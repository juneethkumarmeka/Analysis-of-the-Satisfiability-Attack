module basic_1500_15000_2000_60_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_169,In_129);
nor U1 (N_1,In_481,In_749);
nor U2 (N_2,In_1119,In_159);
nand U3 (N_3,In_50,In_629);
or U4 (N_4,In_820,In_844);
or U5 (N_5,In_176,In_236);
nand U6 (N_6,In_177,In_367);
nand U7 (N_7,In_632,In_317);
nand U8 (N_8,In_153,In_1372);
nand U9 (N_9,In_566,In_1082);
or U10 (N_10,In_433,In_1476);
or U11 (N_11,In_1202,In_982);
or U12 (N_12,In_349,In_826);
xnor U13 (N_13,In_1175,In_1263);
or U14 (N_14,In_376,In_978);
nand U15 (N_15,In_1313,In_1214);
nand U16 (N_16,In_1147,In_1089);
and U17 (N_17,In_839,In_81);
and U18 (N_18,In_797,In_1254);
xor U19 (N_19,In_574,In_567);
nand U20 (N_20,In_54,In_1209);
xnor U21 (N_21,In_1019,In_1468);
or U22 (N_22,In_965,In_1397);
xnor U23 (N_23,In_465,In_833);
and U24 (N_24,In_1279,In_945);
xnor U25 (N_25,In_323,In_843);
nand U26 (N_26,In_1003,In_1422);
nor U27 (N_27,In_411,In_640);
nor U28 (N_28,In_441,In_848);
nor U29 (N_29,In_480,In_538);
nor U30 (N_30,In_908,In_1086);
nor U31 (N_31,In_522,In_36);
or U32 (N_32,In_466,In_1434);
xor U33 (N_33,In_901,In_1233);
or U34 (N_34,In_1290,In_883);
nand U35 (N_35,In_320,In_535);
xor U36 (N_36,In_609,In_943);
or U37 (N_37,In_920,In_1009);
and U38 (N_38,In_489,In_205);
nor U39 (N_39,In_1429,In_836);
xor U40 (N_40,In_854,In_1135);
or U41 (N_41,In_744,In_188);
and U42 (N_42,In_1107,In_1098);
and U43 (N_43,In_692,In_275);
or U44 (N_44,In_456,In_1421);
and U45 (N_45,In_711,In_1469);
nand U46 (N_46,In_1002,In_459);
nand U47 (N_47,In_1121,In_707);
xnor U48 (N_48,In_404,In_1229);
and U49 (N_49,In_1317,In_528);
xor U50 (N_50,In_450,In_703);
and U51 (N_51,In_520,In_336);
xor U52 (N_52,In_1159,In_880);
xor U53 (N_53,In_1172,In_1428);
and U54 (N_54,In_789,In_1287);
xor U55 (N_55,In_612,In_95);
xor U56 (N_56,In_56,In_951);
nand U57 (N_57,In_1437,In_1387);
nor U58 (N_58,In_1327,In_1430);
xor U59 (N_59,In_669,In_577);
and U60 (N_60,In_38,In_948);
xor U61 (N_61,In_1194,In_407);
nor U62 (N_62,In_286,In_333);
and U63 (N_63,In_495,In_135);
and U64 (N_64,In_1027,In_1017);
or U65 (N_65,In_858,In_718);
or U66 (N_66,In_655,In_545);
xor U67 (N_67,In_397,In_1099);
and U68 (N_68,In_351,In_1111);
nor U69 (N_69,In_1205,In_1376);
and U70 (N_70,In_925,In_1261);
or U71 (N_71,In_1226,In_121);
nand U72 (N_72,In_1120,In_1459);
xnor U73 (N_73,In_537,In_1191);
or U74 (N_74,In_1173,In_1222);
nand U75 (N_75,In_1289,In_675);
nand U76 (N_76,In_379,In_1143);
xnor U77 (N_77,In_746,In_1303);
xor U78 (N_78,In_136,In_686);
nand U79 (N_79,In_105,In_932);
nor U80 (N_80,In_97,In_953);
xnor U81 (N_81,In_1240,In_904);
or U82 (N_82,In_1338,In_735);
xnor U83 (N_83,In_506,In_6);
and U84 (N_84,In_147,In_164);
and U85 (N_85,In_521,In_776);
or U86 (N_86,In_621,In_579);
or U87 (N_87,In_699,In_671);
xor U88 (N_88,In_610,In_238);
nand U89 (N_89,In_1088,In_788);
and U90 (N_90,In_467,In_190);
nor U91 (N_91,In_192,In_946);
or U92 (N_92,In_479,In_1127);
xnor U93 (N_93,In_1132,In_1249);
and U94 (N_94,In_391,In_1040);
xnor U95 (N_95,In_1420,In_60);
and U96 (N_96,In_700,In_1235);
xnor U97 (N_97,In_1139,In_211);
nand U98 (N_98,In_1217,In_1395);
nand U99 (N_99,In_791,In_1371);
or U100 (N_100,In_879,In_1273);
and U101 (N_101,In_209,In_1238);
nand U102 (N_102,In_674,In_305);
nor U103 (N_103,In_261,In_794);
and U104 (N_104,In_175,In_1031);
and U105 (N_105,In_432,In_19);
xor U106 (N_106,In_603,In_1267);
xnor U107 (N_107,In_1131,In_738);
or U108 (N_108,In_1444,In_98);
nor U109 (N_109,In_65,In_1188);
or U110 (N_110,In_654,In_770);
xnor U111 (N_111,In_39,In_831);
and U112 (N_112,In_853,In_445);
nor U113 (N_113,In_322,In_48);
or U114 (N_114,In_751,In_146);
and U115 (N_115,In_1025,In_203);
nand U116 (N_116,In_607,In_1396);
xnor U117 (N_117,In_1315,In_386);
xnor U118 (N_118,In_499,In_431);
nor U119 (N_119,In_1283,In_130);
or U120 (N_120,In_548,In_841);
xor U121 (N_121,In_1299,In_464);
or U122 (N_122,In_1304,In_393);
nor U123 (N_123,In_334,In_846);
nand U124 (N_124,In_1220,In_1087);
nor U125 (N_125,In_424,In_102);
and U126 (N_126,In_174,In_315);
xor U127 (N_127,In_570,In_55);
nor U128 (N_128,In_817,In_240);
and U129 (N_129,In_387,In_444);
nor U130 (N_130,In_716,In_1265);
nor U131 (N_131,In_1018,In_1481);
nand U132 (N_132,In_1416,In_443);
and U133 (N_133,In_1309,In_1130);
or U134 (N_134,In_62,In_803);
or U135 (N_135,In_768,In_217);
nand U136 (N_136,In_808,In_111);
and U137 (N_137,In_819,In_1195);
or U138 (N_138,In_1340,In_1016);
or U139 (N_139,In_891,In_1106);
nand U140 (N_140,In_394,In_872);
nand U141 (N_141,In_878,In_1065);
or U142 (N_142,In_1206,In_1180);
and U143 (N_143,In_440,In_1403);
or U144 (N_144,In_42,In_257);
xnor U145 (N_145,In_723,In_357);
xor U146 (N_146,In_611,In_1163);
and U147 (N_147,In_1433,In_596);
or U148 (N_148,In_952,In_1271);
or U149 (N_149,In_682,In_701);
nor U150 (N_150,In_1241,In_270);
nand U151 (N_151,In_578,In_1346);
nand U152 (N_152,In_643,In_1436);
and U153 (N_153,In_77,In_656);
nand U154 (N_154,In_1140,In_1350);
xnor U155 (N_155,In_1490,In_985);
nor U156 (N_156,In_1208,In_714);
nand U157 (N_157,In_668,In_156);
and U158 (N_158,In_615,In_970);
nand U159 (N_159,In_1394,In_933);
nor U160 (N_160,In_99,In_900);
nand U161 (N_161,In_672,In_1076);
and U162 (N_162,In_267,In_804);
nand U163 (N_163,In_491,In_1248);
nor U164 (N_164,In_1015,In_868);
xnor U165 (N_165,In_204,In_1224);
or U166 (N_166,In_902,In_1473);
and U167 (N_167,In_488,In_1198);
nor U168 (N_168,In_116,In_1496);
xor U169 (N_169,In_1186,In_928);
and U170 (N_170,In_760,In_273);
and U171 (N_171,In_995,In_594);
or U172 (N_172,In_1440,In_127);
or U173 (N_173,In_106,In_1013);
nor U174 (N_174,In_182,In_743);
or U175 (N_175,In_131,In_123);
or U176 (N_176,In_1487,In_1425);
xnor U177 (N_177,In_1041,In_758);
nor U178 (N_178,In_696,In_592);
nor U179 (N_179,In_899,In_79);
or U180 (N_180,In_328,In_892);
nor U181 (N_181,In_1413,In_1442);
or U182 (N_182,In_335,In_597);
or U183 (N_183,In_677,In_1390);
or U184 (N_184,In_608,In_547);
nand U185 (N_185,In_816,In_867);
nand U186 (N_186,In_1184,In_490);
xnor U187 (N_187,In_581,In_416);
nor U188 (N_188,In_454,In_1407);
nor U189 (N_189,In_1161,In_1453);
and U190 (N_190,In_1204,In_500);
nand U191 (N_191,In_777,In_893);
nand U192 (N_192,In_828,In_926);
xor U193 (N_193,In_229,In_341);
nand U194 (N_194,In_1492,In_1200);
xor U195 (N_195,In_231,In_1450);
nand U196 (N_196,In_825,In_1439);
or U197 (N_197,In_120,In_967);
or U198 (N_198,In_691,In_365);
and U199 (N_199,In_565,In_1028);
and U200 (N_200,In_1103,In_258);
and U201 (N_201,In_142,In_401);
and U202 (N_202,In_1477,In_207);
nand U203 (N_203,In_830,In_991);
and U204 (N_204,In_1034,In_245);
nor U205 (N_205,In_1068,In_425);
or U206 (N_206,In_1322,In_278);
nand U207 (N_207,In_75,In_251);
xor U208 (N_208,In_216,In_1007);
or U209 (N_209,In_719,In_1398);
or U210 (N_210,In_1149,In_307);
or U211 (N_211,In_1314,In_929);
xor U212 (N_212,In_637,In_1320);
xnor U213 (N_213,In_318,In_1457);
nor U214 (N_214,In_999,In_802);
or U215 (N_215,In_1482,In_1153);
xnor U216 (N_216,In_252,In_1443);
xor U217 (N_217,In_1093,In_1237);
nor U218 (N_218,In_230,In_300);
nand U219 (N_219,In_755,In_1032);
nor U220 (N_220,In_296,In_327);
nor U221 (N_221,In_1069,In_697);
or U222 (N_222,In_473,In_171);
nor U223 (N_223,In_1334,In_223);
xor U224 (N_224,In_96,In_1293);
nand U225 (N_225,In_587,In_745);
or U226 (N_226,In_882,In_14);
nor U227 (N_227,In_232,In_224);
nand U228 (N_228,In_1047,In_189);
and U229 (N_229,In_1268,In_160);
nand U230 (N_230,In_126,In_453);
nand U231 (N_231,In_717,In_1344);
xor U232 (N_232,In_1242,In_362);
or U233 (N_233,In_779,In_1401);
nand U234 (N_234,In_646,In_1102);
nor U235 (N_235,In_875,In_1022);
xor U236 (N_236,In_344,In_364);
or U237 (N_237,In_255,In_1004);
xor U238 (N_238,In_1369,In_818);
nand U239 (N_239,In_811,In_927);
nand U240 (N_240,In_1014,In_477);
or U241 (N_241,In_1462,In_361);
xnor U242 (N_242,In_100,In_1185);
xnor U243 (N_243,In_666,In_782);
and U244 (N_244,In_526,In_731);
xnor U245 (N_245,In_931,In_475);
nand U246 (N_246,In_748,In_753);
and U247 (N_247,In_1187,In_213);
or U248 (N_248,In_1272,In_447);
xor U249 (N_249,In_516,In_468);
or U250 (N_250,In_599,In_604);
nand U251 (N_251,In_1419,N_110);
xor U252 (N_252,In_1495,In_630);
or U253 (N_253,In_876,In_101);
nand U254 (N_254,In_856,N_237);
nor U255 (N_255,In_1463,In_1389);
nor U256 (N_256,In_76,In_180);
xnor U257 (N_257,In_863,In_486);
or U258 (N_258,In_1405,In_1499);
nand U259 (N_259,N_66,In_4);
nand U260 (N_260,In_1228,In_1382);
or U261 (N_261,In_837,In_134);
and U262 (N_262,In_1251,In_256);
nor U263 (N_263,In_1232,In_747);
nor U264 (N_264,N_107,In_63);
nor U265 (N_265,In_527,In_1005);
nand U266 (N_266,In_137,In_984);
nor U267 (N_267,In_72,In_981);
nand U268 (N_268,In_874,In_415);
nor U269 (N_269,In_138,In_128);
xnor U270 (N_270,In_685,In_451);
or U271 (N_271,In_993,In_990);
nor U272 (N_272,In_304,In_469);
xor U273 (N_273,N_94,In_253);
nor U274 (N_274,N_159,In_1213);
nor U275 (N_275,In_762,In_822);
nor U276 (N_276,In_1400,In_268);
nand U277 (N_277,In_800,In_530);
xor U278 (N_278,In_898,In_237);
nand U279 (N_279,In_1308,In_83);
or U280 (N_280,N_135,N_34);
xor U281 (N_281,N_147,In_613);
and U282 (N_282,N_62,N_52);
xnor U283 (N_283,In_1292,In_1033);
nor U284 (N_284,In_695,In_1455);
and U285 (N_285,In_1277,In_1138);
xor U286 (N_286,In_556,In_555);
and U287 (N_287,In_657,In_403);
and U288 (N_288,In_678,N_55);
nand U289 (N_289,N_198,In_264);
nand U290 (N_290,In_661,In_702);
or U291 (N_291,In_1115,In_271);
or U292 (N_292,In_940,N_132);
xnor U293 (N_293,In_1052,In_1438);
nor U294 (N_294,In_954,In_1474);
or U295 (N_295,N_223,In_40);
nor U296 (N_296,In_560,N_56);
nand U297 (N_297,In_1297,In_600);
xor U298 (N_298,N_57,In_1449);
or U299 (N_299,In_312,In_266);
or U300 (N_300,N_42,In_1423);
and U301 (N_301,N_178,N_152);
xnor U302 (N_302,In_618,In_1286);
or U303 (N_303,In_684,In_504);
and U304 (N_304,N_32,In_68);
nor U305 (N_305,N_170,In_324);
nor U306 (N_306,In_647,In_793);
or U307 (N_307,N_74,In_1255);
and U308 (N_308,In_1178,In_569);
xor U309 (N_309,In_482,In_293);
xor U310 (N_310,In_25,N_114);
xor U311 (N_311,In_1046,In_616);
and U312 (N_312,In_1116,N_99);
and U313 (N_313,In_992,In_122);
nor U314 (N_314,In_653,In_1036);
nand U315 (N_315,In_154,In_80);
or U316 (N_316,In_1456,N_122);
and U317 (N_317,In_420,In_413);
nor U318 (N_318,In_774,In_704);
nand U319 (N_319,In_887,In_1260);
or U320 (N_320,In_90,In_82);
nand U321 (N_321,In_1037,In_325);
or U322 (N_322,N_164,In_15);
or U323 (N_323,In_438,In_1384);
xnor U324 (N_324,In_1417,In_1243);
and U325 (N_325,In_601,In_1108);
xor U326 (N_326,In_241,In_358);
nor U327 (N_327,In_29,In_452);
nand U328 (N_328,In_370,In_114);
xor U329 (N_329,In_1152,In_173);
nand U330 (N_330,N_91,In_886);
or U331 (N_331,In_792,In_107);
nand U332 (N_332,In_1051,In_140);
nor U333 (N_333,In_1458,N_240);
nand U334 (N_334,In_1104,In_1259);
xnor U335 (N_335,N_234,N_150);
or U336 (N_336,In_249,In_476);
and U337 (N_337,In_20,In_92);
and U338 (N_338,In_834,N_28);
xnor U339 (N_339,In_1321,In_859);
xnor U340 (N_340,In_149,In_460);
or U341 (N_341,In_119,N_156);
nor U342 (N_342,N_127,In_1060);
xor U343 (N_343,In_561,In_551);
xor U344 (N_344,In_1118,In_1262);
nor U345 (N_345,In_557,In_1083);
nand U346 (N_346,In_124,In_484);
nand U347 (N_347,N_137,In_340);
nand U348 (N_348,In_1181,In_503);
or U349 (N_349,In_225,In_780);
or U350 (N_350,In_956,In_923);
nor U351 (N_351,In_912,N_165);
and U352 (N_352,In_1381,N_65);
nor U353 (N_353,In_1480,In_1276);
nand U354 (N_354,In_191,In_1168);
or U355 (N_355,N_0,N_85);
nand U356 (N_356,In_1300,N_199);
and U357 (N_357,In_442,In_1049);
nand U358 (N_358,In_1472,In_568);
and U359 (N_359,In_1353,In_2);
nand U360 (N_360,N_43,N_11);
xnor U361 (N_361,In_785,In_513);
xor U362 (N_362,In_22,In_645);
and U363 (N_363,N_44,N_160);
and U364 (N_364,N_14,In_588);
nor U365 (N_365,In_517,In_64);
nor U366 (N_366,N_195,N_131);
nand U367 (N_367,N_49,In_247);
nor U368 (N_368,In_32,In_950);
nor U369 (N_369,In_890,In_1427);
nand U370 (N_370,In_1144,N_202);
xor U371 (N_371,N_50,In_771);
and U372 (N_372,N_88,In_91);
nand U373 (N_373,In_812,N_196);
or U374 (N_374,In_761,In_11);
xor U375 (N_375,In_742,N_16);
or U376 (N_376,N_17,In_352);
and U377 (N_377,In_497,In_1001);
nor U378 (N_378,In_418,In_409);
or U379 (N_379,In_961,N_182);
nor U380 (N_380,In_732,In_69);
nor U381 (N_381,In_463,In_1404);
and U382 (N_382,In_110,In_1365);
and U383 (N_383,In_1484,In_881);
or U384 (N_384,In_1329,In_784);
and U385 (N_385,In_103,In_1162);
or U386 (N_386,In_1445,N_133);
nor U387 (N_387,In_642,N_232);
or U388 (N_388,N_245,In_509);
and U389 (N_389,In_221,N_70);
and U390 (N_390,In_41,N_116);
and U391 (N_391,In_1351,In_1364);
and U392 (N_392,In_44,In_1377);
or U393 (N_393,In_1379,N_244);
nand U394 (N_394,N_181,In_1325);
nand U395 (N_395,In_455,In_1171);
xnor U396 (N_396,In_319,In_806);
xor U397 (N_397,In_1335,N_3);
xor U398 (N_398,N_15,In_1045);
xnor U399 (N_399,In_977,In_783);
nand U400 (N_400,In_1418,In_373);
or U401 (N_401,In_542,In_829);
nor U402 (N_402,In_1091,In_1446);
or U403 (N_403,In_243,In_1124);
nand U404 (N_404,In_814,In_641);
xnor U405 (N_405,In_421,In_515);
nor U406 (N_406,In_1,In_824);
nor U407 (N_407,In_550,N_126);
nand U408 (N_408,N_4,In_1101);
nand U409 (N_409,In_1141,In_583);
or U410 (N_410,In_1337,N_38);
nand U411 (N_411,N_25,In_860);
nor U412 (N_412,In_45,In_877);
and U413 (N_413,In_59,In_924);
xnor U414 (N_414,In_1062,In_638);
or U415 (N_415,In_219,In_1012);
or U416 (N_416,In_888,In_385);
nand U417 (N_417,In_576,In_966);
nand U418 (N_418,In_1189,N_228);
nor U419 (N_419,In_28,N_151);
nand U420 (N_420,N_77,In_586);
or U421 (N_421,In_295,N_247);
or U422 (N_422,In_861,In_400);
nand U423 (N_423,In_690,In_781);
or U424 (N_424,In_1385,In_1134);
xor U425 (N_425,In_786,In_1183);
and U426 (N_426,In_1154,In_619);
nand U427 (N_427,In_1368,N_75);
nor U428 (N_428,N_73,In_58);
nor U429 (N_429,In_360,In_1230);
nor U430 (N_430,In_93,In_301);
nor U431 (N_431,In_1215,N_226);
xnor U432 (N_432,N_96,N_138);
nor U433 (N_433,N_171,In_1170);
xor U434 (N_434,In_302,In_1231);
nand U435 (N_435,In_562,In_1146);
and U436 (N_436,In_754,N_142);
xnor U437 (N_437,In_1157,N_189);
xor U438 (N_438,In_85,In_964);
and U439 (N_439,In_390,In_185);
and U440 (N_440,In_1478,In_1362);
nand U441 (N_441,N_201,In_265);
nor U442 (N_442,In_787,In_572);
nor U443 (N_443,In_673,N_30);
or U444 (N_444,N_162,In_329);
or U445 (N_445,In_290,N_174);
nor U446 (N_446,In_331,N_145);
nand U447 (N_447,N_89,In_84);
xor U448 (N_448,In_429,In_614);
and U449 (N_449,N_184,N_105);
xor U450 (N_450,In_809,In_272);
nor U451 (N_451,In_620,N_194);
or U452 (N_452,In_889,N_168);
or U453 (N_453,In_683,N_141);
or U454 (N_454,N_37,In_1498);
or U455 (N_455,In_847,In_1126);
nand U456 (N_456,In_326,In_382);
xnor U457 (N_457,N_153,In_1406);
nor U458 (N_458,In_1466,In_492);
and U459 (N_459,In_531,N_54);
and U460 (N_460,In_573,In_33);
xnor U461 (N_461,In_435,In_470);
or U462 (N_462,N_1,N_120);
nand U463 (N_463,In_9,In_1448);
nor U464 (N_464,In_1029,In_845);
and U465 (N_465,In_355,In_410);
nand U466 (N_466,In_549,In_1288);
nand U467 (N_467,In_197,In_1465);
or U468 (N_468,N_224,In_1079);
nor U469 (N_469,In_795,In_502);
or U470 (N_470,N_108,In_1359);
and U471 (N_471,In_380,In_869);
and U472 (N_472,N_59,N_112);
nor U473 (N_473,In_1113,In_1447);
xnor U474 (N_474,N_61,In_46);
and U475 (N_475,In_388,In_282);
or U476 (N_476,In_1485,In_35);
or U477 (N_477,In_752,In_1212);
nor U478 (N_478,In_449,In_915);
and U479 (N_479,In_1136,In_917);
or U480 (N_480,In_832,In_763);
xor U481 (N_481,N_41,In_728);
or U482 (N_482,In_1123,In_870);
nand U483 (N_483,In_1285,N_193);
nor U484 (N_484,N_179,In_448);
nand U485 (N_485,In_941,In_1316);
xor U486 (N_486,In_1302,In_838);
nand U487 (N_487,In_18,In_1333);
or U488 (N_488,In_1301,In_494);
and U489 (N_489,In_523,In_1030);
nor U490 (N_490,N_212,In_26);
nand U491 (N_491,In_61,In_1479);
or U492 (N_492,In_766,In_417);
and U493 (N_493,In_938,N_104);
and U494 (N_494,In_1408,In_698);
or U495 (N_495,N_233,In_1071);
xor U496 (N_496,In_1190,In_1244);
nor U497 (N_497,In_478,In_143);
xor U498 (N_498,In_1151,In_1169);
xnor U499 (N_499,In_172,In_1460);
and U500 (N_500,In_212,N_436);
nor U501 (N_501,In_636,N_238);
nand U502 (N_502,In_1357,In_162);
nor U503 (N_503,In_342,In_206);
nand U504 (N_504,N_251,N_287);
nand U505 (N_505,N_230,In_215);
xor U506 (N_506,In_125,N_470);
nand U507 (N_507,In_399,In_118);
xor U508 (N_508,N_420,N_190);
or U509 (N_509,In_263,In_897);
and U510 (N_510,N_465,N_403);
xnor U511 (N_511,In_835,In_1216);
or U512 (N_512,In_1039,In_593);
nor U513 (N_513,N_488,In_733);
nand U514 (N_514,In_726,In_906);
nand U515 (N_515,N_314,In_1192);
xor U516 (N_516,N_98,N_321);
and U517 (N_517,In_1343,In_885);
or U518 (N_518,In_1218,N_483);
nor U519 (N_519,N_119,In_884);
xor U520 (N_520,N_33,N_329);
nand U521 (N_521,In_582,In_1061);
or U522 (N_522,In_759,In_815);
nor U523 (N_523,In_181,In_740);
nand U524 (N_524,In_1275,N_29);
nor U525 (N_525,In_648,In_1392);
xnor U526 (N_526,In_1166,In_345);
or U527 (N_527,N_291,In_1258);
nor U528 (N_528,In_756,In_396);
or U529 (N_529,In_1057,In_163);
nand U530 (N_530,N_395,N_39);
or U531 (N_531,In_485,N_315);
xnor U532 (N_532,In_1239,In_337);
xnor U533 (N_533,N_426,In_617);
nand U534 (N_534,In_1278,N_454);
or U535 (N_535,N_274,N_296);
nor U536 (N_536,In_729,N_469);
nor U537 (N_537,In_1158,N_6);
nor U538 (N_538,In_178,In_1486);
and U539 (N_539,N_47,N_266);
or U540 (N_540,In_919,In_1210);
and U541 (N_541,In_974,In_406);
xor U542 (N_542,In_1328,In_1145);
nor U543 (N_543,In_117,In_1182);
nor U544 (N_544,In_983,N_23);
xnor U545 (N_545,In_1280,N_373);
nor U546 (N_546,In_168,In_1035);
nand U547 (N_547,In_372,In_1354);
nor U548 (N_548,In_1080,In_235);
and U549 (N_549,In_152,In_259);
nand U550 (N_550,In_1373,In_827);
and U551 (N_551,In_1411,N_197);
nor U552 (N_552,N_412,In_1264);
xor U553 (N_553,In_540,N_326);
and U554 (N_554,N_388,N_9);
nor U555 (N_555,In_939,N_111);
and U556 (N_556,N_468,In_43);
xnor U557 (N_557,In_13,In_710);
or U558 (N_558,N_496,N_269);
and U559 (N_559,N_18,N_379);
nand U560 (N_560,In_1042,In_662);
nand U561 (N_561,In_1305,N_21);
xnor U562 (N_562,N_338,In_930);
nor U563 (N_563,In_622,In_348);
and U564 (N_564,N_235,N_279);
nand U565 (N_565,N_248,In_947);
nor U566 (N_566,N_271,In_313);
nand U567 (N_567,N_441,N_290);
nor U568 (N_568,In_1410,N_313);
or U569 (N_569,In_1077,In_254);
and U570 (N_570,N_414,In_1094);
nand U571 (N_571,In_546,N_167);
nand U572 (N_572,In_1330,N_437);
or U573 (N_573,In_1341,In_676);
or U574 (N_574,In_1281,N_183);
nor U575 (N_575,In_658,In_969);
xnor U576 (N_576,In_1043,In_1375);
nor U577 (N_577,N_19,N_71);
nand U578 (N_578,N_87,In_1227);
xor U579 (N_579,In_1399,N_413);
xor U580 (N_580,In_74,In_730);
and U581 (N_581,N_451,N_217);
nor U582 (N_582,N_487,N_5);
or U583 (N_583,In_419,In_659);
nand U584 (N_584,In_725,In_292);
xnor U585 (N_585,In_1073,In_715);
or U586 (N_586,N_374,N_166);
or U587 (N_587,In_228,In_487);
and U588 (N_588,In_591,In_306);
nor U589 (N_589,In_155,In_375);
and U590 (N_590,N_316,N_270);
nor U591 (N_591,N_173,N_227);
or U592 (N_592,In_1252,N_434);
and U593 (N_593,N_79,In_1020);
or U594 (N_594,N_443,N_163);
or U595 (N_595,In_1000,In_849);
xnor U596 (N_596,In_505,In_1058);
or U597 (N_597,In_554,N_439);
and U598 (N_598,In_89,N_448);
nor U599 (N_599,N_67,In_519);
or U600 (N_600,N_333,In_598);
and U601 (N_601,In_736,In_558);
and U602 (N_602,N_7,In_1360);
nor U603 (N_603,In_458,In_427);
and U604 (N_604,N_433,In_986);
nand U605 (N_605,In_1038,In_1174);
nor U606 (N_606,In_1125,In_381);
or U607 (N_607,N_347,In_979);
and U608 (N_608,In_1349,In_165);
nor U609 (N_609,N_423,In_532);
nor U610 (N_610,N_380,In_1110);
nor U611 (N_611,In_1269,N_10);
or U612 (N_612,N_298,In_687);
or U613 (N_613,In_706,In_712);
xor U614 (N_614,N_268,N_396);
and U615 (N_615,In_1312,N_486);
or U616 (N_616,In_132,N_429);
xor U617 (N_617,In_807,In_553);
nor U618 (N_618,N_304,N_339);
nor U619 (N_619,In_210,In_667);
nand U620 (N_620,In_144,N_489);
or U621 (N_621,N_331,N_458);
xor U622 (N_622,N_12,In_790);
nor U623 (N_623,In_1493,In_963);
and U624 (N_624,N_356,In_741);
and U625 (N_625,N_72,N_214);
xor U626 (N_626,In_1055,N_250);
nand U627 (N_627,In_1483,In_279);
xor U628 (N_628,In_474,In_356);
or U629 (N_629,In_511,In_1105);
xnor U630 (N_630,In_1008,N_325);
xor U631 (N_631,In_628,N_13);
and U632 (N_632,N_282,N_130);
xor U633 (N_633,N_300,In_193);
xor U634 (N_634,N_421,In_508);
and U635 (N_635,In_1295,In_1246);
xor U636 (N_636,N_490,In_778);
xor U637 (N_637,In_308,N_491);
or U638 (N_638,In_705,N_422);
nor U639 (N_639,In_1415,N_80);
or U640 (N_640,In_821,In_737);
xnor U641 (N_641,In_0,N_272);
and U642 (N_642,N_376,N_352);
xnor U643 (N_643,N_260,N_479);
or U644 (N_644,N_208,In_8);
xnor U645 (N_645,N_215,In_595);
or U646 (N_646,N_364,In_1414);
nor U647 (N_647,In_1488,In_1156);
or U648 (N_648,N_319,In_727);
nor U649 (N_649,In_1177,N_341);
nand U650 (N_650,N_115,In_1494);
and U651 (N_651,N_146,In_757);
xnor U652 (N_652,In_294,N_450);
xor U653 (N_653,N_340,N_424);
or U654 (N_654,N_95,N_209);
xnor U655 (N_655,In_1137,In_1096);
xnor U656 (N_656,In_86,N_385);
xnor U657 (N_657,In_47,In_1196);
or U658 (N_658,N_58,In_1201);
xnor U659 (N_659,N_481,N_359);
xnor U660 (N_660,In_1355,In_383);
and U661 (N_661,In_1050,N_474);
nand U662 (N_662,In_775,N_493);
or U663 (N_663,In_1356,N_323);
nor U664 (N_664,N_348,N_264);
nand U665 (N_665,In_274,N_457);
nor U666 (N_666,In_430,N_461);
nand U667 (N_667,In_1374,N_68);
nand U668 (N_668,N_308,N_447);
and U669 (N_669,In_670,In_525);
nor U670 (N_670,In_31,In_1363);
and U671 (N_671,In_765,In_631);
and U672 (N_672,In_1461,N_206);
or U673 (N_673,In_1342,N_53);
nand U674 (N_674,In_650,N_499);
and U675 (N_675,N_464,In_1176);
nor U676 (N_676,In_585,In_1165);
xor U677 (N_677,N_497,In_1225);
and U678 (N_678,In_354,In_493);
or U679 (N_679,In_720,N_295);
and U680 (N_680,N_303,In_1253);
nor U681 (N_681,In_1307,N_459);
xor U682 (N_682,In_1072,In_1367);
nand U683 (N_683,In_496,N_117);
nand U684 (N_684,In_1179,In_303);
nor U685 (N_685,In_321,In_66);
and U686 (N_686,N_309,In_851);
or U687 (N_687,N_344,In_1431);
or U688 (N_688,N_20,In_1409);
xnor U689 (N_689,N_498,In_1270);
or U690 (N_690,In_510,N_123);
and U691 (N_691,N_176,N_350);
nor U692 (N_692,In_246,In_694);
nor U693 (N_693,In_434,In_12);
or U694 (N_694,N_97,In_289);
xnor U695 (N_695,In_1024,N_361);
nor U696 (N_696,In_1282,In_1245);
and U697 (N_697,In_1336,In_810);
xnor U698 (N_698,In_284,N_252);
nor U699 (N_699,In_1059,N_273);
or U700 (N_700,N_106,In_260);
xor U701 (N_701,In_639,N_328);
and U702 (N_702,In_1310,In_108);
nor U703 (N_703,N_431,N_349);
and U704 (N_704,In_1348,In_208);
nand U705 (N_705,In_1053,N_369);
nand U706 (N_706,N_229,In_1211);
nand U707 (N_707,In_71,In_199);
nand U708 (N_708,N_203,In_864);
nand U709 (N_709,N_192,In_49);
nor U710 (N_710,In_437,N_255);
and U711 (N_711,In_51,In_428);
nand U712 (N_712,In_571,In_145);
and U713 (N_713,N_299,In_739);
and U714 (N_714,N_31,N_257);
nor U715 (N_715,In_862,N_456);
and U716 (N_716,N_261,In_625);
nor U717 (N_717,In_141,N_121);
xor U718 (N_718,N_406,In_1084);
xor U719 (N_719,N_204,In_813);
and U720 (N_720,N_210,In_1221);
xnor U721 (N_721,N_154,N_337);
nand U722 (N_722,N_35,N_382);
xor U723 (N_723,N_430,In_971);
and U724 (N_724,In_1133,In_1067);
xnor U725 (N_725,N_124,In_989);
nor U726 (N_726,In_626,In_347);
and U727 (N_727,N_219,In_34);
nor U728 (N_728,N_2,In_242);
nand U729 (N_729,N_259,In_183);
nor U730 (N_730,N_311,N_418);
nand U731 (N_731,In_1274,In_994);
or U732 (N_732,In_297,N_317);
nor U733 (N_733,N_327,In_1100);
nand U734 (N_734,In_1266,In_1366);
nand U735 (N_735,N_307,N_372);
xor U736 (N_736,N_363,N_370);
nand U737 (N_737,N_297,In_799);
and U738 (N_738,N_267,In_280);
xnor U739 (N_739,In_436,In_529);
xnor U740 (N_740,N_410,In_10);
nor U741 (N_741,N_139,In_187);
and U742 (N_742,In_363,N_22);
nand U743 (N_743,N_249,In_944);
xnor U744 (N_744,In_801,In_405);
nand U745 (N_745,In_514,N_51);
xnor U746 (N_746,In_291,N_281);
nand U747 (N_747,In_1339,In_378);
xor U748 (N_748,N_367,N_289);
nand U749 (N_749,N_478,In_895);
or U750 (N_750,In_709,In_559);
nand U751 (N_751,N_158,N_666);
nor U752 (N_752,In_457,In_1306);
or U753 (N_753,N_473,N_471);
nor U754 (N_754,N_276,N_646);
or U755 (N_755,N_543,N_482);
xor U756 (N_756,N_129,In_412);
nor U757 (N_757,In_972,N_393);
or U758 (N_758,In_17,N_546);
xnor U759 (N_759,In_823,In_57);
nand U760 (N_760,N_686,In_1155);
nor U761 (N_761,In_563,In_934);
and U762 (N_762,In_909,In_1081);
nor U763 (N_763,In_1435,In_606);
nor U764 (N_764,N_571,In_439);
nor U765 (N_765,In_196,N_650);
or U766 (N_766,N_405,N_712);
xor U767 (N_767,N_324,N_90);
nand U768 (N_768,N_216,N_501);
nor U769 (N_769,N_143,In_1426);
xor U770 (N_770,N_632,In_772);
or U771 (N_771,In_350,In_894);
or U772 (N_772,In_635,N_647);
and U773 (N_773,N_662,N_607);
or U774 (N_774,N_665,In_624);
or U775 (N_775,N_627,N_207);
and U776 (N_776,N_351,N_649);
nor U777 (N_777,In_767,N_185);
and U778 (N_778,In_30,N_618);
nor U779 (N_779,In_52,In_366);
xnor U780 (N_780,N_368,N_221);
and U781 (N_781,In_976,N_528);
nor U782 (N_782,N_582,N_577);
or U783 (N_783,N_449,N_444);
nor U784 (N_784,In_959,N_655);
xnor U785 (N_785,N_318,N_394);
and U786 (N_786,In_644,In_589);
and U787 (N_787,N_617,N_705);
or U788 (N_788,N_508,N_504);
or U789 (N_789,N_552,In_1386);
or U790 (N_790,In_330,In_214);
or U791 (N_791,In_53,N_541);
or U792 (N_792,N_566,N_626);
or U793 (N_793,N_572,In_871);
nor U794 (N_794,N_463,N_453);
and U795 (N_795,N_730,In_239);
and U796 (N_796,N_644,N_715);
nand U797 (N_797,N_494,N_84);
xnor U798 (N_798,N_693,N_125);
and U799 (N_799,N_397,N_696);
nor U800 (N_800,N_749,N_518);
nor U801 (N_801,N_664,N_467);
and U802 (N_802,N_222,N_428);
or U803 (N_803,In_713,N_708);
nor U804 (N_804,N_681,N_731);
nor U805 (N_805,In_518,In_907);
xnor U806 (N_806,In_1109,In_359);
or U807 (N_807,In_1491,N_719);
nor U808 (N_808,In_166,In_903);
nand U809 (N_809,In_688,In_1451);
xor U810 (N_810,In_660,In_133);
xnor U811 (N_811,In_534,In_220);
and U812 (N_812,N_254,N_375);
xor U813 (N_813,In_1128,N_220);
and U814 (N_814,N_477,N_522);
xnor U815 (N_815,N_524,In_314);
xnor U816 (N_816,In_1378,In_1074);
nor U817 (N_817,In_988,N_728);
nor U818 (N_818,N_435,In_1223);
or U819 (N_819,N_677,N_625);
and U820 (N_820,In_805,In_369);
nor U821 (N_821,In_921,In_461);
and U822 (N_822,In_652,In_1010);
nor U823 (N_823,N_113,In_408);
or U824 (N_824,In_368,In_507);
xnor U825 (N_825,In_1464,In_922);
and U826 (N_826,N_511,In_1412);
nand U827 (N_827,In_769,N_265);
or U828 (N_828,N_415,N_604);
nor U829 (N_829,In_850,N_599);
and U830 (N_830,N_678,N_231);
or U831 (N_831,In_1219,N_515);
nand U832 (N_832,N_455,N_694);
nand U833 (N_833,N_633,In_1284);
nor U834 (N_834,N_614,N_400);
xor U835 (N_835,N_535,N_452);
xor U836 (N_836,N_657,In_262);
nand U837 (N_837,N_398,N_243);
nand U838 (N_838,N_673,N_583);
nor U839 (N_839,N_672,N_623);
and U840 (N_840,N_674,In_1291);
and U841 (N_841,In_269,N_688);
nand U842 (N_842,In_840,In_1054);
nor U843 (N_843,N_134,N_140);
and U844 (N_844,In_1092,In_1326);
nor U845 (N_845,In_299,In_910);
xor U846 (N_846,N_531,N_741);
and U847 (N_847,N_69,N_722);
nor U848 (N_848,N_567,N_258);
nor U849 (N_849,In_285,In_564);
nand U850 (N_850,In_244,N_263);
xor U851 (N_851,In_462,In_1471);
or U852 (N_852,N_520,In_1026);
nand U853 (N_853,In_936,In_1203);
and U854 (N_854,N_36,In_1234);
or U855 (N_855,In_472,In_623);
and U856 (N_856,N_660,In_158);
and U857 (N_857,N_586,In_1298);
nand U858 (N_858,In_958,In_151);
xnor U859 (N_859,In_423,N_46);
or U860 (N_860,N_579,N_485);
or U861 (N_861,In_1311,In_1475);
xor U862 (N_862,N_606,In_842);
xor U863 (N_863,N_527,N_442);
and U864 (N_864,N_559,In_309);
or U865 (N_865,In_1075,N_390);
or U866 (N_866,In_633,N_191);
nor U867 (N_867,N_371,N_747);
xor U868 (N_868,N_149,N_354);
xnor U869 (N_869,N_732,N_615);
xor U870 (N_870,In_250,In_973);
nand U871 (N_871,N_399,In_5);
xnor U872 (N_872,N_48,In_471);
xnor U873 (N_873,N_507,N_517);
nor U874 (N_874,N_695,In_580);
nand U875 (N_875,N_389,In_605);
or U876 (N_876,In_184,N_542);
xnor U877 (N_877,In_426,N_416);
or U878 (N_878,In_584,N_691);
nor U879 (N_879,In_311,In_398);
or U880 (N_880,In_773,In_283);
or U881 (N_881,In_16,N_602);
nand U882 (N_882,N_81,N_480);
nand U883 (N_883,In_316,In_1250);
and U884 (N_884,N_102,N_312);
and U885 (N_885,N_613,N_500);
xnor U886 (N_886,N_534,N_332);
nor U887 (N_887,In_1090,N_659);
or U888 (N_888,In_935,N_570);
xor U889 (N_889,N_701,In_1070);
xnor U890 (N_890,In_281,N_305);
nor U891 (N_891,N_86,N_172);
nor U892 (N_892,N_180,N_539);
xor U893 (N_893,In_1150,N_334);
nor U894 (N_894,In_997,N_663);
or U895 (N_895,In_1112,N_440);
xnor U896 (N_896,In_371,In_501);
xor U897 (N_897,N_603,N_560);
nand U898 (N_898,In_24,In_873);
or U899 (N_899,N_549,N_596);
nor U900 (N_900,N_510,In_201);
xnor U901 (N_901,N_157,In_1023);
and U902 (N_902,N_253,In_298);
and U903 (N_903,N_721,N_60);
nand U904 (N_904,In_1148,N_554);
nor U905 (N_905,N_322,N_432);
and U906 (N_906,N_684,In_1078);
and U907 (N_907,In_112,In_987);
nor U908 (N_908,In_942,In_7);
nand U909 (N_909,In_680,N_611);
xor U910 (N_910,In_708,In_796);
or U911 (N_911,N_636,N_136);
nand U912 (N_912,In_170,N_366);
xnor U913 (N_913,N_144,In_905);
and U914 (N_914,In_913,N_651);
nor U915 (N_915,N_744,In_1021);
xnor U916 (N_916,N_568,In_1324);
nand U917 (N_917,N_360,In_148);
or U918 (N_918,In_1319,In_1296);
xnor U919 (N_919,In_1056,N_652);
nor U920 (N_920,In_218,In_194);
nand U921 (N_921,N_620,N_64);
xor U922 (N_922,In_1391,In_353);
nor U923 (N_923,In_70,In_483);
and U924 (N_924,N_557,N_600);
xor U925 (N_925,In_1402,N_537);
xor U926 (N_926,N_392,N_648);
and U927 (N_927,In_865,In_1380);
nand U928 (N_928,N_357,In_949);
nor U929 (N_929,In_722,N_419);
nand U930 (N_930,In_1048,N_676);
xor U931 (N_931,N_578,In_186);
and U932 (N_932,N_8,N_492);
nand U933 (N_933,In_27,In_94);
xnor U934 (N_934,N_565,In_627);
or U935 (N_935,In_1358,N_538);
and U936 (N_936,N_345,In_649);
nor U937 (N_937,N_362,In_1331);
nor U938 (N_938,In_998,N_532);
xor U939 (N_939,N_573,N_742);
nor U940 (N_940,In_1383,N_225);
or U941 (N_941,In_1294,N_641);
xor U942 (N_942,In_852,N_736);
nand U943 (N_943,In_1063,N_387);
and U944 (N_944,In_1236,In_414);
nand U945 (N_945,N_598,N_280);
nor U946 (N_946,N_525,N_616);
and U947 (N_947,N_355,N_720);
and U948 (N_948,N_161,N_734);
or U949 (N_949,In_1361,N_92);
nand U950 (N_950,N_246,N_735);
nand U951 (N_951,N_169,N_128);
or U952 (N_952,In_346,N_671);
nand U953 (N_953,In_937,In_918);
nand U954 (N_954,In_1117,N_475);
nor U955 (N_955,In_962,N_26);
xnor U956 (N_956,N_188,In_1197);
xor U957 (N_957,N_301,N_292);
or U958 (N_958,N_729,N_306);
xnor U959 (N_959,N_622,N_409);
and U960 (N_960,N_40,N_718);
xnor U961 (N_961,In_960,In_1467);
nand U962 (N_962,In_721,N_612);
nor U963 (N_963,N_460,N_175);
xnor U964 (N_964,N_533,N_585);
nand U965 (N_965,In_1470,N_726);
xnor U966 (N_966,N_689,N_484);
xnor U967 (N_967,N_343,In_602);
nand U968 (N_968,In_67,N_700);
and U969 (N_969,N_682,N_679);
xor U970 (N_970,N_628,N_592);
nand U971 (N_971,N_704,In_1323);
nand U972 (N_972,In_157,In_87);
and U973 (N_973,N_330,N_505);
nor U974 (N_974,In_104,In_1256);
nor U975 (N_975,N_404,In_764);
or U976 (N_976,In_980,In_1167);
or U977 (N_977,In_896,N_310);
nand U978 (N_978,N_526,N_588);
or U979 (N_979,N_278,N_702);
or U980 (N_980,In_1085,N_407);
nand U981 (N_981,N_590,In_389);
and U982 (N_982,In_1164,N_27);
nor U983 (N_983,N_608,N_476);
or U984 (N_984,N_548,In_88);
xnor U985 (N_985,N_503,N_148);
and U986 (N_986,In_590,In_78);
nor U987 (N_987,N_509,In_1388);
or U988 (N_988,In_689,In_374);
nand U989 (N_989,In_1129,In_23);
nand U990 (N_990,In_161,In_968);
xor U991 (N_991,In_1497,N_286);
nor U992 (N_992,In_198,N_716);
or U993 (N_993,N_637,In_1011);
xnor U994 (N_994,In_446,N_384);
nand U995 (N_995,In_855,N_581);
xor U996 (N_996,N_658,N_118);
xnor U997 (N_997,In_1441,N_377);
xor U998 (N_998,In_395,N_562);
nor U999 (N_999,N_502,In_139);
or U1000 (N_1000,N_882,N_985);
xor U1001 (N_1001,N_697,N_675);
nand U1002 (N_1002,In_195,In_150);
xor U1003 (N_1003,N_909,In_287);
nor U1004 (N_1004,In_1345,N_777);
nor U1005 (N_1005,N_796,N_844);
or U1006 (N_1006,N_948,N_834);
nor U1007 (N_1007,N_989,N_772);
and U1008 (N_1008,N_516,N_893);
nor U1009 (N_1009,N_580,N_963);
nor U1010 (N_1010,N_944,In_109);
and U1011 (N_1011,N_987,N_883);
nor U1012 (N_1012,N_758,In_651);
nand U1013 (N_1013,N_920,N_472);
nand U1014 (N_1014,N_901,N_801);
nand U1015 (N_1015,N_896,N_576);
and U1016 (N_1016,N_764,N_819);
and U1017 (N_1017,N_714,N_187);
xor U1018 (N_1018,In_1142,N_745);
xor U1019 (N_1019,N_462,In_1370);
xnor U1020 (N_1020,N_974,N_792);
xor U1021 (N_1021,N_904,In_1393);
nand U1022 (N_1022,N_957,N_845);
nor U1023 (N_1023,N_564,N_786);
xor U1024 (N_1024,N_670,N_855);
or U1025 (N_1025,N_980,In_167);
nand U1026 (N_1026,N_943,In_955);
nor U1027 (N_1027,In_693,N_837);
nand U1028 (N_1028,N_544,N_890);
nor U1029 (N_1029,N_954,N_610);
or U1030 (N_1030,N_848,N_861);
and U1031 (N_1031,N_365,N_767);
and U1032 (N_1032,N_561,N_942);
nor U1033 (N_1033,In_200,In_338);
or U1034 (N_1034,N_401,N_869);
xnor U1035 (N_1035,N_100,N_236);
or U1036 (N_1036,N_294,N_791);
nand U1037 (N_1037,N_894,N_914);
nand U1038 (N_1038,N_551,N_667);
and U1039 (N_1039,N_750,N_838);
and U1040 (N_1040,N_438,N_806);
xor U1041 (N_1041,N_302,N_748);
nand U1042 (N_1042,N_242,N_63);
xor U1043 (N_1043,N_683,In_1066);
xor U1044 (N_1044,N_540,N_594);
and U1045 (N_1045,N_798,N_770);
or U1046 (N_1046,N_555,In_533);
xnor U1047 (N_1047,N_907,In_226);
nor U1048 (N_1048,N_998,N_723);
or U1049 (N_1049,N_601,N_774);
or U1050 (N_1050,In_1193,In_665);
or U1051 (N_1051,N_427,N_917);
or U1052 (N_1052,N_574,N_872);
xor U1053 (N_1053,N_342,N_811);
or U1054 (N_1054,N_680,N_828);
nor U1055 (N_1055,In_498,In_21);
nor U1056 (N_1056,N_739,N_699);
nand U1057 (N_1057,N_793,N_865);
or U1058 (N_1058,N_445,In_541);
nand U1059 (N_1059,N_784,N_898);
xnor U1060 (N_1060,N_922,N_840);
nor U1061 (N_1061,In_276,N_990);
and U1062 (N_1062,N_879,N_808);
or U1063 (N_1063,N_962,N_24);
xnor U1064 (N_1064,In_1432,N_769);
or U1065 (N_1065,N_737,N_771);
xnor U1066 (N_1066,N_986,In_857);
nand U1067 (N_1067,N_905,N_155);
xnor U1068 (N_1068,N_863,N_529);
xor U1069 (N_1069,N_884,N_335);
or U1070 (N_1070,N_213,N_411);
nand U1071 (N_1071,In_1006,N_935);
nor U1072 (N_1072,N_746,N_624);
nand U1073 (N_1073,N_858,N_654);
nor U1074 (N_1074,N_970,N_978);
nor U1075 (N_1075,N_773,N_983);
xor U1076 (N_1076,N_558,N_466);
xnor U1077 (N_1077,N_851,In_115);
nor U1078 (N_1078,In_339,N_743);
nand U1079 (N_1079,In_1199,N_827);
nand U1080 (N_1080,N_906,N_759);
or U1081 (N_1081,In_996,N_575);
nor U1082 (N_1082,N_584,N_724);
xnor U1083 (N_1083,N_895,N_919);
and U1084 (N_1084,N_866,N_717);
xor U1085 (N_1085,N_710,N_768);
xnor U1086 (N_1086,N_857,N_911);
or U1087 (N_1087,N_283,N_619);
nor U1088 (N_1088,N_386,N_929);
or U1089 (N_1089,N_669,N_874);
nor U1090 (N_1090,N_913,N_975);
nor U1091 (N_1091,N_690,N_733);
or U1092 (N_1092,N_656,N_928);
xnor U1093 (N_1093,In_634,N_591);
nand U1094 (N_1094,N_803,In_1347);
nand U1095 (N_1095,N_947,N_800);
nand U1096 (N_1096,N_45,N_936);
or U1097 (N_1097,N_921,In_543);
or U1098 (N_1098,N_864,In_1097);
or U1099 (N_1099,N_877,N_910);
and U1100 (N_1100,N_814,N_999);
xnor U1101 (N_1101,N_831,N_262);
nor U1102 (N_1102,In_392,N_880);
nand U1103 (N_1103,N_284,N_653);
and U1104 (N_1104,N_886,N_756);
nor U1105 (N_1105,N_821,N_932);
xnor U1106 (N_1106,N_186,N_995);
nand U1107 (N_1107,N_818,N_82);
or U1108 (N_1108,N_495,N_83);
xnor U1109 (N_1109,N_523,N_103);
and U1110 (N_1110,N_417,In_422);
or U1111 (N_1111,In_1489,In_1044);
nand U1112 (N_1112,N_997,N_994);
xor U1113 (N_1113,In_911,N_996);
xor U1114 (N_1114,N_829,N_766);
xnor U1115 (N_1115,N_639,In_512);
and U1116 (N_1116,N_293,In_1114);
or U1117 (N_1117,N_854,In_681);
and U1118 (N_1118,In_1247,N_934);
nor U1119 (N_1119,N_938,N_842);
nand U1120 (N_1120,N_939,In_724);
nand U1121 (N_1121,In_3,N_812);
xnor U1122 (N_1122,In_234,N_727);
or U1123 (N_1123,N_878,N_876);
nor U1124 (N_1124,N_809,N_797);
nor U1125 (N_1125,N_763,N_826);
and U1126 (N_1126,N_871,N_506);
or U1127 (N_1127,N_738,N_973);
nor U1128 (N_1128,N_621,N_790);
nand U1129 (N_1129,N_976,N_916);
xnor U1130 (N_1130,In_539,N_949);
xnor U1131 (N_1131,N_707,N_873);
and U1132 (N_1132,In_679,N_288);
xor U1133 (N_1133,N_593,In_663);
or U1134 (N_1134,N_959,N_241);
or U1135 (N_1135,N_629,In_1257);
and U1136 (N_1136,In_1122,N_824);
or U1137 (N_1137,N_899,N_703);
nand U1138 (N_1138,In_384,N_867);
nand U1139 (N_1139,N_765,N_946);
or U1140 (N_1140,N_940,N_425);
nor U1141 (N_1141,N_200,N_988);
nor U1142 (N_1142,N_569,N_830);
or U1143 (N_1143,N_897,N_981);
xor U1144 (N_1144,N_277,N_383);
and U1145 (N_1145,In_536,N_903);
and U1146 (N_1146,N_862,N_692);
and U1147 (N_1147,N_711,N_761);
nor U1148 (N_1148,N_836,N_810);
nor U1149 (N_1149,N_902,N_953);
nor U1150 (N_1150,N_950,In_914);
and U1151 (N_1151,N_977,In_524);
nor U1152 (N_1152,N_76,N_706);
and U1153 (N_1153,N_982,N_631);
xor U1154 (N_1154,N_984,In_1207);
xor U1155 (N_1155,N_101,N_807);
nor U1156 (N_1156,In_750,N_888);
nand U1157 (N_1157,N_933,N_780);
nor U1158 (N_1158,N_887,N_587);
nor U1159 (N_1159,N_927,N_446);
nor U1160 (N_1160,N_545,N_930);
nor U1161 (N_1161,N_852,N_937);
nor U1162 (N_1162,N_782,N_755);
xor U1163 (N_1163,In_222,In_798);
nor U1164 (N_1164,N_972,N_941);
xnor U1165 (N_1165,N_820,N_788);
nor U1166 (N_1166,N_918,N_713);
or U1167 (N_1167,N_965,In_544);
nand U1168 (N_1168,In_866,N_992);
or U1169 (N_1169,N_968,N_892);
nor U1170 (N_1170,N_709,N_971);
nor U1171 (N_1171,N_881,N_960);
or U1172 (N_1172,N_550,N_634);
nor U1173 (N_1173,N_835,N_378);
nor U1174 (N_1174,N_408,N_951);
nor U1175 (N_1175,N_336,N_783);
and U1176 (N_1176,N_752,N_78);
xor U1177 (N_1177,N_969,N_961);
and U1178 (N_1178,N_320,N_875);
or U1179 (N_1179,N_785,N_211);
xor U1180 (N_1180,In_1318,N_813);
or U1181 (N_1181,In_957,N_595);
nor U1182 (N_1182,N_923,N_239);
xor U1183 (N_1183,N_816,N_860);
xor U1184 (N_1184,In_1452,In_113);
and U1185 (N_1185,N_924,In_734);
nand U1186 (N_1186,N_638,N_945);
and U1187 (N_1187,In_975,N_687);
nand U1188 (N_1188,N_753,N_853);
nand U1189 (N_1189,In_233,In_1454);
xnor U1190 (N_1190,N_519,N_815);
xnor U1191 (N_1191,In_575,N_964);
xnor U1192 (N_1192,N_760,N_850);
or U1193 (N_1193,N_885,N_109);
or U1194 (N_1194,N_605,In_552);
xnor U1195 (N_1195,N_891,N_781);
nand U1196 (N_1196,N_402,N_846);
nor U1197 (N_1197,N_889,N_177);
or U1198 (N_1198,N_868,N_779);
xor U1199 (N_1199,N_513,N_795);
and U1200 (N_1200,N_822,N_563);
xnor U1201 (N_1201,N_609,N_536);
and U1202 (N_1202,N_841,N_775);
nor U1203 (N_1203,In_1095,N_856);
nor U1204 (N_1204,N_740,In_1424);
or U1205 (N_1205,In_227,N_832);
or U1206 (N_1206,N_776,In_664);
nor U1207 (N_1207,In_1352,N_958);
nor U1208 (N_1208,N_794,N_804);
xnor U1209 (N_1209,N_908,N_955);
nand U1210 (N_1210,N_751,N_778);
xor U1211 (N_1211,N_275,N_381);
xor U1212 (N_1212,N_789,N_833);
xnor U1213 (N_1213,N_967,N_353);
nand U1214 (N_1214,N_645,N_635);
or U1215 (N_1215,In_1160,N_93);
nor U1216 (N_1216,N_530,N_966);
and U1217 (N_1217,N_847,N_802);
nor U1218 (N_1218,N_521,N_993);
and U1219 (N_1219,In_402,N_553);
xor U1220 (N_1220,N_931,In_1064);
xnor U1221 (N_1221,N_642,N_661);
nor U1222 (N_1222,N_817,N_839);
nand U1223 (N_1223,In_73,N_956);
or U1224 (N_1224,In_332,N_346);
nand U1225 (N_1225,N_912,N_589);
nor U1226 (N_1226,N_205,N_391);
nand U1227 (N_1227,In_37,N_925);
or U1228 (N_1228,N_685,In_202);
nor U1229 (N_1229,N_597,N_979);
xnor U1230 (N_1230,N_870,N_698);
or U1231 (N_1231,In_377,N_926);
and U1232 (N_1232,N_823,In_310);
and U1233 (N_1233,In_277,In_248);
or U1234 (N_1234,N_762,N_285);
nand U1235 (N_1235,In_288,N_843);
nor U1236 (N_1236,N_787,N_547);
and U1237 (N_1237,In_343,In_916);
xnor U1238 (N_1238,N_630,N_514);
or U1239 (N_1239,N_512,In_179);
nor U1240 (N_1240,N_900,N_218);
xnor U1241 (N_1241,N_952,N_754);
xor U1242 (N_1242,N_991,N_668);
xnor U1243 (N_1243,N_757,In_1332);
nor U1244 (N_1244,N_825,N_556);
or U1245 (N_1245,N_643,N_849);
or U1246 (N_1246,N_799,N_725);
or U1247 (N_1247,N_915,N_805);
or U1248 (N_1248,N_256,N_358);
and U1249 (N_1249,N_640,N_859);
nor U1250 (N_1250,N_1172,N_1183);
and U1251 (N_1251,N_1152,N_1014);
or U1252 (N_1252,N_1055,N_1191);
nor U1253 (N_1253,N_1121,N_1189);
xnor U1254 (N_1254,N_1165,N_1168);
and U1255 (N_1255,N_1115,N_1213);
xnor U1256 (N_1256,N_1156,N_1018);
nor U1257 (N_1257,N_1111,N_1202);
xnor U1258 (N_1258,N_1206,N_1036);
nor U1259 (N_1259,N_1056,N_1131);
xnor U1260 (N_1260,N_1242,N_1114);
nor U1261 (N_1261,N_1231,N_1057);
and U1262 (N_1262,N_1042,N_1052);
and U1263 (N_1263,N_1110,N_1001);
xor U1264 (N_1264,N_1070,N_1095);
xnor U1265 (N_1265,N_1178,N_1100);
and U1266 (N_1266,N_1162,N_1039);
nand U1267 (N_1267,N_1151,N_1120);
nand U1268 (N_1268,N_1236,N_1140);
nor U1269 (N_1269,N_1104,N_1022);
nand U1270 (N_1270,N_1196,N_1179);
xnor U1271 (N_1271,N_1221,N_1240);
nand U1272 (N_1272,N_1145,N_1082);
nand U1273 (N_1273,N_1048,N_1008);
xnor U1274 (N_1274,N_1085,N_1103);
and U1275 (N_1275,N_1109,N_1139);
xnor U1276 (N_1276,N_1074,N_1123);
nor U1277 (N_1277,N_1235,N_1245);
nor U1278 (N_1278,N_1164,N_1160);
nor U1279 (N_1279,N_1154,N_1031);
nor U1280 (N_1280,N_1169,N_1177);
and U1281 (N_1281,N_1180,N_1117);
nand U1282 (N_1282,N_1025,N_1066);
and U1283 (N_1283,N_1105,N_1144);
nor U1284 (N_1284,N_1079,N_1034);
nor U1285 (N_1285,N_1155,N_1166);
and U1286 (N_1286,N_1194,N_1219);
or U1287 (N_1287,N_1050,N_1138);
nand U1288 (N_1288,N_1116,N_1005);
nor U1289 (N_1289,N_1086,N_1107);
or U1290 (N_1290,N_1217,N_1244);
and U1291 (N_1291,N_1112,N_1043);
and U1292 (N_1292,N_1125,N_1149);
xor U1293 (N_1293,N_1075,N_1247);
and U1294 (N_1294,N_1032,N_1146);
nand U1295 (N_1295,N_1096,N_1068);
nor U1296 (N_1296,N_1176,N_1019);
xor U1297 (N_1297,N_1136,N_1137);
or U1298 (N_1298,N_1218,N_1241);
nor U1299 (N_1299,N_1119,N_1201);
nor U1300 (N_1300,N_1076,N_1186);
xor U1301 (N_1301,N_1197,N_1141);
nor U1302 (N_1302,N_1227,N_1159);
nor U1303 (N_1303,N_1143,N_1220);
and U1304 (N_1304,N_1098,N_1228);
xnor U1305 (N_1305,N_1239,N_1080);
and U1306 (N_1306,N_1013,N_1062);
nor U1307 (N_1307,N_1028,N_1071);
and U1308 (N_1308,N_1187,N_1044);
nand U1309 (N_1309,N_1003,N_1210);
xnor U1310 (N_1310,N_1006,N_1222);
or U1311 (N_1311,N_1148,N_1053);
xnor U1312 (N_1312,N_1170,N_1040);
nor U1313 (N_1313,N_1161,N_1246);
and U1314 (N_1314,N_1113,N_1163);
or U1315 (N_1315,N_1058,N_1203);
and U1316 (N_1316,N_1090,N_1015);
xnor U1317 (N_1317,N_1078,N_1016);
nand U1318 (N_1318,N_1030,N_1041);
xnor U1319 (N_1319,N_1094,N_1069);
nor U1320 (N_1320,N_1190,N_1249);
xnor U1321 (N_1321,N_1046,N_1195);
xor U1322 (N_1322,N_1212,N_1065);
nor U1323 (N_1323,N_1207,N_1226);
and U1324 (N_1324,N_1216,N_1193);
nor U1325 (N_1325,N_1127,N_1229);
or U1326 (N_1326,N_1126,N_1214);
or U1327 (N_1327,N_1158,N_1004);
or U1328 (N_1328,N_1063,N_1153);
or U1329 (N_1329,N_1029,N_1089);
nor U1330 (N_1330,N_1185,N_1208);
nand U1331 (N_1331,N_1097,N_1174);
or U1332 (N_1332,N_1188,N_1130);
nand U1333 (N_1333,N_1184,N_1128);
nor U1334 (N_1334,N_1064,N_1059);
nand U1335 (N_1335,N_1088,N_1087);
nand U1336 (N_1336,N_1233,N_1000);
xor U1337 (N_1337,N_1045,N_1173);
nand U1338 (N_1338,N_1023,N_1175);
or U1339 (N_1339,N_1225,N_1230);
nand U1340 (N_1340,N_1021,N_1101);
xor U1341 (N_1341,N_1204,N_1135);
xor U1342 (N_1342,N_1072,N_1108);
and U1343 (N_1343,N_1092,N_1009);
xor U1344 (N_1344,N_1051,N_1234);
and U1345 (N_1345,N_1238,N_1083);
xnor U1346 (N_1346,N_1133,N_1060);
xnor U1347 (N_1347,N_1017,N_1223);
nand U1348 (N_1348,N_1106,N_1038);
xor U1349 (N_1349,N_1012,N_1200);
xnor U1350 (N_1350,N_1102,N_1002);
xnor U1351 (N_1351,N_1224,N_1198);
nand U1352 (N_1352,N_1054,N_1199);
or U1353 (N_1353,N_1209,N_1134);
nor U1354 (N_1354,N_1091,N_1211);
nor U1355 (N_1355,N_1215,N_1118);
nand U1356 (N_1356,N_1033,N_1007);
nand U1357 (N_1357,N_1037,N_1020);
or U1358 (N_1358,N_1093,N_1171);
xnor U1359 (N_1359,N_1248,N_1243);
or U1360 (N_1360,N_1122,N_1024);
and U1361 (N_1361,N_1157,N_1181);
and U1362 (N_1362,N_1129,N_1077);
nor U1363 (N_1363,N_1084,N_1205);
xor U1364 (N_1364,N_1061,N_1132);
and U1365 (N_1365,N_1081,N_1150);
nor U1366 (N_1366,N_1067,N_1142);
nor U1367 (N_1367,N_1027,N_1192);
nor U1368 (N_1368,N_1047,N_1026);
xor U1369 (N_1369,N_1011,N_1237);
xnor U1370 (N_1370,N_1035,N_1010);
or U1371 (N_1371,N_1232,N_1049);
nand U1372 (N_1372,N_1182,N_1073);
xnor U1373 (N_1373,N_1167,N_1099);
nand U1374 (N_1374,N_1124,N_1147);
nand U1375 (N_1375,N_1075,N_1015);
nor U1376 (N_1376,N_1029,N_1033);
xnor U1377 (N_1377,N_1138,N_1110);
xnor U1378 (N_1378,N_1230,N_1065);
or U1379 (N_1379,N_1014,N_1050);
and U1380 (N_1380,N_1097,N_1090);
nor U1381 (N_1381,N_1044,N_1022);
and U1382 (N_1382,N_1064,N_1099);
and U1383 (N_1383,N_1024,N_1095);
or U1384 (N_1384,N_1179,N_1224);
nor U1385 (N_1385,N_1147,N_1180);
and U1386 (N_1386,N_1189,N_1195);
xnor U1387 (N_1387,N_1217,N_1223);
xnor U1388 (N_1388,N_1197,N_1234);
nand U1389 (N_1389,N_1122,N_1195);
nor U1390 (N_1390,N_1071,N_1184);
nand U1391 (N_1391,N_1157,N_1133);
and U1392 (N_1392,N_1000,N_1051);
nor U1393 (N_1393,N_1203,N_1174);
nand U1394 (N_1394,N_1172,N_1035);
or U1395 (N_1395,N_1079,N_1026);
or U1396 (N_1396,N_1111,N_1048);
xor U1397 (N_1397,N_1141,N_1135);
nor U1398 (N_1398,N_1168,N_1139);
xnor U1399 (N_1399,N_1248,N_1108);
xor U1400 (N_1400,N_1194,N_1190);
and U1401 (N_1401,N_1190,N_1093);
or U1402 (N_1402,N_1072,N_1012);
nor U1403 (N_1403,N_1241,N_1119);
xor U1404 (N_1404,N_1199,N_1149);
nand U1405 (N_1405,N_1202,N_1142);
nand U1406 (N_1406,N_1124,N_1100);
xnor U1407 (N_1407,N_1120,N_1066);
xnor U1408 (N_1408,N_1140,N_1072);
and U1409 (N_1409,N_1135,N_1220);
and U1410 (N_1410,N_1059,N_1145);
or U1411 (N_1411,N_1062,N_1008);
nor U1412 (N_1412,N_1120,N_1209);
and U1413 (N_1413,N_1170,N_1165);
nand U1414 (N_1414,N_1061,N_1113);
nand U1415 (N_1415,N_1043,N_1174);
nor U1416 (N_1416,N_1235,N_1072);
or U1417 (N_1417,N_1072,N_1214);
nor U1418 (N_1418,N_1034,N_1159);
nor U1419 (N_1419,N_1044,N_1228);
or U1420 (N_1420,N_1024,N_1235);
nand U1421 (N_1421,N_1225,N_1169);
and U1422 (N_1422,N_1041,N_1212);
xnor U1423 (N_1423,N_1194,N_1137);
nand U1424 (N_1424,N_1114,N_1031);
xnor U1425 (N_1425,N_1207,N_1041);
and U1426 (N_1426,N_1130,N_1145);
nand U1427 (N_1427,N_1146,N_1157);
xor U1428 (N_1428,N_1030,N_1132);
nand U1429 (N_1429,N_1105,N_1209);
xnor U1430 (N_1430,N_1236,N_1151);
nand U1431 (N_1431,N_1086,N_1162);
nand U1432 (N_1432,N_1043,N_1072);
and U1433 (N_1433,N_1186,N_1115);
and U1434 (N_1434,N_1211,N_1110);
or U1435 (N_1435,N_1226,N_1183);
xor U1436 (N_1436,N_1046,N_1187);
xor U1437 (N_1437,N_1011,N_1226);
and U1438 (N_1438,N_1223,N_1039);
and U1439 (N_1439,N_1073,N_1129);
nand U1440 (N_1440,N_1067,N_1007);
nand U1441 (N_1441,N_1183,N_1189);
or U1442 (N_1442,N_1186,N_1095);
nor U1443 (N_1443,N_1004,N_1089);
or U1444 (N_1444,N_1033,N_1052);
nor U1445 (N_1445,N_1236,N_1137);
nand U1446 (N_1446,N_1064,N_1030);
nor U1447 (N_1447,N_1107,N_1054);
xnor U1448 (N_1448,N_1090,N_1137);
nor U1449 (N_1449,N_1040,N_1133);
nor U1450 (N_1450,N_1051,N_1155);
and U1451 (N_1451,N_1147,N_1051);
nand U1452 (N_1452,N_1061,N_1172);
xnor U1453 (N_1453,N_1070,N_1180);
or U1454 (N_1454,N_1178,N_1119);
nor U1455 (N_1455,N_1005,N_1081);
nand U1456 (N_1456,N_1043,N_1145);
nand U1457 (N_1457,N_1069,N_1048);
nor U1458 (N_1458,N_1090,N_1053);
and U1459 (N_1459,N_1038,N_1210);
and U1460 (N_1460,N_1164,N_1131);
nand U1461 (N_1461,N_1212,N_1150);
nor U1462 (N_1462,N_1185,N_1128);
xnor U1463 (N_1463,N_1183,N_1223);
nor U1464 (N_1464,N_1123,N_1073);
nand U1465 (N_1465,N_1048,N_1125);
nand U1466 (N_1466,N_1112,N_1210);
nor U1467 (N_1467,N_1199,N_1172);
and U1468 (N_1468,N_1173,N_1143);
and U1469 (N_1469,N_1006,N_1209);
nor U1470 (N_1470,N_1004,N_1091);
and U1471 (N_1471,N_1008,N_1022);
and U1472 (N_1472,N_1225,N_1151);
or U1473 (N_1473,N_1127,N_1090);
nand U1474 (N_1474,N_1062,N_1082);
and U1475 (N_1475,N_1036,N_1046);
or U1476 (N_1476,N_1085,N_1094);
and U1477 (N_1477,N_1026,N_1206);
xor U1478 (N_1478,N_1168,N_1159);
xnor U1479 (N_1479,N_1061,N_1009);
nor U1480 (N_1480,N_1117,N_1050);
nor U1481 (N_1481,N_1211,N_1112);
and U1482 (N_1482,N_1186,N_1180);
and U1483 (N_1483,N_1074,N_1085);
nor U1484 (N_1484,N_1074,N_1116);
xor U1485 (N_1485,N_1122,N_1059);
nand U1486 (N_1486,N_1044,N_1097);
xor U1487 (N_1487,N_1182,N_1181);
xnor U1488 (N_1488,N_1027,N_1187);
nor U1489 (N_1489,N_1102,N_1034);
and U1490 (N_1490,N_1133,N_1222);
nand U1491 (N_1491,N_1096,N_1170);
and U1492 (N_1492,N_1159,N_1115);
nor U1493 (N_1493,N_1221,N_1090);
or U1494 (N_1494,N_1158,N_1039);
xnor U1495 (N_1495,N_1161,N_1065);
nor U1496 (N_1496,N_1074,N_1137);
nand U1497 (N_1497,N_1109,N_1191);
or U1498 (N_1498,N_1119,N_1011);
nand U1499 (N_1499,N_1040,N_1244);
nor U1500 (N_1500,N_1297,N_1475);
xnor U1501 (N_1501,N_1413,N_1323);
xnor U1502 (N_1502,N_1259,N_1453);
nor U1503 (N_1503,N_1472,N_1425);
nor U1504 (N_1504,N_1456,N_1484);
xor U1505 (N_1505,N_1277,N_1424);
nor U1506 (N_1506,N_1345,N_1333);
or U1507 (N_1507,N_1418,N_1481);
or U1508 (N_1508,N_1359,N_1258);
and U1509 (N_1509,N_1463,N_1421);
and U1510 (N_1510,N_1386,N_1433);
nor U1511 (N_1511,N_1315,N_1497);
nand U1512 (N_1512,N_1492,N_1283);
xnor U1513 (N_1513,N_1488,N_1266);
xor U1514 (N_1514,N_1379,N_1401);
or U1515 (N_1515,N_1302,N_1293);
or U1516 (N_1516,N_1402,N_1473);
nand U1517 (N_1517,N_1321,N_1465);
nor U1518 (N_1518,N_1372,N_1408);
xor U1519 (N_1519,N_1252,N_1311);
or U1520 (N_1520,N_1279,N_1368);
xnor U1521 (N_1521,N_1385,N_1255);
and U1522 (N_1522,N_1287,N_1480);
xnor U1523 (N_1523,N_1328,N_1457);
nand U1524 (N_1524,N_1291,N_1367);
xor U1525 (N_1525,N_1330,N_1254);
nor U1526 (N_1526,N_1347,N_1343);
xnor U1527 (N_1527,N_1409,N_1290);
or U1528 (N_1528,N_1319,N_1441);
and U1529 (N_1529,N_1495,N_1431);
nand U1530 (N_1530,N_1439,N_1419);
xor U1531 (N_1531,N_1286,N_1373);
and U1532 (N_1532,N_1435,N_1332);
or U1533 (N_1533,N_1407,N_1427);
or U1534 (N_1534,N_1423,N_1309);
and U1535 (N_1535,N_1442,N_1436);
xnor U1536 (N_1536,N_1483,N_1262);
xnor U1537 (N_1537,N_1305,N_1256);
nand U1538 (N_1538,N_1468,N_1449);
or U1539 (N_1539,N_1351,N_1422);
and U1540 (N_1540,N_1316,N_1461);
nand U1541 (N_1541,N_1400,N_1467);
or U1542 (N_1542,N_1493,N_1393);
xnor U1543 (N_1543,N_1378,N_1337);
nor U1544 (N_1544,N_1296,N_1406);
and U1545 (N_1545,N_1490,N_1295);
and U1546 (N_1546,N_1250,N_1269);
nand U1547 (N_1547,N_1450,N_1358);
nor U1548 (N_1548,N_1395,N_1324);
nor U1549 (N_1549,N_1459,N_1273);
xnor U1550 (N_1550,N_1460,N_1380);
nor U1551 (N_1551,N_1491,N_1346);
and U1552 (N_1552,N_1394,N_1479);
nor U1553 (N_1553,N_1498,N_1284);
or U1554 (N_1554,N_1478,N_1445);
nor U1555 (N_1555,N_1257,N_1403);
xor U1556 (N_1556,N_1384,N_1381);
nor U1557 (N_1557,N_1253,N_1398);
xor U1558 (N_1558,N_1455,N_1350);
xor U1559 (N_1559,N_1298,N_1348);
or U1560 (N_1560,N_1338,N_1251);
and U1561 (N_1561,N_1264,N_1272);
nand U1562 (N_1562,N_1270,N_1308);
or U1563 (N_1563,N_1438,N_1494);
xor U1564 (N_1564,N_1443,N_1451);
and U1565 (N_1565,N_1322,N_1454);
nor U1566 (N_1566,N_1356,N_1404);
nand U1567 (N_1567,N_1278,N_1260);
xnor U1568 (N_1568,N_1434,N_1437);
nand U1569 (N_1569,N_1353,N_1271);
nor U1570 (N_1570,N_1362,N_1375);
and U1571 (N_1571,N_1444,N_1417);
xnor U1572 (N_1572,N_1392,N_1469);
nand U1573 (N_1573,N_1383,N_1313);
or U1574 (N_1574,N_1341,N_1477);
or U1575 (N_1575,N_1429,N_1352);
and U1576 (N_1576,N_1331,N_1304);
nor U1577 (N_1577,N_1446,N_1363);
nand U1578 (N_1578,N_1334,N_1397);
xnor U1579 (N_1579,N_1452,N_1292);
nor U1580 (N_1580,N_1399,N_1405);
nor U1581 (N_1581,N_1389,N_1416);
or U1582 (N_1582,N_1336,N_1325);
nand U1583 (N_1583,N_1275,N_1349);
xor U1584 (N_1584,N_1448,N_1354);
xnor U1585 (N_1585,N_1382,N_1474);
and U1586 (N_1586,N_1280,N_1268);
nor U1587 (N_1587,N_1428,N_1471);
nand U1588 (N_1588,N_1282,N_1329);
nor U1589 (N_1589,N_1320,N_1299);
xor U1590 (N_1590,N_1371,N_1388);
nor U1591 (N_1591,N_1289,N_1489);
or U1592 (N_1592,N_1327,N_1374);
xnor U1593 (N_1593,N_1306,N_1387);
or U1594 (N_1594,N_1391,N_1300);
xnor U1595 (N_1595,N_1344,N_1307);
nand U1596 (N_1596,N_1340,N_1415);
nand U1597 (N_1597,N_1281,N_1360);
nand U1598 (N_1598,N_1318,N_1364);
xnor U1599 (N_1599,N_1496,N_1261);
nor U1600 (N_1600,N_1294,N_1411);
nand U1601 (N_1601,N_1440,N_1263);
xor U1602 (N_1602,N_1303,N_1276);
nand U1603 (N_1603,N_1487,N_1342);
or U1604 (N_1604,N_1390,N_1361);
nor U1605 (N_1605,N_1462,N_1366);
xnor U1606 (N_1606,N_1466,N_1370);
xor U1607 (N_1607,N_1267,N_1447);
or U1608 (N_1608,N_1414,N_1396);
xnor U1609 (N_1609,N_1339,N_1485);
xnor U1610 (N_1610,N_1326,N_1335);
nor U1611 (N_1611,N_1412,N_1432);
and U1612 (N_1612,N_1301,N_1420);
or U1613 (N_1613,N_1464,N_1310);
xnor U1614 (N_1614,N_1470,N_1476);
nand U1615 (N_1615,N_1410,N_1486);
nand U1616 (N_1616,N_1426,N_1499);
or U1617 (N_1617,N_1377,N_1357);
nand U1618 (N_1618,N_1312,N_1288);
nor U1619 (N_1619,N_1355,N_1317);
xor U1620 (N_1620,N_1458,N_1274);
or U1621 (N_1621,N_1365,N_1285);
xor U1622 (N_1622,N_1430,N_1369);
nand U1623 (N_1623,N_1376,N_1265);
nand U1624 (N_1624,N_1482,N_1314);
xor U1625 (N_1625,N_1416,N_1269);
nor U1626 (N_1626,N_1318,N_1305);
xnor U1627 (N_1627,N_1351,N_1427);
or U1628 (N_1628,N_1364,N_1282);
xnor U1629 (N_1629,N_1367,N_1483);
xor U1630 (N_1630,N_1437,N_1419);
nand U1631 (N_1631,N_1301,N_1304);
or U1632 (N_1632,N_1309,N_1485);
xor U1633 (N_1633,N_1282,N_1331);
or U1634 (N_1634,N_1455,N_1346);
or U1635 (N_1635,N_1290,N_1451);
nor U1636 (N_1636,N_1448,N_1301);
xnor U1637 (N_1637,N_1386,N_1447);
xor U1638 (N_1638,N_1334,N_1301);
nand U1639 (N_1639,N_1450,N_1342);
nand U1640 (N_1640,N_1412,N_1303);
nor U1641 (N_1641,N_1476,N_1267);
nand U1642 (N_1642,N_1279,N_1322);
and U1643 (N_1643,N_1498,N_1290);
xnor U1644 (N_1644,N_1336,N_1494);
nor U1645 (N_1645,N_1398,N_1397);
xnor U1646 (N_1646,N_1295,N_1298);
or U1647 (N_1647,N_1291,N_1491);
and U1648 (N_1648,N_1316,N_1390);
and U1649 (N_1649,N_1467,N_1408);
and U1650 (N_1650,N_1491,N_1266);
nor U1651 (N_1651,N_1341,N_1427);
or U1652 (N_1652,N_1463,N_1419);
nor U1653 (N_1653,N_1331,N_1371);
nand U1654 (N_1654,N_1297,N_1427);
and U1655 (N_1655,N_1490,N_1250);
xor U1656 (N_1656,N_1372,N_1289);
nand U1657 (N_1657,N_1366,N_1467);
and U1658 (N_1658,N_1452,N_1291);
nor U1659 (N_1659,N_1381,N_1342);
or U1660 (N_1660,N_1464,N_1399);
nand U1661 (N_1661,N_1373,N_1377);
xnor U1662 (N_1662,N_1313,N_1376);
xor U1663 (N_1663,N_1312,N_1292);
and U1664 (N_1664,N_1301,N_1478);
or U1665 (N_1665,N_1388,N_1288);
nor U1666 (N_1666,N_1379,N_1342);
nor U1667 (N_1667,N_1453,N_1300);
nor U1668 (N_1668,N_1484,N_1332);
xor U1669 (N_1669,N_1394,N_1399);
nand U1670 (N_1670,N_1388,N_1417);
and U1671 (N_1671,N_1266,N_1397);
and U1672 (N_1672,N_1498,N_1283);
or U1673 (N_1673,N_1358,N_1293);
or U1674 (N_1674,N_1415,N_1326);
and U1675 (N_1675,N_1323,N_1284);
and U1676 (N_1676,N_1467,N_1415);
nor U1677 (N_1677,N_1338,N_1295);
and U1678 (N_1678,N_1326,N_1385);
and U1679 (N_1679,N_1483,N_1298);
nand U1680 (N_1680,N_1389,N_1317);
nand U1681 (N_1681,N_1377,N_1407);
nand U1682 (N_1682,N_1428,N_1383);
or U1683 (N_1683,N_1255,N_1497);
or U1684 (N_1684,N_1254,N_1495);
and U1685 (N_1685,N_1460,N_1332);
nor U1686 (N_1686,N_1445,N_1415);
xor U1687 (N_1687,N_1343,N_1377);
nand U1688 (N_1688,N_1431,N_1338);
nor U1689 (N_1689,N_1455,N_1313);
xor U1690 (N_1690,N_1300,N_1435);
or U1691 (N_1691,N_1408,N_1399);
or U1692 (N_1692,N_1468,N_1428);
or U1693 (N_1693,N_1262,N_1382);
xor U1694 (N_1694,N_1277,N_1355);
xnor U1695 (N_1695,N_1427,N_1332);
xor U1696 (N_1696,N_1496,N_1274);
nand U1697 (N_1697,N_1284,N_1353);
and U1698 (N_1698,N_1362,N_1389);
nand U1699 (N_1699,N_1428,N_1311);
and U1700 (N_1700,N_1294,N_1322);
and U1701 (N_1701,N_1291,N_1405);
and U1702 (N_1702,N_1399,N_1349);
or U1703 (N_1703,N_1431,N_1372);
and U1704 (N_1704,N_1272,N_1330);
or U1705 (N_1705,N_1356,N_1426);
xor U1706 (N_1706,N_1308,N_1483);
nand U1707 (N_1707,N_1285,N_1464);
xor U1708 (N_1708,N_1377,N_1385);
and U1709 (N_1709,N_1313,N_1464);
nor U1710 (N_1710,N_1497,N_1301);
and U1711 (N_1711,N_1253,N_1329);
or U1712 (N_1712,N_1267,N_1348);
nor U1713 (N_1713,N_1354,N_1459);
nand U1714 (N_1714,N_1423,N_1476);
nand U1715 (N_1715,N_1279,N_1276);
or U1716 (N_1716,N_1259,N_1322);
and U1717 (N_1717,N_1310,N_1431);
and U1718 (N_1718,N_1493,N_1275);
or U1719 (N_1719,N_1343,N_1254);
nand U1720 (N_1720,N_1262,N_1366);
nor U1721 (N_1721,N_1374,N_1338);
or U1722 (N_1722,N_1480,N_1387);
nor U1723 (N_1723,N_1285,N_1382);
or U1724 (N_1724,N_1432,N_1311);
nand U1725 (N_1725,N_1415,N_1293);
and U1726 (N_1726,N_1422,N_1430);
or U1727 (N_1727,N_1393,N_1429);
xnor U1728 (N_1728,N_1447,N_1356);
and U1729 (N_1729,N_1461,N_1448);
and U1730 (N_1730,N_1400,N_1253);
nand U1731 (N_1731,N_1481,N_1287);
nor U1732 (N_1732,N_1335,N_1359);
xor U1733 (N_1733,N_1359,N_1345);
and U1734 (N_1734,N_1494,N_1398);
nand U1735 (N_1735,N_1302,N_1420);
nor U1736 (N_1736,N_1353,N_1293);
xor U1737 (N_1737,N_1276,N_1404);
nand U1738 (N_1738,N_1298,N_1342);
or U1739 (N_1739,N_1414,N_1429);
nor U1740 (N_1740,N_1461,N_1279);
nor U1741 (N_1741,N_1483,N_1414);
or U1742 (N_1742,N_1402,N_1264);
xor U1743 (N_1743,N_1326,N_1419);
xnor U1744 (N_1744,N_1352,N_1354);
or U1745 (N_1745,N_1385,N_1412);
nand U1746 (N_1746,N_1388,N_1406);
or U1747 (N_1747,N_1464,N_1250);
nor U1748 (N_1748,N_1360,N_1493);
nand U1749 (N_1749,N_1340,N_1397);
nand U1750 (N_1750,N_1568,N_1635);
nand U1751 (N_1751,N_1626,N_1560);
nor U1752 (N_1752,N_1703,N_1532);
and U1753 (N_1753,N_1653,N_1527);
and U1754 (N_1754,N_1526,N_1590);
nor U1755 (N_1755,N_1574,N_1596);
nor U1756 (N_1756,N_1600,N_1510);
nand U1757 (N_1757,N_1674,N_1639);
and U1758 (N_1758,N_1732,N_1717);
nand U1759 (N_1759,N_1671,N_1669);
or U1760 (N_1760,N_1530,N_1629);
and U1761 (N_1761,N_1556,N_1707);
and U1762 (N_1762,N_1744,N_1567);
or U1763 (N_1763,N_1644,N_1615);
and U1764 (N_1764,N_1578,N_1617);
nor U1765 (N_1765,N_1517,N_1519);
nand U1766 (N_1766,N_1749,N_1677);
xor U1767 (N_1767,N_1603,N_1702);
nand U1768 (N_1768,N_1662,N_1518);
nor U1769 (N_1769,N_1588,N_1610);
or U1770 (N_1770,N_1746,N_1569);
or U1771 (N_1771,N_1681,N_1656);
nand U1772 (N_1772,N_1724,N_1535);
xnor U1773 (N_1773,N_1505,N_1718);
or U1774 (N_1774,N_1570,N_1747);
nand U1775 (N_1775,N_1745,N_1733);
and U1776 (N_1776,N_1507,N_1711);
nor U1777 (N_1777,N_1604,N_1516);
or U1778 (N_1778,N_1704,N_1624);
xnor U1779 (N_1779,N_1719,N_1739);
and U1780 (N_1780,N_1571,N_1658);
or U1781 (N_1781,N_1661,N_1619);
or U1782 (N_1782,N_1665,N_1506);
nor U1783 (N_1783,N_1728,N_1737);
or U1784 (N_1784,N_1691,N_1651);
and U1785 (N_1785,N_1508,N_1502);
and U1786 (N_1786,N_1742,N_1633);
or U1787 (N_1787,N_1553,N_1642);
xnor U1788 (N_1788,N_1537,N_1706);
and U1789 (N_1789,N_1521,N_1566);
xnor U1790 (N_1790,N_1585,N_1544);
nand U1791 (N_1791,N_1673,N_1735);
nor U1792 (N_1792,N_1562,N_1623);
xor U1793 (N_1793,N_1545,N_1637);
xor U1794 (N_1794,N_1701,N_1589);
nor U1795 (N_1795,N_1705,N_1727);
nand U1796 (N_1796,N_1551,N_1602);
nor U1797 (N_1797,N_1734,N_1688);
xnor U1798 (N_1798,N_1664,N_1687);
or U1799 (N_1799,N_1700,N_1743);
nand U1800 (N_1800,N_1698,N_1685);
or U1801 (N_1801,N_1559,N_1652);
or U1802 (N_1802,N_1631,N_1609);
nand U1803 (N_1803,N_1680,N_1646);
xnor U1804 (N_1804,N_1641,N_1572);
xor U1805 (N_1805,N_1523,N_1621);
or U1806 (N_1806,N_1586,N_1540);
nor U1807 (N_1807,N_1686,N_1618);
or U1808 (N_1808,N_1670,N_1693);
and U1809 (N_1809,N_1716,N_1663);
nor U1810 (N_1810,N_1533,N_1584);
nor U1811 (N_1811,N_1666,N_1607);
nand U1812 (N_1812,N_1645,N_1576);
nand U1813 (N_1813,N_1547,N_1543);
nor U1814 (N_1814,N_1606,N_1729);
nand U1815 (N_1815,N_1573,N_1723);
nor U1816 (N_1816,N_1557,N_1689);
xor U1817 (N_1817,N_1640,N_1672);
or U1818 (N_1818,N_1726,N_1622);
nor U1819 (N_1819,N_1713,N_1536);
or U1820 (N_1820,N_1612,N_1512);
or U1821 (N_1821,N_1504,N_1613);
nand U1822 (N_1822,N_1528,N_1509);
and U1823 (N_1823,N_1592,N_1740);
and U1824 (N_1824,N_1614,N_1599);
nand U1825 (N_1825,N_1524,N_1534);
and U1826 (N_1826,N_1643,N_1683);
nand U1827 (N_1827,N_1655,N_1679);
xnor U1828 (N_1828,N_1684,N_1514);
nor U1829 (N_1829,N_1668,N_1546);
nor U1830 (N_1830,N_1577,N_1697);
xnor U1831 (N_1831,N_1736,N_1725);
and U1832 (N_1832,N_1548,N_1594);
or U1833 (N_1833,N_1579,N_1538);
and U1834 (N_1834,N_1541,N_1748);
or U1835 (N_1835,N_1676,N_1625);
xnor U1836 (N_1836,N_1649,N_1565);
and U1837 (N_1837,N_1598,N_1708);
and U1838 (N_1838,N_1709,N_1738);
or U1839 (N_1839,N_1501,N_1582);
nor U1840 (N_1840,N_1531,N_1611);
or U1841 (N_1841,N_1710,N_1678);
xor U1842 (N_1842,N_1587,N_1715);
nor U1843 (N_1843,N_1522,N_1520);
xor U1844 (N_1844,N_1561,N_1682);
xnor U1845 (N_1845,N_1675,N_1692);
nand U1846 (N_1846,N_1714,N_1581);
xor U1847 (N_1847,N_1593,N_1542);
and U1848 (N_1848,N_1564,N_1634);
xor U1849 (N_1849,N_1647,N_1741);
nand U1850 (N_1850,N_1597,N_1591);
and U1851 (N_1851,N_1515,N_1638);
and U1852 (N_1852,N_1549,N_1627);
nor U1853 (N_1853,N_1659,N_1630);
xor U1854 (N_1854,N_1595,N_1500);
and U1855 (N_1855,N_1580,N_1654);
or U1856 (N_1856,N_1636,N_1712);
nand U1857 (N_1857,N_1722,N_1632);
and U1858 (N_1858,N_1503,N_1605);
nand U1859 (N_1859,N_1730,N_1563);
and U1860 (N_1860,N_1513,N_1695);
nand U1861 (N_1861,N_1648,N_1601);
xor U1862 (N_1862,N_1660,N_1583);
nor U1863 (N_1863,N_1550,N_1731);
nor U1864 (N_1864,N_1529,N_1525);
nand U1865 (N_1865,N_1690,N_1616);
nor U1866 (N_1866,N_1650,N_1694);
nand U1867 (N_1867,N_1608,N_1699);
and U1868 (N_1868,N_1539,N_1575);
nor U1869 (N_1869,N_1628,N_1720);
or U1870 (N_1870,N_1511,N_1620);
nand U1871 (N_1871,N_1555,N_1667);
and U1872 (N_1872,N_1558,N_1721);
nand U1873 (N_1873,N_1657,N_1554);
nor U1874 (N_1874,N_1552,N_1696);
and U1875 (N_1875,N_1737,N_1739);
or U1876 (N_1876,N_1691,N_1609);
nor U1877 (N_1877,N_1557,N_1534);
nor U1878 (N_1878,N_1515,N_1633);
xor U1879 (N_1879,N_1709,N_1689);
or U1880 (N_1880,N_1692,N_1557);
nor U1881 (N_1881,N_1598,N_1583);
or U1882 (N_1882,N_1668,N_1679);
xor U1883 (N_1883,N_1584,N_1628);
nor U1884 (N_1884,N_1572,N_1658);
xor U1885 (N_1885,N_1733,N_1637);
nor U1886 (N_1886,N_1614,N_1693);
or U1887 (N_1887,N_1739,N_1647);
nand U1888 (N_1888,N_1662,N_1520);
nand U1889 (N_1889,N_1580,N_1561);
xnor U1890 (N_1890,N_1727,N_1680);
nor U1891 (N_1891,N_1505,N_1652);
or U1892 (N_1892,N_1517,N_1677);
and U1893 (N_1893,N_1658,N_1690);
nand U1894 (N_1894,N_1523,N_1581);
nand U1895 (N_1895,N_1648,N_1687);
or U1896 (N_1896,N_1545,N_1625);
nand U1897 (N_1897,N_1596,N_1568);
and U1898 (N_1898,N_1552,N_1516);
or U1899 (N_1899,N_1501,N_1605);
or U1900 (N_1900,N_1525,N_1514);
and U1901 (N_1901,N_1642,N_1586);
and U1902 (N_1902,N_1738,N_1619);
nand U1903 (N_1903,N_1637,N_1528);
nand U1904 (N_1904,N_1684,N_1617);
nor U1905 (N_1905,N_1543,N_1657);
and U1906 (N_1906,N_1598,N_1608);
nor U1907 (N_1907,N_1708,N_1568);
or U1908 (N_1908,N_1601,N_1703);
and U1909 (N_1909,N_1502,N_1641);
nor U1910 (N_1910,N_1617,N_1643);
nand U1911 (N_1911,N_1680,N_1616);
or U1912 (N_1912,N_1624,N_1649);
nand U1913 (N_1913,N_1656,N_1510);
nor U1914 (N_1914,N_1546,N_1611);
nor U1915 (N_1915,N_1629,N_1697);
xnor U1916 (N_1916,N_1522,N_1708);
and U1917 (N_1917,N_1599,N_1701);
or U1918 (N_1918,N_1557,N_1539);
or U1919 (N_1919,N_1593,N_1612);
nor U1920 (N_1920,N_1602,N_1727);
nor U1921 (N_1921,N_1688,N_1510);
or U1922 (N_1922,N_1508,N_1724);
xor U1923 (N_1923,N_1695,N_1634);
nand U1924 (N_1924,N_1524,N_1563);
xor U1925 (N_1925,N_1575,N_1657);
or U1926 (N_1926,N_1743,N_1537);
nor U1927 (N_1927,N_1728,N_1707);
and U1928 (N_1928,N_1712,N_1527);
or U1929 (N_1929,N_1664,N_1688);
xor U1930 (N_1930,N_1620,N_1738);
nand U1931 (N_1931,N_1614,N_1695);
xnor U1932 (N_1932,N_1616,N_1536);
or U1933 (N_1933,N_1535,N_1713);
nand U1934 (N_1934,N_1643,N_1668);
or U1935 (N_1935,N_1746,N_1521);
or U1936 (N_1936,N_1646,N_1661);
xor U1937 (N_1937,N_1661,N_1731);
nor U1938 (N_1938,N_1668,N_1727);
nor U1939 (N_1939,N_1509,N_1740);
and U1940 (N_1940,N_1546,N_1574);
or U1941 (N_1941,N_1749,N_1650);
and U1942 (N_1942,N_1717,N_1563);
nand U1943 (N_1943,N_1624,N_1625);
nor U1944 (N_1944,N_1553,N_1651);
xor U1945 (N_1945,N_1656,N_1560);
xnor U1946 (N_1946,N_1625,N_1667);
or U1947 (N_1947,N_1646,N_1727);
nand U1948 (N_1948,N_1582,N_1670);
nand U1949 (N_1949,N_1601,N_1745);
and U1950 (N_1950,N_1507,N_1630);
or U1951 (N_1951,N_1701,N_1702);
nand U1952 (N_1952,N_1613,N_1645);
nor U1953 (N_1953,N_1656,N_1703);
nor U1954 (N_1954,N_1545,N_1514);
xnor U1955 (N_1955,N_1667,N_1637);
nand U1956 (N_1956,N_1612,N_1537);
nand U1957 (N_1957,N_1596,N_1689);
nand U1958 (N_1958,N_1559,N_1730);
xnor U1959 (N_1959,N_1717,N_1747);
nand U1960 (N_1960,N_1683,N_1558);
xnor U1961 (N_1961,N_1527,N_1564);
or U1962 (N_1962,N_1505,N_1579);
nand U1963 (N_1963,N_1696,N_1589);
nand U1964 (N_1964,N_1541,N_1708);
nor U1965 (N_1965,N_1595,N_1531);
and U1966 (N_1966,N_1698,N_1626);
nand U1967 (N_1967,N_1591,N_1634);
and U1968 (N_1968,N_1712,N_1745);
nor U1969 (N_1969,N_1551,N_1597);
or U1970 (N_1970,N_1629,N_1621);
xnor U1971 (N_1971,N_1574,N_1669);
or U1972 (N_1972,N_1712,N_1535);
and U1973 (N_1973,N_1514,N_1637);
nor U1974 (N_1974,N_1519,N_1733);
xor U1975 (N_1975,N_1515,N_1634);
nand U1976 (N_1976,N_1731,N_1669);
or U1977 (N_1977,N_1558,N_1607);
nand U1978 (N_1978,N_1582,N_1728);
nand U1979 (N_1979,N_1679,N_1697);
and U1980 (N_1980,N_1725,N_1585);
nand U1981 (N_1981,N_1731,N_1665);
and U1982 (N_1982,N_1687,N_1532);
nand U1983 (N_1983,N_1614,N_1682);
or U1984 (N_1984,N_1564,N_1503);
xnor U1985 (N_1985,N_1701,N_1533);
nor U1986 (N_1986,N_1595,N_1532);
or U1987 (N_1987,N_1668,N_1519);
or U1988 (N_1988,N_1723,N_1665);
xor U1989 (N_1989,N_1704,N_1662);
xnor U1990 (N_1990,N_1574,N_1506);
or U1991 (N_1991,N_1629,N_1618);
nand U1992 (N_1992,N_1658,N_1585);
or U1993 (N_1993,N_1556,N_1565);
xnor U1994 (N_1994,N_1560,N_1609);
and U1995 (N_1995,N_1647,N_1745);
nor U1996 (N_1996,N_1525,N_1594);
or U1997 (N_1997,N_1647,N_1708);
nand U1998 (N_1998,N_1674,N_1543);
xor U1999 (N_1999,N_1701,N_1530);
and U2000 (N_2000,N_1964,N_1810);
xnor U2001 (N_2001,N_1985,N_1843);
nand U2002 (N_2002,N_1910,N_1992);
nor U2003 (N_2003,N_1962,N_1833);
and U2004 (N_2004,N_1914,N_1872);
nor U2005 (N_2005,N_1887,N_1926);
and U2006 (N_2006,N_1867,N_1956);
nand U2007 (N_2007,N_1850,N_1915);
nand U2008 (N_2008,N_1870,N_1827);
xor U2009 (N_2009,N_1883,N_1969);
nand U2010 (N_2010,N_1873,N_1800);
and U2011 (N_2011,N_1788,N_1866);
and U2012 (N_2012,N_1756,N_1909);
or U2013 (N_2013,N_1903,N_1752);
or U2014 (N_2014,N_1841,N_1812);
nand U2015 (N_2015,N_1929,N_1894);
and U2016 (N_2016,N_1899,N_1967);
and U2017 (N_2017,N_1806,N_1973);
and U2018 (N_2018,N_1905,N_1759);
or U2019 (N_2019,N_1983,N_1953);
xnor U2020 (N_2020,N_1977,N_1880);
nand U2021 (N_2021,N_1842,N_1796);
or U2022 (N_2022,N_1837,N_1943);
nor U2023 (N_2023,N_1978,N_1811);
and U2024 (N_2024,N_1789,N_1881);
or U2025 (N_2025,N_1922,N_1911);
nand U2026 (N_2026,N_1938,N_1819);
xor U2027 (N_2027,N_1888,N_1805);
xor U2028 (N_2028,N_1890,N_1908);
or U2029 (N_2029,N_1774,N_1942);
xor U2030 (N_2030,N_1767,N_1856);
nand U2031 (N_2031,N_1944,N_1802);
and U2032 (N_2032,N_1982,N_1923);
nand U2033 (N_2033,N_1885,N_1831);
nand U2034 (N_2034,N_1772,N_1935);
nand U2035 (N_2035,N_1751,N_1766);
nor U2036 (N_2036,N_1879,N_1989);
nor U2037 (N_2037,N_1927,N_1864);
or U2038 (N_2038,N_1886,N_1750);
nor U2039 (N_2039,N_1844,N_1892);
and U2040 (N_2040,N_1994,N_1845);
or U2041 (N_2041,N_1853,N_1839);
or U2042 (N_2042,N_1986,N_1959);
and U2043 (N_2043,N_1895,N_1787);
nand U2044 (N_2044,N_1778,N_1808);
and U2045 (N_2045,N_1893,N_1999);
nor U2046 (N_2046,N_1835,N_1768);
nand U2047 (N_2047,N_1813,N_1777);
nand U2048 (N_2048,N_1821,N_1940);
nor U2049 (N_2049,N_1794,N_1945);
and U2050 (N_2050,N_1975,N_1960);
or U2051 (N_2051,N_1901,N_1939);
nand U2052 (N_2052,N_1790,N_1784);
nor U2053 (N_2053,N_1814,N_1912);
nand U2054 (N_2054,N_1775,N_1776);
or U2055 (N_2055,N_1980,N_1990);
or U2056 (N_2056,N_1884,N_1765);
nand U2057 (N_2057,N_1902,N_1852);
nand U2058 (N_2058,N_1836,N_1921);
xor U2059 (N_2059,N_1848,N_1898);
nand U2060 (N_2060,N_1861,N_1770);
xor U2061 (N_2061,N_1854,N_1987);
nor U2062 (N_2062,N_1968,N_1906);
nor U2063 (N_2063,N_1920,N_1809);
nor U2064 (N_2064,N_1930,N_1860);
or U2065 (N_2065,N_1838,N_1798);
and U2066 (N_2066,N_1760,N_1781);
nor U2067 (N_2067,N_1971,N_1807);
nor U2068 (N_2068,N_1791,N_1993);
nand U2069 (N_2069,N_1826,N_1937);
and U2070 (N_2070,N_1928,N_1825);
xnor U2071 (N_2071,N_1823,N_1782);
nor U2072 (N_2072,N_1761,N_1851);
and U2073 (N_2073,N_1830,N_1769);
xor U2074 (N_2074,N_1995,N_1832);
and U2075 (N_2075,N_1965,N_1828);
and U2076 (N_2076,N_1780,N_1869);
xor U2077 (N_2077,N_1815,N_1816);
and U2078 (N_2078,N_1952,N_1981);
xor U2079 (N_2079,N_1858,N_1803);
nor U2080 (N_2080,N_1896,N_1755);
and U2081 (N_2081,N_1931,N_1984);
nor U2082 (N_2082,N_1793,N_1829);
nor U2083 (N_2083,N_1855,N_1795);
or U2084 (N_2084,N_1877,N_1916);
xor U2085 (N_2085,N_1865,N_1979);
xnor U2086 (N_2086,N_1868,N_1950);
nand U2087 (N_2087,N_1785,N_1976);
xnor U2088 (N_2088,N_1941,N_1924);
xnor U2089 (N_2089,N_1970,N_1773);
or U2090 (N_2090,N_1919,N_1949);
xnor U2091 (N_2091,N_1801,N_1817);
nand U2092 (N_2092,N_1972,N_1988);
or U2093 (N_2093,N_1934,N_1834);
and U2094 (N_2094,N_1840,N_1786);
nand U2095 (N_2095,N_1974,N_1875);
and U2096 (N_2096,N_1997,N_1862);
nand U2097 (N_2097,N_1783,N_1996);
nor U2098 (N_2098,N_1925,N_1891);
nor U2099 (N_2099,N_1753,N_1900);
xnor U2100 (N_2100,N_1889,N_1874);
and U2101 (N_2101,N_1792,N_1754);
nand U2102 (N_2102,N_1932,N_1824);
nand U2103 (N_2103,N_1918,N_1955);
and U2104 (N_2104,N_1913,N_1762);
or U2105 (N_2105,N_1863,N_1820);
or U2106 (N_2106,N_1946,N_1882);
or U2107 (N_2107,N_1763,N_1947);
and U2108 (N_2108,N_1779,N_1847);
nor U2109 (N_2109,N_1871,N_1958);
xnor U2110 (N_2110,N_1917,N_1991);
nand U2111 (N_2111,N_1936,N_1878);
or U2112 (N_2112,N_1897,N_1876);
xnor U2113 (N_2113,N_1907,N_1857);
nor U2114 (N_2114,N_1966,N_1764);
or U2115 (N_2115,N_1757,N_1963);
or U2116 (N_2116,N_1951,N_1933);
and U2117 (N_2117,N_1758,N_1957);
and U2118 (N_2118,N_1948,N_1771);
nand U2119 (N_2119,N_1954,N_1799);
and U2120 (N_2120,N_1961,N_1822);
and U2121 (N_2121,N_1849,N_1998);
xor U2122 (N_2122,N_1846,N_1797);
and U2123 (N_2123,N_1804,N_1859);
nand U2124 (N_2124,N_1818,N_1904);
xnor U2125 (N_2125,N_1906,N_1964);
or U2126 (N_2126,N_1893,N_1796);
xor U2127 (N_2127,N_1867,N_1852);
nor U2128 (N_2128,N_1752,N_1921);
xor U2129 (N_2129,N_1767,N_1925);
nand U2130 (N_2130,N_1797,N_1813);
nor U2131 (N_2131,N_1951,N_1786);
or U2132 (N_2132,N_1754,N_1918);
or U2133 (N_2133,N_1791,N_1876);
xor U2134 (N_2134,N_1912,N_1913);
xor U2135 (N_2135,N_1985,N_1917);
and U2136 (N_2136,N_1971,N_1954);
nor U2137 (N_2137,N_1953,N_1820);
nor U2138 (N_2138,N_1785,N_1884);
nand U2139 (N_2139,N_1790,N_1909);
or U2140 (N_2140,N_1756,N_1802);
xnor U2141 (N_2141,N_1828,N_1796);
xnor U2142 (N_2142,N_1766,N_1783);
or U2143 (N_2143,N_1887,N_1888);
or U2144 (N_2144,N_1815,N_1870);
nor U2145 (N_2145,N_1950,N_1770);
nor U2146 (N_2146,N_1915,N_1819);
nand U2147 (N_2147,N_1762,N_1962);
xor U2148 (N_2148,N_1812,N_1967);
xnor U2149 (N_2149,N_1801,N_1887);
nand U2150 (N_2150,N_1804,N_1974);
nor U2151 (N_2151,N_1909,N_1936);
nand U2152 (N_2152,N_1942,N_1854);
nor U2153 (N_2153,N_1938,N_1931);
nor U2154 (N_2154,N_1822,N_1984);
xor U2155 (N_2155,N_1809,N_1885);
nand U2156 (N_2156,N_1932,N_1843);
xor U2157 (N_2157,N_1794,N_1871);
and U2158 (N_2158,N_1942,N_1821);
nand U2159 (N_2159,N_1828,N_1916);
nand U2160 (N_2160,N_1817,N_1891);
or U2161 (N_2161,N_1908,N_1800);
or U2162 (N_2162,N_1918,N_1803);
or U2163 (N_2163,N_1947,N_1942);
and U2164 (N_2164,N_1791,N_1917);
and U2165 (N_2165,N_1761,N_1821);
xnor U2166 (N_2166,N_1802,N_1892);
nand U2167 (N_2167,N_1778,N_1871);
nand U2168 (N_2168,N_1830,N_1773);
nor U2169 (N_2169,N_1860,N_1911);
or U2170 (N_2170,N_1999,N_1986);
xor U2171 (N_2171,N_1932,N_1835);
and U2172 (N_2172,N_1907,N_1848);
nand U2173 (N_2173,N_1885,N_1882);
nand U2174 (N_2174,N_1778,N_1955);
or U2175 (N_2175,N_1912,N_1966);
nand U2176 (N_2176,N_1758,N_1903);
nor U2177 (N_2177,N_1891,N_1800);
nand U2178 (N_2178,N_1805,N_1860);
or U2179 (N_2179,N_1760,N_1787);
nand U2180 (N_2180,N_1865,N_1802);
nor U2181 (N_2181,N_1796,N_1752);
xnor U2182 (N_2182,N_1821,N_1772);
xor U2183 (N_2183,N_1833,N_1906);
xnor U2184 (N_2184,N_1969,N_1934);
or U2185 (N_2185,N_1765,N_1825);
or U2186 (N_2186,N_1853,N_1775);
xor U2187 (N_2187,N_1777,N_1984);
nor U2188 (N_2188,N_1841,N_1969);
or U2189 (N_2189,N_1945,N_1813);
xnor U2190 (N_2190,N_1819,N_1870);
nor U2191 (N_2191,N_1962,N_1924);
xnor U2192 (N_2192,N_1750,N_1903);
nor U2193 (N_2193,N_1989,N_1853);
nor U2194 (N_2194,N_1767,N_1878);
nand U2195 (N_2195,N_1854,N_1943);
or U2196 (N_2196,N_1832,N_1782);
xor U2197 (N_2197,N_1902,N_1790);
and U2198 (N_2198,N_1848,N_1962);
nor U2199 (N_2199,N_1911,N_1811);
nand U2200 (N_2200,N_1978,N_1850);
or U2201 (N_2201,N_1816,N_1840);
nor U2202 (N_2202,N_1853,N_1822);
nand U2203 (N_2203,N_1974,N_1836);
nor U2204 (N_2204,N_1924,N_1930);
or U2205 (N_2205,N_1829,N_1889);
xnor U2206 (N_2206,N_1820,N_1847);
or U2207 (N_2207,N_1919,N_1787);
nor U2208 (N_2208,N_1762,N_1971);
or U2209 (N_2209,N_1877,N_1948);
or U2210 (N_2210,N_1782,N_1921);
or U2211 (N_2211,N_1867,N_1954);
nand U2212 (N_2212,N_1855,N_1802);
nand U2213 (N_2213,N_1768,N_1986);
nand U2214 (N_2214,N_1771,N_1990);
nor U2215 (N_2215,N_1851,N_1962);
or U2216 (N_2216,N_1994,N_1892);
xnor U2217 (N_2217,N_1877,N_1801);
nor U2218 (N_2218,N_1868,N_1954);
and U2219 (N_2219,N_1894,N_1858);
nand U2220 (N_2220,N_1861,N_1790);
nand U2221 (N_2221,N_1971,N_1784);
and U2222 (N_2222,N_1903,N_1960);
or U2223 (N_2223,N_1896,N_1821);
nor U2224 (N_2224,N_1947,N_1757);
nor U2225 (N_2225,N_1897,N_1880);
nand U2226 (N_2226,N_1837,N_1978);
and U2227 (N_2227,N_1834,N_1803);
or U2228 (N_2228,N_1900,N_1928);
or U2229 (N_2229,N_1908,N_1874);
and U2230 (N_2230,N_1897,N_1756);
or U2231 (N_2231,N_1779,N_1767);
nand U2232 (N_2232,N_1809,N_1807);
nor U2233 (N_2233,N_1758,N_1765);
or U2234 (N_2234,N_1866,N_1776);
nand U2235 (N_2235,N_1757,N_1821);
and U2236 (N_2236,N_1807,N_1850);
xnor U2237 (N_2237,N_1935,N_1883);
xnor U2238 (N_2238,N_1993,N_1806);
and U2239 (N_2239,N_1760,N_1932);
nand U2240 (N_2240,N_1947,N_1937);
and U2241 (N_2241,N_1875,N_1835);
and U2242 (N_2242,N_1912,N_1842);
xnor U2243 (N_2243,N_1803,N_1924);
or U2244 (N_2244,N_1892,N_1846);
nor U2245 (N_2245,N_1935,N_1869);
or U2246 (N_2246,N_1966,N_1798);
and U2247 (N_2247,N_1903,N_1893);
nand U2248 (N_2248,N_1939,N_1944);
nand U2249 (N_2249,N_1810,N_1995);
xnor U2250 (N_2250,N_2187,N_2195);
nor U2251 (N_2251,N_2207,N_2124);
nand U2252 (N_2252,N_2192,N_2050);
nor U2253 (N_2253,N_2115,N_2020);
or U2254 (N_2254,N_2044,N_2132);
nand U2255 (N_2255,N_2019,N_2218);
and U2256 (N_2256,N_2016,N_2228);
and U2257 (N_2257,N_2152,N_2085);
nor U2258 (N_2258,N_2236,N_2137);
and U2259 (N_2259,N_2076,N_2173);
and U2260 (N_2260,N_2186,N_2081);
and U2261 (N_2261,N_2133,N_2119);
and U2262 (N_2262,N_2143,N_2015);
or U2263 (N_2263,N_2047,N_2151);
nand U2264 (N_2264,N_2175,N_2042);
xnor U2265 (N_2265,N_2178,N_2031);
nor U2266 (N_2266,N_2247,N_2083);
xor U2267 (N_2267,N_2208,N_2048);
nand U2268 (N_2268,N_2161,N_2017);
and U2269 (N_2269,N_2146,N_2136);
nand U2270 (N_2270,N_2166,N_2026);
nand U2271 (N_2271,N_2204,N_2191);
or U2272 (N_2272,N_2174,N_2006);
and U2273 (N_2273,N_2172,N_2093);
or U2274 (N_2274,N_2056,N_2153);
nand U2275 (N_2275,N_2231,N_2002);
and U2276 (N_2276,N_2025,N_2205);
nor U2277 (N_2277,N_2194,N_2011);
or U2278 (N_2278,N_2080,N_2127);
or U2279 (N_2279,N_2176,N_2032);
or U2280 (N_2280,N_2033,N_2067);
nand U2281 (N_2281,N_2165,N_2149);
nand U2282 (N_2282,N_2217,N_2230);
xor U2283 (N_2283,N_2206,N_2144);
nor U2284 (N_2284,N_2224,N_2053);
or U2285 (N_2285,N_2037,N_2167);
nor U2286 (N_2286,N_2180,N_2227);
nor U2287 (N_2287,N_2241,N_2156);
or U2288 (N_2288,N_2084,N_2128);
xnor U2289 (N_2289,N_2045,N_2116);
or U2290 (N_2290,N_2125,N_2014);
nand U2291 (N_2291,N_2065,N_2185);
xor U2292 (N_2292,N_2160,N_2063);
xor U2293 (N_2293,N_2130,N_2069);
and U2294 (N_2294,N_2029,N_2100);
nand U2295 (N_2295,N_2052,N_2216);
nand U2296 (N_2296,N_2072,N_2077);
or U2297 (N_2297,N_2070,N_2009);
or U2298 (N_2298,N_2121,N_2196);
xor U2299 (N_2299,N_2079,N_2168);
nand U2300 (N_2300,N_2066,N_2030);
nor U2301 (N_2301,N_2117,N_2169);
or U2302 (N_2302,N_2007,N_2041);
xor U2303 (N_2303,N_2222,N_2059);
xor U2304 (N_2304,N_2145,N_2091);
xor U2305 (N_2305,N_2107,N_2110);
and U2306 (N_2306,N_2109,N_2181);
or U2307 (N_2307,N_2098,N_2082);
nor U2308 (N_2308,N_2162,N_2104);
xnor U2309 (N_2309,N_2038,N_2234);
and U2310 (N_2310,N_2183,N_2113);
or U2311 (N_2311,N_2164,N_2012);
nor U2312 (N_2312,N_2068,N_2248);
or U2313 (N_2313,N_2190,N_2213);
nand U2314 (N_2314,N_2086,N_2158);
nand U2315 (N_2315,N_2060,N_2090);
nand U2316 (N_2316,N_2058,N_2154);
or U2317 (N_2317,N_2046,N_2106);
or U2318 (N_2318,N_2170,N_2103);
nor U2319 (N_2319,N_2035,N_2078);
or U2320 (N_2320,N_2142,N_2123);
nand U2321 (N_2321,N_2022,N_2120);
or U2322 (N_2322,N_2099,N_2000);
and U2323 (N_2323,N_2075,N_2027);
and U2324 (N_2324,N_2220,N_2249);
nand U2325 (N_2325,N_2242,N_2126);
nor U2326 (N_2326,N_2232,N_2102);
xor U2327 (N_2327,N_2157,N_2054);
xor U2328 (N_2328,N_2237,N_2193);
xor U2329 (N_2329,N_2214,N_2074);
nor U2330 (N_2330,N_2159,N_2095);
xnor U2331 (N_2331,N_2004,N_2049);
and U2332 (N_2332,N_2036,N_2182);
and U2333 (N_2333,N_2163,N_2094);
and U2334 (N_2334,N_2245,N_2171);
nand U2335 (N_2335,N_2051,N_2097);
nand U2336 (N_2336,N_2088,N_2219);
xor U2337 (N_2337,N_2221,N_2005);
nand U2338 (N_2338,N_2062,N_2189);
nor U2339 (N_2339,N_2039,N_2118);
xor U2340 (N_2340,N_2010,N_2024);
or U2341 (N_2341,N_2210,N_2244);
nand U2342 (N_2342,N_2135,N_2021);
or U2343 (N_2343,N_2089,N_2003);
and U2344 (N_2344,N_2018,N_2223);
nand U2345 (N_2345,N_2071,N_2229);
nand U2346 (N_2346,N_2201,N_2200);
nand U2347 (N_2347,N_2243,N_2246);
xnor U2348 (N_2348,N_2202,N_2138);
xor U2349 (N_2349,N_2199,N_2105);
nand U2350 (N_2350,N_2008,N_2134);
and U2351 (N_2351,N_2238,N_2028);
nor U2352 (N_2352,N_2096,N_2226);
and U2353 (N_2353,N_2055,N_2212);
and U2354 (N_2354,N_2139,N_2179);
nand U2355 (N_2355,N_2203,N_2155);
xor U2356 (N_2356,N_2073,N_2197);
nor U2357 (N_2357,N_2188,N_2064);
and U2358 (N_2358,N_2225,N_2112);
nand U2359 (N_2359,N_2215,N_2147);
nand U2360 (N_2360,N_2040,N_2184);
or U2361 (N_2361,N_2023,N_2092);
xnor U2362 (N_2362,N_2061,N_2240);
and U2363 (N_2363,N_2239,N_2198);
nor U2364 (N_2364,N_2108,N_2101);
nand U2365 (N_2365,N_2087,N_2114);
or U2366 (N_2366,N_2129,N_2122);
xnor U2367 (N_2367,N_2235,N_2150);
nor U2368 (N_2368,N_2233,N_2057);
or U2369 (N_2369,N_2034,N_2209);
or U2370 (N_2370,N_2013,N_2043);
nand U2371 (N_2371,N_2141,N_2177);
and U2372 (N_2372,N_2131,N_2001);
nor U2373 (N_2373,N_2111,N_2211);
nor U2374 (N_2374,N_2140,N_2148);
or U2375 (N_2375,N_2194,N_2242);
or U2376 (N_2376,N_2029,N_2197);
xor U2377 (N_2377,N_2123,N_2235);
nand U2378 (N_2378,N_2210,N_2184);
xor U2379 (N_2379,N_2113,N_2073);
nor U2380 (N_2380,N_2011,N_2036);
and U2381 (N_2381,N_2211,N_2219);
xnor U2382 (N_2382,N_2174,N_2177);
nand U2383 (N_2383,N_2047,N_2061);
xor U2384 (N_2384,N_2109,N_2171);
or U2385 (N_2385,N_2192,N_2241);
or U2386 (N_2386,N_2177,N_2180);
nand U2387 (N_2387,N_2244,N_2046);
nand U2388 (N_2388,N_2017,N_2041);
nor U2389 (N_2389,N_2010,N_2055);
and U2390 (N_2390,N_2182,N_2228);
or U2391 (N_2391,N_2205,N_2186);
and U2392 (N_2392,N_2206,N_2075);
nor U2393 (N_2393,N_2120,N_2204);
or U2394 (N_2394,N_2040,N_2135);
xor U2395 (N_2395,N_2043,N_2091);
and U2396 (N_2396,N_2132,N_2151);
or U2397 (N_2397,N_2120,N_2207);
or U2398 (N_2398,N_2063,N_2078);
nor U2399 (N_2399,N_2054,N_2194);
nand U2400 (N_2400,N_2180,N_2182);
and U2401 (N_2401,N_2228,N_2086);
and U2402 (N_2402,N_2205,N_2160);
nor U2403 (N_2403,N_2180,N_2150);
nor U2404 (N_2404,N_2189,N_2035);
xor U2405 (N_2405,N_2241,N_2174);
nand U2406 (N_2406,N_2156,N_2140);
or U2407 (N_2407,N_2160,N_2234);
nand U2408 (N_2408,N_2049,N_2245);
xor U2409 (N_2409,N_2214,N_2152);
nand U2410 (N_2410,N_2056,N_2221);
and U2411 (N_2411,N_2145,N_2138);
and U2412 (N_2412,N_2230,N_2215);
xnor U2413 (N_2413,N_2010,N_2072);
nor U2414 (N_2414,N_2009,N_2127);
xor U2415 (N_2415,N_2006,N_2100);
or U2416 (N_2416,N_2004,N_2178);
or U2417 (N_2417,N_2228,N_2024);
nand U2418 (N_2418,N_2192,N_2122);
xnor U2419 (N_2419,N_2122,N_2184);
nor U2420 (N_2420,N_2134,N_2024);
or U2421 (N_2421,N_2187,N_2208);
nand U2422 (N_2422,N_2042,N_2170);
nor U2423 (N_2423,N_2024,N_2218);
and U2424 (N_2424,N_2223,N_2147);
xor U2425 (N_2425,N_2219,N_2163);
and U2426 (N_2426,N_2161,N_2228);
or U2427 (N_2427,N_2010,N_2126);
or U2428 (N_2428,N_2023,N_2037);
xor U2429 (N_2429,N_2080,N_2148);
or U2430 (N_2430,N_2183,N_2046);
nand U2431 (N_2431,N_2099,N_2032);
or U2432 (N_2432,N_2123,N_2000);
nand U2433 (N_2433,N_2193,N_2057);
xnor U2434 (N_2434,N_2168,N_2023);
xnor U2435 (N_2435,N_2120,N_2115);
nand U2436 (N_2436,N_2230,N_2114);
nand U2437 (N_2437,N_2110,N_2051);
and U2438 (N_2438,N_2215,N_2154);
and U2439 (N_2439,N_2195,N_2176);
nand U2440 (N_2440,N_2238,N_2075);
and U2441 (N_2441,N_2163,N_2147);
or U2442 (N_2442,N_2094,N_2014);
nor U2443 (N_2443,N_2242,N_2074);
nand U2444 (N_2444,N_2076,N_2095);
xnor U2445 (N_2445,N_2143,N_2044);
nand U2446 (N_2446,N_2203,N_2114);
and U2447 (N_2447,N_2181,N_2122);
nor U2448 (N_2448,N_2152,N_2105);
or U2449 (N_2449,N_2234,N_2217);
or U2450 (N_2450,N_2015,N_2219);
or U2451 (N_2451,N_2067,N_2051);
nor U2452 (N_2452,N_2019,N_2234);
nand U2453 (N_2453,N_2224,N_2136);
xor U2454 (N_2454,N_2105,N_2040);
nand U2455 (N_2455,N_2097,N_2090);
and U2456 (N_2456,N_2017,N_2163);
nor U2457 (N_2457,N_2234,N_2064);
or U2458 (N_2458,N_2081,N_2049);
nor U2459 (N_2459,N_2128,N_2094);
and U2460 (N_2460,N_2018,N_2033);
or U2461 (N_2461,N_2066,N_2147);
xor U2462 (N_2462,N_2246,N_2186);
and U2463 (N_2463,N_2190,N_2237);
and U2464 (N_2464,N_2150,N_2073);
nand U2465 (N_2465,N_2116,N_2041);
and U2466 (N_2466,N_2197,N_2142);
and U2467 (N_2467,N_2195,N_2026);
nor U2468 (N_2468,N_2137,N_2117);
nand U2469 (N_2469,N_2079,N_2189);
or U2470 (N_2470,N_2134,N_2139);
or U2471 (N_2471,N_2167,N_2090);
and U2472 (N_2472,N_2086,N_2171);
or U2473 (N_2473,N_2240,N_2225);
nor U2474 (N_2474,N_2158,N_2209);
nand U2475 (N_2475,N_2188,N_2138);
xnor U2476 (N_2476,N_2003,N_2186);
or U2477 (N_2477,N_2178,N_2179);
or U2478 (N_2478,N_2197,N_2085);
nand U2479 (N_2479,N_2230,N_2111);
and U2480 (N_2480,N_2113,N_2236);
xor U2481 (N_2481,N_2025,N_2096);
and U2482 (N_2482,N_2083,N_2209);
nor U2483 (N_2483,N_2095,N_2183);
nand U2484 (N_2484,N_2011,N_2097);
nor U2485 (N_2485,N_2231,N_2075);
or U2486 (N_2486,N_2057,N_2128);
nor U2487 (N_2487,N_2211,N_2204);
or U2488 (N_2488,N_2231,N_2086);
and U2489 (N_2489,N_2116,N_2098);
and U2490 (N_2490,N_2152,N_2176);
nor U2491 (N_2491,N_2187,N_2221);
nor U2492 (N_2492,N_2106,N_2103);
xnor U2493 (N_2493,N_2021,N_2110);
xor U2494 (N_2494,N_2009,N_2063);
xnor U2495 (N_2495,N_2123,N_2003);
xnor U2496 (N_2496,N_2066,N_2198);
xor U2497 (N_2497,N_2074,N_2227);
xor U2498 (N_2498,N_2217,N_2086);
nand U2499 (N_2499,N_2220,N_2080);
nand U2500 (N_2500,N_2471,N_2287);
nor U2501 (N_2501,N_2261,N_2340);
nand U2502 (N_2502,N_2482,N_2290);
and U2503 (N_2503,N_2251,N_2385);
or U2504 (N_2504,N_2318,N_2322);
and U2505 (N_2505,N_2352,N_2497);
xnor U2506 (N_2506,N_2462,N_2461);
nor U2507 (N_2507,N_2275,N_2380);
nand U2508 (N_2508,N_2400,N_2439);
nor U2509 (N_2509,N_2425,N_2337);
or U2510 (N_2510,N_2296,N_2323);
nor U2511 (N_2511,N_2445,N_2263);
and U2512 (N_2512,N_2386,N_2269);
nand U2513 (N_2513,N_2257,N_2405);
or U2514 (N_2514,N_2419,N_2272);
and U2515 (N_2515,N_2343,N_2372);
and U2516 (N_2516,N_2452,N_2265);
nor U2517 (N_2517,N_2448,N_2442);
nand U2518 (N_2518,N_2381,N_2331);
nand U2519 (N_2519,N_2488,N_2361);
and U2520 (N_2520,N_2390,N_2464);
nand U2521 (N_2521,N_2431,N_2324);
and U2522 (N_2522,N_2301,N_2481);
or U2523 (N_2523,N_2271,N_2449);
nor U2524 (N_2524,N_2313,N_2455);
and U2525 (N_2525,N_2289,N_2293);
nand U2526 (N_2526,N_2438,N_2491);
and U2527 (N_2527,N_2451,N_2432);
xnor U2528 (N_2528,N_2256,N_2463);
or U2529 (N_2529,N_2410,N_2396);
xor U2530 (N_2530,N_2260,N_2298);
nor U2531 (N_2531,N_2268,N_2344);
nor U2532 (N_2532,N_2255,N_2294);
nand U2533 (N_2533,N_2364,N_2387);
xnor U2534 (N_2534,N_2404,N_2474);
nor U2535 (N_2535,N_2466,N_2366);
nor U2536 (N_2536,N_2490,N_2310);
nand U2537 (N_2537,N_2341,N_2330);
and U2538 (N_2538,N_2456,N_2435);
and U2539 (N_2539,N_2373,N_2424);
or U2540 (N_2540,N_2311,N_2370);
xor U2541 (N_2541,N_2300,N_2483);
nor U2542 (N_2542,N_2325,N_2258);
and U2543 (N_2543,N_2351,N_2363);
xnor U2544 (N_2544,N_2430,N_2412);
nor U2545 (N_2545,N_2409,N_2327);
nand U2546 (N_2546,N_2468,N_2357);
and U2547 (N_2547,N_2349,N_2414);
and U2548 (N_2548,N_2319,N_2437);
nand U2549 (N_2549,N_2486,N_2411);
nor U2550 (N_2550,N_2353,N_2454);
xnor U2551 (N_2551,N_2374,N_2329);
xnor U2552 (N_2552,N_2338,N_2479);
or U2553 (N_2553,N_2378,N_2460);
nor U2554 (N_2554,N_2458,N_2253);
nor U2555 (N_2555,N_2434,N_2436);
and U2556 (N_2556,N_2383,N_2484);
nor U2557 (N_2557,N_2459,N_2403);
nor U2558 (N_2558,N_2284,N_2264);
xnor U2559 (N_2559,N_2358,N_2450);
nor U2560 (N_2560,N_2393,N_2391);
xnor U2561 (N_2561,N_2326,N_2428);
nor U2562 (N_2562,N_2427,N_2371);
nor U2563 (N_2563,N_2429,N_2280);
nor U2564 (N_2564,N_2397,N_2346);
xor U2565 (N_2565,N_2467,N_2423);
or U2566 (N_2566,N_2406,N_2274);
nor U2567 (N_2567,N_2267,N_2398);
nor U2568 (N_2568,N_2279,N_2440);
nor U2569 (N_2569,N_2335,N_2498);
and U2570 (N_2570,N_2375,N_2392);
nor U2571 (N_2571,N_2476,N_2312);
xor U2572 (N_2572,N_2288,N_2252);
xor U2573 (N_2573,N_2447,N_2377);
nor U2574 (N_2574,N_2336,N_2356);
nor U2575 (N_2575,N_2382,N_2302);
xor U2576 (N_2576,N_2291,N_2444);
nor U2577 (N_2577,N_2407,N_2369);
or U2578 (N_2578,N_2345,N_2399);
xor U2579 (N_2579,N_2270,N_2266);
nor U2580 (N_2580,N_2443,N_2416);
and U2581 (N_2581,N_2485,N_2250);
nor U2582 (N_2582,N_2283,N_2303);
nand U2583 (N_2583,N_2415,N_2334);
and U2584 (N_2584,N_2295,N_2495);
nor U2585 (N_2585,N_2333,N_2342);
and U2586 (N_2586,N_2308,N_2402);
or U2587 (N_2587,N_2478,N_2394);
nor U2588 (N_2588,N_2388,N_2367);
or U2589 (N_2589,N_2350,N_2473);
or U2590 (N_2590,N_2365,N_2315);
nor U2591 (N_2591,N_2457,N_2305);
nand U2592 (N_2592,N_2276,N_2328);
xor U2593 (N_2593,N_2408,N_2320);
nor U2594 (N_2594,N_2339,N_2332);
nand U2595 (N_2595,N_2477,N_2254);
nor U2596 (N_2596,N_2355,N_2379);
nor U2597 (N_2597,N_2420,N_2489);
nand U2598 (N_2598,N_2306,N_2499);
and U2599 (N_2599,N_2422,N_2309);
nand U2600 (N_2600,N_2354,N_2494);
xor U2601 (N_2601,N_2496,N_2304);
nand U2602 (N_2602,N_2321,N_2472);
nand U2603 (N_2603,N_2465,N_2426);
or U2604 (N_2604,N_2470,N_2384);
nor U2605 (N_2605,N_2389,N_2317);
and U2606 (N_2606,N_2314,N_2347);
xor U2607 (N_2607,N_2273,N_2487);
and U2608 (N_2608,N_2299,N_2259);
or U2609 (N_2609,N_2281,N_2441);
or U2610 (N_2610,N_2446,N_2433);
nor U2611 (N_2611,N_2297,N_2469);
or U2612 (N_2612,N_2316,N_2453);
xnor U2613 (N_2613,N_2307,N_2492);
and U2614 (N_2614,N_2359,N_2262);
xor U2615 (N_2615,N_2421,N_2368);
nor U2616 (N_2616,N_2475,N_2417);
xnor U2617 (N_2617,N_2418,N_2395);
and U2618 (N_2618,N_2278,N_2362);
and U2619 (N_2619,N_2360,N_2480);
and U2620 (N_2620,N_2285,N_2348);
and U2621 (N_2621,N_2376,N_2282);
and U2622 (N_2622,N_2493,N_2286);
nand U2623 (N_2623,N_2413,N_2401);
or U2624 (N_2624,N_2277,N_2292);
and U2625 (N_2625,N_2381,N_2316);
nor U2626 (N_2626,N_2401,N_2488);
and U2627 (N_2627,N_2370,N_2484);
or U2628 (N_2628,N_2415,N_2445);
nor U2629 (N_2629,N_2411,N_2459);
nand U2630 (N_2630,N_2446,N_2418);
xnor U2631 (N_2631,N_2364,N_2457);
or U2632 (N_2632,N_2472,N_2394);
nor U2633 (N_2633,N_2391,N_2273);
nand U2634 (N_2634,N_2483,N_2415);
nor U2635 (N_2635,N_2374,N_2427);
or U2636 (N_2636,N_2251,N_2401);
nor U2637 (N_2637,N_2374,N_2349);
xor U2638 (N_2638,N_2271,N_2313);
or U2639 (N_2639,N_2489,N_2347);
or U2640 (N_2640,N_2275,N_2332);
nor U2641 (N_2641,N_2363,N_2416);
and U2642 (N_2642,N_2355,N_2347);
or U2643 (N_2643,N_2331,N_2444);
or U2644 (N_2644,N_2327,N_2383);
and U2645 (N_2645,N_2406,N_2305);
or U2646 (N_2646,N_2320,N_2309);
xnor U2647 (N_2647,N_2429,N_2455);
and U2648 (N_2648,N_2392,N_2474);
xnor U2649 (N_2649,N_2308,N_2254);
nor U2650 (N_2650,N_2363,N_2274);
nand U2651 (N_2651,N_2257,N_2415);
xnor U2652 (N_2652,N_2308,N_2251);
nor U2653 (N_2653,N_2486,N_2492);
or U2654 (N_2654,N_2410,N_2438);
or U2655 (N_2655,N_2354,N_2370);
xor U2656 (N_2656,N_2312,N_2403);
nand U2657 (N_2657,N_2453,N_2299);
xor U2658 (N_2658,N_2275,N_2295);
and U2659 (N_2659,N_2354,N_2478);
or U2660 (N_2660,N_2408,N_2255);
or U2661 (N_2661,N_2419,N_2447);
nor U2662 (N_2662,N_2340,N_2297);
or U2663 (N_2663,N_2443,N_2331);
or U2664 (N_2664,N_2279,N_2331);
nor U2665 (N_2665,N_2433,N_2498);
xor U2666 (N_2666,N_2371,N_2328);
nand U2667 (N_2667,N_2356,N_2297);
nand U2668 (N_2668,N_2462,N_2403);
and U2669 (N_2669,N_2417,N_2455);
and U2670 (N_2670,N_2479,N_2284);
nor U2671 (N_2671,N_2327,N_2447);
or U2672 (N_2672,N_2391,N_2296);
xor U2673 (N_2673,N_2293,N_2375);
nand U2674 (N_2674,N_2440,N_2338);
or U2675 (N_2675,N_2425,N_2275);
nor U2676 (N_2676,N_2277,N_2498);
xnor U2677 (N_2677,N_2304,N_2297);
and U2678 (N_2678,N_2462,N_2275);
xor U2679 (N_2679,N_2346,N_2466);
xnor U2680 (N_2680,N_2287,N_2332);
nand U2681 (N_2681,N_2491,N_2268);
and U2682 (N_2682,N_2457,N_2324);
xor U2683 (N_2683,N_2406,N_2373);
nand U2684 (N_2684,N_2288,N_2328);
nor U2685 (N_2685,N_2310,N_2415);
or U2686 (N_2686,N_2348,N_2467);
xnor U2687 (N_2687,N_2307,N_2489);
nand U2688 (N_2688,N_2378,N_2300);
xor U2689 (N_2689,N_2405,N_2479);
xnor U2690 (N_2690,N_2398,N_2385);
and U2691 (N_2691,N_2433,N_2479);
nand U2692 (N_2692,N_2270,N_2475);
nand U2693 (N_2693,N_2288,N_2270);
and U2694 (N_2694,N_2376,N_2498);
and U2695 (N_2695,N_2269,N_2319);
xnor U2696 (N_2696,N_2315,N_2361);
and U2697 (N_2697,N_2480,N_2486);
xnor U2698 (N_2698,N_2256,N_2389);
and U2699 (N_2699,N_2384,N_2344);
xnor U2700 (N_2700,N_2274,N_2287);
and U2701 (N_2701,N_2298,N_2262);
nand U2702 (N_2702,N_2320,N_2354);
and U2703 (N_2703,N_2420,N_2358);
or U2704 (N_2704,N_2483,N_2441);
xor U2705 (N_2705,N_2390,N_2403);
nand U2706 (N_2706,N_2466,N_2311);
and U2707 (N_2707,N_2427,N_2327);
nor U2708 (N_2708,N_2476,N_2315);
or U2709 (N_2709,N_2274,N_2318);
or U2710 (N_2710,N_2399,N_2392);
xor U2711 (N_2711,N_2329,N_2469);
nor U2712 (N_2712,N_2428,N_2261);
xor U2713 (N_2713,N_2370,N_2296);
nand U2714 (N_2714,N_2334,N_2489);
nor U2715 (N_2715,N_2275,N_2362);
xor U2716 (N_2716,N_2252,N_2271);
nor U2717 (N_2717,N_2473,N_2302);
xor U2718 (N_2718,N_2490,N_2387);
and U2719 (N_2719,N_2455,N_2369);
or U2720 (N_2720,N_2365,N_2468);
nand U2721 (N_2721,N_2436,N_2425);
and U2722 (N_2722,N_2414,N_2268);
nor U2723 (N_2723,N_2309,N_2296);
or U2724 (N_2724,N_2496,N_2300);
or U2725 (N_2725,N_2470,N_2407);
or U2726 (N_2726,N_2289,N_2281);
xnor U2727 (N_2727,N_2460,N_2390);
nand U2728 (N_2728,N_2290,N_2329);
nor U2729 (N_2729,N_2259,N_2257);
nand U2730 (N_2730,N_2455,N_2305);
xnor U2731 (N_2731,N_2479,N_2259);
or U2732 (N_2732,N_2327,N_2318);
nor U2733 (N_2733,N_2360,N_2478);
or U2734 (N_2734,N_2342,N_2424);
or U2735 (N_2735,N_2473,N_2296);
nor U2736 (N_2736,N_2442,N_2337);
nor U2737 (N_2737,N_2416,N_2470);
or U2738 (N_2738,N_2329,N_2410);
and U2739 (N_2739,N_2295,N_2492);
nand U2740 (N_2740,N_2307,N_2253);
nor U2741 (N_2741,N_2499,N_2475);
nor U2742 (N_2742,N_2255,N_2326);
nand U2743 (N_2743,N_2266,N_2488);
and U2744 (N_2744,N_2419,N_2498);
and U2745 (N_2745,N_2452,N_2475);
nand U2746 (N_2746,N_2479,N_2341);
nand U2747 (N_2747,N_2370,N_2476);
or U2748 (N_2748,N_2299,N_2317);
or U2749 (N_2749,N_2261,N_2293);
nor U2750 (N_2750,N_2524,N_2550);
xnor U2751 (N_2751,N_2596,N_2713);
nand U2752 (N_2752,N_2599,N_2581);
or U2753 (N_2753,N_2576,N_2526);
and U2754 (N_2754,N_2548,N_2665);
or U2755 (N_2755,N_2538,N_2572);
nand U2756 (N_2756,N_2544,N_2556);
and U2757 (N_2757,N_2689,N_2533);
and U2758 (N_2758,N_2681,N_2652);
and U2759 (N_2759,N_2644,N_2687);
and U2760 (N_2760,N_2531,N_2619);
or U2761 (N_2761,N_2563,N_2589);
nand U2762 (N_2762,N_2664,N_2719);
nand U2763 (N_2763,N_2542,N_2701);
nor U2764 (N_2764,N_2568,N_2574);
nor U2765 (N_2765,N_2691,N_2671);
nor U2766 (N_2766,N_2724,N_2547);
xor U2767 (N_2767,N_2677,N_2582);
nand U2768 (N_2768,N_2562,N_2702);
nor U2769 (N_2769,N_2700,N_2735);
or U2770 (N_2770,N_2520,N_2516);
or U2771 (N_2771,N_2670,N_2728);
nor U2772 (N_2772,N_2669,N_2712);
xnor U2773 (N_2773,N_2586,N_2505);
nor U2774 (N_2774,N_2616,N_2660);
nor U2775 (N_2775,N_2668,N_2584);
and U2776 (N_2776,N_2507,N_2674);
or U2777 (N_2777,N_2605,N_2537);
nand U2778 (N_2778,N_2553,N_2588);
nor U2779 (N_2779,N_2529,N_2650);
nand U2780 (N_2780,N_2643,N_2692);
and U2781 (N_2781,N_2680,N_2571);
and U2782 (N_2782,N_2500,N_2679);
and U2783 (N_2783,N_2593,N_2527);
nor U2784 (N_2784,N_2578,N_2733);
xor U2785 (N_2785,N_2512,N_2651);
xor U2786 (N_2786,N_2626,N_2631);
xor U2787 (N_2787,N_2502,N_2704);
nor U2788 (N_2788,N_2630,N_2504);
nor U2789 (N_2789,N_2693,N_2648);
xor U2790 (N_2790,N_2602,N_2698);
nand U2791 (N_2791,N_2746,N_2570);
or U2792 (N_2792,N_2645,N_2590);
xnor U2793 (N_2793,N_2716,N_2506);
and U2794 (N_2794,N_2717,N_2729);
or U2795 (N_2795,N_2723,N_2612);
nor U2796 (N_2796,N_2627,N_2573);
and U2797 (N_2797,N_2708,N_2628);
xor U2798 (N_2798,N_2647,N_2711);
and U2799 (N_2799,N_2560,N_2513);
or U2800 (N_2800,N_2667,N_2609);
xnor U2801 (N_2801,N_2747,N_2549);
and U2802 (N_2802,N_2532,N_2743);
nor U2803 (N_2803,N_2515,N_2684);
and U2804 (N_2804,N_2678,N_2511);
xnor U2805 (N_2805,N_2567,N_2591);
or U2806 (N_2806,N_2718,N_2551);
nor U2807 (N_2807,N_2534,N_2579);
or U2808 (N_2808,N_2682,N_2694);
nor U2809 (N_2809,N_2510,N_2638);
nand U2810 (N_2810,N_2696,N_2725);
or U2811 (N_2811,N_2597,N_2720);
nand U2812 (N_2812,N_2539,N_2623);
and U2813 (N_2813,N_2501,N_2583);
xnor U2814 (N_2814,N_2654,N_2649);
and U2815 (N_2815,N_2714,N_2634);
nor U2816 (N_2816,N_2614,N_2595);
or U2817 (N_2817,N_2639,N_2697);
nand U2818 (N_2818,N_2709,N_2690);
xnor U2819 (N_2819,N_2740,N_2528);
nor U2820 (N_2820,N_2530,N_2726);
and U2821 (N_2821,N_2686,N_2657);
or U2822 (N_2822,N_2519,N_2736);
nor U2823 (N_2823,N_2517,N_2662);
and U2824 (N_2824,N_2732,N_2554);
xnor U2825 (N_2825,N_2521,N_2561);
or U2826 (N_2826,N_2545,N_2536);
or U2827 (N_2827,N_2575,N_2587);
or U2828 (N_2828,N_2508,N_2683);
nor U2829 (N_2829,N_2566,N_2640);
nand U2830 (N_2830,N_2675,N_2565);
xnor U2831 (N_2831,N_2632,N_2540);
nor U2832 (N_2832,N_2555,N_2624);
xor U2833 (N_2833,N_2688,N_2592);
or U2834 (N_2834,N_2727,N_2585);
xnor U2835 (N_2835,N_2601,N_2706);
or U2836 (N_2836,N_2738,N_2636);
and U2837 (N_2837,N_2705,N_2594);
nand U2838 (N_2838,N_2722,N_2621);
xor U2839 (N_2839,N_2559,N_2633);
xor U2840 (N_2840,N_2734,N_2695);
or U2841 (N_2841,N_2629,N_2741);
nand U2842 (N_2842,N_2710,N_2600);
and U2843 (N_2843,N_2731,N_2685);
xor U2844 (N_2844,N_2699,N_2635);
xnor U2845 (N_2845,N_2598,N_2666);
or U2846 (N_2846,N_2661,N_2622);
nand U2847 (N_2847,N_2715,N_2658);
and U2848 (N_2848,N_2672,N_2577);
or U2849 (N_2849,N_2611,N_2509);
nor U2850 (N_2850,N_2604,N_2625);
xor U2851 (N_2851,N_2558,N_2637);
and U2852 (N_2852,N_2739,N_2503);
nor U2853 (N_2853,N_2610,N_2620);
or U2854 (N_2854,N_2656,N_2707);
nand U2855 (N_2855,N_2744,N_2745);
or U2856 (N_2856,N_2721,N_2742);
or U2857 (N_2857,N_2749,N_2673);
xnor U2858 (N_2858,N_2676,N_2603);
nand U2859 (N_2859,N_2618,N_2564);
xnor U2860 (N_2860,N_2703,N_2535);
nand U2861 (N_2861,N_2525,N_2557);
nand U2862 (N_2862,N_2552,N_2641);
or U2863 (N_2863,N_2569,N_2615);
xor U2864 (N_2864,N_2522,N_2646);
and U2865 (N_2865,N_2606,N_2514);
xnor U2866 (N_2866,N_2663,N_2748);
or U2867 (N_2867,N_2617,N_2655);
nor U2868 (N_2868,N_2608,N_2523);
xnor U2869 (N_2869,N_2518,N_2607);
nor U2870 (N_2870,N_2541,N_2543);
or U2871 (N_2871,N_2653,N_2737);
or U2872 (N_2872,N_2546,N_2659);
or U2873 (N_2873,N_2642,N_2730);
xnor U2874 (N_2874,N_2580,N_2613);
nand U2875 (N_2875,N_2631,N_2527);
nor U2876 (N_2876,N_2625,N_2719);
xnor U2877 (N_2877,N_2676,N_2608);
nor U2878 (N_2878,N_2725,N_2557);
or U2879 (N_2879,N_2527,N_2602);
or U2880 (N_2880,N_2735,N_2730);
or U2881 (N_2881,N_2553,N_2668);
nand U2882 (N_2882,N_2565,N_2560);
nor U2883 (N_2883,N_2618,N_2693);
xnor U2884 (N_2884,N_2731,N_2697);
xnor U2885 (N_2885,N_2667,N_2679);
xor U2886 (N_2886,N_2522,N_2551);
nand U2887 (N_2887,N_2674,N_2740);
and U2888 (N_2888,N_2676,N_2600);
and U2889 (N_2889,N_2699,N_2647);
and U2890 (N_2890,N_2604,N_2596);
and U2891 (N_2891,N_2640,N_2584);
and U2892 (N_2892,N_2680,N_2608);
nand U2893 (N_2893,N_2604,N_2519);
and U2894 (N_2894,N_2654,N_2720);
or U2895 (N_2895,N_2594,N_2619);
or U2896 (N_2896,N_2648,N_2511);
xor U2897 (N_2897,N_2602,N_2665);
xor U2898 (N_2898,N_2722,N_2602);
nand U2899 (N_2899,N_2665,N_2637);
nor U2900 (N_2900,N_2719,N_2621);
xnor U2901 (N_2901,N_2597,N_2692);
nor U2902 (N_2902,N_2732,N_2572);
or U2903 (N_2903,N_2716,N_2646);
and U2904 (N_2904,N_2683,N_2575);
and U2905 (N_2905,N_2588,N_2565);
and U2906 (N_2906,N_2634,N_2519);
nor U2907 (N_2907,N_2588,N_2673);
xnor U2908 (N_2908,N_2623,N_2614);
nor U2909 (N_2909,N_2629,N_2585);
nor U2910 (N_2910,N_2627,N_2696);
nor U2911 (N_2911,N_2674,N_2690);
nand U2912 (N_2912,N_2666,N_2704);
xnor U2913 (N_2913,N_2548,N_2596);
or U2914 (N_2914,N_2638,N_2551);
nor U2915 (N_2915,N_2569,N_2688);
nand U2916 (N_2916,N_2708,N_2589);
nor U2917 (N_2917,N_2559,N_2651);
nand U2918 (N_2918,N_2582,N_2554);
or U2919 (N_2919,N_2532,N_2609);
xor U2920 (N_2920,N_2704,N_2636);
nand U2921 (N_2921,N_2568,N_2509);
xnor U2922 (N_2922,N_2622,N_2583);
and U2923 (N_2923,N_2522,N_2547);
xor U2924 (N_2924,N_2548,N_2678);
xor U2925 (N_2925,N_2528,N_2619);
and U2926 (N_2926,N_2560,N_2619);
and U2927 (N_2927,N_2680,N_2705);
nand U2928 (N_2928,N_2508,N_2734);
and U2929 (N_2929,N_2543,N_2662);
or U2930 (N_2930,N_2525,N_2558);
xor U2931 (N_2931,N_2645,N_2501);
nand U2932 (N_2932,N_2620,N_2525);
xor U2933 (N_2933,N_2608,N_2530);
xnor U2934 (N_2934,N_2632,N_2695);
nand U2935 (N_2935,N_2585,N_2746);
nor U2936 (N_2936,N_2571,N_2598);
or U2937 (N_2937,N_2739,N_2607);
and U2938 (N_2938,N_2624,N_2712);
nand U2939 (N_2939,N_2560,N_2579);
nor U2940 (N_2940,N_2724,N_2727);
or U2941 (N_2941,N_2566,N_2564);
nor U2942 (N_2942,N_2731,N_2702);
or U2943 (N_2943,N_2724,N_2533);
xnor U2944 (N_2944,N_2729,N_2714);
nand U2945 (N_2945,N_2641,N_2620);
nand U2946 (N_2946,N_2645,N_2726);
or U2947 (N_2947,N_2591,N_2550);
xor U2948 (N_2948,N_2555,N_2557);
xnor U2949 (N_2949,N_2565,N_2524);
or U2950 (N_2950,N_2671,N_2605);
nor U2951 (N_2951,N_2549,N_2593);
nor U2952 (N_2952,N_2694,N_2667);
xnor U2953 (N_2953,N_2730,N_2524);
nand U2954 (N_2954,N_2632,N_2657);
nor U2955 (N_2955,N_2634,N_2582);
nand U2956 (N_2956,N_2584,N_2533);
nor U2957 (N_2957,N_2740,N_2586);
nor U2958 (N_2958,N_2704,N_2669);
nor U2959 (N_2959,N_2746,N_2686);
or U2960 (N_2960,N_2712,N_2709);
nor U2961 (N_2961,N_2716,N_2612);
nor U2962 (N_2962,N_2664,N_2652);
and U2963 (N_2963,N_2608,N_2536);
xnor U2964 (N_2964,N_2565,N_2512);
or U2965 (N_2965,N_2694,N_2585);
nor U2966 (N_2966,N_2560,N_2650);
nand U2967 (N_2967,N_2535,N_2528);
nand U2968 (N_2968,N_2696,N_2558);
xor U2969 (N_2969,N_2511,N_2546);
nand U2970 (N_2970,N_2684,N_2546);
xnor U2971 (N_2971,N_2697,N_2687);
and U2972 (N_2972,N_2660,N_2505);
or U2973 (N_2973,N_2720,N_2593);
nor U2974 (N_2974,N_2730,N_2580);
nor U2975 (N_2975,N_2590,N_2556);
and U2976 (N_2976,N_2637,N_2566);
and U2977 (N_2977,N_2697,N_2595);
nor U2978 (N_2978,N_2552,N_2518);
or U2979 (N_2979,N_2518,N_2622);
nor U2980 (N_2980,N_2537,N_2667);
nor U2981 (N_2981,N_2705,N_2587);
or U2982 (N_2982,N_2639,N_2581);
nand U2983 (N_2983,N_2655,N_2709);
and U2984 (N_2984,N_2668,N_2529);
or U2985 (N_2985,N_2670,N_2660);
and U2986 (N_2986,N_2721,N_2698);
nor U2987 (N_2987,N_2677,N_2526);
nor U2988 (N_2988,N_2738,N_2511);
or U2989 (N_2989,N_2597,N_2561);
nor U2990 (N_2990,N_2692,N_2609);
or U2991 (N_2991,N_2636,N_2745);
or U2992 (N_2992,N_2620,N_2706);
nor U2993 (N_2993,N_2537,N_2718);
nand U2994 (N_2994,N_2608,N_2556);
or U2995 (N_2995,N_2581,N_2675);
nor U2996 (N_2996,N_2582,N_2695);
xor U2997 (N_2997,N_2654,N_2668);
and U2998 (N_2998,N_2608,N_2667);
and U2999 (N_2999,N_2510,N_2547);
nor U3000 (N_3000,N_2887,N_2905);
and U3001 (N_3001,N_2805,N_2890);
nor U3002 (N_3002,N_2756,N_2788);
or U3003 (N_3003,N_2778,N_2791);
nor U3004 (N_3004,N_2884,N_2949);
xnor U3005 (N_3005,N_2812,N_2866);
or U3006 (N_3006,N_2961,N_2888);
nand U3007 (N_3007,N_2984,N_2762);
or U3008 (N_3008,N_2899,N_2840);
nor U3009 (N_3009,N_2754,N_2996);
nand U3010 (N_3010,N_2814,N_2808);
nor U3011 (N_3011,N_2842,N_2940);
nand U3012 (N_3012,N_2944,N_2848);
nand U3013 (N_3013,N_2894,N_2925);
or U3014 (N_3014,N_2864,N_2986);
or U3015 (N_3015,N_2943,N_2836);
nand U3016 (N_3016,N_2911,N_2983);
and U3017 (N_3017,N_2909,N_2912);
nor U3018 (N_3018,N_2766,N_2845);
xnor U3019 (N_3019,N_2868,N_2908);
and U3020 (N_3020,N_2967,N_2898);
nand U3021 (N_3021,N_2981,N_2871);
and U3022 (N_3022,N_2797,N_2819);
nor U3023 (N_3023,N_2763,N_2801);
xor U3024 (N_3024,N_2950,N_2968);
xnor U3025 (N_3025,N_2767,N_2793);
nand U3026 (N_3026,N_2902,N_2773);
or U3027 (N_3027,N_2859,N_2904);
and U3028 (N_3028,N_2844,N_2951);
nor U3029 (N_3029,N_2958,N_2969);
and U3030 (N_3030,N_2772,N_2799);
or U3031 (N_3031,N_2807,N_2930);
and U3032 (N_3032,N_2921,N_2851);
or U3033 (N_3033,N_2988,N_2960);
xnor U3034 (N_3034,N_2815,N_2975);
or U3035 (N_3035,N_2946,N_2832);
nor U3036 (N_3036,N_2897,N_2831);
xor U3037 (N_3037,N_2913,N_2833);
nor U3038 (N_3038,N_2976,N_2796);
nor U3039 (N_3039,N_2769,N_2985);
nor U3040 (N_3040,N_2900,N_2818);
nor U3041 (N_3041,N_2876,N_2910);
or U3042 (N_3042,N_2809,N_2823);
nand U3043 (N_3043,N_2811,N_2835);
or U3044 (N_3044,N_2760,N_2953);
nand U3045 (N_3045,N_2777,N_2813);
nand U3046 (N_3046,N_2874,N_2834);
nor U3047 (N_3047,N_2952,N_2820);
xor U3048 (N_3048,N_2880,N_2794);
nor U3049 (N_3049,N_2750,N_2990);
or U3050 (N_3050,N_2856,N_2989);
or U3051 (N_3051,N_2783,N_2924);
xnor U3052 (N_3052,N_2790,N_2916);
nor U3053 (N_3053,N_2895,N_2903);
and U3054 (N_3054,N_2860,N_2886);
and U3055 (N_3055,N_2915,N_2802);
or U3056 (N_3056,N_2929,N_2945);
nand U3057 (N_3057,N_2992,N_2974);
xnor U3058 (N_3058,N_2828,N_2971);
xnor U3059 (N_3059,N_2928,N_2873);
or U3060 (N_3060,N_2926,N_2784);
nand U3061 (N_3061,N_2979,N_2954);
nor U3062 (N_3062,N_2917,N_2978);
and U3063 (N_3063,N_2935,N_2998);
nand U3064 (N_3064,N_2972,N_2765);
or U3065 (N_3065,N_2837,N_2795);
xor U3066 (N_3066,N_2780,N_2907);
nor U3067 (N_3067,N_2885,N_2821);
nand U3068 (N_3068,N_2798,N_2948);
xnor U3069 (N_3069,N_2931,N_2785);
and U3070 (N_3070,N_2761,N_2982);
or U3071 (N_3071,N_2938,N_2934);
xor U3072 (N_3072,N_2770,N_2824);
nand U3073 (N_3073,N_2841,N_2955);
xnor U3074 (N_3074,N_2869,N_2867);
nand U3075 (N_3075,N_2774,N_2987);
or U3076 (N_3076,N_2927,N_2829);
and U3077 (N_3077,N_2937,N_2786);
nor U3078 (N_3078,N_2826,N_2965);
nand U3079 (N_3079,N_2933,N_2906);
or U3080 (N_3080,N_2771,N_2816);
and U3081 (N_3081,N_2957,N_2849);
xnor U3082 (N_3082,N_2922,N_2995);
nand U3083 (N_3083,N_2855,N_2962);
or U3084 (N_3084,N_2932,N_2920);
or U3085 (N_3085,N_2843,N_2879);
nand U3086 (N_3086,N_2991,N_2964);
xnor U3087 (N_3087,N_2817,N_2959);
nor U3088 (N_3088,N_2993,N_2839);
and U3089 (N_3089,N_2861,N_2980);
xnor U3090 (N_3090,N_2792,N_2936);
xnor U3091 (N_3091,N_2914,N_2857);
or U3092 (N_3092,N_2764,N_2999);
nor U3093 (N_3093,N_2896,N_2782);
nand U3094 (N_3094,N_2883,N_2942);
nor U3095 (N_3095,N_2755,N_2977);
xnor U3096 (N_3096,N_2752,N_2901);
nand U3097 (N_3097,N_2822,N_2827);
nand U3098 (N_3098,N_2779,N_2753);
or U3099 (N_3099,N_2956,N_2847);
xnor U3100 (N_3100,N_2804,N_2781);
and U3101 (N_3101,N_2882,N_2825);
nor U3102 (N_3102,N_2850,N_2789);
nor U3103 (N_3103,N_2941,N_2862);
or U3104 (N_3104,N_2846,N_2758);
xnor U3105 (N_3105,N_2970,N_2800);
or U3106 (N_3106,N_2878,N_2810);
nor U3107 (N_3107,N_2854,N_2973);
or U3108 (N_3108,N_2852,N_2870);
nor U3109 (N_3109,N_2966,N_2853);
nand U3110 (N_3110,N_2891,N_2892);
and U3111 (N_3111,N_2963,N_2757);
nand U3112 (N_3112,N_2863,N_2889);
nand U3113 (N_3113,N_2830,N_2947);
and U3114 (N_3114,N_2893,N_2751);
nor U3115 (N_3115,N_2787,N_2919);
and U3116 (N_3116,N_2918,N_2997);
or U3117 (N_3117,N_2775,N_2875);
xnor U3118 (N_3118,N_2865,N_2939);
xnor U3119 (N_3119,N_2858,N_2872);
and U3120 (N_3120,N_2881,N_2838);
nor U3121 (N_3121,N_2768,N_2994);
or U3122 (N_3122,N_2803,N_2806);
or U3123 (N_3123,N_2776,N_2759);
xor U3124 (N_3124,N_2923,N_2877);
xnor U3125 (N_3125,N_2973,N_2781);
xor U3126 (N_3126,N_2793,N_2842);
xnor U3127 (N_3127,N_2992,N_2955);
nand U3128 (N_3128,N_2813,N_2864);
or U3129 (N_3129,N_2842,N_2816);
or U3130 (N_3130,N_2904,N_2947);
nor U3131 (N_3131,N_2926,N_2988);
nand U3132 (N_3132,N_2910,N_2983);
nor U3133 (N_3133,N_2828,N_2907);
xor U3134 (N_3134,N_2825,N_2754);
nor U3135 (N_3135,N_2799,N_2807);
and U3136 (N_3136,N_2988,N_2782);
and U3137 (N_3137,N_2873,N_2945);
nor U3138 (N_3138,N_2961,N_2758);
nor U3139 (N_3139,N_2972,N_2914);
nor U3140 (N_3140,N_2776,N_2991);
or U3141 (N_3141,N_2806,N_2808);
and U3142 (N_3142,N_2932,N_2875);
nor U3143 (N_3143,N_2781,N_2799);
and U3144 (N_3144,N_2796,N_2916);
nand U3145 (N_3145,N_2875,N_2855);
and U3146 (N_3146,N_2795,N_2850);
nor U3147 (N_3147,N_2822,N_2962);
nand U3148 (N_3148,N_2986,N_2991);
nand U3149 (N_3149,N_2971,N_2931);
nor U3150 (N_3150,N_2920,N_2870);
or U3151 (N_3151,N_2850,N_2939);
nand U3152 (N_3152,N_2838,N_2859);
xnor U3153 (N_3153,N_2989,N_2826);
and U3154 (N_3154,N_2923,N_2989);
xor U3155 (N_3155,N_2932,N_2919);
nor U3156 (N_3156,N_2909,N_2898);
nor U3157 (N_3157,N_2837,N_2963);
xnor U3158 (N_3158,N_2890,N_2791);
xnor U3159 (N_3159,N_2900,N_2910);
or U3160 (N_3160,N_2855,N_2964);
and U3161 (N_3161,N_2895,N_2977);
xor U3162 (N_3162,N_2922,N_2868);
nand U3163 (N_3163,N_2933,N_2798);
nor U3164 (N_3164,N_2920,N_2882);
and U3165 (N_3165,N_2943,N_2775);
nor U3166 (N_3166,N_2868,N_2762);
nand U3167 (N_3167,N_2772,N_2851);
xnor U3168 (N_3168,N_2837,N_2995);
xnor U3169 (N_3169,N_2991,N_2838);
nand U3170 (N_3170,N_2869,N_2991);
nand U3171 (N_3171,N_2849,N_2813);
or U3172 (N_3172,N_2913,N_2793);
nand U3173 (N_3173,N_2918,N_2983);
nor U3174 (N_3174,N_2825,N_2897);
nand U3175 (N_3175,N_2973,N_2809);
and U3176 (N_3176,N_2772,N_2871);
or U3177 (N_3177,N_2881,N_2804);
nand U3178 (N_3178,N_2854,N_2950);
or U3179 (N_3179,N_2830,N_2945);
nand U3180 (N_3180,N_2806,N_2931);
xnor U3181 (N_3181,N_2809,N_2875);
or U3182 (N_3182,N_2837,N_2891);
or U3183 (N_3183,N_2772,N_2948);
nor U3184 (N_3184,N_2959,N_2962);
nand U3185 (N_3185,N_2955,N_2987);
nor U3186 (N_3186,N_2854,N_2844);
and U3187 (N_3187,N_2771,N_2836);
nor U3188 (N_3188,N_2896,N_2949);
nand U3189 (N_3189,N_2891,N_2879);
nand U3190 (N_3190,N_2884,N_2777);
or U3191 (N_3191,N_2973,N_2927);
and U3192 (N_3192,N_2907,N_2767);
and U3193 (N_3193,N_2790,N_2924);
nor U3194 (N_3194,N_2926,N_2960);
nor U3195 (N_3195,N_2918,N_2872);
xor U3196 (N_3196,N_2992,N_2885);
or U3197 (N_3197,N_2945,N_2843);
or U3198 (N_3198,N_2763,N_2931);
or U3199 (N_3199,N_2935,N_2763);
xor U3200 (N_3200,N_2809,N_2821);
or U3201 (N_3201,N_2752,N_2831);
nand U3202 (N_3202,N_2936,N_2954);
or U3203 (N_3203,N_2935,N_2866);
and U3204 (N_3204,N_2902,N_2878);
and U3205 (N_3205,N_2975,N_2851);
nand U3206 (N_3206,N_2752,N_2888);
xor U3207 (N_3207,N_2988,N_2937);
or U3208 (N_3208,N_2875,N_2804);
nor U3209 (N_3209,N_2996,N_2750);
and U3210 (N_3210,N_2919,N_2914);
nor U3211 (N_3211,N_2791,N_2758);
nand U3212 (N_3212,N_2836,N_2792);
nor U3213 (N_3213,N_2779,N_2959);
xor U3214 (N_3214,N_2823,N_2815);
nor U3215 (N_3215,N_2870,N_2863);
and U3216 (N_3216,N_2871,N_2858);
nand U3217 (N_3217,N_2965,N_2985);
and U3218 (N_3218,N_2840,N_2864);
nor U3219 (N_3219,N_2989,N_2799);
xnor U3220 (N_3220,N_2784,N_2850);
nand U3221 (N_3221,N_2896,N_2764);
nand U3222 (N_3222,N_2870,N_2884);
or U3223 (N_3223,N_2755,N_2857);
nand U3224 (N_3224,N_2784,N_2810);
or U3225 (N_3225,N_2794,N_2939);
and U3226 (N_3226,N_2998,N_2895);
nor U3227 (N_3227,N_2910,N_2831);
nand U3228 (N_3228,N_2786,N_2861);
xnor U3229 (N_3229,N_2973,N_2786);
xnor U3230 (N_3230,N_2768,N_2956);
nand U3231 (N_3231,N_2802,N_2974);
nand U3232 (N_3232,N_2870,N_2875);
nor U3233 (N_3233,N_2876,N_2917);
nor U3234 (N_3234,N_2925,N_2758);
nor U3235 (N_3235,N_2949,N_2954);
or U3236 (N_3236,N_2976,N_2754);
xnor U3237 (N_3237,N_2786,N_2945);
or U3238 (N_3238,N_2752,N_2860);
and U3239 (N_3239,N_2870,N_2955);
xnor U3240 (N_3240,N_2873,N_2821);
and U3241 (N_3241,N_2884,N_2975);
nor U3242 (N_3242,N_2896,N_2846);
nor U3243 (N_3243,N_2772,N_2919);
or U3244 (N_3244,N_2928,N_2837);
nor U3245 (N_3245,N_2997,N_2783);
xor U3246 (N_3246,N_2986,N_2777);
nor U3247 (N_3247,N_2936,N_2834);
nor U3248 (N_3248,N_2889,N_2990);
or U3249 (N_3249,N_2844,N_2753);
and U3250 (N_3250,N_3048,N_3106);
and U3251 (N_3251,N_3021,N_3069);
nand U3252 (N_3252,N_3092,N_3065);
nand U3253 (N_3253,N_3130,N_3140);
nand U3254 (N_3254,N_3053,N_3055);
or U3255 (N_3255,N_3093,N_3166);
xor U3256 (N_3256,N_3020,N_3017);
or U3257 (N_3257,N_3153,N_3104);
or U3258 (N_3258,N_3002,N_3082);
nor U3259 (N_3259,N_3072,N_3212);
nor U3260 (N_3260,N_3137,N_3011);
nor U3261 (N_3261,N_3000,N_3059);
nor U3262 (N_3262,N_3161,N_3223);
xnor U3263 (N_3263,N_3085,N_3242);
nand U3264 (N_3264,N_3236,N_3240);
nand U3265 (N_3265,N_3045,N_3219);
or U3266 (N_3266,N_3148,N_3225);
nor U3267 (N_3267,N_3139,N_3136);
or U3268 (N_3268,N_3118,N_3127);
or U3269 (N_3269,N_3133,N_3041);
nand U3270 (N_3270,N_3229,N_3080);
nor U3271 (N_3271,N_3076,N_3138);
or U3272 (N_3272,N_3012,N_3235);
nor U3273 (N_3273,N_3099,N_3026);
and U3274 (N_3274,N_3015,N_3014);
xor U3275 (N_3275,N_3063,N_3191);
or U3276 (N_3276,N_3102,N_3052);
nand U3277 (N_3277,N_3169,N_3158);
or U3278 (N_3278,N_3019,N_3058);
or U3279 (N_3279,N_3211,N_3246);
nor U3280 (N_3280,N_3183,N_3215);
or U3281 (N_3281,N_3200,N_3206);
nand U3282 (N_3282,N_3234,N_3054);
xor U3283 (N_3283,N_3168,N_3146);
and U3284 (N_3284,N_3221,N_3196);
nand U3285 (N_3285,N_3067,N_3199);
nor U3286 (N_3286,N_3018,N_3034);
xnor U3287 (N_3287,N_3064,N_3023);
nand U3288 (N_3288,N_3079,N_3029);
or U3289 (N_3289,N_3124,N_3167);
nand U3290 (N_3290,N_3004,N_3181);
or U3291 (N_3291,N_3237,N_3134);
and U3292 (N_3292,N_3033,N_3036);
and U3293 (N_3293,N_3180,N_3193);
nand U3294 (N_3294,N_3081,N_3131);
and U3295 (N_3295,N_3224,N_3113);
nand U3296 (N_3296,N_3205,N_3051);
xnor U3297 (N_3297,N_3078,N_3057);
nand U3298 (N_3298,N_3032,N_3097);
nand U3299 (N_3299,N_3024,N_3088);
nor U3300 (N_3300,N_3145,N_3143);
xor U3301 (N_3301,N_3141,N_3202);
nor U3302 (N_3302,N_3144,N_3003);
xor U3303 (N_3303,N_3165,N_3050);
nand U3304 (N_3304,N_3109,N_3117);
and U3305 (N_3305,N_3178,N_3031);
nand U3306 (N_3306,N_3094,N_3123);
xor U3307 (N_3307,N_3101,N_3039);
nand U3308 (N_3308,N_3009,N_3096);
and U3309 (N_3309,N_3037,N_3070);
xnor U3310 (N_3310,N_3120,N_3112);
nand U3311 (N_3311,N_3174,N_3013);
or U3312 (N_3312,N_3244,N_3089);
xnor U3313 (N_3313,N_3160,N_3185);
or U3314 (N_3314,N_3044,N_3245);
or U3315 (N_3315,N_3091,N_3111);
nor U3316 (N_3316,N_3187,N_3061);
nand U3317 (N_3317,N_3149,N_3100);
nand U3318 (N_3318,N_3025,N_3201);
or U3319 (N_3319,N_3232,N_3084);
xor U3320 (N_3320,N_3074,N_3098);
xnor U3321 (N_3321,N_3164,N_3090);
nand U3322 (N_3322,N_3230,N_3142);
and U3323 (N_3323,N_3121,N_3049);
and U3324 (N_3324,N_3056,N_3207);
xnor U3325 (N_3325,N_3126,N_3108);
xnor U3326 (N_3326,N_3075,N_3046);
or U3327 (N_3327,N_3198,N_3177);
nor U3328 (N_3328,N_3114,N_3190);
nand U3329 (N_3329,N_3008,N_3086);
nand U3330 (N_3330,N_3083,N_3233);
nor U3331 (N_3331,N_3095,N_3071);
xnor U3332 (N_3332,N_3001,N_3125);
or U3333 (N_3333,N_3239,N_3103);
or U3334 (N_3334,N_3171,N_3155);
xor U3335 (N_3335,N_3179,N_3173);
nor U3336 (N_3336,N_3062,N_3204);
nor U3337 (N_3337,N_3110,N_3042);
nand U3338 (N_3338,N_3105,N_3213);
and U3339 (N_3339,N_3188,N_3040);
nand U3340 (N_3340,N_3043,N_3154);
and U3341 (N_3341,N_3247,N_3231);
and U3342 (N_3342,N_3132,N_3227);
or U3343 (N_3343,N_3068,N_3016);
nand U3344 (N_3344,N_3077,N_3214);
and U3345 (N_3345,N_3107,N_3218);
nor U3346 (N_3346,N_3226,N_3010);
and U3347 (N_3347,N_3241,N_3157);
and U3348 (N_3348,N_3152,N_3194);
nand U3349 (N_3349,N_3119,N_3248);
and U3350 (N_3350,N_3115,N_3022);
nand U3351 (N_3351,N_3243,N_3116);
or U3352 (N_3352,N_3249,N_3170);
nor U3353 (N_3353,N_3197,N_3217);
or U3354 (N_3354,N_3238,N_3195);
and U3355 (N_3355,N_3060,N_3163);
and U3356 (N_3356,N_3028,N_3129);
or U3357 (N_3357,N_3038,N_3006);
nor U3358 (N_3358,N_3186,N_3027);
nand U3359 (N_3359,N_3172,N_3035);
nand U3360 (N_3360,N_3184,N_3150);
nand U3361 (N_3361,N_3047,N_3176);
or U3362 (N_3362,N_3220,N_3005);
nor U3363 (N_3363,N_3216,N_3073);
or U3364 (N_3364,N_3147,N_3135);
and U3365 (N_3365,N_3222,N_3210);
nor U3366 (N_3366,N_3122,N_3156);
nand U3367 (N_3367,N_3189,N_3087);
xnor U3368 (N_3368,N_3066,N_3175);
nand U3369 (N_3369,N_3209,N_3192);
and U3370 (N_3370,N_3128,N_3228);
or U3371 (N_3371,N_3030,N_3162);
or U3372 (N_3372,N_3208,N_3203);
nor U3373 (N_3373,N_3182,N_3007);
xnor U3374 (N_3374,N_3151,N_3159);
xor U3375 (N_3375,N_3089,N_3158);
nand U3376 (N_3376,N_3086,N_3057);
nor U3377 (N_3377,N_3221,N_3074);
nand U3378 (N_3378,N_3172,N_3200);
nor U3379 (N_3379,N_3015,N_3130);
nand U3380 (N_3380,N_3022,N_3181);
nand U3381 (N_3381,N_3218,N_3136);
nor U3382 (N_3382,N_3002,N_3145);
xnor U3383 (N_3383,N_3222,N_3229);
nor U3384 (N_3384,N_3042,N_3191);
nand U3385 (N_3385,N_3213,N_3038);
nand U3386 (N_3386,N_3144,N_3174);
nand U3387 (N_3387,N_3051,N_3113);
or U3388 (N_3388,N_3174,N_3239);
nand U3389 (N_3389,N_3167,N_3100);
xor U3390 (N_3390,N_3147,N_3226);
or U3391 (N_3391,N_3084,N_3214);
xor U3392 (N_3392,N_3126,N_3077);
and U3393 (N_3393,N_3102,N_3177);
xor U3394 (N_3394,N_3097,N_3080);
nor U3395 (N_3395,N_3249,N_3101);
nand U3396 (N_3396,N_3009,N_3228);
or U3397 (N_3397,N_3168,N_3172);
nand U3398 (N_3398,N_3221,N_3194);
and U3399 (N_3399,N_3040,N_3132);
and U3400 (N_3400,N_3083,N_3032);
nor U3401 (N_3401,N_3087,N_3149);
xor U3402 (N_3402,N_3186,N_3196);
xor U3403 (N_3403,N_3214,N_3235);
nor U3404 (N_3404,N_3048,N_3148);
nor U3405 (N_3405,N_3135,N_3217);
nor U3406 (N_3406,N_3204,N_3229);
or U3407 (N_3407,N_3114,N_3211);
or U3408 (N_3408,N_3110,N_3188);
and U3409 (N_3409,N_3156,N_3219);
or U3410 (N_3410,N_3136,N_3172);
or U3411 (N_3411,N_3237,N_3153);
or U3412 (N_3412,N_3056,N_3042);
and U3413 (N_3413,N_3064,N_3141);
nand U3414 (N_3414,N_3168,N_3020);
or U3415 (N_3415,N_3065,N_3016);
and U3416 (N_3416,N_3134,N_3059);
nor U3417 (N_3417,N_3026,N_3245);
xor U3418 (N_3418,N_3083,N_3039);
nor U3419 (N_3419,N_3031,N_3209);
nand U3420 (N_3420,N_3070,N_3086);
xor U3421 (N_3421,N_3185,N_3034);
xor U3422 (N_3422,N_3031,N_3086);
nor U3423 (N_3423,N_3224,N_3123);
and U3424 (N_3424,N_3216,N_3003);
nor U3425 (N_3425,N_3050,N_3178);
nand U3426 (N_3426,N_3248,N_3136);
and U3427 (N_3427,N_3090,N_3173);
nor U3428 (N_3428,N_3160,N_3132);
xnor U3429 (N_3429,N_3065,N_3009);
nor U3430 (N_3430,N_3110,N_3151);
xnor U3431 (N_3431,N_3151,N_3005);
xnor U3432 (N_3432,N_3110,N_3097);
or U3433 (N_3433,N_3072,N_3114);
and U3434 (N_3434,N_3117,N_3019);
nand U3435 (N_3435,N_3098,N_3109);
nor U3436 (N_3436,N_3247,N_3118);
nor U3437 (N_3437,N_3172,N_3216);
nand U3438 (N_3438,N_3048,N_3133);
nor U3439 (N_3439,N_3198,N_3191);
or U3440 (N_3440,N_3069,N_3105);
xnor U3441 (N_3441,N_3045,N_3096);
xnor U3442 (N_3442,N_3123,N_3065);
or U3443 (N_3443,N_3170,N_3199);
nand U3444 (N_3444,N_3227,N_3125);
and U3445 (N_3445,N_3008,N_3216);
nor U3446 (N_3446,N_3152,N_3017);
nand U3447 (N_3447,N_3184,N_3248);
nand U3448 (N_3448,N_3005,N_3234);
or U3449 (N_3449,N_3047,N_3233);
xnor U3450 (N_3450,N_3235,N_3029);
nor U3451 (N_3451,N_3059,N_3049);
and U3452 (N_3452,N_3028,N_3230);
nor U3453 (N_3453,N_3240,N_3235);
nand U3454 (N_3454,N_3175,N_3225);
and U3455 (N_3455,N_3056,N_3145);
and U3456 (N_3456,N_3175,N_3119);
nand U3457 (N_3457,N_3152,N_3239);
and U3458 (N_3458,N_3046,N_3168);
nor U3459 (N_3459,N_3001,N_3144);
nor U3460 (N_3460,N_3168,N_3151);
nor U3461 (N_3461,N_3196,N_3064);
or U3462 (N_3462,N_3226,N_3005);
and U3463 (N_3463,N_3235,N_3095);
xor U3464 (N_3464,N_3038,N_3080);
nor U3465 (N_3465,N_3001,N_3149);
nor U3466 (N_3466,N_3228,N_3147);
nor U3467 (N_3467,N_3200,N_3106);
xor U3468 (N_3468,N_3230,N_3017);
xnor U3469 (N_3469,N_3153,N_3009);
or U3470 (N_3470,N_3167,N_3150);
or U3471 (N_3471,N_3219,N_3104);
nor U3472 (N_3472,N_3214,N_3040);
and U3473 (N_3473,N_3183,N_3021);
and U3474 (N_3474,N_3205,N_3146);
nor U3475 (N_3475,N_3194,N_3033);
xnor U3476 (N_3476,N_3183,N_3129);
xor U3477 (N_3477,N_3155,N_3168);
xnor U3478 (N_3478,N_3144,N_3013);
nor U3479 (N_3479,N_3118,N_3007);
and U3480 (N_3480,N_3071,N_3098);
nor U3481 (N_3481,N_3096,N_3055);
xnor U3482 (N_3482,N_3061,N_3067);
nand U3483 (N_3483,N_3124,N_3098);
or U3484 (N_3484,N_3092,N_3010);
nor U3485 (N_3485,N_3049,N_3210);
nand U3486 (N_3486,N_3138,N_3048);
or U3487 (N_3487,N_3089,N_3029);
nor U3488 (N_3488,N_3002,N_3095);
xor U3489 (N_3489,N_3100,N_3037);
xor U3490 (N_3490,N_3057,N_3089);
or U3491 (N_3491,N_3009,N_3117);
and U3492 (N_3492,N_3145,N_3057);
and U3493 (N_3493,N_3049,N_3007);
xor U3494 (N_3494,N_3084,N_3180);
nand U3495 (N_3495,N_3063,N_3107);
nor U3496 (N_3496,N_3132,N_3229);
nand U3497 (N_3497,N_3193,N_3241);
xor U3498 (N_3498,N_3093,N_3187);
or U3499 (N_3499,N_3086,N_3053);
xnor U3500 (N_3500,N_3421,N_3264);
nand U3501 (N_3501,N_3383,N_3450);
and U3502 (N_3502,N_3476,N_3466);
and U3503 (N_3503,N_3467,N_3358);
and U3504 (N_3504,N_3377,N_3257);
nor U3505 (N_3505,N_3389,N_3255);
nand U3506 (N_3506,N_3302,N_3371);
and U3507 (N_3507,N_3492,N_3369);
and U3508 (N_3508,N_3381,N_3309);
nor U3509 (N_3509,N_3442,N_3418);
or U3510 (N_3510,N_3499,N_3354);
and U3511 (N_3511,N_3333,N_3472);
or U3512 (N_3512,N_3431,N_3307);
xnor U3513 (N_3513,N_3471,N_3464);
nand U3514 (N_3514,N_3347,N_3409);
or U3515 (N_3515,N_3490,N_3289);
nand U3516 (N_3516,N_3391,N_3335);
nor U3517 (N_3517,N_3411,N_3488);
nand U3518 (N_3518,N_3328,N_3373);
or U3519 (N_3519,N_3429,N_3412);
nand U3520 (N_3520,N_3286,N_3493);
or U3521 (N_3521,N_3375,N_3362);
nor U3522 (N_3522,N_3420,N_3292);
or U3523 (N_3523,N_3465,N_3387);
and U3524 (N_3524,N_3285,N_3337);
nand U3525 (N_3525,N_3306,N_3366);
xor U3526 (N_3526,N_3269,N_3460);
nand U3527 (N_3527,N_3270,N_3274);
nor U3528 (N_3528,N_3267,N_3395);
and U3529 (N_3529,N_3479,N_3384);
or U3530 (N_3530,N_3296,N_3338);
or U3531 (N_3531,N_3363,N_3339);
xor U3532 (N_3532,N_3253,N_3319);
and U3533 (N_3533,N_3297,N_3298);
xor U3534 (N_3534,N_3324,N_3305);
nand U3535 (N_3535,N_3397,N_3413);
xor U3536 (N_3536,N_3326,N_3321);
nor U3537 (N_3537,N_3315,N_3344);
nand U3538 (N_3538,N_3399,N_3407);
nand U3539 (N_3539,N_3468,N_3393);
nand U3540 (N_3540,N_3251,N_3279);
nor U3541 (N_3541,N_3386,N_3341);
nand U3542 (N_3542,N_3470,N_3382);
nor U3543 (N_3543,N_3353,N_3443);
nor U3544 (N_3544,N_3474,N_3317);
and U3545 (N_3545,N_3497,N_3480);
and U3546 (N_3546,N_3435,N_3262);
nor U3547 (N_3547,N_3331,N_3401);
nor U3548 (N_3548,N_3436,N_3355);
xor U3549 (N_3549,N_3446,N_3459);
nor U3550 (N_3550,N_3327,N_3405);
or U3551 (N_3551,N_3275,N_3304);
xnor U3552 (N_3552,N_3287,N_3364);
nand U3553 (N_3553,N_3430,N_3408);
and U3554 (N_3554,N_3404,N_3276);
nand U3555 (N_3555,N_3416,N_3433);
xor U3556 (N_3556,N_3496,N_3308);
xor U3557 (N_3557,N_3489,N_3498);
nor U3558 (N_3558,N_3441,N_3437);
xor U3559 (N_3559,N_3481,N_3448);
or U3560 (N_3560,N_3314,N_3424);
nor U3561 (N_3561,N_3390,N_3477);
xor U3562 (N_3562,N_3372,N_3281);
or U3563 (N_3563,N_3343,N_3311);
nand U3564 (N_3564,N_3402,N_3340);
and U3565 (N_3565,N_3438,N_3290);
xnor U3566 (N_3566,N_3398,N_3392);
xor U3567 (N_3567,N_3434,N_3361);
nor U3568 (N_3568,N_3425,N_3440);
nand U3569 (N_3569,N_3414,N_3428);
nor U3570 (N_3570,N_3380,N_3365);
xor U3571 (N_3571,N_3280,N_3449);
nand U3572 (N_3572,N_3310,N_3445);
nor U3573 (N_3573,N_3427,N_3359);
and U3574 (N_3574,N_3318,N_3417);
nor U3575 (N_3575,N_3334,N_3288);
and U3576 (N_3576,N_3301,N_3379);
xor U3577 (N_3577,N_3284,N_3293);
nand U3578 (N_3578,N_3478,N_3266);
and U3579 (N_3579,N_3348,N_3403);
nand U3580 (N_3580,N_3378,N_3273);
or U3581 (N_3581,N_3320,N_3444);
nor U3582 (N_3582,N_3332,N_3261);
nor U3583 (N_3583,N_3463,N_3439);
and U3584 (N_3584,N_3323,N_3316);
nand U3585 (N_3585,N_3396,N_3495);
xnor U3586 (N_3586,N_3491,N_3350);
nand U3587 (N_3587,N_3455,N_3277);
and U3588 (N_3588,N_3299,N_3356);
and U3589 (N_3589,N_3283,N_3268);
nand U3590 (N_3590,N_3325,N_3454);
nor U3591 (N_3591,N_3447,N_3294);
nor U3592 (N_3592,N_3473,N_3259);
and U3593 (N_3593,N_3475,N_3345);
and U3594 (N_3594,N_3456,N_3352);
or U3595 (N_3595,N_3374,N_3388);
xnor U3596 (N_3596,N_3370,N_3303);
nor U3597 (N_3597,N_3254,N_3263);
and U3598 (N_3598,N_3485,N_3342);
and U3599 (N_3599,N_3432,N_3271);
nand U3600 (N_3600,N_3312,N_3300);
xor U3601 (N_3601,N_3360,N_3295);
and U3602 (N_3602,N_3368,N_3400);
nand U3603 (N_3603,N_3349,N_3313);
nand U3604 (N_3604,N_3452,N_3367);
xnor U3605 (N_3605,N_3252,N_3451);
and U3606 (N_3606,N_3376,N_3336);
and U3607 (N_3607,N_3256,N_3462);
or U3608 (N_3608,N_3482,N_3330);
or U3609 (N_3609,N_3487,N_3250);
or U3610 (N_3610,N_3410,N_3415);
xor U3611 (N_3611,N_3291,N_3329);
and U3612 (N_3612,N_3322,N_3458);
nor U3613 (N_3613,N_3426,N_3272);
nor U3614 (N_3614,N_3494,N_3278);
nand U3615 (N_3615,N_3419,N_3483);
and U3616 (N_3616,N_3260,N_3484);
nand U3617 (N_3617,N_3265,N_3457);
and U3618 (N_3618,N_3357,N_3406);
and U3619 (N_3619,N_3346,N_3351);
nor U3620 (N_3620,N_3394,N_3385);
and U3621 (N_3621,N_3469,N_3258);
and U3622 (N_3622,N_3453,N_3461);
xnor U3623 (N_3623,N_3282,N_3422);
nor U3624 (N_3624,N_3423,N_3486);
and U3625 (N_3625,N_3327,N_3345);
and U3626 (N_3626,N_3464,N_3426);
xnor U3627 (N_3627,N_3381,N_3360);
or U3628 (N_3628,N_3328,N_3476);
or U3629 (N_3629,N_3273,N_3387);
nor U3630 (N_3630,N_3310,N_3385);
and U3631 (N_3631,N_3292,N_3301);
nor U3632 (N_3632,N_3255,N_3339);
xnor U3633 (N_3633,N_3426,N_3419);
xor U3634 (N_3634,N_3414,N_3288);
nand U3635 (N_3635,N_3377,N_3282);
nand U3636 (N_3636,N_3484,N_3333);
xor U3637 (N_3637,N_3452,N_3322);
and U3638 (N_3638,N_3336,N_3351);
xnor U3639 (N_3639,N_3364,N_3288);
and U3640 (N_3640,N_3336,N_3449);
nor U3641 (N_3641,N_3422,N_3272);
or U3642 (N_3642,N_3384,N_3311);
nor U3643 (N_3643,N_3418,N_3349);
and U3644 (N_3644,N_3495,N_3363);
nor U3645 (N_3645,N_3484,N_3270);
nand U3646 (N_3646,N_3404,N_3497);
nor U3647 (N_3647,N_3431,N_3479);
and U3648 (N_3648,N_3293,N_3318);
nor U3649 (N_3649,N_3438,N_3370);
nand U3650 (N_3650,N_3389,N_3250);
or U3651 (N_3651,N_3333,N_3371);
xor U3652 (N_3652,N_3496,N_3321);
nor U3653 (N_3653,N_3378,N_3348);
or U3654 (N_3654,N_3294,N_3344);
and U3655 (N_3655,N_3487,N_3307);
nor U3656 (N_3656,N_3324,N_3487);
nor U3657 (N_3657,N_3295,N_3276);
nand U3658 (N_3658,N_3439,N_3256);
nand U3659 (N_3659,N_3424,N_3252);
nand U3660 (N_3660,N_3491,N_3475);
nor U3661 (N_3661,N_3430,N_3468);
or U3662 (N_3662,N_3348,N_3376);
nand U3663 (N_3663,N_3478,N_3442);
and U3664 (N_3664,N_3467,N_3378);
and U3665 (N_3665,N_3299,N_3460);
and U3666 (N_3666,N_3397,N_3478);
xor U3667 (N_3667,N_3288,N_3337);
xnor U3668 (N_3668,N_3424,N_3383);
nand U3669 (N_3669,N_3323,N_3336);
and U3670 (N_3670,N_3334,N_3426);
or U3671 (N_3671,N_3256,N_3370);
nand U3672 (N_3672,N_3348,N_3356);
or U3673 (N_3673,N_3366,N_3496);
and U3674 (N_3674,N_3319,N_3291);
and U3675 (N_3675,N_3406,N_3328);
nor U3676 (N_3676,N_3322,N_3330);
xor U3677 (N_3677,N_3357,N_3269);
or U3678 (N_3678,N_3329,N_3368);
xnor U3679 (N_3679,N_3380,N_3359);
nand U3680 (N_3680,N_3300,N_3321);
or U3681 (N_3681,N_3499,N_3259);
nand U3682 (N_3682,N_3352,N_3493);
and U3683 (N_3683,N_3287,N_3393);
or U3684 (N_3684,N_3313,N_3253);
xor U3685 (N_3685,N_3484,N_3300);
or U3686 (N_3686,N_3354,N_3452);
nor U3687 (N_3687,N_3412,N_3485);
nand U3688 (N_3688,N_3470,N_3426);
xor U3689 (N_3689,N_3374,N_3310);
or U3690 (N_3690,N_3424,N_3401);
or U3691 (N_3691,N_3259,N_3417);
nor U3692 (N_3692,N_3496,N_3250);
xor U3693 (N_3693,N_3368,N_3261);
xor U3694 (N_3694,N_3435,N_3490);
or U3695 (N_3695,N_3313,N_3415);
nand U3696 (N_3696,N_3448,N_3394);
or U3697 (N_3697,N_3364,N_3455);
nand U3698 (N_3698,N_3477,N_3412);
nor U3699 (N_3699,N_3318,N_3358);
nand U3700 (N_3700,N_3467,N_3274);
or U3701 (N_3701,N_3270,N_3403);
nor U3702 (N_3702,N_3284,N_3310);
nor U3703 (N_3703,N_3353,N_3433);
or U3704 (N_3704,N_3303,N_3304);
nand U3705 (N_3705,N_3412,N_3356);
and U3706 (N_3706,N_3347,N_3429);
xor U3707 (N_3707,N_3381,N_3421);
nor U3708 (N_3708,N_3465,N_3399);
nand U3709 (N_3709,N_3316,N_3307);
nand U3710 (N_3710,N_3284,N_3361);
nand U3711 (N_3711,N_3353,N_3279);
or U3712 (N_3712,N_3369,N_3399);
nor U3713 (N_3713,N_3263,N_3489);
nor U3714 (N_3714,N_3325,N_3350);
nor U3715 (N_3715,N_3269,N_3351);
nand U3716 (N_3716,N_3494,N_3475);
nand U3717 (N_3717,N_3314,N_3291);
xor U3718 (N_3718,N_3489,N_3338);
xor U3719 (N_3719,N_3425,N_3480);
nand U3720 (N_3720,N_3298,N_3257);
or U3721 (N_3721,N_3286,N_3464);
xnor U3722 (N_3722,N_3427,N_3490);
or U3723 (N_3723,N_3375,N_3338);
xnor U3724 (N_3724,N_3327,N_3466);
nand U3725 (N_3725,N_3266,N_3437);
nand U3726 (N_3726,N_3490,N_3378);
and U3727 (N_3727,N_3414,N_3354);
or U3728 (N_3728,N_3388,N_3408);
nor U3729 (N_3729,N_3359,N_3373);
xnor U3730 (N_3730,N_3481,N_3494);
and U3731 (N_3731,N_3439,N_3485);
nand U3732 (N_3732,N_3391,N_3373);
or U3733 (N_3733,N_3290,N_3388);
or U3734 (N_3734,N_3413,N_3289);
nand U3735 (N_3735,N_3275,N_3482);
nand U3736 (N_3736,N_3431,N_3390);
and U3737 (N_3737,N_3429,N_3332);
nor U3738 (N_3738,N_3391,N_3448);
nor U3739 (N_3739,N_3457,N_3373);
nor U3740 (N_3740,N_3461,N_3488);
xor U3741 (N_3741,N_3262,N_3255);
xor U3742 (N_3742,N_3343,N_3340);
xor U3743 (N_3743,N_3403,N_3387);
nand U3744 (N_3744,N_3280,N_3427);
or U3745 (N_3745,N_3374,N_3289);
nor U3746 (N_3746,N_3383,N_3329);
nand U3747 (N_3747,N_3399,N_3323);
nand U3748 (N_3748,N_3444,N_3372);
nand U3749 (N_3749,N_3484,N_3406);
nor U3750 (N_3750,N_3733,N_3588);
xnor U3751 (N_3751,N_3660,N_3609);
and U3752 (N_3752,N_3611,N_3629);
and U3753 (N_3753,N_3627,N_3618);
and U3754 (N_3754,N_3632,N_3625);
nand U3755 (N_3755,N_3593,N_3692);
and U3756 (N_3756,N_3713,N_3650);
nor U3757 (N_3757,N_3623,N_3649);
or U3758 (N_3758,N_3705,N_3718);
or U3759 (N_3759,N_3570,N_3691);
or U3760 (N_3760,N_3523,N_3507);
or U3761 (N_3761,N_3518,N_3529);
nor U3762 (N_3762,N_3734,N_3622);
nor U3763 (N_3763,N_3655,N_3509);
xor U3764 (N_3764,N_3582,N_3737);
and U3765 (N_3765,N_3602,N_3645);
xnor U3766 (N_3766,N_3574,N_3740);
nor U3767 (N_3767,N_3659,N_3682);
or U3768 (N_3768,N_3633,N_3578);
nand U3769 (N_3769,N_3741,N_3634);
xnor U3770 (N_3770,N_3666,N_3550);
nand U3771 (N_3771,N_3693,N_3505);
and U3772 (N_3772,N_3712,N_3603);
and U3773 (N_3773,N_3553,N_3576);
or U3774 (N_3774,N_3548,N_3558);
and U3775 (N_3775,N_3624,N_3644);
and U3776 (N_3776,N_3688,N_3663);
and U3777 (N_3777,N_3561,N_3555);
nand U3778 (N_3778,N_3689,N_3512);
nand U3779 (N_3779,N_3596,N_3665);
or U3780 (N_3780,N_3677,N_3566);
or U3781 (N_3781,N_3584,N_3711);
nand U3782 (N_3782,N_3641,N_3679);
and U3783 (N_3783,N_3717,N_3569);
xnor U3784 (N_3784,N_3654,N_3510);
or U3785 (N_3785,N_3703,N_3695);
or U3786 (N_3786,N_3540,N_3522);
xnor U3787 (N_3787,N_3556,N_3539);
nor U3788 (N_3788,N_3729,N_3652);
xor U3789 (N_3789,N_3552,N_3544);
or U3790 (N_3790,N_3606,N_3565);
nor U3791 (N_3791,N_3575,N_3564);
or U3792 (N_3792,N_3563,N_3668);
xnor U3793 (N_3793,N_3700,N_3516);
nor U3794 (N_3794,N_3626,N_3651);
and U3795 (N_3795,N_3736,N_3714);
or U3796 (N_3796,N_3551,N_3690);
and U3797 (N_3797,N_3701,N_3513);
nand U3798 (N_3798,N_3722,N_3676);
xor U3799 (N_3799,N_3735,N_3600);
nand U3800 (N_3800,N_3587,N_3662);
or U3801 (N_3801,N_3738,N_3685);
and U3802 (N_3802,N_3543,N_3630);
nor U3803 (N_3803,N_3560,N_3595);
nand U3804 (N_3804,N_3608,N_3694);
nor U3805 (N_3805,N_3646,N_3520);
and U3806 (N_3806,N_3669,N_3557);
nand U3807 (N_3807,N_3541,N_3657);
nor U3808 (N_3808,N_3672,N_3726);
xnor U3809 (N_3809,N_3573,N_3667);
nor U3810 (N_3810,N_3591,N_3580);
nor U3811 (N_3811,N_3579,N_3610);
nand U3812 (N_3812,N_3592,N_3501);
xnor U3813 (N_3813,N_3528,N_3581);
nor U3814 (N_3814,N_3656,N_3613);
or U3815 (N_3815,N_3533,N_3707);
nand U3816 (N_3816,N_3607,N_3614);
and U3817 (N_3817,N_3612,N_3537);
and U3818 (N_3818,N_3716,N_3597);
and U3819 (N_3819,N_3631,N_3728);
or U3820 (N_3820,N_3704,N_3601);
xnor U3821 (N_3821,N_3747,N_3643);
nor U3822 (N_3822,N_3742,N_3671);
and U3823 (N_3823,N_3661,N_3594);
nand U3824 (N_3824,N_3635,N_3532);
nand U3825 (N_3825,N_3583,N_3708);
and U3826 (N_3826,N_3673,N_3619);
nand U3827 (N_3827,N_3559,N_3658);
xor U3828 (N_3828,N_3664,N_3521);
nand U3829 (N_3829,N_3604,N_3542);
nor U3830 (N_3830,N_3525,N_3549);
or U3831 (N_3831,N_3589,N_3545);
nor U3832 (N_3832,N_3647,N_3506);
nand U3833 (N_3833,N_3680,N_3515);
xnor U3834 (N_3834,N_3547,N_3710);
nor U3835 (N_3835,N_3621,N_3577);
nor U3836 (N_3836,N_3730,N_3698);
xnor U3837 (N_3837,N_3511,N_3536);
nor U3838 (N_3838,N_3743,N_3674);
nand U3839 (N_3839,N_3720,N_3620);
xnor U3840 (N_3840,N_3670,N_3715);
xor U3841 (N_3841,N_3684,N_3653);
nor U3842 (N_3842,N_3502,N_3723);
nand U3843 (N_3843,N_3616,N_3534);
nor U3844 (N_3844,N_3719,N_3709);
xnor U3845 (N_3845,N_3727,N_3749);
nand U3846 (N_3846,N_3686,N_3503);
xor U3847 (N_3847,N_3514,N_3731);
and U3848 (N_3848,N_3568,N_3744);
xor U3849 (N_3849,N_3526,N_3732);
and U3850 (N_3850,N_3640,N_3599);
and U3851 (N_3851,N_3598,N_3527);
nand U3852 (N_3852,N_3562,N_3724);
nand U3853 (N_3853,N_3586,N_3697);
nand U3854 (N_3854,N_3531,N_3567);
and U3855 (N_3855,N_3678,N_3681);
and U3856 (N_3856,N_3615,N_3590);
nor U3857 (N_3857,N_3636,N_3585);
nand U3858 (N_3858,N_3508,N_3605);
and U3859 (N_3859,N_3721,N_3746);
or U3860 (N_3860,N_3675,N_3745);
or U3861 (N_3861,N_3696,N_3546);
nor U3862 (N_3862,N_3571,N_3530);
or U3863 (N_3863,N_3517,N_3535);
nand U3864 (N_3864,N_3702,N_3642);
and U3865 (N_3865,N_3500,N_3706);
and U3866 (N_3866,N_3524,N_3683);
or U3867 (N_3867,N_3748,N_3504);
nand U3868 (N_3868,N_3554,N_3699);
xnor U3869 (N_3869,N_3648,N_3538);
or U3870 (N_3870,N_3638,N_3687);
nand U3871 (N_3871,N_3639,N_3628);
xor U3872 (N_3872,N_3617,N_3725);
nand U3873 (N_3873,N_3519,N_3637);
nor U3874 (N_3874,N_3572,N_3739);
or U3875 (N_3875,N_3722,N_3520);
or U3876 (N_3876,N_3610,N_3607);
xor U3877 (N_3877,N_3749,N_3530);
xor U3878 (N_3878,N_3577,N_3531);
xor U3879 (N_3879,N_3746,N_3508);
nand U3880 (N_3880,N_3541,N_3723);
nor U3881 (N_3881,N_3522,N_3524);
and U3882 (N_3882,N_3570,N_3528);
or U3883 (N_3883,N_3694,N_3600);
or U3884 (N_3884,N_3538,N_3618);
nor U3885 (N_3885,N_3705,N_3744);
xnor U3886 (N_3886,N_3659,N_3661);
xor U3887 (N_3887,N_3644,N_3524);
xor U3888 (N_3888,N_3588,N_3543);
and U3889 (N_3889,N_3729,N_3587);
xor U3890 (N_3890,N_3621,N_3610);
xor U3891 (N_3891,N_3582,N_3535);
and U3892 (N_3892,N_3652,N_3629);
or U3893 (N_3893,N_3600,N_3552);
xnor U3894 (N_3894,N_3586,N_3708);
and U3895 (N_3895,N_3577,N_3658);
nand U3896 (N_3896,N_3564,N_3697);
nor U3897 (N_3897,N_3620,N_3680);
nor U3898 (N_3898,N_3697,N_3556);
xor U3899 (N_3899,N_3688,N_3736);
or U3900 (N_3900,N_3708,N_3506);
nor U3901 (N_3901,N_3560,N_3548);
nor U3902 (N_3902,N_3567,N_3706);
or U3903 (N_3903,N_3702,N_3705);
or U3904 (N_3904,N_3652,N_3674);
nor U3905 (N_3905,N_3646,N_3587);
and U3906 (N_3906,N_3730,N_3565);
or U3907 (N_3907,N_3715,N_3737);
xor U3908 (N_3908,N_3743,N_3689);
xnor U3909 (N_3909,N_3510,N_3698);
nor U3910 (N_3910,N_3605,N_3733);
nand U3911 (N_3911,N_3578,N_3536);
nor U3912 (N_3912,N_3528,N_3553);
nor U3913 (N_3913,N_3732,N_3717);
xor U3914 (N_3914,N_3544,N_3728);
xnor U3915 (N_3915,N_3699,N_3596);
nor U3916 (N_3916,N_3530,N_3617);
or U3917 (N_3917,N_3622,N_3553);
nor U3918 (N_3918,N_3714,N_3539);
xnor U3919 (N_3919,N_3661,N_3608);
nand U3920 (N_3920,N_3557,N_3551);
xnor U3921 (N_3921,N_3533,N_3523);
or U3922 (N_3922,N_3626,N_3627);
or U3923 (N_3923,N_3568,N_3562);
nand U3924 (N_3924,N_3711,N_3631);
and U3925 (N_3925,N_3591,N_3712);
nor U3926 (N_3926,N_3741,N_3592);
nand U3927 (N_3927,N_3640,N_3558);
xnor U3928 (N_3928,N_3653,N_3729);
or U3929 (N_3929,N_3699,N_3597);
nand U3930 (N_3930,N_3738,N_3552);
and U3931 (N_3931,N_3673,N_3632);
and U3932 (N_3932,N_3658,N_3536);
or U3933 (N_3933,N_3573,N_3605);
nor U3934 (N_3934,N_3542,N_3609);
nor U3935 (N_3935,N_3511,N_3639);
nand U3936 (N_3936,N_3747,N_3548);
nand U3937 (N_3937,N_3583,N_3684);
or U3938 (N_3938,N_3513,N_3542);
or U3939 (N_3939,N_3640,N_3660);
nand U3940 (N_3940,N_3527,N_3663);
nor U3941 (N_3941,N_3563,N_3602);
or U3942 (N_3942,N_3519,N_3739);
or U3943 (N_3943,N_3684,N_3564);
nand U3944 (N_3944,N_3722,N_3588);
nor U3945 (N_3945,N_3612,N_3614);
nand U3946 (N_3946,N_3721,N_3688);
xnor U3947 (N_3947,N_3742,N_3630);
or U3948 (N_3948,N_3663,N_3673);
xnor U3949 (N_3949,N_3638,N_3607);
or U3950 (N_3950,N_3563,N_3625);
or U3951 (N_3951,N_3539,N_3625);
or U3952 (N_3952,N_3706,N_3539);
xnor U3953 (N_3953,N_3561,N_3578);
nand U3954 (N_3954,N_3581,N_3634);
xnor U3955 (N_3955,N_3699,N_3555);
or U3956 (N_3956,N_3508,N_3521);
nand U3957 (N_3957,N_3653,N_3607);
nand U3958 (N_3958,N_3666,N_3646);
or U3959 (N_3959,N_3607,N_3509);
nor U3960 (N_3960,N_3532,N_3609);
xor U3961 (N_3961,N_3676,N_3653);
nand U3962 (N_3962,N_3673,N_3729);
and U3963 (N_3963,N_3648,N_3705);
xor U3964 (N_3964,N_3632,N_3604);
nor U3965 (N_3965,N_3677,N_3536);
xor U3966 (N_3966,N_3653,N_3544);
xor U3967 (N_3967,N_3655,N_3570);
or U3968 (N_3968,N_3512,N_3584);
nand U3969 (N_3969,N_3554,N_3667);
nand U3970 (N_3970,N_3640,N_3623);
xnor U3971 (N_3971,N_3730,N_3567);
xnor U3972 (N_3972,N_3685,N_3741);
xor U3973 (N_3973,N_3672,N_3617);
and U3974 (N_3974,N_3706,N_3538);
or U3975 (N_3975,N_3604,N_3656);
and U3976 (N_3976,N_3625,N_3619);
nor U3977 (N_3977,N_3674,N_3682);
nor U3978 (N_3978,N_3723,N_3605);
nand U3979 (N_3979,N_3624,N_3693);
xnor U3980 (N_3980,N_3600,N_3709);
or U3981 (N_3981,N_3701,N_3608);
nand U3982 (N_3982,N_3617,N_3618);
nor U3983 (N_3983,N_3547,N_3581);
nor U3984 (N_3984,N_3620,N_3590);
and U3985 (N_3985,N_3629,N_3677);
xnor U3986 (N_3986,N_3713,N_3697);
and U3987 (N_3987,N_3736,N_3502);
nor U3988 (N_3988,N_3707,N_3638);
xnor U3989 (N_3989,N_3703,N_3675);
or U3990 (N_3990,N_3590,N_3654);
and U3991 (N_3991,N_3617,N_3682);
nand U3992 (N_3992,N_3719,N_3514);
nand U3993 (N_3993,N_3662,N_3630);
nand U3994 (N_3994,N_3579,N_3594);
nor U3995 (N_3995,N_3514,N_3699);
and U3996 (N_3996,N_3511,N_3532);
xor U3997 (N_3997,N_3562,N_3548);
nand U3998 (N_3998,N_3539,N_3564);
and U3999 (N_3999,N_3679,N_3715);
nand U4000 (N_4000,N_3879,N_3862);
xor U4001 (N_4001,N_3857,N_3877);
nand U4002 (N_4002,N_3967,N_3897);
or U4003 (N_4003,N_3902,N_3886);
nand U4004 (N_4004,N_3943,N_3942);
xnor U4005 (N_4005,N_3973,N_3842);
xnor U4006 (N_4006,N_3888,N_3776);
nor U4007 (N_4007,N_3946,N_3751);
nor U4008 (N_4008,N_3851,N_3763);
or U4009 (N_4009,N_3969,N_3872);
nand U4010 (N_4010,N_3951,N_3750);
nor U4011 (N_4011,N_3808,N_3914);
xor U4012 (N_4012,N_3976,N_3994);
xnor U4013 (N_4013,N_3850,N_3871);
nor U4014 (N_4014,N_3950,N_3796);
nand U4015 (N_4015,N_3865,N_3873);
xnor U4016 (N_4016,N_3800,N_3819);
nand U4017 (N_4017,N_3835,N_3775);
nand U4018 (N_4018,N_3810,N_3966);
and U4019 (N_4019,N_3794,N_3923);
or U4020 (N_4020,N_3880,N_3814);
and U4021 (N_4021,N_3958,N_3766);
nor U4022 (N_4022,N_3761,N_3961);
and U4023 (N_4023,N_3990,N_3982);
or U4024 (N_4024,N_3968,N_3759);
nand U4025 (N_4025,N_3824,N_3828);
xnor U4026 (N_4026,N_3997,N_3986);
nor U4027 (N_4027,N_3786,N_3908);
and U4028 (N_4028,N_3853,N_3875);
and U4029 (N_4029,N_3930,N_3785);
xnor U4030 (N_4030,N_3895,N_3983);
xnor U4031 (N_4031,N_3753,N_3783);
and U4032 (N_4032,N_3841,N_3878);
nor U4033 (N_4033,N_3787,N_3803);
nand U4034 (N_4034,N_3899,N_3805);
and U4035 (N_4035,N_3768,N_3834);
nor U4036 (N_4036,N_3876,N_3840);
or U4037 (N_4037,N_3778,N_3993);
nand U4038 (N_4038,N_3770,N_3954);
and U4039 (N_4039,N_3821,N_3991);
and U4040 (N_4040,N_3891,N_3765);
nand U4041 (N_4041,N_3779,N_3965);
nand U4042 (N_4042,N_3844,N_3910);
or U4043 (N_4043,N_3827,N_3826);
xnor U4044 (N_4044,N_3836,N_3864);
and U4045 (N_4045,N_3911,N_3758);
xnor U4046 (N_4046,N_3929,N_3846);
xnor U4047 (N_4047,N_3843,N_3798);
and U4048 (N_4048,N_3964,N_3859);
xnor U4049 (N_4049,N_3855,N_3935);
xnor U4050 (N_4050,N_3801,N_3949);
nor U4051 (N_4051,N_3782,N_3934);
nand U4052 (N_4052,N_3863,N_3944);
xnor U4053 (N_4053,N_3815,N_3984);
nand U4054 (N_4054,N_3833,N_3909);
xnor U4055 (N_4055,N_3963,N_3870);
and U4056 (N_4056,N_3938,N_3913);
xnor U4057 (N_4057,N_3874,N_3988);
or U4058 (N_4058,N_3922,N_3989);
xnor U4059 (N_4059,N_3959,N_3777);
nor U4060 (N_4060,N_3974,N_3883);
nand U4061 (N_4061,N_3892,N_3987);
nor U4062 (N_4062,N_3767,N_3854);
and U4063 (N_4063,N_3957,N_3893);
or U4064 (N_4064,N_3918,N_3795);
xnor U4065 (N_4065,N_3978,N_3797);
nor U4066 (N_4066,N_3928,N_3894);
xnor U4067 (N_4067,N_3941,N_3849);
nand U4068 (N_4068,N_3868,N_3816);
or U4069 (N_4069,N_3769,N_3904);
xor U4070 (N_4070,N_3998,N_3939);
xnor U4071 (N_4071,N_3975,N_3948);
nor U4072 (N_4072,N_3900,N_3885);
or U4073 (N_4073,N_3804,N_3784);
or U4074 (N_4074,N_3757,N_3907);
xnor U4075 (N_4075,N_3809,N_3756);
nand U4076 (N_4076,N_3896,N_3831);
or U4077 (N_4077,N_3752,N_3890);
and U4078 (N_4078,N_3829,N_3817);
xor U4079 (N_4079,N_3999,N_3867);
and U4080 (N_4080,N_3755,N_3953);
and U4081 (N_4081,N_3932,N_3856);
nor U4082 (N_4082,N_3771,N_3995);
nand U4083 (N_4083,N_3789,N_3860);
and U4084 (N_4084,N_3773,N_3917);
and U4085 (N_4085,N_3980,N_3981);
nand U4086 (N_4086,N_3839,N_3952);
and U4087 (N_4087,N_3848,N_3920);
xor U4088 (N_4088,N_3881,N_3972);
xor U4089 (N_4089,N_3882,N_3780);
and U4090 (N_4090,N_3919,N_3781);
xor U4091 (N_4091,N_3985,N_3916);
and U4092 (N_4092,N_3992,N_3772);
or U4093 (N_4093,N_3921,N_3936);
and U4094 (N_4094,N_3811,N_3903);
nand U4095 (N_4095,N_3764,N_3956);
xnor U4096 (N_4096,N_3820,N_3937);
xnor U4097 (N_4097,N_3979,N_3793);
or U4098 (N_4098,N_3905,N_3818);
xnor U4099 (N_4099,N_3847,N_3925);
or U4100 (N_4100,N_3837,N_3926);
and U4101 (N_4101,N_3760,N_3887);
or U4102 (N_4102,N_3754,N_3792);
and U4103 (N_4103,N_3977,N_3813);
nand U4104 (N_4104,N_3852,N_3901);
or U4105 (N_4105,N_3955,N_3906);
nor U4106 (N_4106,N_3924,N_3845);
or U4107 (N_4107,N_3861,N_3799);
nand U4108 (N_4108,N_3884,N_3869);
nor U4109 (N_4109,N_3940,N_3915);
and U4110 (N_4110,N_3971,N_3788);
or U4111 (N_4111,N_3806,N_3931);
nand U4112 (N_4112,N_3812,N_3898);
or U4113 (N_4113,N_3790,N_3822);
or U4114 (N_4114,N_3832,N_3889);
or U4115 (N_4115,N_3774,N_3830);
xnor U4116 (N_4116,N_3838,N_3970);
nand U4117 (N_4117,N_3962,N_3791);
or U4118 (N_4118,N_3960,N_3933);
or U4119 (N_4119,N_3823,N_3762);
nand U4120 (N_4120,N_3912,N_3927);
xor U4121 (N_4121,N_3807,N_3858);
and U4122 (N_4122,N_3825,N_3947);
nand U4123 (N_4123,N_3802,N_3866);
nor U4124 (N_4124,N_3996,N_3945);
or U4125 (N_4125,N_3867,N_3783);
nand U4126 (N_4126,N_3960,N_3969);
nand U4127 (N_4127,N_3911,N_3982);
nand U4128 (N_4128,N_3954,N_3896);
xnor U4129 (N_4129,N_3867,N_3895);
xor U4130 (N_4130,N_3762,N_3787);
nor U4131 (N_4131,N_3909,N_3991);
nor U4132 (N_4132,N_3886,N_3990);
nor U4133 (N_4133,N_3928,N_3797);
nor U4134 (N_4134,N_3993,N_3785);
nand U4135 (N_4135,N_3981,N_3910);
and U4136 (N_4136,N_3902,N_3752);
and U4137 (N_4137,N_3887,N_3803);
nor U4138 (N_4138,N_3937,N_3916);
nor U4139 (N_4139,N_3840,N_3763);
and U4140 (N_4140,N_3984,N_3777);
xor U4141 (N_4141,N_3762,N_3972);
xor U4142 (N_4142,N_3756,N_3962);
and U4143 (N_4143,N_3830,N_3769);
or U4144 (N_4144,N_3810,N_3799);
and U4145 (N_4145,N_3799,N_3961);
or U4146 (N_4146,N_3992,N_3878);
and U4147 (N_4147,N_3759,N_3792);
xor U4148 (N_4148,N_3962,N_3970);
or U4149 (N_4149,N_3948,N_3875);
and U4150 (N_4150,N_3942,N_3806);
or U4151 (N_4151,N_3825,N_3830);
nand U4152 (N_4152,N_3775,N_3884);
nor U4153 (N_4153,N_3961,N_3954);
or U4154 (N_4154,N_3974,N_3794);
nor U4155 (N_4155,N_3848,N_3983);
nand U4156 (N_4156,N_3939,N_3830);
xnor U4157 (N_4157,N_3846,N_3754);
xor U4158 (N_4158,N_3887,N_3967);
nand U4159 (N_4159,N_3962,N_3841);
xor U4160 (N_4160,N_3816,N_3931);
xnor U4161 (N_4161,N_3993,N_3759);
and U4162 (N_4162,N_3929,N_3997);
or U4163 (N_4163,N_3797,N_3782);
xor U4164 (N_4164,N_3776,N_3807);
nor U4165 (N_4165,N_3863,N_3945);
nand U4166 (N_4166,N_3985,N_3804);
nor U4167 (N_4167,N_3910,N_3752);
or U4168 (N_4168,N_3929,N_3874);
and U4169 (N_4169,N_3914,N_3895);
or U4170 (N_4170,N_3838,N_3938);
and U4171 (N_4171,N_3910,N_3956);
nor U4172 (N_4172,N_3800,N_3760);
or U4173 (N_4173,N_3774,N_3789);
xnor U4174 (N_4174,N_3948,N_3985);
nor U4175 (N_4175,N_3994,N_3786);
nand U4176 (N_4176,N_3772,N_3944);
xnor U4177 (N_4177,N_3790,N_3968);
nor U4178 (N_4178,N_3830,N_3928);
nand U4179 (N_4179,N_3927,N_3793);
or U4180 (N_4180,N_3846,N_3951);
or U4181 (N_4181,N_3884,N_3954);
and U4182 (N_4182,N_3952,N_3895);
xnor U4183 (N_4183,N_3871,N_3925);
nor U4184 (N_4184,N_3905,N_3808);
nor U4185 (N_4185,N_3783,N_3916);
or U4186 (N_4186,N_3827,N_3879);
nand U4187 (N_4187,N_3771,N_3883);
nor U4188 (N_4188,N_3769,N_3782);
xnor U4189 (N_4189,N_3987,N_3860);
or U4190 (N_4190,N_3897,N_3791);
xor U4191 (N_4191,N_3953,N_3869);
xor U4192 (N_4192,N_3913,N_3917);
xnor U4193 (N_4193,N_3787,N_3870);
or U4194 (N_4194,N_3935,N_3958);
nor U4195 (N_4195,N_3974,N_3975);
xor U4196 (N_4196,N_3976,N_3982);
xor U4197 (N_4197,N_3998,N_3795);
and U4198 (N_4198,N_3752,N_3833);
nor U4199 (N_4199,N_3826,N_3944);
and U4200 (N_4200,N_3868,N_3947);
nor U4201 (N_4201,N_3763,N_3916);
xnor U4202 (N_4202,N_3912,N_3938);
or U4203 (N_4203,N_3815,N_3844);
xor U4204 (N_4204,N_3942,N_3764);
or U4205 (N_4205,N_3752,N_3886);
xor U4206 (N_4206,N_3771,N_3824);
xor U4207 (N_4207,N_3838,N_3827);
nand U4208 (N_4208,N_3868,N_3762);
xor U4209 (N_4209,N_3907,N_3807);
nand U4210 (N_4210,N_3799,N_3793);
xor U4211 (N_4211,N_3950,N_3836);
nand U4212 (N_4212,N_3797,N_3967);
and U4213 (N_4213,N_3754,N_3824);
nand U4214 (N_4214,N_3822,N_3983);
or U4215 (N_4215,N_3837,N_3839);
nand U4216 (N_4216,N_3993,N_3935);
xor U4217 (N_4217,N_3933,N_3964);
and U4218 (N_4218,N_3892,N_3950);
nand U4219 (N_4219,N_3849,N_3942);
nand U4220 (N_4220,N_3755,N_3872);
and U4221 (N_4221,N_3804,N_3956);
xor U4222 (N_4222,N_3855,N_3794);
or U4223 (N_4223,N_3843,N_3813);
nand U4224 (N_4224,N_3889,N_3783);
and U4225 (N_4225,N_3838,N_3899);
nor U4226 (N_4226,N_3965,N_3876);
xnor U4227 (N_4227,N_3862,N_3907);
xor U4228 (N_4228,N_3917,N_3751);
nand U4229 (N_4229,N_3809,N_3966);
and U4230 (N_4230,N_3881,N_3802);
nand U4231 (N_4231,N_3933,N_3883);
or U4232 (N_4232,N_3823,N_3787);
and U4233 (N_4233,N_3788,N_3882);
and U4234 (N_4234,N_3769,N_3844);
or U4235 (N_4235,N_3869,N_3983);
nand U4236 (N_4236,N_3945,N_3904);
xnor U4237 (N_4237,N_3999,N_3897);
nor U4238 (N_4238,N_3864,N_3878);
nor U4239 (N_4239,N_3750,N_3977);
nor U4240 (N_4240,N_3967,N_3995);
xnor U4241 (N_4241,N_3897,N_3856);
or U4242 (N_4242,N_3956,N_3937);
nor U4243 (N_4243,N_3908,N_3921);
xnor U4244 (N_4244,N_3981,N_3868);
xor U4245 (N_4245,N_3787,N_3779);
and U4246 (N_4246,N_3832,N_3783);
and U4247 (N_4247,N_3965,N_3961);
and U4248 (N_4248,N_3899,N_3820);
and U4249 (N_4249,N_3773,N_3805);
nand U4250 (N_4250,N_4047,N_4104);
nor U4251 (N_4251,N_4083,N_4182);
xor U4252 (N_4252,N_4185,N_4155);
xnor U4253 (N_4253,N_4124,N_4049);
nand U4254 (N_4254,N_4168,N_4203);
or U4255 (N_4255,N_4048,N_4023);
nand U4256 (N_4256,N_4019,N_4022);
xnor U4257 (N_4257,N_4177,N_4077);
and U4258 (N_4258,N_4141,N_4127);
and U4259 (N_4259,N_4175,N_4070);
nand U4260 (N_4260,N_4113,N_4016);
xnor U4261 (N_4261,N_4025,N_4217);
xor U4262 (N_4262,N_4146,N_4190);
xnor U4263 (N_4263,N_4241,N_4086);
xor U4264 (N_4264,N_4001,N_4231);
or U4265 (N_4265,N_4050,N_4209);
and U4266 (N_4266,N_4053,N_4243);
and U4267 (N_4267,N_4199,N_4205);
or U4268 (N_4268,N_4198,N_4115);
and U4269 (N_4269,N_4108,N_4102);
xor U4270 (N_4270,N_4100,N_4240);
nor U4271 (N_4271,N_4043,N_4040);
and U4272 (N_4272,N_4161,N_4044);
and U4273 (N_4273,N_4066,N_4029);
and U4274 (N_4274,N_4026,N_4009);
nand U4275 (N_4275,N_4105,N_4162);
xnor U4276 (N_4276,N_4111,N_4238);
nor U4277 (N_4277,N_4027,N_4193);
or U4278 (N_4278,N_4246,N_4219);
nor U4279 (N_4279,N_4008,N_4035);
xnor U4280 (N_4280,N_4129,N_4020);
xnor U4281 (N_4281,N_4189,N_4148);
or U4282 (N_4282,N_4072,N_4153);
nand U4283 (N_4283,N_4125,N_4114);
xor U4284 (N_4284,N_4051,N_4180);
nand U4285 (N_4285,N_4091,N_4166);
xnor U4286 (N_4286,N_4229,N_4096);
xnor U4287 (N_4287,N_4159,N_4173);
xnor U4288 (N_4288,N_4112,N_4076);
and U4289 (N_4289,N_4227,N_4233);
nand U4290 (N_4290,N_4088,N_4082);
nor U4291 (N_4291,N_4015,N_4164);
or U4292 (N_4292,N_4158,N_4207);
nor U4293 (N_4293,N_4143,N_4000);
or U4294 (N_4294,N_4041,N_4014);
or U4295 (N_4295,N_4213,N_4081);
xnor U4296 (N_4296,N_4117,N_4031);
nand U4297 (N_4297,N_4210,N_4071);
xor U4298 (N_4298,N_4055,N_4201);
xnor U4299 (N_4299,N_4157,N_4073);
xor U4300 (N_4300,N_4131,N_4099);
nor U4301 (N_4301,N_4140,N_4184);
nor U4302 (N_4302,N_4191,N_4196);
xnor U4303 (N_4303,N_4062,N_4216);
and U4304 (N_4304,N_4174,N_4080);
nand U4305 (N_4305,N_4060,N_4248);
xor U4306 (N_4306,N_4017,N_4186);
or U4307 (N_4307,N_4172,N_4065);
xnor U4308 (N_4308,N_4171,N_4085);
or U4309 (N_4309,N_4154,N_4002);
nor U4310 (N_4310,N_4068,N_4084);
or U4311 (N_4311,N_4223,N_4200);
nor U4312 (N_4312,N_4144,N_4107);
xnor U4313 (N_4313,N_4061,N_4003);
and U4314 (N_4314,N_4123,N_4024);
and U4315 (N_4315,N_4239,N_4006);
nor U4316 (N_4316,N_4056,N_4188);
nand U4317 (N_4317,N_4220,N_4206);
or U4318 (N_4318,N_4119,N_4244);
xor U4319 (N_4319,N_4093,N_4092);
nand U4320 (N_4320,N_4089,N_4110);
nor U4321 (N_4321,N_4234,N_4195);
or U4322 (N_4322,N_4042,N_4245);
xnor U4323 (N_4323,N_4218,N_4152);
and U4324 (N_4324,N_4018,N_4036);
or U4325 (N_4325,N_4067,N_4128);
or U4326 (N_4326,N_4054,N_4126);
nand U4327 (N_4327,N_4136,N_4121);
nor U4328 (N_4328,N_4098,N_4187);
nand U4329 (N_4329,N_4038,N_4212);
or U4330 (N_4330,N_4079,N_4087);
and U4331 (N_4331,N_4090,N_4074);
nand U4332 (N_4332,N_4028,N_4197);
xnor U4333 (N_4333,N_4094,N_4170);
and U4334 (N_4334,N_4147,N_4004);
nand U4335 (N_4335,N_4011,N_4075);
nor U4336 (N_4336,N_4134,N_4179);
xnor U4337 (N_4337,N_4225,N_4169);
or U4338 (N_4338,N_4010,N_4228);
nor U4339 (N_4339,N_4215,N_4226);
xor U4340 (N_4340,N_4192,N_4101);
nand U4341 (N_4341,N_4063,N_4237);
xor U4342 (N_4342,N_4130,N_4204);
or U4343 (N_4343,N_4052,N_4214);
and U4344 (N_4344,N_4142,N_4012);
and U4345 (N_4345,N_4135,N_4034);
or U4346 (N_4346,N_4167,N_4160);
and U4347 (N_4347,N_4005,N_4202);
or U4348 (N_4348,N_4097,N_4095);
and U4349 (N_4349,N_4132,N_4059);
nand U4350 (N_4350,N_4211,N_4194);
xor U4351 (N_4351,N_4176,N_4120);
and U4352 (N_4352,N_4138,N_4183);
nor U4353 (N_4353,N_4247,N_4178);
nand U4354 (N_4354,N_4030,N_4137);
or U4355 (N_4355,N_4116,N_4045);
xnor U4356 (N_4356,N_4232,N_4230);
nand U4357 (N_4357,N_4145,N_4133);
xor U4358 (N_4358,N_4069,N_4078);
and U4359 (N_4359,N_4222,N_4037);
xor U4360 (N_4360,N_4149,N_4032);
nand U4361 (N_4361,N_4165,N_4057);
and U4362 (N_4362,N_4007,N_4106);
nor U4363 (N_4363,N_4013,N_4208);
and U4364 (N_4364,N_4139,N_4221);
xor U4365 (N_4365,N_4236,N_4151);
and U4366 (N_4366,N_4242,N_4109);
nand U4367 (N_4367,N_4039,N_4058);
nand U4368 (N_4368,N_4249,N_4224);
xnor U4369 (N_4369,N_4118,N_4163);
nor U4370 (N_4370,N_4122,N_4033);
or U4371 (N_4371,N_4156,N_4103);
or U4372 (N_4372,N_4181,N_4046);
and U4373 (N_4373,N_4021,N_4235);
nand U4374 (N_4374,N_4064,N_4150);
nand U4375 (N_4375,N_4189,N_4193);
or U4376 (N_4376,N_4186,N_4022);
xor U4377 (N_4377,N_4193,N_4085);
nor U4378 (N_4378,N_4162,N_4066);
nand U4379 (N_4379,N_4210,N_4104);
and U4380 (N_4380,N_4012,N_4067);
and U4381 (N_4381,N_4052,N_4059);
nand U4382 (N_4382,N_4009,N_4205);
or U4383 (N_4383,N_4010,N_4022);
nand U4384 (N_4384,N_4190,N_4249);
nand U4385 (N_4385,N_4017,N_4078);
nor U4386 (N_4386,N_4054,N_4222);
and U4387 (N_4387,N_4113,N_4077);
or U4388 (N_4388,N_4195,N_4164);
nor U4389 (N_4389,N_4141,N_4022);
and U4390 (N_4390,N_4230,N_4018);
and U4391 (N_4391,N_4109,N_4238);
nand U4392 (N_4392,N_4170,N_4131);
nor U4393 (N_4393,N_4068,N_4046);
xor U4394 (N_4394,N_4186,N_4233);
xor U4395 (N_4395,N_4123,N_4179);
nand U4396 (N_4396,N_4117,N_4178);
nand U4397 (N_4397,N_4163,N_4222);
nand U4398 (N_4398,N_4200,N_4114);
nor U4399 (N_4399,N_4109,N_4110);
nand U4400 (N_4400,N_4108,N_4152);
xor U4401 (N_4401,N_4096,N_4054);
xor U4402 (N_4402,N_4027,N_4070);
nand U4403 (N_4403,N_4221,N_4070);
nor U4404 (N_4404,N_4131,N_4026);
xnor U4405 (N_4405,N_4248,N_4155);
xor U4406 (N_4406,N_4016,N_4028);
and U4407 (N_4407,N_4164,N_4004);
xnor U4408 (N_4408,N_4151,N_4094);
and U4409 (N_4409,N_4016,N_4112);
and U4410 (N_4410,N_4206,N_4145);
xnor U4411 (N_4411,N_4111,N_4149);
nand U4412 (N_4412,N_4045,N_4214);
and U4413 (N_4413,N_4117,N_4097);
xnor U4414 (N_4414,N_4020,N_4204);
nor U4415 (N_4415,N_4197,N_4099);
and U4416 (N_4416,N_4166,N_4036);
and U4417 (N_4417,N_4170,N_4114);
nand U4418 (N_4418,N_4003,N_4002);
nor U4419 (N_4419,N_4069,N_4157);
nor U4420 (N_4420,N_4203,N_4034);
nor U4421 (N_4421,N_4202,N_4131);
nand U4422 (N_4422,N_4096,N_4099);
or U4423 (N_4423,N_4232,N_4226);
and U4424 (N_4424,N_4093,N_4119);
xnor U4425 (N_4425,N_4038,N_4158);
or U4426 (N_4426,N_4131,N_4081);
or U4427 (N_4427,N_4126,N_4087);
and U4428 (N_4428,N_4185,N_4142);
xnor U4429 (N_4429,N_4197,N_4190);
and U4430 (N_4430,N_4073,N_4094);
nor U4431 (N_4431,N_4158,N_4063);
nor U4432 (N_4432,N_4132,N_4035);
or U4433 (N_4433,N_4191,N_4061);
or U4434 (N_4434,N_4209,N_4006);
and U4435 (N_4435,N_4219,N_4004);
nor U4436 (N_4436,N_4154,N_4006);
xor U4437 (N_4437,N_4009,N_4116);
nor U4438 (N_4438,N_4050,N_4105);
xnor U4439 (N_4439,N_4051,N_4005);
and U4440 (N_4440,N_4078,N_4056);
or U4441 (N_4441,N_4000,N_4128);
xnor U4442 (N_4442,N_4092,N_4142);
or U4443 (N_4443,N_4146,N_4020);
nand U4444 (N_4444,N_4064,N_4151);
nand U4445 (N_4445,N_4218,N_4177);
and U4446 (N_4446,N_4193,N_4190);
nor U4447 (N_4447,N_4158,N_4013);
nand U4448 (N_4448,N_4185,N_4229);
nor U4449 (N_4449,N_4201,N_4131);
or U4450 (N_4450,N_4197,N_4206);
and U4451 (N_4451,N_4145,N_4172);
nand U4452 (N_4452,N_4131,N_4236);
nor U4453 (N_4453,N_4095,N_4118);
and U4454 (N_4454,N_4176,N_4077);
nand U4455 (N_4455,N_4138,N_4206);
and U4456 (N_4456,N_4100,N_4112);
xor U4457 (N_4457,N_4245,N_4249);
or U4458 (N_4458,N_4207,N_4049);
xor U4459 (N_4459,N_4078,N_4049);
nand U4460 (N_4460,N_4093,N_4207);
and U4461 (N_4461,N_4001,N_4166);
nor U4462 (N_4462,N_4206,N_4234);
nor U4463 (N_4463,N_4231,N_4150);
or U4464 (N_4464,N_4000,N_4058);
and U4465 (N_4465,N_4005,N_4249);
nor U4466 (N_4466,N_4036,N_4059);
nand U4467 (N_4467,N_4239,N_4109);
xnor U4468 (N_4468,N_4123,N_4011);
nor U4469 (N_4469,N_4107,N_4103);
nor U4470 (N_4470,N_4152,N_4060);
or U4471 (N_4471,N_4230,N_4058);
nand U4472 (N_4472,N_4016,N_4171);
and U4473 (N_4473,N_4150,N_4157);
or U4474 (N_4474,N_4242,N_4233);
nor U4475 (N_4475,N_4023,N_4123);
xnor U4476 (N_4476,N_4080,N_4118);
and U4477 (N_4477,N_4103,N_4203);
nor U4478 (N_4478,N_4059,N_4207);
nor U4479 (N_4479,N_4055,N_4086);
nor U4480 (N_4480,N_4204,N_4015);
xor U4481 (N_4481,N_4241,N_4110);
or U4482 (N_4482,N_4074,N_4196);
nor U4483 (N_4483,N_4194,N_4119);
nor U4484 (N_4484,N_4209,N_4068);
nor U4485 (N_4485,N_4060,N_4007);
nor U4486 (N_4486,N_4026,N_4016);
nand U4487 (N_4487,N_4131,N_4180);
nand U4488 (N_4488,N_4066,N_4013);
xnor U4489 (N_4489,N_4133,N_4244);
nand U4490 (N_4490,N_4214,N_4123);
xnor U4491 (N_4491,N_4129,N_4196);
or U4492 (N_4492,N_4014,N_4102);
or U4493 (N_4493,N_4129,N_4092);
or U4494 (N_4494,N_4119,N_4086);
nand U4495 (N_4495,N_4129,N_4014);
nor U4496 (N_4496,N_4089,N_4209);
or U4497 (N_4497,N_4128,N_4031);
and U4498 (N_4498,N_4113,N_4187);
or U4499 (N_4499,N_4201,N_4128);
or U4500 (N_4500,N_4484,N_4342);
or U4501 (N_4501,N_4489,N_4469);
nand U4502 (N_4502,N_4452,N_4471);
nand U4503 (N_4503,N_4395,N_4426);
nor U4504 (N_4504,N_4305,N_4450);
and U4505 (N_4505,N_4329,N_4333);
and U4506 (N_4506,N_4390,N_4495);
nand U4507 (N_4507,N_4366,N_4492);
or U4508 (N_4508,N_4257,N_4465);
nand U4509 (N_4509,N_4360,N_4377);
xnor U4510 (N_4510,N_4434,N_4293);
and U4511 (N_4511,N_4253,N_4481);
and U4512 (N_4512,N_4255,N_4267);
and U4513 (N_4513,N_4499,N_4336);
and U4514 (N_4514,N_4361,N_4449);
nor U4515 (N_4515,N_4472,N_4440);
nand U4516 (N_4516,N_4370,N_4418);
nor U4517 (N_4517,N_4467,N_4468);
xor U4518 (N_4518,N_4381,N_4261);
xor U4519 (N_4519,N_4274,N_4455);
nor U4520 (N_4520,N_4308,N_4345);
nand U4521 (N_4521,N_4337,N_4362);
xor U4522 (N_4522,N_4463,N_4276);
nor U4523 (N_4523,N_4351,N_4436);
or U4524 (N_4524,N_4454,N_4414);
nor U4525 (N_4525,N_4421,N_4363);
xnor U4526 (N_4526,N_4392,N_4335);
xnor U4527 (N_4527,N_4283,N_4396);
xor U4528 (N_4528,N_4314,N_4427);
and U4529 (N_4529,N_4394,N_4376);
nand U4530 (N_4530,N_4411,N_4295);
xor U4531 (N_4531,N_4324,N_4288);
xnor U4532 (N_4532,N_4493,N_4458);
nor U4533 (N_4533,N_4358,N_4278);
and U4534 (N_4534,N_4289,N_4309);
nor U4535 (N_4535,N_4425,N_4387);
or U4536 (N_4536,N_4321,N_4432);
nand U4537 (N_4537,N_4483,N_4316);
xnor U4538 (N_4538,N_4273,N_4339);
and U4539 (N_4539,N_4397,N_4413);
nor U4540 (N_4540,N_4400,N_4490);
or U4541 (N_4541,N_4447,N_4417);
xor U4542 (N_4542,N_4429,N_4422);
or U4543 (N_4543,N_4254,N_4457);
or U4544 (N_4544,N_4344,N_4486);
or U4545 (N_4545,N_4343,N_4444);
nor U4546 (N_4546,N_4372,N_4327);
and U4547 (N_4547,N_4439,N_4476);
xnor U4548 (N_4548,N_4350,N_4258);
nand U4549 (N_4549,N_4298,N_4412);
nor U4550 (N_4550,N_4431,N_4306);
xor U4551 (N_4551,N_4252,N_4259);
or U4552 (N_4552,N_4389,N_4250);
nor U4553 (N_4553,N_4386,N_4275);
nand U4554 (N_4554,N_4485,N_4368);
or U4555 (N_4555,N_4263,N_4311);
nand U4556 (N_4556,N_4374,N_4369);
xnor U4557 (N_4557,N_4320,N_4357);
nor U4558 (N_4558,N_4364,N_4460);
nor U4559 (N_4559,N_4367,N_4302);
nand U4560 (N_4560,N_4494,N_4262);
and U4561 (N_4561,N_4282,N_4317);
nor U4562 (N_4562,N_4496,N_4269);
or U4563 (N_4563,N_4281,N_4319);
nand U4564 (N_4564,N_4433,N_4446);
and U4565 (N_4565,N_4488,N_4297);
nor U4566 (N_4566,N_4409,N_4277);
or U4567 (N_4567,N_4478,N_4470);
nand U4568 (N_4568,N_4415,N_4286);
or U4569 (N_4569,N_4264,N_4299);
and U4570 (N_4570,N_4294,N_4430);
nor U4571 (N_4571,N_4420,N_4441);
nand U4572 (N_4572,N_4371,N_4315);
nor U4573 (N_4573,N_4466,N_4325);
or U4574 (N_4574,N_4338,N_4428);
nand U4575 (N_4575,N_4347,N_4323);
xor U4576 (N_4576,N_4405,N_4380);
or U4577 (N_4577,N_4328,N_4379);
xnor U4578 (N_4578,N_4391,N_4353);
xor U4579 (N_4579,N_4475,N_4408);
nand U4580 (N_4580,N_4419,N_4404);
xor U4581 (N_4581,N_4318,N_4473);
nor U4582 (N_4582,N_4416,N_4442);
nor U4583 (N_4583,N_4385,N_4406);
or U4584 (N_4584,N_4340,N_4291);
and U4585 (N_4585,N_4296,N_4453);
nand U4586 (N_4586,N_4352,N_4266);
or U4587 (N_4587,N_4498,N_4304);
nand U4588 (N_4588,N_4355,N_4265);
xor U4589 (N_4589,N_4334,N_4497);
nor U4590 (N_4590,N_4410,N_4349);
nand U4591 (N_4591,N_4402,N_4407);
and U4592 (N_4592,N_4383,N_4403);
xnor U4593 (N_4593,N_4401,N_4456);
nand U4594 (N_4594,N_4326,N_4399);
or U4595 (N_4595,N_4365,N_4448);
and U4596 (N_4596,N_4443,N_4310);
xor U4597 (N_4597,N_4346,N_4437);
xor U4598 (N_4598,N_4331,N_4307);
or U4599 (N_4599,N_4279,N_4424);
xnor U4600 (N_4600,N_4375,N_4312);
nor U4601 (N_4601,N_4445,N_4271);
xnor U4602 (N_4602,N_4303,N_4341);
nor U4603 (N_4603,N_4354,N_4474);
nor U4604 (N_4604,N_4462,N_4251);
nor U4605 (N_4605,N_4459,N_4464);
nor U4606 (N_4606,N_4268,N_4348);
nor U4607 (N_4607,N_4270,N_4290);
nand U4608 (N_4608,N_4287,N_4256);
or U4609 (N_4609,N_4480,N_4332);
and U4610 (N_4610,N_4451,N_4435);
and U4611 (N_4611,N_4313,N_4322);
nor U4612 (N_4612,N_4285,N_4482);
nand U4613 (N_4613,N_4260,N_4423);
nand U4614 (N_4614,N_4284,N_4292);
or U4615 (N_4615,N_4388,N_4438);
or U4616 (N_4616,N_4301,N_4356);
nor U4617 (N_4617,N_4378,N_4398);
nand U4618 (N_4618,N_4393,N_4300);
xnor U4619 (N_4619,N_4373,N_4384);
or U4620 (N_4620,N_4382,N_4461);
nand U4621 (N_4621,N_4359,N_4491);
nand U4622 (N_4622,N_4272,N_4479);
or U4623 (N_4623,N_4330,N_4280);
nor U4624 (N_4624,N_4477,N_4487);
xor U4625 (N_4625,N_4409,N_4297);
nor U4626 (N_4626,N_4271,N_4402);
nor U4627 (N_4627,N_4494,N_4253);
nand U4628 (N_4628,N_4489,N_4397);
nand U4629 (N_4629,N_4447,N_4299);
and U4630 (N_4630,N_4476,N_4462);
nor U4631 (N_4631,N_4412,N_4497);
or U4632 (N_4632,N_4487,N_4316);
or U4633 (N_4633,N_4324,N_4365);
nand U4634 (N_4634,N_4273,N_4487);
nor U4635 (N_4635,N_4475,N_4343);
nand U4636 (N_4636,N_4342,N_4278);
xnor U4637 (N_4637,N_4368,N_4289);
nor U4638 (N_4638,N_4296,N_4256);
and U4639 (N_4639,N_4359,N_4317);
or U4640 (N_4640,N_4350,N_4486);
xor U4641 (N_4641,N_4475,N_4332);
and U4642 (N_4642,N_4398,N_4329);
xnor U4643 (N_4643,N_4407,N_4436);
or U4644 (N_4644,N_4263,N_4488);
or U4645 (N_4645,N_4417,N_4319);
xnor U4646 (N_4646,N_4459,N_4331);
nand U4647 (N_4647,N_4391,N_4259);
xor U4648 (N_4648,N_4365,N_4412);
or U4649 (N_4649,N_4322,N_4403);
nor U4650 (N_4650,N_4305,N_4270);
xnor U4651 (N_4651,N_4490,N_4300);
nor U4652 (N_4652,N_4270,N_4325);
xnor U4653 (N_4653,N_4396,N_4355);
or U4654 (N_4654,N_4367,N_4370);
nor U4655 (N_4655,N_4411,N_4328);
xnor U4656 (N_4656,N_4337,N_4348);
nand U4657 (N_4657,N_4352,N_4357);
nand U4658 (N_4658,N_4413,N_4298);
and U4659 (N_4659,N_4256,N_4273);
or U4660 (N_4660,N_4307,N_4482);
xor U4661 (N_4661,N_4378,N_4346);
nor U4662 (N_4662,N_4363,N_4418);
and U4663 (N_4663,N_4259,N_4452);
nor U4664 (N_4664,N_4489,N_4442);
xnor U4665 (N_4665,N_4272,N_4384);
nor U4666 (N_4666,N_4253,N_4406);
or U4667 (N_4667,N_4293,N_4289);
or U4668 (N_4668,N_4283,N_4398);
and U4669 (N_4669,N_4276,N_4330);
nand U4670 (N_4670,N_4491,N_4494);
nor U4671 (N_4671,N_4458,N_4416);
nor U4672 (N_4672,N_4375,N_4351);
and U4673 (N_4673,N_4398,N_4438);
xor U4674 (N_4674,N_4306,N_4398);
and U4675 (N_4675,N_4336,N_4304);
nor U4676 (N_4676,N_4499,N_4274);
nand U4677 (N_4677,N_4281,N_4296);
and U4678 (N_4678,N_4493,N_4367);
nand U4679 (N_4679,N_4387,N_4436);
xnor U4680 (N_4680,N_4271,N_4332);
nor U4681 (N_4681,N_4372,N_4319);
nand U4682 (N_4682,N_4308,N_4417);
nor U4683 (N_4683,N_4311,N_4497);
xnor U4684 (N_4684,N_4469,N_4415);
and U4685 (N_4685,N_4435,N_4453);
and U4686 (N_4686,N_4419,N_4254);
and U4687 (N_4687,N_4334,N_4255);
nand U4688 (N_4688,N_4412,N_4438);
or U4689 (N_4689,N_4335,N_4311);
or U4690 (N_4690,N_4329,N_4480);
xor U4691 (N_4691,N_4364,N_4499);
nand U4692 (N_4692,N_4482,N_4463);
nor U4693 (N_4693,N_4499,N_4467);
or U4694 (N_4694,N_4350,N_4389);
nand U4695 (N_4695,N_4496,N_4388);
or U4696 (N_4696,N_4318,N_4257);
nor U4697 (N_4697,N_4324,N_4494);
nor U4698 (N_4698,N_4405,N_4404);
nand U4699 (N_4699,N_4442,N_4456);
and U4700 (N_4700,N_4293,N_4416);
nor U4701 (N_4701,N_4454,N_4482);
nand U4702 (N_4702,N_4411,N_4282);
or U4703 (N_4703,N_4373,N_4446);
and U4704 (N_4704,N_4286,N_4450);
and U4705 (N_4705,N_4406,N_4431);
nand U4706 (N_4706,N_4340,N_4383);
nand U4707 (N_4707,N_4432,N_4437);
nand U4708 (N_4708,N_4313,N_4433);
nor U4709 (N_4709,N_4356,N_4458);
or U4710 (N_4710,N_4319,N_4460);
nor U4711 (N_4711,N_4451,N_4364);
xnor U4712 (N_4712,N_4384,N_4381);
or U4713 (N_4713,N_4298,N_4447);
or U4714 (N_4714,N_4366,N_4430);
nand U4715 (N_4715,N_4272,N_4473);
or U4716 (N_4716,N_4401,N_4361);
nor U4717 (N_4717,N_4393,N_4258);
nor U4718 (N_4718,N_4287,N_4343);
and U4719 (N_4719,N_4264,N_4411);
nand U4720 (N_4720,N_4493,N_4313);
xor U4721 (N_4721,N_4349,N_4451);
and U4722 (N_4722,N_4441,N_4439);
nand U4723 (N_4723,N_4450,N_4304);
nand U4724 (N_4724,N_4397,N_4456);
xnor U4725 (N_4725,N_4263,N_4270);
or U4726 (N_4726,N_4491,N_4326);
nor U4727 (N_4727,N_4354,N_4430);
and U4728 (N_4728,N_4378,N_4431);
and U4729 (N_4729,N_4364,N_4430);
or U4730 (N_4730,N_4337,N_4285);
or U4731 (N_4731,N_4485,N_4371);
and U4732 (N_4732,N_4282,N_4492);
or U4733 (N_4733,N_4433,N_4481);
nor U4734 (N_4734,N_4345,N_4266);
or U4735 (N_4735,N_4475,N_4349);
and U4736 (N_4736,N_4435,N_4395);
nand U4737 (N_4737,N_4317,N_4394);
nor U4738 (N_4738,N_4310,N_4378);
nand U4739 (N_4739,N_4382,N_4276);
or U4740 (N_4740,N_4465,N_4453);
nor U4741 (N_4741,N_4339,N_4375);
and U4742 (N_4742,N_4364,N_4377);
nor U4743 (N_4743,N_4316,N_4369);
or U4744 (N_4744,N_4250,N_4253);
or U4745 (N_4745,N_4465,N_4254);
nand U4746 (N_4746,N_4327,N_4484);
nor U4747 (N_4747,N_4422,N_4277);
nand U4748 (N_4748,N_4472,N_4417);
nand U4749 (N_4749,N_4292,N_4465);
xnor U4750 (N_4750,N_4707,N_4675);
or U4751 (N_4751,N_4689,N_4506);
or U4752 (N_4752,N_4623,N_4664);
nor U4753 (N_4753,N_4740,N_4609);
nand U4754 (N_4754,N_4570,N_4644);
and U4755 (N_4755,N_4723,N_4586);
or U4756 (N_4756,N_4666,N_4731);
nor U4757 (N_4757,N_4631,N_4533);
nand U4758 (N_4758,N_4507,N_4656);
or U4759 (N_4759,N_4538,N_4571);
nand U4760 (N_4760,N_4554,N_4640);
xnor U4761 (N_4761,N_4677,N_4564);
nand U4762 (N_4762,N_4706,N_4509);
and U4763 (N_4763,N_4648,N_4712);
xor U4764 (N_4764,N_4622,N_4702);
xor U4765 (N_4765,N_4526,N_4663);
nor U4766 (N_4766,N_4659,N_4651);
nor U4767 (N_4767,N_4693,N_4572);
xnor U4768 (N_4768,N_4634,N_4715);
and U4769 (N_4769,N_4713,N_4661);
xnor U4770 (N_4770,N_4552,N_4558);
and U4771 (N_4771,N_4515,N_4510);
nand U4772 (N_4772,N_4624,N_4735);
nand U4773 (N_4773,N_4670,N_4620);
nand U4774 (N_4774,N_4692,N_4699);
or U4775 (N_4775,N_4589,N_4512);
or U4776 (N_4776,N_4528,N_4744);
and U4777 (N_4777,N_4683,N_4685);
or U4778 (N_4778,N_4690,N_4592);
nand U4779 (N_4779,N_4732,N_4601);
xor U4780 (N_4780,N_4652,N_4730);
and U4781 (N_4781,N_4700,N_4544);
and U4782 (N_4782,N_4524,N_4567);
xnor U4783 (N_4783,N_4614,N_4579);
nor U4784 (N_4784,N_4698,N_4657);
nor U4785 (N_4785,N_4696,N_4574);
nor U4786 (N_4786,N_4518,N_4610);
or U4787 (N_4787,N_4514,N_4697);
or U4788 (N_4788,N_4537,N_4674);
nand U4789 (N_4789,N_4708,N_4501);
or U4790 (N_4790,N_4709,N_4569);
and U4791 (N_4791,N_4637,N_4555);
or U4792 (N_4792,N_4695,N_4556);
or U4793 (N_4793,N_4549,N_4653);
xor U4794 (N_4794,N_4673,N_4546);
xor U4795 (N_4795,N_4517,N_4676);
nor U4796 (N_4796,N_4655,N_4600);
and U4797 (N_4797,N_4604,N_4545);
xnor U4798 (N_4798,N_4532,N_4523);
nand U4799 (N_4799,N_4606,N_4611);
and U4800 (N_4800,N_4626,N_4748);
nand U4801 (N_4801,N_4503,N_4671);
xor U4802 (N_4802,N_4553,N_4627);
xor U4803 (N_4803,N_4691,N_4582);
nor U4804 (N_4804,N_4585,N_4703);
nand U4805 (N_4805,N_4728,N_4565);
xnor U4806 (N_4806,N_4628,N_4743);
and U4807 (N_4807,N_4568,N_4608);
xnor U4808 (N_4808,N_4649,N_4688);
or U4809 (N_4809,N_4590,N_4641);
xor U4810 (N_4810,N_4662,N_4660);
xor U4811 (N_4811,N_4531,N_4643);
nand U4812 (N_4812,N_4529,N_4605);
nor U4813 (N_4813,N_4629,N_4535);
nand U4814 (N_4814,N_4591,N_4642);
or U4815 (N_4815,N_4513,N_4598);
nand U4816 (N_4816,N_4678,N_4504);
xnor U4817 (N_4817,N_4551,N_4541);
xor U4818 (N_4818,N_4741,N_4718);
xnor U4819 (N_4819,N_4632,N_4701);
nor U4820 (N_4820,N_4733,N_4502);
xnor U4821 (N_4821,N_4746,N_4617);
nand U4822 (N_4822,N_4658,N_4596);
and U4823 (N_4823,N_4527,N_4505);
nor U4824 (N_4824,N_4667,N_4520);
and U4825 (N_4825,N_4721,N_4516);
and U4826 (N_4826,N_4542,N_4638);
nand U4827 (N_4827,N_4665,N_4588);
and U4828 (N_4828,N_4540,N_4563);
or U4829 (N_4829,N_4726,N_4684);
or U4830 (N_4830,N_4716,N_4580);
nor U4831 (N_4831,N_4749,N_4725);
or U4832 (N_4832,N_4560,N_4704);
xor U4833 (N_4833,N_4602,N_4714);
nand U4834 (N_4834,N_4736,N_4584);
and U4835 (N_4835,N_4550,N_4742);
or U4836 (N_4836,N_4682,N_4630);
nor U4837 (N_4837,N_4561,N_4616);
xor U4838 (N_4838,N_4615,N_4687);
and U4839 (N_4839,N_4508,N_4668);
nor U4840 (N_4840,N_4686,N_4747);
or U4841 (N_4841,N_4633,N_4647);
or U4842 (N_4842,N_4618,N_4521);
xnor U4843 (N_4843,N_4619,N_4672);
and U4844 (N_4844,N_4737,N_4650);
nor U4845 (N_4845,N_4621,N_4613);
and U4846 (N_4846,N_4727,N_4511);
xnor U4847 (N_4847,N_4625,N_4587);
and U4848 (N_4848,N_4680,N_4557);
and U4849 (N_4849,N_4578,N_4738);
and U4850 (N_4850,N_4577,N_4519);
or U4851 (N_4851,N_4681,N_4720);
xnor U4852 (N_4852,N_4562,N_4539);
nor U4853 (N_4853,N_4534,N_4612);
nor U4854 (N_4854,N_4581,N_4724);
and U4855 (N_4855,N_4593,N_4635);
or U4856 (N_4856,N_4729,N_4717);
nor U4857 (N_4857,N_4710,N_4575);
xor U4858 (N_4858,N_4603,N_4719);
nand U4859 (N_4859,N_4576,N_4694);
nor U4860 (N_4860,N_4745,N_4734);
or U4861 (N_4861,N_4522,N_4500);
nor U4862 (N_4862,N_4711,N_4594);
and U4863 (N_4863,N_4646,N_4645);
nor U4864 (N_4864,N_4530,N_4525);
xnor U4865 (N_4865,N_4599,N_4583);
nand U4866 (N_4866,N_4597,N_4595);
nor U4867 (N_4867,N_4536,N_4636);
or U4868 (N_4868,N_4654,N_4639);
or U4869 (N_4869,N_4679,N_4547);
xnor U4870 (N_4870,N_4543,N_4607);
nor U4871 (N_4871,N_4573,N_4722);
xnor U4872 (N_4872,N_4739,N_4669);
xnor U4873 (N_4873,N_4559,N_4705);
and U4874 (N_4874,N_4566,N_4548);
nor U4875 (N_4875,N_4555,N_4700);
and U4876 (N_4876,N_4549,N_4658);
or U4877 (N_4877,N_4528,N_4735);
xor U4878 (N_4878,N_4576,N_4658);
or U4879 (N_4879,N_4632,N_4630);
and U4880 (N_4880,N_4731,N_4558);
xnor U4881 (N_4881,N_4507,N_4532);
nor U4882 (N_4882,N_4502,N_4674);
nor U4883 (N_4883,N_4528,N_4521);
and U4884 (N_4884,N_4505,N_4730);
and U4885 (N_4885,N_4652,N_4595);
and U4886 (N_4886,N_4660,N_4686);
nor U4887 (N_4887,N_4658,N_4749);
nand U4888 (N_4888,N_4667,N_4690);
and U4889 (N_4889,N_4621,N_4638);
or U4890 (N_4890,N_4511,N_4546);
xnor U4891 (N_4891,N_4619,N_4595);
and U4892 (N_4892,N_4651,N_4664);
nand U4893 (N_4893,N_4606,N_4600);
or U4894 (N_4894,N_4587,N_4624);
or U4895 (N_4895,N_4585,N_4506);
nor U4896 (N_4896,N_4511,N_4506);
nand U4897 (N_4897,N_4572,N_4698);
xnor U4898 (N_4898,N_4623,N_4579);
and U4899 (N_4899,N_4558,N_4631);
or U4900 (N_4900,N_4502,N_4520);
xor U4901 (N_4901,N_4680,N_4672);
nor U4902 (N_4902,N_4538,N_4505);
xor U4903 (N_4903,N_4735,N_4663);
nand U4904 (N_4904,N_4731,N_4703);
nand U4905 (N_4905,N_4687,N_4731);
nor U4906 (N_4906,N_4719,N_4665);
nor U4907 (N_4907,N_4593,N_4597);
or U4908 (N_4908,N_4706,N_4671);
nand U4909 (N_4909,N_4690,N_4550);
xor U4910 (N_4910,N_4655,N_4537);
or U4911 (N_4911,N_4703,N_4663);
or U4912 (N_4912,N_4745,N_4609);
or U4913 (N_4913,N_4690,N_4653);
nor U4914 (N_4914,N_4737,N_4581);
nand U4915 (N_4915,N_4515,N_4627);
or U4916 (N_4916,N_4520,N_4728);
nor U4917 (N_4917,N_4659,N_4693);
nor U4918 (N_4918,N_4677,N_4603);
nor U4919 (N_4919,N_4625,N_4686);
or U4920 (N_4920,N_4542,N_4703);
nand U4921 (N_4921,N_4547,N_4732);
nor U4922 (N_4922,N_4510,N_4530);
nand U4923 (N_4923,N_4721,N_4540);
nand U4924 (N_4924,N_4588,N_4708);
nand U4925 (N_4925,N_4639,N_4540);
xor U4926 (N_4926,N_4545,N_4637);
or U4927 (N_4927,N_4518,N_4532);
xor U4928 (N_4928,N_4737,N_4613);
and U4929 (N_4929,N_4553,N_4524);
or U4930 (N_4930,N_4609,N_4730);
xor U4931 (N_4931,N_4644,N_4623);
or U4932 (N_4932,N_4725,N_4640);
and U4933 (N_4933,N_4672,N_4616);
nand U4934 (N_4934,N_4602,N_4729);
xnor U4935 (N_4935,N_4739,N_4636);
nand U4936 (N_4936,N_4700,N_4643);
and U4937 (N_4937,N_4652,N_4617);
and U4938 (N_4938,N_4623,N_4611);
nand U4939 (N_4939,N_4702,N_4577);
nand U4940 (N_4940,N_4667,N_4688);
nor U4941 (N_4941,N_4621,N_4603);
nor U4942 (N_4942,N_4568,N_4746);
or U4943 (N_4943,N_4711,N_4661);
nor U4944 (N_4944,N_4516,N_4593);
nand U4945 (N_4945,N_4529,N_4597);
xnor U4946 (N_4946,N_4616,N_4607);
and U4947 (N_4947,N_4703,N_4584);
nor U4948 (N_4948,N_4625,N_4629);
or U4949 (N_4949,N_4591,N_4698);
nor U4950 (N_4950,N_4738,N_4748);
or U4951 (N_4951,N_4632,N_4697);
xor U4952 (N_4952,N_4711,N_4663);
and U4953 (N_4953,N_4541,N_4554);
xnor U4954 (N_4954,N_4705,N_4723);
nor U4955 (N_4955,N_4714,N_4640);
xor U4956 (N_4956,N_4501,N_4722);
xnor U4957 (N_4957,N_4660,N_4628);
and U4958 (N_4958,N_4547,N_4610);
or U4959 (N_4959,N_4748,N_4647);
and U4960 (N_4960,N_4683,N_4640);
and U4961 (N_4961,N_4524,N_4612);
nor U4962 (N_4962,N_4648,N_4735);
nor U4963 (N_4963,N_4509,N_4679);
nand U4964 (N_4964,N_4537,N_4721);
or U4965 (N_4965,N_4545,N_4523);
nand U4966 (N_4966,N_4587,N_4567);
nor U4967 (N_4967,N_4507,N_4598);
and U4968 (N_4968,N_4561,N_4579);
and U4969 (N_4969,N_4742,N_4609);
nand U4970 (N_4970,N_4680,N_4594);
and U4971 (N_4971,N_4653,N_4517);
xor U4972 (N_4972,N_4657,N_4633);
or U4973 (N_4973,N_4689,N_4647);
or U4974 (N_4974,N_4683,N_4665);
nand U4975 (N_4975,N_4596,N_4720);
or U4976 (N_4976,N_4681,N_4524);
or U4977 (N_4977,N_4716,N_4637);
and U4978 (N_4978,N_4510,N_4685);
xnor U4979 (N_4979,N_4748,N_4637);
and U4980 (N_4980,N_4676,N_4526);
xor U4981 (N_4981,N_4510,N_4527);
or U4982 (N_4982,N_4586,N_4634);
xor U4983 (N_4983,N_4569,N_4651);
nor U4984 (N_4984,N_4713,N_4620);
nor U4985 (N_4985,N_4644,N_4689);
xor U4986 (N_4986,N_4582,N_4679);
nand U4987 (N_4987,N_4506,N_4561);
nand U4988 (N_4988,N_4665,N_4618);
or U4989 (N_4989,N_4714,N_4707);
and U4990 (N_4990,N_4622,N_4663);
xnor U4991 (N_4991,N_4744,N_4663);
nor U4992 (N_4992,N_4502,N_4663);
xor U4993 (N_4993,N_4621,N_4668);
nor U4994 (N_4994,N_4692,N_4727);
and U4995 (N_4995,N_4548,N_4746);
or U4996 (N_4996,N_4538,N_4568);
or U4997 (N_4997,N_4671,N_4743);
nor U4998 (N_4998,N_4588,N_4582);
xnor U4999 (N_4999,N_4612,N_4642);
and U5000 (N_5000,N_4785,N_4877);
and U5001 (N_5001,N_4885,N_4818);
and U5002 (N_5002,N_4899,N_4850);
nand U5003 (N_5003,N_4772,N_4894);
nor U5004 (N_5004,N_4790,N_4838);
xor U5005 (N_5005,N_4960,N_4854);
nor U5006 (N_5006,N_4799,N_4876);
or U5007 (N_5007,N_4886,N_4862);
or U5008 (N_5008,N_4989,N_4828);
xnor U5009 (N_5009,N_4815,N_4856);
nor U5010 (N_5010,N_4996,N_4895);
and U5011 (N_5011,N_4773,N_4827);
or U5012 (N_5012,N_4811,N_4927);
nor U5013 (N_5013,N_4978,N_4820);
nor U5014 (N_5014,N_4931,N_4756);
xnor U5015 (N_5015,N_4921,N_4997);
and U5016 (N_5016,N_4831,N_4963);
xnor U5017 (N_5017,N_4757,N_4884);
nand U5018 (N_5018,N_4900,N_4910);
or U5019 (N_5019,N_4936,N_4958);
and U5020 (N_5020,N_4941,N_4792);
and U5021 (N_5021,N_4979,N_4986);
nand U5022 (N_5022,N_4806,N_4925);
nor U5023 (N_5023,N_4801,N_4949);
xor U5024 (N_5024,N_4964,N_4858);
nor U5025 (N_5025,N_4967,N_4852);
and U5026 (N_5026,N_4980,N_4882);
nor U5027 (N_5027,N_4912,N_4945);
xnor U5028 (N_5028,N_4883,N_4871);
or U5029 (N_5029,N_4789,N_4798);
xor U5030 (N_5030,N_4847,N_4846);
or U5031 (N_5031,N_4843,N_4771);
xor U5032 (N_5032,N_4870,N_4962);
nand U5033 (N_5033,N_4873,N_4922);
and U5034 (N_5034,N_4944,N_4926);
nand U5035 (N_5035,N_4840,N_4754);
nand U5036 (N_5036,N_4794,N_4923);
nor U5037 (N_5037,N_4928,N_4954);
nor U5038 (N_5038,N_4763,N_4890);
or U5039 (N_5039,N_4988,N_4867);
and U5040 (N_5040,N_4764,N_4803);
nor U5041 (N_5041,N_4902,N_4888);
nand U5042 (N_5042,N_4943,N_4880);
and U5043 (N_5043,N_4836,N_4913);
nand U5044 (N_5044,N_4950,N_4968);
nand U5045 (N_5045,N_4819,N_4752);
xnor U5046 (N_5046,N_4791,N_4977);
and U5047 (N_5047,N_4875,N_4999);
and U5048 (N_5048,N_4804,N_4774);
and U5049 (N_5049,N_4783,N_4842);
or U5050 (N_5050,N_4879,N_4830);
or U5051 (N_5051,N_4932,N_4861);
and U5052 (N_5052,N_4955,N_4829);
or U5053 (N_5053,N_4930,N_4768);
nor U5054 (N_5054,N_4959,N_4957);
xor U5055 (N_5055,N_4758,N_4812);
or U5056 (N_5056,N_4788,N_4837);
or U5057 (N_5057,N_4821,N_4981);
and U5058 (N_5058,N_4841,N_4918);
nand U5059 (N_5059,N_4907,N_4793);
nor U5060 (N_5060,N_4809,N_4975);
and U5061 (N_5061,N_4807,N_4782);
nand U5062 (N_5062,N_4753,N_4851);
xnor U5063 (N_5063,N_4786,N_4937);
or U5064 (N_5064,N_4951,N_4859);
nand U5065 (N_5065,N_4965,N_4755);
nand U5066 (N_5066,N_4776,N_4972);
and U5067 (N_5067,N_4935,N_4770);
nor U5068 (N_5068,N_4984,N_4919);
or U5069 (N_5069,N_4761,N_4853);
or U5070 (N_5070,N_4929,N_4952);
nor U5071 (N_5071,N_4874,N_4866);
and U5072 (N_5072,N_4973,N_4780);
or U5073 (N_5073,N_4933,N_4868);
nand U5074 (N_5074,N_4924,N_4849);
nand U5075 (N_5075,N_4982,N_4947);
and U5076 (N_5076,N_4992,N_4891);
nor U5077 (N_5077,N_4825,N_4816);
and U5078 (N_5078,N_4760,N_4908);
or U5079 (N_5079,N_4946,N_4869);
or U5080 (N_5080,N_4860,N_4775);
xnor U5081 (N_5081,N_4857,N_4762);
nor U5082 (N_5082,N_4814,N_4904);
xor U5083 (N_5083,N_4994,N_4844);
nor U5084 (N_5084,N_4795,N_4845);
nand U5085 (N_5085,N_4892,N_4961);
or U5086 (N_5086,N_4787,N_4833);
nand U5087 (N_5087,N_4934,N_4878);
xor U5088 (N_5088,N_4948,N_4805);
nor U5089 (N_5089,N_4766,N_4839);
or U5090 (N_5090,N_4916,N_4767);
xnor U5091 (N_5091,N_4864,N_4897);
nor U5092 (N_5092,N_4779,N_4881);
xor U5093 (N_5093,N_4769,N_4993);
or U5094 (N_5094,N_4810,N_4808);
xor U5095 (N_5095,N_4985,N_4911);
nand U5096 (N_5096,N_4966,N_4887);
nand U5097 (N_5097,N_4990,N_4872);
nand U5098 (N_5098,N_4906,N_4898);
xor U5099 (N_5099,N_4995,N_4956);
xnor U5100 (N_5100,N_4751,N_4823);
nor U5101 (N_5101,N_4991,N_4765);
and U5102 (N_5102,N_4802,N_4778);
xor U5103 (N_5103,N_4822,N_4974);
nand U5104 (N_5104,N_4903,N_4750);
xnor U5105 (N_5105,N_4971,N_4983);
and U5106 (N_5106,N_4835,N_4800);
nand U5107 (N_5107,N_4938,N_4940);
nor U5108 (N_5108,N_4796,N_4969);
and U5109 (N_5109,N_4953,N_4797);
nor U5110 (N_5110,N_4901,N_4909);
and U5111 (N_5111,N_4942,N_4784);
nor U5112 (N_5112,N_4813,N_4855);
xnor U5113 (N_5113,N_4863,N_4905);
and U5114 (N_5114,N_4915,N_4824);
and U5115 (N_5115,N_4865,N_4889);
and U5116 (N_5116,N_4848,N_4832);
nand U5117 (N_5117,N_4920,N_4759);
or U5118 (N_5118,N_4893,N_4998);
or U5119 (N_5119,N_4914,N_4970);
or U5120 (N_5120,N_4834,N_4781);
nand U5121 (N_5121,N_4917,N_4976);
or U5122 (N_5122,N_4987,N_4939);
or U5123 (N_5123,N_4896,N_4826);
nand U5124 (N_5124,N_4817,N_4777);
nor U5125 (N_5125,N_4795,N_4957);
xnor U5126 (N_5126,N_4966,N_4856);
nor U5127 (N_5127,N_4887,N_4987);
xnor U5128 (N_5128,N_4823,N_4969);
xnor U5129 (N_5129,N_4884,N_4980);
and U5130 (N_5130,N_4862,N_4995);
and U5131 (N_5131,N_4996,N_4838);
or U5132 (N_5132,N_4954,N_4793);
or U5133 (N_5133,N_4936,N_4817);
nor U5134 (N_5134,N_4889,N_4821);
and U5135 (N_5135,N_4953,N_4901);
nand U5136 (N_5136,N_4878,N_4810);
xnor U5137 (N_5137,N_4862,N_4892);
xnor U5138 (N_5138,N_4791,N_4858);
nor U5139 (N_5139,N_4977,N_4811);
or U5140 (N_5140,N_4833,N_4774);
nand U5141 (N_5141,N_4989,N_4819);
xnor U5142 (N_5142,N_4867,N_4767);
xnor U5143 (N_5143,N_4814,N_4872);
xnor U5144 (N_5144,N_4826,N_4907);
or U5145 (N_5145,N_4806,N_4980);
or U5146 (N_5146,N_4844,N_4974);
nor U5147 (N_5147,N_4949,N_4863);
and U5148 (N_5148,N_4867,N_4797);
xor U5149 (N_5149,N_4946,N_4860);
or U5150 (N_5150,N_4767,N_4880);
and U5151 (N_5151,N_4954,N_4803);
or U5152 (N_5152,N_4843,N_4896);
nor U5153 (N_5153,N_4810,N_4817);
and U5154 (N_5154,N_4823,N_4973);
or U5155 (N_5155,N_4979,N_4881);
xor U5156 (N_5156,N_4772,N_4880);
or U5157 (N_5157,N_4833,N_4981);
nand U5158 (N_5158,N_4794,N_4797);
nor U5159 (N_5159,N_4906,N_4850);
nor U5160 (N_5160,N_4763,N_4797);
and U5161 (N_5161,N_4911,N_4777);
and U5162 (N_5162,N_4935,N_4753);
xnor U5163 (N_5163,N_4792,N_4942);
xnor U5164 (N_5164,N_4892,N_4925);
or U5165 (N_5165,N_4977,N_4959);
or U5166 (N_5166,N_4914,N_4780);
xnor U5167 (N_5167,N_4875,N_4993);
xnor U5168 (N_5168,N_4847,N_4900);
nor U5169 (N_5169,N_4927,N_4926);
xor U5170 (N_5170,N_4752,N_4972);
nand U5171 (N_5171,N_4909,N_4893);
and U5172 (N_5172,N_4806,N_4763);
nand U5173 (N_5173,N_4847,N_4875);
nand U5174 (N_5174,N_4806,N_4829);
or U5175 (N_5175,N_4750,N_4980);
or U5176 (N_5176,N_4839,N_4985);
or U5177 (N_5177,N_4964,N_4932);
or U5178 (N_5178,N_4831,N_4756);
nand U5179 (N_5179,N_4830,N_4798);
nand U5180 (N_5180,N_4839,N_4765);
or U5181 (N_5181,N_4811,N_4784);
nand U5182 (N_5182,N_4927,N_4838);
nand U5183 (N_5183,N_4773,N_4938);
and U5184 (N_5184,N_4786,N_4983);
xnor U5185 (N_5185,N_4958,N_4974);
xnor U5186 (N_5186,N_4814,N_4941);
xnor U5187 (N_5187,N_4872,N_4798);
nor U5188 (N_5188,N_4911,N_4901);
nand U5189 (N_5189,N_4893,N_4835);
xor U5190 (N_5190,N_4762,N_4893);
xor U5191 (N_5191,N_4831,N_4931);
nand U5192 (N_5192,N_4980,N_4755);
xnor U5193 (N_5193,N_4912,N_4755);
and U5194 (N_5194,N_4882,N_4912);
nand U5195 (N_5195,N_4834,N_4979);
or U5196 (N_5196,N_4966,N_4984);
and U5197 (N_5197,N_4767,N_4884);
xor U5198 (N_5198,N_4889,N_4837);
or U5199 (N_5199,N_4995,N_4993);
or U5200 (N_5200,N_4754,N_4907);
and U5201 (N_5201,N_4992,N_4988);
xor U5202 (N_5202,N_4915,N_4954);
or U5203 (N_5203,N_4827,N_4801);
xor U5204 (N_5204,N_4953,N_4952);
and U5205 (N_5205,N_4759,N_4841);
xnor U5206 (N_5206,N_4778,N_4962);
and U5207 (N_5207,N_4947,N_4954);
and U5208 (N_5208,N_4824,N_4829);
nor U5209 (N_5209,N_4918,N_4771);
and U5210 (N_5210,N_4790,N_4988);
xnor U5211 (N_5211,N_4902,N_4977);
and U5212 (N_5212,N_4862,N_4911);
or U5213 (N_5213,N_4762,N_4856);
and U5214 (N_5214,N_4944,N_4870);
xnor U5215 (N_5215,N_4825,N_4991);
nor U5216 (N_5216,N_4783,N_4923);
nor U5217 (N_5217,N_4902,N_4838);
and U5218 (N_5218,N_4964,N_4924);
xnor U5219 (N_5219,N_4802,N_4971);
or U5220 (N_5220,N_4754,N_4908);
xor U5221 (N_5221,N_4888,N_4996);
nor U5222 (N_5222,N_4840,N_4947);
nand U5223 (N_5223,N_4990,N_4950);
and U5224 (N_5224,N_4946,N_4780);
xnor U5225 (N_5225,N_4947,N_4981);
and U5226 (N_5226,N_4938,N_4914);
xnor U5227 (N_5227,N_4838,N_4986);
xor U5228 (N_5228,N_4889,N_4973);
nor U5229 (N_5229,N_4806,N_4996);
nand U5230 (N_5230,N_4878,N_4969);
xor U5231 (N_5231,N_4785,N_4935);
nor U5232 (N_5232,N_4770,N_4903);
or U5233 (N_5233,N_4866,N_4850);
nand U5234 (N_5234,N_4825,N_4797);
xor U5235 (N_5235,N_4843,N_4827);
and U5236 (N_5236,N_4911,N_4856);
xor U5237 (N_5237,N_4895,N_4839);
and U5238 (N_5238,N_4896,N_4753);
xnor U5239 (N_5239,N_4942,N_4905);
or U5240 (N_5240,N_4949,N_4939);
or U5241 (N_5241,N_4758,N_4981);
and U5242 (N_5242,N_4801,N_4769);
nor U5243 (N_5243,N_4939,N_4848);
nor U5244 (N_5244,N_4866,N_4793);
xnor U5245 (N_5245,N_4955,N_4925);
nand U5246 (N_5246,N_4814,N_4838);
and U5247 (N_5247,N_4871,N_4890);
nand U5248 (N_5248,N_4859,N_4920);
or U5249 (N_5249,N_4805,N_4826);
xor U5250 (N_5250,N_5164,N_5186);
xnor U5251 (N_5251,N_5205,N_5121);
nand U5252 (N_5252,N_5128,N_5022);
xnor U5253 (N_5253,N_5013,N_5061);
nor U5254 (N_5254,N_5188,N_5001);
or U5255 (N_5255,N_5249,N_5191);
and U5256 (N_5256,N_5209,N_5005);
nand U5257 (N_5257,N_5032,N_5217);
nor U5258 (N_5258,N_5154,N_5090);
and U5259 (N_5259,N_5099,N_5212);
xnor U5260 (N_5260,N_5236,N_5073);
nand U5261 (N_5261,N_5101,N_5181);
and U5262 (N_5262,N_5214,N_5148);
xor U5263 (N_5263,N_5177,N_5114);
nand U5264 (N_5264,N_5056,N_5016);
nand U5265 (N_5265,N_5126,N_5058);
nand U5266 (N_5266,N_5033,N_5132);
and U5267 (N_5267,N_5144,N_5149);
nor U5268 (N_5268,N_5194,N_5244);
nor U5269 (N_5269,N_5012,N_5136);
nor U5270 (N_5270,N_5167,N_5196);
and U5271 (N_5271,N_5072,N_5047);
nor U5272 (N_5272,N_5108,N_5075);
and U5273 (N_5273,N_5054,N_5003);
nor U5274 (N_5274,N_5153,N_5037);
and U5275 (N_5275,N_5215,N_5112);
nand U5276 (N_5276,N_5046,N_5239);
or U5277 (N_5277,N_5100,N_5222);
xor U5278 (N_5278,N_5208,N_5009);
or U5279 (N_5279,N_5116,N_5086);
and U5280 (N_5280,N_5179,N_5227);
xnor U5281 (N_5281,N_5130,N_5050);
or U5282 (N_5282,N_5057,N_5125);
or U5283 (N_5283,N_5064,N_5048);
or U5284 (N_5284,N_5074,N_5183);
or U5285 (N_5285,N_5105,N_5135);
xnor U5286 (N_5286,N_5229,N_5141);
and U5287 (N_5287,N_5044,N_5143);
or U5288 (N_5288,N_5137,N_5223);
xor U5289 (N_5289,N_5080,N_5202);
nand U5290 (N_5290,N_5083,N_5010);
and U5291 (N_5291,N_5241,N_5119);
or U5292 (N_5292,N_5192,N_5020);
and U5293 (N_5293,N_5242,N_5038);
xnor U5294 (N_5294,N_5059,N_5028);
and U5295 (N_5295,N_5138,N_5157);
or U5296 (N_5296,N_5200,N_5007);
and U5297 (N_5297,N_5066,N_5160);
nand U5298 (N_5298,N_5049,N_5139);
xor U5299 (N_5299,N_5173,N_5067);
nand U5300 (N_5300,N_5078,N_5129);
xnor U5301 (N_5301,N_5146,N_5127);
or U5302 (N_5302,N_5107,N_5204);
nor U5303 (N_5303,N_5238,N_5095);
xor U5304 (N_5304,N_5004,N_5026);
or U5305 (N_5305,N_5069,N_5220);
or U5306 (N_5306,N_5002,N_5079);
nor U5307 (N_5307,N_5062,N_5060);
or U5308 (N_5308,N_5023,N_5096);
and U5309 (N_5309,N_5187,N_5133);
xor U5310 (N_5310,N_5140,N_5025);
xor U5311 (N_5311,N_5030,N_5093);
or U5312 (N_5312,N_5055,N_5159);
nor U5313 (N_5313,N_5034,N_5199);
and U5314 (N_5314,N_5039,N_5195);
nor U5315 (N_5315,N_5006,N_5162);
xnor U5316 (N_5316,N_5156,N_5243);
nand U5317 (N_5317,N_5169,N_5185);
nand U5318 (N_5318,N_5092,N_5225);
or U5319 (N_5319,N_5221,N_5216);
nand U5320 (N_5320,N_5098,N_5068);
or U5321 (N_5321,N_5245,N_5029);
nor U5322 (N_5322,N_5088,N_5234);
and U5323 (N_5323,N_5158,N_5247);
or U5324 (N_5324,N_5166,N_5071);
or U5325 (N_5325,N_5015,N_5031);
nand U5326 (N_5326,N_5197,N_5176);
xor U5327 (N_5327,N_5065,N_5134);
xnor U5328 (N_5328,N_5000,N_5226);
and U5329 (N_5329,N_5237,N_5165);
xnor U5330 (N_5330,N_5168,N_5207);
nor U5331 (N_5331,N_5218,N_5152);
nor U5332 (N_5332,N_5109,N_5171);
nand U5333 (N_5333,N_5102,N_5018);
or U5334 (N_5334,N_5211,N_5027);
nor U5335 (N_5335,N_5070,N_5063);
xnor U5336 (N_5336,N_5190,N_5201);
and U5337 (N_5337,N_5122,N_5240);
xor U5338 (N_5338,N_5189,N_5228);
and U5339 (N_5339,N_5089,N_5097);
nand U5340 (N_5340,N_5087,N_5091);
nand U5341 (N_5341,N_5131,N_5142);
and U5342 (N_5342,N_5219,N_5120);
nand U5343 (N_5343,N_5051,N_5117);
nor U5344 (N_5344,N_5076,N_5017);
nor U5345 (N_5345,N_5113,N_5145);
nor U5346 (N_5346,N_5150,N_5115);
nand U5347 (N_5347,N_5172,N_5045);
and U5348 (N_5348,N_5206,N_5008);
and U5349 (N_5349,N_5184,N_5110);
xor U5350 (N_5350,N_5042,N_5021);
and U5351 (N_5351,N_5235,N_5011);
xor U5352 (N_5352,N_5036,N_5224);
nor U5353 (N_5353,N_5155,N_5085);
xnor U5354 (N_5354,N_5111,N_5182);
xnor U5355 (N_5355,N_5233,N_5246);
or U5356 (N_5356,N_5104,N_5178);
or U5357 (N_5357,N_5231,N_5248);
nand U5358 (N_5358,N_5193,N_5147);
or U5359 (N_5359,N_5180,N_5014);
nor U5360 (N_5360,N_5203,N_5213);
or U5361 (N_5361,N_5163,N_5118);
nor U5362 (N_5362,N_5103,N_5040);
xnor U5363 (N_5363,N_5024,N_5094);
xor U5364 (N_5364,N_5124,N_5174);
nand U5365 (N_5365,N_5151,N_5052);
or U5366 (N_5366,N_5106,N_5053);
xor U5367 (N_5367,N_5035,N_5082);
nand U5368 (N_5368,N_5043,N_5084);
xnor U5369 (N_5369,N_5123,N_5161);
or U5370 (N_5370,N_5232,N_5198);
nand U5371 (N_5371,N_5175,N_5210);
or U5372 (N_5372,N_5170,N_5230);
nor U5373 (N_5373,N_5081,N_5041);
xor U5374 (N_5374,N_5077,N_5019);
nor U5375 (N_5375,N_5004,N_5043);
nor U5376 (N_5376,N_5118,N_5015);
nand U5377 (N_5377,N_5190,N_5199);
nand U5378 (N_5378,N_5136,N_5089);
and U5379 (N_5379,N_5014,N_5081);
xnor U5380 (N_5380,N_5242,N_5107);
nor U5381 (N_5381,N_5095,N_5240);
xnor U5382 (N_5382,N_5102,N_5055);
nand U5383 (N_5383,N_5086,N_5066);
and U5384 (N_5384,N_5102,N_5075);
nor U5385 (N_5385,N_5200,N_5182);
nor U5386 (N_5386,N_5207,N_5225);
nand U5387 (N_5387,N_5216,N_5152);
nor U5388 (N_5388,N_5240,N_5068);
and U5389 (N_5389,N_5211,N_5115);
xor U5390 (N_5390,N_5175,N_5230);
xnor U5391 (N_5391,N_5154,N_5077);
or U5392 (N_5392,N_5051,N_5155);
xnor U5393 (N_5393,N_5216,N_5157);
nand U5394 (N_5394,N_5053,N_5229);
xnor U5395 (N_5395,N_5120,N_5034);
nand U5396 (N_5396,N_5093,N_5071);
nor U5397 (N_5397,N_5143,N_5014);
nand U5398 (N_5398,N_5230,N_5065);
xnor U5399 (N_5399,N_5228,N_5076);
nor U5400 (N_5400,N_5245,N_5068);
and U5401 (N_5401,N_5184,N_5071);
and U5402 (N_5402,N_5105,N_5106);
or U5403 (N_5403,N_5057,N_5095);
nand U5404 (N_5404,N_5146,N_5192);
and U5405 (N_5405,N_5085,N_5201);
nand U5406 (N_5406,N_5090,N_5047);
xor U5407 (N_5407,N_5228,N_5065);
xnor U5408 (N_5408,N_5249,N_5147);
nand U5409 (N_5409,N_5087,N_5153);
nand U5410 (N_5410,N_5062,N_5004);
nand U5411 (N_5411,N_5237,N_5188);
xnor U5412 (N_5412,N_5199,N_5054);
and U5413 (N_5413,N_5080,N_5239);
or U5414 (N_5414,N_5147,N_5113);
nor U5415 (N_5415,N_5177,N_5173);
or U5416 (N_5416,N_5025,N_5036);
or U5417 (N_5417,N_5076,N_5157);
nand U5418 (N_5418,N_5049,N_5137);
and U5419 (N_5419,N_5159,N_5082);
or U5420 (N_5420,N_5017,N_5203);
nand U5421 (N_5421,N_5012,N_5045);
nand U5422 (N_5422,N_5173,N_5207);
nand U5423 (N_5423,N_5113,N_5239);
or U5424 (N_5424,N_5141,N_5228);
nor U5425 (N_5425,N_5133,N_5216);
or U5426 (N_5426,N_5245,N_5164);
and U5427 (N_5427,N_5206,N_5133);
or U5428 (N_5428,N_5201,N_5042);
and U5429 (N_5429,N_5214,N_5022);
xor U5430 (N_5430,N_5216,N_5180);
xor U5431 (N_5431,N_5111,N_5196);
and U5432 (N_5432,N_5193,N_5241);
and U5433 (N_5433,N_5064,N_5151);
xor U5434 (N_5434,N_5182,N_5164);
xnor U5435 (N_5435,N_5157,N_5217);
nor U5436 (N_5436,N_5133,N_5083);
nand U5437 (N_5437,N_5179,N_5214);
nor U5438 (N_5438,N_5149,N_5100);
nor U5439 (N_5439,N_5179,N_5006);
nor U5440 (N_5440,N_5023,N_5076);
nor U5441 (N_5441,N_5029,N_5004);
nor U5442 (N_5442,N_5244,N_5032);
and U5443 (N_5443,N_5091,N_5037);
nand U5444 (N_5444,N_5062,N_5196);
and U5445 (N_5445,N_5236,N_5132);
and U5446 (N_5446,N_5225,N_5112);
nand U5447 (N_5447,N_5096,N_5065);
xor U5448 (N_5448,N_5205,N_5231);
xor U5449 (N_5449,N_5063,N_5074);
nor U5450 (N_5450,N_5062,N_5219);
nand U5451 (N_5451,N_5201,N_5213);
or U5452 (N_5452,N_5153,N_5088);
xnor U5453 (N_5453,N_5021,N_5124);
nor U5454 (N_5454,N_5140,N_5205);
nand U5455 (N_5455,N_5125,N_5052);
nor U5456 (N_5456,N_5049,N_5116);
nor U5457 (N_5457,N_5103,N_5217);
xor U5458 (N_5458,N_5101,N_5029);
nand U5459 (N_5459,N_5071,N_5212);
or U5460 (N_5460,N_5245,N_5090);
nand U5461 (N_5461,N_5083,N_5039);
nor U5462 (N_5462,N_5143,N_5190);
and U5463 (N_5463,N_5170,N_5161);
or U5464 (N_5464,N_5138,N_5180);
nor U5465 (N_5465,N_5026,N_5089);
nor U5466 (N_5466,N_5015,N_5196);
or U5467 (N_5467,N_5039,N_5079);
and U5468 (N_5468,N_5070,N_5230);
nand U5469 (N_5469,N_5239,N_5249);
nand U5470 (N_5470,N_5019,N_5182);
xnor U5471 (N_5471,N_5143,N_5202);
nor U5472 (N_5472,N_5143,N_5129);
xor U5473 (N_5473,N_5129,N_5049);
nor U5474 (N_5474,N_5057,N_5040);
xor U5475 (N_5475,N_5139,N_5194);
nand U5476 (N_5476,N_5001,N_5217);
and U5477 (N_5477,N_5190,N_5086);
xnor U5478 (N_5478,N_5232,N_5126);
xor U5479 (N_5479,N_5090,N_5084);
nor U5480 (N_5480,N_5199,N_5048);
or U5481 (N_5481,N_5191,N_5012);
nand U5482 (N_5482,N_5099,N_5179);
or U5483 (N_5483,N_5110,N_5100);
or U5484 (N_5484,N_5212,N_5037);
nor U5485 (N_5485,N_5212,N_5220);
or U5486 (N_5486,N_5243,N_5224);
and U5487 (N_5487,N_5088,N_5039);
and U5488 (N_5488,N_5186,N_5224);
or U5489 (N_5489,N_5055,N_5144);
nor U5490 (N_5490,N_5119,N_5038);
nand U5491 (N_5491,N_5033,N_5068);
and U5492 (N_5492,N_5170,N_5054);
or U5493 (N_5493,N_5025,N_5143);
or U5494 (N_5494,N_5050,N_5056);
nor U5495 (N_5495,N_5042,N_5087);
or U5496 (N_5496,N_5078,N_5239);
nand U5497 (N_5497,N_5237,N_5219);
or U5498 (N_5498,N_5246,N_5148);
xor U5499 (N_5499,N_5127,N_5005);
nand U5500 (N_5500,N_5274,N_5323);
nand U5501 (N_5501,N_5410,N_5431);
nand U5502 (N_5502,N_5307,N_5265);
nor U5503 (N_5503,N_5476,N_5260);
or U5504 (N_5504,N_5273,N_5498);
and U5505 (N_5505,N_5312,N_5438);
nor U5506 (N_5506,N_5390,N_5373);
nand U5507 (N_5507,N_5456,N_5442);
xnor U5508 (N_5508,N_5435,N_5464);
and U5509 (N_5509,N_5400,N_5282);
xor U5510 (N_5510,N_5360,N_5475);
or U5511 (N_5511,N_5327,N_5259);
xor U5512 (N_5512,N_5301,N_5277);
xor U5513 (N_5513,N_5384,N_5361);
or U5514 (N_5514,N_5430,N_5446);
nor U5515 (N_5515,N_5377,N_5401);
and U5516 (N_5516,N_5492,N_5291);
xor U5517 (N_5517,N_5445,N_5457);
nand U5518 (N_5518,N_5349,N_5402);
xor U5519 (N_5519,N_5350,N_5276);
nor U5520 (N_5520,N_5294,N_5329);
or U5521 (N_5521,N_5394,N_5316);
nand U5522 (N_5522,N_5451,N_5321);
nor U5523 (N_5523,N_5486,N_5279);
xor U5524 (N_5524,N_5280,N_5336);
nor U5525 (N_5525,N_5449,N_5258);
nand U5526 (N_5526,N_5396,N_5302);
and U5527 (N_5527,N_5426,N_5416);
or U5528 (N_5528,N_5345,N_5458);
nand U5529 (N_5529,N_5419,N_5309);
nand U5530 (N_5530,N_5412,N_5285);
nand U5531 (N_5531,N_5303,N_5363);
or U5532 (N_5532,N_5351,N_5403);
nor U5533 (N_5533,N_5368,N_5364);
and U5534 (N_5534,N_5346,N_5432);
nand U5535 (N_5535,N_5481,N_5489);
nand U5536 (N_5536,N_5487,N_5341);
nand U5537 (N_5537,N_5315,N_5469);
or U5538 (N_5538,N_5310,N_5452);
xnor U5539 (N_5539,N_5287,N_5304);
and U5540 (N_5540,N_5472,N_5497);
nand U5541 (N_5541,N_5459,N_5494);
nor U5542 (N_5542,N_5496,N_5284);
nand U5543 (N_5543,N_5328,N_5275);
or U5544 (N_5544,N_5293,N_5369);
and U5545 (N_5545,N_5439,N_5420);
and U5546 (N_5546,N_5331,N_5334);
and U5547 (N_5547,N_5257,N_5447);
nor U5548 (N_5548,N_5450,N_5256);
or U5549 (N_5549,N_5366,N_5385);
xnor U5550 (N_5550,N_5437,N_5371);
nand U5551 (N_5551,N_5397,N_5393);
xnor U5552 (N_5552,N_5281,N_5297);
nor U5553 (N_5553,N_5320,N_5478);
and U5554 (N_5554,N_5295,N_5250);
nand U5555 (N_5555,N_5324,N_5343);
nand U5556 (N_5556,N_5424,N_5264);
nor U5557 (N_5557,N_5415,N_5335);
nor U5558 (N_5558,N_5380,N_5375);
xor U5559 (N_5559,N_5367,N_5399);
and U5560 (N_5560,N_5465,N_5460);
nand U5561 (N_5561,N_5300,N_5339);
xor U5562 (N_5562,N_5383,N_5386);
nor U5563 (N_5563,N_5255,N_5443);
nor U5564 (N_5564,N_5296,N_5357);
xnor U5565 (N_5565,N_5395,N_5358);
nand U5566 (N_5566,N_5330,N_5425);
nand U5567 (N_5567,N_5466,N_5359);
nand U5568 (N_5568,N_5499,N_5338);
and U5569 (N_5569,N_5421,N_5267);
xor U5570 (N_5570,N_5290,N_5470);
xor U5571 (N_5571,N_5408,N_5326);
or U5572 (N_5572,N_5271,N_5354);
nand U5573 (N_5573,N_5461,N_5379);
nand U5574 (N_5574,N_5305,N_5352);
or U5575 (N_5575,N_5333,N_5391);
nand U5576 (N_5576,N_5266,N_5306);
or U5577 (N_5577,N_5283,N_5453);
xor U5578 (N_5578,N_5422,N_5436);
nand U5579 (N_5579,N_5491,N_5387);
and U5580 (N_5580,N_5471,N_5268);
and U5581 (N_5581,N_5405,N_5298);
or U5582 (N_5582,N_5253,N_5289);
nand U5583 (N_5583,N_5370,N_5314);
and U5584 (N_5584,N_5374,N_5355);
xnor U5585 (N_5585,N_5313,N_5372);
nand U5586 (N_5586,N_5428,N_5454);
xnor U5587 (N_5587,N_5474,N_5477);
xor U5588 (N_5588,N_5440,N_5462);
and U5589 (N_5589,N_5490,N_5406);
nor U5590 (N_5590,N_5407,N_5473);
nor U5591 (N_5591,N_5311,N_5365);
nor U5592 (N_5592,N_5493,N_5463);
and U5593 (N_5593,N_5272,N_5299);
or U5594 (N_5594,N_5417,N_5348);
and U5595 (N_5595,N_5353,N_5318);
xnor U5596 (N_5596,N_5468,N_5411);
nand U5597 (N_5597,N_5434,N_5429);
nand U5598 (N_5598,N_5392,N_5262);
or U5599 (N_5599,N_5444,N_5278);
or U5600 (N_5600,N_5332,N_5378);
and U5601 (N_5601,N_5484,N_5482);
nor U5602 (N_5602,N_5376,N_5347);
and U5603 (N_5603,N_5288,N_5261);
or U5604 (N_5604,N_5423,N_5441);
and U5605 (N_5605,N_5388,N_5413);
nand U5606 (N_5606,N_5344,N_5398);
nor U5607 (N_5607,N_5337,N_5254);
nor U5608 (N_5608,N_5252,N_5263);
and U5609 (N_5609,N_5381,N_5418);
xor U5610 (N_5610,N_5427,N_5270);
xnor U5611 (N_5611,N_5389,N_5404);
nor U5612 (N_5612,N_5483,N_5409);
or U5613 (N_5613,N_5356,N_5342);
xor U5614 (N_5614,N_5362,N_5455);
and U5615 (N_5615,N_5286,N_5308);
xnor U5616 (N_5616,N_5319,N_5251);
and U5617 (N_5617,N_5495,N_5467);
and U5618 (N_5618,N_5414,N_5479);
nor U5619 (N_5619,N_5480,N_5485);
nor U5620 (N_5620,N_5269,N_5317);
xor U5621 (N_5621,N_5322,N_5292);
and U5622 (N_5622,N_5325,N_5448);
or U5623 (N_5623,N_5340,N_5382);
nor U5624 (N_5624,N_5488,N_5433);
or U5625 (N_5625,N_5331,N_5298);
and U5626 (N_5626,N_5338,N_5280);
xnor U5627 (N_5627,N_5254,N_5432);
and U5628 (N_5628,N_5360,N_5321);
xor U5629 (N_5629,N_5276,N_5481);
xnor U5630 (N_5630,N_5443,N_5417);
or U5631 (N_5631,N_5286,N_5356);
nor U5632 (N_5632,N_5398,N_5365);
and U5633 (N_5633,N_5257,N_5305);
nand U5634 (N_5634,N_5311,N_5326);
nor U5635 (N_5635,N_5294,N_5381);
and U5636 (N_5636,N_5355,N_5321);
xnor U5637 (N_5637,N_5299,N_5437);
and U5638 (N_5638,N_5404,N_5463);
nand U5639 (N_5639,N_5263,N_5343);
xor U5640 (N_5640,N_5319,N_5312);
or U5641 (N_5641,N_5458,N_5414);
nor U5642 (N_5642,N_5484,N_5336);
xor U5643 (N_5643,N_5453,N_5472);
or U5644 (N_5644,N_5349,N_5293);
nor U5645 (N_5645,N_5397,N_5308);
nor U5646 (N_5646,N_5445,N_5395);
nand U5647 (N_5647,N_5391,N_5285);
and U5648 (N_5648,N_5291,N_5331);
or U5649 (N_5649,N_5421,N_5499);
and U5650 (N_5650,N_5350,N_5423);
and U5651 (N_5651,N_5286,N_5447);
or U5652 (N_5652,N_5402,N_5317);
xor U5653 (N_5653,N_5343,N_5327);
and U5654 (N_5654,N_5304,N_5325);
nand U5655 (N_5655,N_5377,N_5360);
nor U5656 (N_5656,N_5285,N_5254);
and U5657 (N_5657,N_5381,N_5254);
and U5658 (N_5658,N_5364,N_5333);
and U5659 (N_5659,N_5263,N_5382);
and U5660 (N_5660,N_5273,N_5395);
xnor U5661 (N_5661,N_5370,N_5293);
xor U5662 (N_5662,N_5498,N_5319);
nor U5663 (N_5663,N_5357,N_5454);
nor U5664 (N_5664,N_5446,N_5286);
and U5665 (N_5665,N_5288,N_5458);
or U5666 (N_5666,N_5414,N_5422);
nand U5667 (N_5667,N_5414,N_5336);
or U5668 (N_5668,N_5368,N_5309);
nor U5669 (N_5669,N_5349,N_5280);
nand U5670 (N_5670,N_5459,N_5376);
xnor U5671 (N_5671,N_5382,N_5252);
nor U5672 (N_5672,N_5374,N_5434);
nor U5673 (N_5673,N_5322,N_5400);
xnor U5674 (N_5674,N_5389,N_5280);
xnor U5675 (N_5675,N_5328,N_5407);
and U5676 (N_5676,N_5456,N_5377);
nand U5677 (N_5677,N_5487,N_5291);
nor U5678 (N_5678,N_5311,N_5288);
xor U5679 (N_5679,N_5411,N_5420);
or U5680 (N_5680,N_5267,N_5256);
xor U5681 (N_5681,N_5417,N_5369);
nor U5682 (N_5682,N_5282,N_5374);
and U5683 (N_5683,N_5391,N_5432);
nand U5684 (N_5684,N_5461,N_5405);
xor U5685 (N_5685,N_5401,N_5250);
or U5686 (N_5686,N_5280,N_5333);
or U5687 (N_5687,N_5441,N_5417);
and U5688 (N_5688,N_5483,N_5374);
or U5689 (N_5689,N_5336,N_5349);
nor U5690 (N_5690,N_5256,N_5446);
or U5691 (N_5691,N_5319,N_5310);
nand U5692 (N_5692,N_5298,N_5296);
xor U5693 (N_5693,N_5321,N_5304);
nand U5694 (N_5694,N_5320,N_5369);
and U5695 (N_5695,N_5292,N_5414);
nor U5696 (N_5696,N_5291,N_5429);
or U5697 (N_5697,N_5431,N_5479);
nor U5698 (N_5698,N_5409,N_5428);
nor U5699 (N_5699,N_5388,N_5337);
nor U5700 (N_5700,N_5417,N_5427);
xnor U5701 (N_5701,N_5451,N_5482);
nor U5702 (N_5702,N_5360,N_5432);
xnor U5703 (N_5703,N_5357,N_5369);
nand U5704 (N_5704,N_5268,N_5333);
nand U5705 (N_5705,N_5493,N_5423);
nor U5706 (N_5706,N_5483,N_5381);
xor U5707 (N_5707,N_5347,N_5281);
nand U5708 (N_5708,N_5481,N_5311);
nor U5709 (N_5709,N_5493,N_5271);
nand U5710 (N_5710,N_5378,N_5499);
and U5711 (N_5711,N_5471,N_5357);
and U5712 (N_5712,N_5483,N_5420);
xnor U5713 (N_5713,N_5419,N_5446);
xnor U5714 (N_5714,N_5257,N_5345);
nand U5715 (N_5715,N_5297,N_5383);
nand U5716 (N_5716,N_5385,N_5460);
and U5717 (N_5717,N_5363,N_5479);
and U5718 (N_5718,N_5442,N_5368);
nor U5719 (N_5719,N_5358,N_5270);
xor U5720 (N_5720,N_5311,N_5468);
nor U5721 (N_5721,N_5384,N_5463);
nand U5722 (N_5722,N_5338,N_5441);
nand U5723 (N_5723,N_5256,N_5254);
xor U5724 (N_5724,N_5408,N_5271);
and U5725 (N_5725,N_5406,N_5400);
or U5726 (N_5726,N_5383,N_5315);
nor U5727 (N_5727,N_5453,N_5321);
and U5728 (N_5728,N_5309,N_5496);
nand U5729 (N_5729,N_5307,N_5432);
nor U5730 (N_5730,N_5313,N_5479);
or U5731 (N_5731,N_5250,N_5302);
nor U5732 (N_5732,N_5416,N_5322);
nand U5733 (N_5733,N_5460,N_5345);
xnor U5734 (N_5734,N_5400,N_5274);
nor U5735 (N_5735,N_5394,N_5337);
nand U5736 (N_5736,N_5469,N_5268);
nor U5737 (N_5737,N_5320,N_5405);
or U5738 (N_5738,N_5312,N_5265);
nand U5739 (N_5739,N_5257,N_5359);
nand U5740 (N_5740,N_5257,N_5456);
or U5741 (N_5741,N_5255,N_5420);
or U5742 (N_5742,N_5261,N_5253);
and U5743 (N_5743,N_5279,N_5306);
nor U5744 (N_5744,N_5334,N_5381);
and U5745 (N_5745,N_5282,N_5328);
and U5746 (N_5746,N_5409,N_5455);
nor U5747 (N_5747,N_5477,N_5478);
xor U5748 (N_5748,N_5390,N_5464);
nor U5749 (N_5749,N_5361,N_5430);
nand U5750 (N_5750,N_5718,N_5678);
or U5751 (N_5751,N_5637,N_5578);
or U5752 (N_5752,N_5685,N_5689);
nand U5753 (N_5753,N_5632,N_5663);
and U5754 (N_5754,N_5609,N_5604);
nor U5755 (N_5755,N_5534,N_5684);
and U5756 (N_5756,N_5549,N_5626);
nor U5757 (N_5757,N_5543,N_5621);
nor U5758 (N_5758,N_5680,N_5598);
and U5759 (N_5759,N_5639,N_5638);
or U5760 (N_5760,N_5592,N_5608);
nand U5761 (N_5761,N_5558,N_5739);
and U5762 (N_5762,N_5742,N_5583);
xnor U5763 (N_5763,N_5599,N_5605);
and U5764 (N_5764,N_5597,N_5733);
xor U5765 (N_5765,N_5567,N_5643);
nor U5766 (N_5766,N_5540,N_5631);
or U5767 (N_5767,N_5521,N_5533);
xnor U5768 (N_5768,N_5606,N_5554);
nor U5769 (N_5769,N_5594,N_5587);
nand U5770 (N_5770,N_5525,N_5568);
and U5771 (N_5771,N_5520,N_5664);
nand U5772 (N_5772,N_5641,N_5749);
or U5773 (N_5773,N_5575,N_5528);
nor U5774 (N_5774,N_5555,N_5693);
nor U5775 (N_5775,N_5603,N_5672);
xor U5776 (N_5776,N_5746,N_5618);
xor U5777 (N_5777,N_5705,N_5647);
and U5778 (N_5778,N_5503,N_5610);
xor U5779 (N_5779,N_5624,N_5653);
nor U5780 (N_5780,N_5564,N_5725);
xnor U5781 (N_5781,N_5711,N_5566);
nor U5782 (N_5782,N_5649,N_5539);
nand U5783 (N_5783,N_5629,N_5572);
nand U5784 (N_5784,N_5745,N_5737);
or U5785 (N_5785,N_5524,N_5561);
nor U5786 (N_5786,N_5652,N_5660);
nor U5787 (N_5787,N_5505,N_5508);
or U5788 (N_5788,N_5691,N_5584);
or U5789 (N_5789,N_5613,N_5715);
or U5790 (N_5790,N_5514,N_5612);
nor U5791 (N_5791,N_5547,N_5573);
and U5792 (N_5792,N_5501,N_5602);
and U5793 (N_5793,N_5697,N_5654);
and U5794 (N_5794,N_5551,N_5730);
or U5795 (N_5795,N_5512,N_5601);
and U5796 (N_5796,N_5710,N_5511);
or U5797 (N_5797,N_5617,N_5581);
or U5798 (N_5798,N_5531,N_5698);
nand U5799 (N_5799,N_5513,N_5642);
and U5800 (N_5800,N_5738,N_5545);
nor U5801 (N_5801,N_5559,N_5553);
and U5802 (N_5802,N_5607,N_5735);
and U5803 (N_5803,N_5577,N_5530);
and U5804 (N_5804,N_5668,N_5695);
nor U5805 (N_5805,N_5504,N_5690);
nor U5806 (N_5806,N_5648,N_5667);
nor U5807 (N_5807,N_5728,N_5627);
nand U5808 (N_5808,N_5519,N_5628);
nand U5809 (N_5809,N_5744,N_5517);
nand U5810 (N_5810,N_5717,N_5546);
xor U5811 (N_5811,N_5634,N_5576);
nand U5812 (N_5812,N_5515,N_5523);
nor U5813 (N_5813,N_5719,N_5593);
nand U5814 (N_5814,N_5623,N_5651);
and U5815 (N_5815,N_5633,N_5724);
or U5816 (N_5816,N_5526,N_5707);
and U5817 (N_5817,N_5679,N_5591);
or U5818 (N_5818,N_5644,N_5600);
nor U5819 (N_5819,N_5538,N_5589);
and U5820 (N_5820,N_5692,N_5743);
nand U5821 (N_5821,N_5544,N_5510);
nand U5822 (N_5822,N_5708,N_5736);
nand U5823 (N_5823,N_5506,N_5509);
nand U5824 (N_5824,N_5732,N_5646);
or U5825 (N_5825,N_5703,N_5557);
and U5826 (N_5826,N_5709,N_5579);
nor U5827 (N_5827,N_5671,N_5569);
xor U5828 (N_5828,N_5655,N_5611);
nand U5829 (N_5829,N_5535,N_5681);
or U5830 (N_5830,N_5516,N_5622);
nand U5831 (N_5831,N_5635,N_5748);
nor U5832 (N_5832,N_5688,N_5687);
or U5833 (N_5833,N_5701,N_5726);
xnor U5834 (N_5834,N_5548,N_5676);
nor U5835 (N_5835,N_5675,N_5507);
xnor U5836 (N_5836,N_5723,N_5713);
or U5837 (N_5837,N_5716,N_5500);
nand U5838 (N_5838,N_5630,N_5645);
or U5839 (N_5839,N_5674,N_5590);
nor U5840 (N_5840,N_5574,N_5704);
nor U5841 (N_5841,N_5677,N_5699);
nand U5842 (N_5842,N_5586,N_5683);
nand U5843 (N_5843,N_5616,N_5669);
xnor U5844 (N_5844,N_5502,N_5596);
xnor U5845 (N_5845,N_5585,N_5595);
and U5846 (N_5846,N_5582,N_5556);
or U5847 (N_5847,N_5619,N_5527);
nand U5848 (N_5848,N_5650,N_5706);
nand U5849 (N_5849,N_5560,N_5537);
nor U5850 (N_5850,N_5721,N_5565);
nor U5851 (N_5851,N_5734,N_5666);
nor U5852 (N_5852,N_5747,N_5615);
and U5853 (N_5853,N_5700,N_5536);
and U5854 (N_5854,N_5659,N_5720);
nand U5855 (N_5855,N_5562,N_5532);
xnor U5856 (N_5856,N_5614,N_5673);
nand U5857 (N_5857,N_5731,N_5570);
nor U5858 (N_5858,N_5662,N_5722);
xor U5859 (N_5859,N_5658,N_5712);
and U5860 (N_5860,N_5741,N_5580);
or U5861 (N_5861,N_5661,N_5729);
xor U5862 (N_5862,N_5694,N_5588);
nand U5863 (N_5863,N_5518,N_5550);
nand U5864 (N_5864,N_5522,N_5702);
or U5865 (N_5865,N_5625,N_5542);
xor U5866 (N_5866,N_5541,N_5657);
and U5867 (N_5867,N_5529,N_5682);
and U5868 (N_5868,N_5665,N_5552);
xor U5869 (N_5869,N_5696,N_5714);
nand U5870 (N_5870,N_5656,N_5636);
nand U5871 (N_5871,N_5727,N_5670);
or U5872 (N_5872,N_5571,N_5563);
nor U5873 (N_5873,N_5740,N_5640);
xnor U5874 (N_5874,N_5686,N_5620);
nor U5875 (N_5875,N_5594,N_5578);
nor U5876 (N_5876,N_5542,N_5569);
xor U5877 (N_5877,N_5626,N_5513);
nand U5878 (N_5878,N_5603,N_5585);
and U5879 (N_5879,N_5548,N_5525);
and U5880 (N_5880,N_5566,N_5536);
xnor U5881 (N_5881,N_5677,N_5514);
nor U5882 (N_5882,N_5508,N_5667);
nand U5883 (N_5883,N_5501,N_5592);
nand U5884 (N_5884,N_5734,N_5723);
xnor U5885 (N_5885,N_5609,N_5678);
nor U5886 (N_5886,N_5508,N_5685);
xor U5887 (N_5887,N_5593,N_5638);
xor U5888 (N_5888,N_5659,N_5504);
nand U5889 (N_5889,N_5507,N_5618);
xor U5890 (N_5890,N_5506,N_5738);
or U5891 (N_5891,N_5689,N_5674);
xor U5892 (N_5892,N_5660,N_5566);
or U5893 (N_5893,N_5531,N_5536);
xor U5894 (N_5894,N_5679,N_5523);
nand U5895 (N_5895,N_5720,N_5658);
nor U5896 (N_5896,N_5501,N_5566);
or U5897 (N_5897,N_5682,N_5606);
or U5898 (N_5898,N_5604,N_5623);
nand U5899 (N_5899,N_5624,N_5615);
nor U5900 (N_5900,N_5592,N_5506);
and U5901 (N_5901,N_5664,N_5650);
nor U5902 (N_5902,N_5542,N_5558);
nor U5903 (N_5903,N_5616,N_5688);
and U5904 (N_5904,N_5690,N_5694);
xnor U5905 (N_5905,N_5712,N_5644);
nor U5906 (N_5906,N_5546,N_5510);
or U5907 (N_5907,N_5572,N_5531);
nand U5908 (N_5908,N_5723,N_5698);
xor U5909 (N_5909,N_5646,N_5681);
nor U5910 (N_5910,N_5744,N_5678);
nand U5911 (N_5911,N_5682,N_5660);
or U5912 (N_5912,N_5537,N_5578);
nor U5913 (N_5913,N_5737,N_5546);
xnor U5914 (N_5914,N_5556,N_5694);
nor U5915 (N_5915,N_5722,N_5537);
or U5916 (N_5916,N_5695,N_5593);
or U5917 (N_5917,N_5547,N_5719);
and U5918 (N_5918,N_5548,N_5560);
and U5919 (N_5919,N_5521,N_5514);
xnor U5920 (N_5920,N_5594,N_5732);
nor U5921 (N_5921,N_5571,N_5504);
or U5922 (N_5922,N_5505,N_5606);
nor U5923 (N_5923,N_5737,N_5739);
or U5924 (N_5924,N_5608,N_5713);
nor U5925 (N_5925,N_5715,N_5695);
nand U5926 (N_5926,N_5547,N_5676);
and U5927 (N_5927,N_5597,N_5617);
and U5928 (N_5928,N_5747,N_5631);
nor U5929 (N_5929,N_5536,N_5681);
xor U5930 (N_5930,N_5658,N_5569);
nor U5931 (N_5931,N_5503,N_5533);
xor U5932 (N_5932,N_5668,N_5684);
or U5933 (N_5933,N_5722,N_5518);
or U5934 (N_5934,N_5621,N_5509);
xnor U5935 (N_5935,N_5707,N_5539);
or U5936 (N_5936,N_5561,N_5593);
nand U5937 (N_5937,N_5736,N_5545);
nand U5938 (N_5938,N_5574,N_5735);
nand U5939 (N_5939,N_5739,N_5724);
nor U5940 (N_5940,N_5622,N_5598);
or U5941 (N_5941,N_5566,N_5687);
xnor U5942 (N_5942,N_5603,N_5513);
xor U5943 (N_5943,N_5721,N_5720);
nand U5944 (N_5944,N_5592,N_5582);
xor U5945 (N_5945,N_5686,N_5701);
and U5946 (N_5946,N_5643,N_5665);
xor U5947 (N_5947,N_5619,N_5731);
or U5948 (N_5948,N_5663,N_5615);
nor U5949 (N_5949,N_5643,N_5688);
and U5950 (N_5950,N_5521,N_5653);
or U5951 (N_5951,N_5597,N_5718);
and U5952 (N_5952,N_5574,N_5581);
nand U5953 (N_5953,N_5622,N_5599);
nor U5954 (N_5954,N_5527,N_5608);
nand U5955 (N_5955,N_5652,N_5592);
or U5956 (N_5956,N_5641,N_5549);
nand U5957 (N_5957,N_5620,N_5614);
nor U5958 (N_5958,N_5510,N_5712);
and U5959 (N_5959,N_5592,N_5647);
nor U5960 (N_5960,N_5650,N_5566);
xor U5961 (N_5961,N_5662,N_5736);
or U5962 (N_5962,N_5584,N_5728);
or U5963 (N_5963,N_5531,N_5727);
nand U5964 (N_5964,N_5724,N_5626);
or U5965 (N_5965,N_5577,N_5672);
nor U5966 (N_5966,N_5500,N_5576);
nand U5967 (N_5967,N_5737,N_5637);
xor U5968 (N_5968,N_5571,N_5714);
nor U5969 (N_5969,N_5595,N_5594);
and U5970 (N_5970,N_5562,N_5592);
nor U5971 (N_5971,N_5663,N_5716);
or U5972 (N_5972,N_5539,N_5686);
nor U5973 (N_5973,N_5708,N_5680);
nand U5974 (N_5974,N_5614,N_5652);
nand U5975 (N_5975,N_5721,N_5520);
nor U5976 (N_5976,N_5694,N_5564);
or U5977 (N_5977,N_5521,N_5675);
and U5978 (N_5978,N_5651,N_5598);
or U5979 (N_5979,N_5627,N_5537);
and U5980 (N_5980,N_5719,N_5685);
nor U5981 (N_5981,N_5504,N_5670);
nor U5982 (N_5982,N_5553,N_5745);
or U5983 (N_5983,N_5613,N_5746);
nand U5984 (N_5984,N_5661,N_5627);
xor U5985 (N_5985,N_5534,N_5628);
xor U5986 (N_5986,N_5673,N_5696);
and U5987 (N_5987,N_5583,N_5614);
xnor U5988 (N_5988,N_5502,N_5665);
nor U5989 (N_5989,N_5628,N_5737);
xnor U5990 (N_5990,N_5576,N_5688);
and U5991 (N_5991,N_5549,N_5732);
nand U5992 (N_5992,N_5704,N_5567);
or U5993 (N_5993,N_5510,N_5713);
nor U5994 (N_5994,N_5525,N_5545);
nor U5995 (N_5995,N_5609,N_5530);
xnor U5996 (N_5996,N_5670,N_5577);
nor U5997 (N_5997,N_5739,N_5523);
nand U5998 (N_5998,N_5504,N_5698);
and U5999 (N_5999,N_5560,N_5585);
and U6000 (N_6000,N_5804,N_5785);
or U6001 (N_6001,N_5783,N_5872);
nor U6002 (N_6002,N_5927,N_5854);
nand U6003 (N_6003,N_5974,N_5791);
nor U6004 (N_6004,N_5892,N_5773);
or U6005 (N_6005,N_5751,N_5953);
xor U6006 (N_6006,N_5792,N_5915);
xor U6007 (N_6007,N_5798,N_5830);
and U6008 (N_6008,N_5962,N_5979);
nand U6009 (N_6009,N_5863,N_5985);
nor U6010 (N_6010,N_5754,N_5924);
nor U6011 (N_6011,N_5951,N_5988);
nor U6012 (N_6012,N_5855,N_5813);
or U6013 (N_6013,N_5906,N_5940);
xor U6014 (N_6014,N_5986,N_5797);
nand U6015 (N_6015,N_5905,N_5862);
xor U6016 (N_6016,N_5762,N_5950);
or U6017 (N_6017,N_5822,N_5981);
nand U6018 (N_6018,N_5828,N_5914);
xor U6019 (N_6019,N_5808,N_5760);
and U6020 (N_6020,N_5764,N_5904);
nand U6021 (N_6021,N_5838,N_5810);
nor U6022 (N_6022,N_5834,N_5938);
and U6023 (N_6023,N_5769,N_5923);
and U6024 (N_6024,N_5947,N_5835);
nand U6025 (N_6025,N_5805,N_5993);
nor U6026 (N_6026,N_5917,N_5933);
or U6027 (N_6027,N_5857,N_5870);
and U6028 (N_6028,N_5753,N_5881);
nor U6029 (N_6029,N_5952,N_5864);
xor U6030 (N_6030,N_5861,N_5928);
xnor U6031 (N_6031,N_5941,N_5944);
or U6032 (N_6032,N_5890,N_5829);
nor U6033 (N_6033,N_5989,N_5771);
xor U6034 (N_6034,N_5960,N_5766);
or U6035 (N_6035,N_5982,N_5918);
nor U6036 (N_6036,N_5776,N_5820);
nand U6037 (N_6037,N_5980,N_5803);
nand U6038 (N_6038,N_5759,N_5866);
xor U6039 (N_6039,N_5782,N_5775);
xor U6040 (N_6040,N_5868,N_5873);
nor U6041 (N_6041,N_5883,N_5972);
xnor U6042 (N_6042,N_5877,N_5955);
or U6043 (N_6043,N_5853,N_5837);
xor U6044 (N_6044,N_5945,N_5911);
xor U6045 (N_6045,N_5789,N_5836);
and U6046 (N_6046,N_5875,N_5949);
and U6047 (N_6047,N_5788,N_5990);
nand U6048 (N_6048,N_5765,N_5796);
nor U6049 (N_6049,N_5894,N_5849);
and U6050 (N_6050,N_5846,N_5887);
nor U6051 (N_6051,N_5799,N_5874);
or U6052 (N_6052,N_5984,N_5954);
nor U6053 (N_6053,N_5833,N_5845);
and U6054 (N_6054,N_5856,N_5968);
xor U6055 (N_6055,N_5943,N_5898);
xnor U6056 (N_6056,N_5871,N_5926);
and U6057 (N_6057,N_5876,N_5793);
or U6058 (N_6058,N_5992,N_5889);
nor U6059 (N_6059,N_5959,N_5896);
nor U6060 (N_6060,N_5869,N_5885);
xor U6061 (N_6061,N_5925,N_5816);
or U6062 (N_6062,N_5790,N_5969);
xor U6063 (N_6063,N_5860,N_5922);
nand U6064 (N_6064,N_5910,N_5879);
or U6065 (N_6065,N_5802,N_5995);
nor U6066 (N_6066,N_5916,N_5811);
or U6067 (N_6067,N_5931,N_5821);
or U6068 (N_6068,N_5865,N_5850);
nor U6069 (N_6069,N_5843,N_5975);
nand U6070 (N_6070,N_5919,N_5942);
nand U6071 (N_6071,N_5848,N_5779);
nand U6072 (N_6072,N_5888,N_5971);
nand U6073 (N_6073,N_5761,N_5840);
or U6074 (N_6074,N_5794,N_5755);
or U6075 (N_6075,N_5824,N_5958);
nand U6076 (N_6076,N_5920,N_5978);
xnor U6077 (N_6077,N_5930,N_5756);
nor U6078 (N_6078,N_5763,N_5819);
xnor U6079 (N_6079,N_5806,N_5784);
or U6080 (N_6080,N_5902,N_5977);
or U6081 (N_6081,N_5812,N_5815);
and U6082 (N_6082,N_5913,N_5778);
and U6083 (N_6083,N_5814,N_5961);
or U6084 (N_6084,N_5908,N_5946);
nor U6085 (N_6085,N_5826,N_5770);
nor U6086 (N_6086,N_5809,N_5936);
nor U6087 (N_6087,N_5777,N_5987);
xnor U6088 (N_6088,N_5901,N_5800);
nand U6089 (N_6089,N_5882,N_5963);
nor U6090 (N_6090,N_5893,N_5973);
xor U6091 (N_6091,N_5772,N_5878);
xor U6092 (N_6092,N_5867,N_5891);
or U6093 (N_6093,N_5994,N_5842);
and U6094 (N_6094,N_5965,N_5886);
and U6095 (N_6095,N_5895,N_5847);
nor U6096 (N_6096,N_5932,N_5966);
xor U6097 (N_6097,N_5998,N_5970);
or U6098 (N_6098,N_5851,N_5884);
nand U6099 (N_6099,N_5948,N_5921);
nand U6100 (N_6100,N_5801,N_5858);
xnor U6101 (N_6101,N_5832,N_5823);
or U6102 (N_6102,N_5758,N_5880);
or U6103 (N_6103,N_5956,N_5859);
xor U6104 (N_6104,N_5957,N_5786);
nor U6105 (N_6105,N_5997,N_5752);
nor U6106 (N_6106,N_5817,N_5935);
or U6107 (N_6107,N_5831,N_5912);
nor U6108 (N_6108,N_5991,N_5976);
and U6109 (N_6109,N_5781,N_5768);
nand U6110 (N_6110,N_5996,N_5780);
and U6111 (N_6111,N_5999,N_5839);
or U6112 (N_6112,N_5807,N_5767);
or U6113 (N_6113,N_5841,N_5787);
nor U6114 (N_6114,N_5934,N_5897);
nand U6115 (N_6115,N_5900,N_5852);
or U6116 (N_6116,N_5937,N_5795);
and U6117 (N_6117,N_5909,N_5939);
nor U6118 (N_6118,N_5983,N_5750);
and U6119 (N_6119,N_5899,N_5757);
and U6120 (N_6120,N_5967,N_5774);
nor U6121 (N_6121,N_5907,N_5825);
nand U6122 (N_6122,N_5844,N_5964);
and U6123 (N_6123,N_5818,N_5903);
nor U6124 (N_6124,N_5929,N_5827);
and U6125 (N_6125,N_5933,N_5935);
nor U6126 (N_6126,N_5756,N_5921);
or U6127 (N_6127,N_5948,N_5780);
and U6128 (N_6128,N_5813,N_5810);
and U6129 (N_6129,N_5805,N_5976);
xor U6130 (N_6130,N_5826,N_5780);
and U6131 (N_6131,N_5831,N_5840);
nor U6132 (N_6132,N_5860,N_5783);
nor U6133 (N_6133,N_5795,N_5925);
xnor U6134 (N_6134,N_5831,N_5901);
xnor U6135 (N_6135,N_5997,N_5907);
or U6136 (N_6136,N_5969,N_5956);
nand U6137 (N_6137,N_5801,N_5760);
or U6138 (N_6138,N_5765,N_5953);
nor U6139 (N_6139,N_5875,N_5914);
or U6140 (N_6140,N_5904,N_5951);
and U6141 (N_6141,N_5810,N_5806);
or U6142 (N_6142,N_5923,N_5758);
or U6143 (N_6143,N_5984,N_5903);
nor U6144 (N_6144,N_5890,N_5985);
nand U6145 (N_6145,N_5817,N_5835);
xnor U6146 (N_6146,N_5990,N_5936);
nor U6147 (N_6147,N_5874,N_5809);
nor U6148 (N_6148,N_5964,N_5796);
nand U6149 (N_6149,N_5819,N_5896);
nand U6150 (N_6150,N_5974,N_5848);
nor U6151 (N_6151,N_5824,N_5916);
nand U6152 (N_6152,N_5804,N_5793);
nand U6153 (N_6153,N_5865,N_5963);
xor U6154 (N_6154,N_5868,N_5768);
or U6155 (N_6155,N_5926,N_5852);
nand U6156 (N_6156,N_5851,N_5918);
xor U6157 (N_6157,N_5919,N_5952);
and U6158 (N_6158,N_5785,N_5859);
or U6159 (N_6159,N_5831,N_5769);
or U6160 (N_6160,N_5902,N_5962);
nand U6161 (N_6161,N_5850,N_5806);
nand U6162 (N_6162,N_5878,N_5989);
nor U6163 (N_6163,N_5757,N_5967);
nand U6164 (N_6164,N_5821,N_5783);
xnor U6165 (N_6165,N_5813,N_5894);
nand U6166 (N_6166,N_5868,N_5811);
nor U6167 (N_6167,N_5928,N_5866);
nand U6168 (N_6168,N_5963,N_5935);
or U6169 (N_6169,N_5826,N_5789);
and U6170 (N_6170,N_5766,N_5856);
nand U6171 (N_6171,N_5956,N_5811);
nor U6172 (N_6172,N_5810,N_5837);
nand U6173 (N_6173,N_5861,N_5820);
nor U6174 (N_6174,N_5758,N_5822);
or U6175 (N_6175,N_5929,N_5768);
nand U6176 (N_6176,N_5791,N_5819);
or U6177 (N_6177,N_5960,N_5943);
or U6178 (N_6178,N_5872,N_5875);
nand U6179 (N_6179,N_5912,N_5773);
xor U6180 (N_6180,N_5868,N_5940);
xor U6181 (N_6181,N_5891,N_5838);
and U6182 (N_6182,N_5892,N_5975);
or U6183 (N_6183,N_5855,N_5967);
nand U6184 (N_6184,N_5977,N_5942);
or U6185 (N_6185,N_5820,N_5853);
xor U6186 (N_6186,N_5845,N_5852);
and U6187 (N_6187,N_5824,N_5964);
nor U6188 (N_6188,N_5924,N_5820);
xnor U6189 (N_6189,N_5861,N_5836);
xor U6190 (N_6190,N_5810,N_5882);
or U6191 (N_6191,N_5929,N_5964);
and U6192 (N_6192,N_5850,N_5948);
or U6193 (N_6193,N_5997,N_5821);
nor U6194 (N_6194,N_5869,N_5760);
nor U6195 (N_6195,N_5784,N_5853);
nand U6196 (N_6196,N_5848,N_5989);
and U6197 (N_6197,N_5896,N_5984);
nor U6198 (N_6198,N_5849,N_5886);
nor U6199 (N_6199,N_5864,N_5759);
nand U6200 (N_6200,N_5774,N_5956);
and U6201 (N_6201,N_5762,N_5837);
nor U6202 (N_6202,N_5853,N_5958);
or U6203 (N_6203,N_5778,N_5756);
nand U6204 (N_6204,N_5903,N_5832);
or U6205 (N_6205,N_5903,N_5844);
nor U6206 (N_6206,N_5935,N_5795);
or U6207 (N_6207,N_5919,N_5891);
xnor U6208 (N_6208,N_5949,N_5788);
or U6209 (N_6209,N_5826,N_5876);
or U6210 (N_6210,N_5933,N_5900);
nor U6211 (N_6211,N_5882,N_5996);
and U6212 (N_6212,N_5848,N_5882);
nand U6213 (N_6213,N_5758,N_5766);
xor U6214 (N_6214,N_5953,N_5967);
nand U6215 (N_6215,N_5848,N_5859);
nand U6216 (N_6216,N_5808,N_5819);
nor U6217 (N_6217,N_5932,N_5949);
or U6218 (N_6218,N_5987,N_5791);
or U6219 (N_6219,N_5781,N_5907);
or U6220 (N_6220,N_5852,N_5968);
nor U6221 (N_6221,N_5785,N_5836);
and U6222 (N_6222,N_5846,N_5788);
and U6223 (N_6223,N_5958,N_5906);
nor U6224 (N_6224,N_5868,N_5882);
nand U6225 (N_6225,N_5821,N_5939);
and U6226 (N_6226,N_5806,N_5752);
xor U6227 (N_6227,N_5891,N_5932);
nor U6228 (N_6228,N_5888,N_5754);
xor U6229 (N_6229,N_5826,N_5910);
nor U6230 (N_6230,N_5931,N_5938);
xor U6231 (N_6231,N_5882,N_5877);
xor U6232 (N_6232,N_5807,N_5772);
and U6233 (N_6233,N_5814,N_5946);
nand U6234 (N_6234,N_5982,N_5791);
nand U6235 (N_6235,N_5895,N_5990);
nor U6236 (N_6236,N_5950,N_5922);
nor U6237 (N_6237,N_5780,N_5849);
nor U6238 (N_6238,N_5909,N_5961);
nand U6239 (N_6239,N_5979,N_5762);
nor U6240 (N_6240,N_5755,N_5827);
and U6241 (N_6241,N_5971,N_5857);
or U6242 (N_6242,N_5984,N_5956);
and U6243 (N_6243,N_5818,N_5988);
nor U6244 (N_6244,N_5983,N_5856);
and U6245 (N_6245,N_5974,N_5861);
xnor U6246 (N_6246,N_5963,N_5829);
xnor U6247 (N_6247,N_5864,N_5842);
nor U6248 (N_6248,N_5907,N_5867);
and U6249 (N_6249,N_5796,N_5768);
nor U6250 (N_6250,N_6138,N_6223);
and U6251 (N_6251,N_6199,N_6041);
nor U6252 (N_6252,N_6076,N_6129);
nor U6253 (N_6253,N_6142,N_6144);
xnor U6254 (N_6254,N_6085,N_6044);
nor U6255 (N_6255,N_6237,N_6033);
nand U6256 (N_6256,N_6230,N_6143);
or U6257 (N_6257,N_6080,N_6136);
nor U6258 (N_6258,N_6026,N_6231);
and U6259 (N_6259,N_6115,N_6017);
or U6260 (N_6260,N_6239,N_6028);
and U6261 (N_6261,N_6098,N_6067);
or U6262 (N_6262,N_6013,N_6141);
nand U6263 (N_6263,N_6179,N_6197);
nand U6264 (N_6264,N_6247,N_6075);
or U6265 (N_6265,N_6112,N_6225);
nand U6266 (N_6266,N_6185,N_6158);
or U6267 (N_6267,N_6206,N_6220);
nor U6268 (N_6268,N_6196,N_6228);
nor U6269 (N_6269,N_6042,N_6039);
nand U6270 (N_6270,N_6084,N_6093);
nor U6271 (N_6271,N_6131,N_6148);
nor U6272 (N_6272,N_6047,N_6245);
xor U6273 (N_6273,N_6030,N_6159);
nor U6274 (N_6274,N_6246,N_6011);
and U6275 (N_6275,N_6120,N_6051);
xor U6276 (N_6276,N_6130,N_6006);
nor U6277 (N_6277,N_6069,N_6232);
and U6278 (N_6278,N_6105,N_6053);
nor U6279 (N_6279,N_6204,N_6181);
nor U6280 (N_6280,N_6208,N_6027);
and U6281 (N_6281,N_6107,N_6235);
and U6282 (N_6282,N_6091,N_6116);
nand U6283 (N_6283,N_6173,N_6177);
xnor U6284 (N_6284,N_6032,N_6106);
nand U6285 (N_6285,N_6012,N_6134);
or U6286 (N_6286,N_6149,N_6025);
nor U6287 (N_6287,N_6070,N_6221);
nor U6288 (N_6288,N_6078,N_6122);
xnor U6289 (N_6289,N_6101,N_6203);
nand U6290 (N_6290,N_6156,N_6095);
and U6291 (N_6291,N_6040,N_6238);
nand U6292 (N_6292,N_6043,N_6154);
nand U6293 (N_6293,N_6211,N_6209);
nor U6294 (N_6294,N_6019,N_6077);
xnor U6295 (N_6295,N_6036,N_6088);
xnor U6296 (N_6296,N_6009,N_6083);
and U6297 (N_6297,N_6137,N_6200);
and U6298 (N_6298,N_6218,N_6191);
and U6299 (N_6299,N_6213,N_6065);
xnor U6300 (N_6300,N_6103,N_6180);
nor U6301 (N_6301,N_6187,N_6167);
or U6302 (N_6302,N_6125,N_6219);
nand U6303 (N_6303,N_6074,N_6150);
nand U6304 (N_6304,N_6099,N_6072);
and U6305 (N_6305,N_6233,N_6241);
and U6306 (N_6306,N_6016,N_6100);
xnor U6307 (N_6307,N_6057,N_6210);
nor U6308 (N_6308,N_6201,N_6182);
nand U6309 (N_6309,N_6014,N_6021);
and U6310 (N_6310,N_6198,N_6001);
nor U6311 (N_6311,N_6071,N_6108);
or U6312 (N_6312,N_6121,N_6062);
or U6313 (N_6313,N_6189,N_6104);
and U6314 (N_6314,N_6236,N_6248);
and U6315 (N_6315,N_6061,N_6045);
or U6316 (N_6316,N_6056,N_6176);
nor U6317 (N_6317,N_6094,N_6117);
or U6318 (N_6318,N_6163,N_6068);
and U6319 (N_6319,N_6145,N_6029);
nor U6320 (N_6320,N_6227,N_6217);
nand U6321 (N_6321,N_6073,N_6054);
nor U6322 (N_6322,N_6202,N_6124);
or U6323 (N_6323,N_6242,N_6034);
xnor U6324 (N_6324,N_6022,N_6172);
nand U6325 (N_6325,N_6058,N_6193);
nand U6326 (N_6326,N_6119,N_6166);
xnor U6327 (N_6327,N_6005,N_6055);
and U6328 (N_6328,N_6222,N_6212);
or U6329 (N_6329,N_6018,N_6063);
nor U6330 (N_6330,N_6002,N_6031);
or U6331 (N_6331,N_6089,N_6153);
and U6332 (N_6332,N_6171,N_6000);
xnor U6333 (N_6333,N_6035,N_6126);
and U6334 (N_6334,N_6165,N_6244);
and U6335 (N_6335,N_6090,N_6178);
nand U6336 (N_6336,N_6140,N_6157);
nor U6337 (N_6337,N_6183,N_6170);
xor U6338 (N_6338,N_6109,N_6086);
xnor U6339 (N_6339,N_6060,N_6132);
and U6340 (N_6340,N_6205,N_6234);
xor U6341 (N_6341,N_6139,N_6114);
and U6342 (N_6342,N_6081,N_6240);
xor U6343 (N_6343,N_6050,N_6243);
or U6344 (N_6344,N_6151,N_6037);
and U6345 (N_6345,N_6146,N_6175);
or U6346 (N_6346,N_6155,N_6184);
nor U6347 (N_6347,N_6079,N_6216);
and U6348 (N_6348,N_6066,N_6192);
or U6349 (N_6349,N_6004,N_6174);
xnor U6350 (N_6350,N_6007,N_6188);
nand U6351 (N_6351,N_6087,N_6128);
or U6352 (N_6352,N_6008,N_6038);
nand U6353 (N_6353,N_6195,N_6168);
nand U6354 (N_6354,N_6064,N_6229);
or U6355 (N_6355,N_6249,N_6023);
or U6356 (N_6356,N_6010,N_6152);
xnor U6357 (N_6357,N_6207,N_6015);
nor U6358 (N_6358,N_6133,N_6003);
nand U6359 (N_6359,N_6097,N_6111);
or U6360 (N_6360,N_6214,N_6082);
nor U6361 (N_6361,N_6024,N_6215);
xnor U6362 (N_6362,N_6110,N_6123);
or U6363 (N_6363,N_6135,N_6092);
nor U6364 (N_6364,N_6020,N_6052);
nand U6365 (N_6365,N_6186,N_6161);
and U6366 (N_6366,N_6147,N_6048);
nor U6367 (N_6367,N_6162,N_6194);
and U6368 (N_6368,N_6127,N_6049);
or U6369 (N_6369,N_6160,N_6046);
nand U6370 (N_6370,N_6113,N_6096);
and U6371 (N_6371,N_6224,N_6102);
nand U6372 (N_6372,N_6059,N_6226);
and U6373 (N_6373,N_6169,N_6190);
or U6374 (N_6374,N_6118,N_6164);
xnor U6375 (N_6375,N_6212,N_6072);
and U6376 (N_6376,N_6179,N_6044);
and U6377 (N_6377,N_6235,N_6144);
or U6378 (N_6378,N_6081,N_6010);
or U6379 (N_6379,N_6101,N_6154);
xnor U6380 (N_6380,N_6022,N_6110);
nor U6381 (N_6381,N_6045,N_6012);
or U6382 (N_6382,N_6143,N_6097);
or U6383 (N_6383,N_6138,N_6084);
nor U6384 (N_6384,N_6035,N_6006);
or U6385 (N_6385,N_6158,N_6076);
xor U6386 (N_6386,N_6208,N_6077);
xor U6387 (N_6387,N_6220,N_6185);
xor U6388 (N_6388,N_6227,N_6128);
nor U6389 (N_6389,N_6173,N_6203);
nand U6390 (N_6390,N_6241,N_6062);
nand U6391 (N_6391,N_6181,N_6078);
nand U6392 (N_6392,N_6039,N_6175);
and U6393 (N_6393,N_6057,N_6038);
xor U6394 (N_6394,N_6233,N_6016);
nor U6395 (N_6395,N_6046,N_6042);
nor U6396 (N_6396,N_6022,N_6175);
nor U6397 (N_6397,N_6244,N_6068);
xnor U6398 (N_6398,N_6099,N_6054);
xor U6399 (N_6399,N_6005,N_6193);
nor U6400 (N_6400,N_6124,N_6169);
and U6401 (N_6401,N_6199,N_6168);
or U6402 (N_6402,N_6041,N_6246);
or U6403 (N_6403,N_6172,N_6059);
and U6404 (N_6404,N_6229,N_6199);
and U6405 (N_6405,N_6129,N_6159);
or U6406 (N_6406,N_6149,N_6019);
and U6407 (N_6407,N_6135,N_6248);
nand U6408 (N_6408,N_6139,N_6021);
nor U6409 (N_6409,N_6071,N_6236);
nand U6410 (N_6410,N_6091,N_6113);
xnor U6411 (N_6411,N_6188,N_6208);
nand U6412 (N_6412,N_6040,N_6058);
or U6413 (N_6413,N_6160,N_6017);
or U6414 (N_6414,N_6058,N_6024);
and U6415 (N_6415,N_6125,N_6082);
or U6416 (N_6416,N_6079,N_6154);
nand U6417 (N_6417,N_6124,N_6018);
or U6418 (N_6418,N_6045,N_6228);
nand U6419 (N_6419,N_6098,N_6118);
and U6420 (N_6420,N_6232,N_6117);
or U6421 (N_6421,N_6104,N_6011);
or U6422 (N_6422,N_6056,N_6001);
nor U6423 (N_6423,N_6014,N_6188);
or U6424 (N_6424,N_6071,N_6181);
and U6425 (N_6425,N_6057,N_6108);
and U6426 (N_6426,N_6182,N_6195);
nand U6427 (N_6427,N_6140,N_6075);
and U6428 (N_6428,N_6066,N_6180);
nand U6429 (N_6429,N_6134,N_6017);
and U6430 (N_6430,N_6046,N_6075);
or U6431 (N_6431,N_6054,N_6000);
or U6432 (N_6432,N_6011,N_6215);
xor U6433 (N_6433,N_6130,N_6059);
or U6434 (N_6434,N_6099,N_6137);
and U6435 (N_6435,N_6032,N_6194);
or U6436 (N_6436,N_6195,N_6040);
and U6437 (N_6437,N_6122,N_6007);
xnor U6438 (N_6438,N_6143,N_6117);
and U6439 (N_6439,N_6011,N_6118);
and U6440 (N_6440,N_6118,N_6153);
xor U6441 (N_6441,N_6217,N_6154);
nor U6442 (N_6442,N_6000,N_6150);
nand U6443 (N_6443,N_6089,N_6054);
or U6444 (N_6444,N_6229,N_6164);
xor U6445 (N_6445,N_6226,N_6087);
nand U6446 (N_6446,N_6007,N_6163);
nor U6447 (N_6447,N_6239,N_6220);
or U6448 (N_6448,N_6224,N_6021);
nor U6449 (N_6449,N_6047,N_6219);
nand U6450 (N_6450,N_6184,N_6196);
or U6451 (N_6451,N_6211,N_6060);
and U6452 (N_6452,N_6237,N_6060);
or U6453 (N_6453,N_6187,N_6095);
or U6454 (N_6454,N_6047,N_6111);
nand U6455 (N_6455,N_6090,N_6113);
or U6456 (N_6456,N_6134,N_6069);
xnor U6457 (N_6457,N_6083,N_6160);
xnor U6458 (N_6458,N_6029,N_6175);
nor U6459 (N_6459,N_6179,N_6040);
nand U6460 (N_6460,N_6001,N_6207);
or U6461 (N_6461,N_6249,N_6086);
nand U6462 (N_6462,N_6240,N_6168);
xnor U6463 (N_6463,N_6107,N_6115);
or U6464 (N_6464,N_6114,N_6071);
xnor U6465 (N_6465,N_6214,N_6154);
nand U6466 (N_6466,N_6008,N_6035);
xnor U6467 (N_6467,N_6045,N_6236);
and U6468 (N_6468,N_6086,N_6058);
xor U6469 (N_6469,N_6148,N_6072);
and U6470 (N_6470,N_6211,N_6094);
or U6471 (N_6471,N_6045,N_6152);
xor U6472 (N_6472,N_6054,N_6108);
nand U6473 (N_6473,N_6150,N_6172);
or U6474 (N_6474,N_6178,N_6237);
xor U6475 (N_6475,N_6137,N_6198);
xor U6476 (N_6476,N_6064,N_6026);
and U6477 (N_6477,N_6035,N_6226);
and U6478 (N_6478,N_6161,N_6069);
or U6479 (N_6479,N_6248,N_6097);
or U6480 (N_6480,N_6088,N_6046);
nor U6481 (N_6481,N_6000,N_6249);
nor U6482 (N_6482,N_6027,N_6153);
and U6483 (N_6483,N_6214,N_6195);
nor U6484 (N_6484,N_6016,N_6028);
xnor U6485 (N_6485,N_6017,N_6215);
xnor U6486 (N_6486,N_6239,N_6015);
or U6487 (N_6487,N_6184,N_6120);
nor U6488 (N_6488,N_6127,N_6034);
nand U6489 (N_6489,N_6074,N_6134);
nor U6490 (N_6490,N_6212,N_6018);
nor U6491 (N_6491,N_6064,N_6030);
nor U6492 (N_6492,N_6167,N_6075);
and U6493 (N_6493,N_6125,N_6062);
or U6494 (N_6494,N_6179,N_6222);
and U6495 (N_6495,N_6028,N_6163);
xor U6496 (N_6496,N_6190,N_6062);
and U6497 (N_6497,N_6168,N_6069);
and U6498 (N_6498,N_6136,N_6121);
nor U6499 (N_6499,N_6198,N_6035);
nor U6500 (N_6500,N_6440,N_6376);
nand U6501 (N_6501,N_6448,N_6286);
or U6502 (N_6502,N_6310,N_6273);
nor U6503 (N_6503,N_6406,N_6322);
or U6504 (N_6504,N_6432,N_6267);
nor U6505 (N_6505,N_6383,N_6455);
or U6506 (N_6506,N_6329,N_6372);
xnor U6507 (N_6507,N_6358,N_6494);
nor U6508 (N_6508,N_6497,N_6466);
or U6509 (N_6509,N_6318,N_6435);
nor U6510 (N_6510,N_6446,N_6370);
or U6511 (N_6511,N_6429,N_6407);
nor U6512 (N_6512,N_6436,N_6332);
and U6513 (N_6513,N_6297,N_6315);
or U6514 (N_6514,N_6366,N_6290);
and U6515 (N_6515,N_6388,N_6265);
and U6516 (N_6516,N_6364,N_6454);
nand U6517 (N_6517,N_6387,N_6416);
nand U6518 (N_6518,N_6488,N_6258);
or U6519 (N_6519,N_6324,N_6319);
and U6520 (N_6520,N_6398,N_6452);
or U6521 (N_6521,N_6414,N_6347);
nand U6522 (N_6522,N_6447,N_6333);
nand U6523 (N_6523,N_6392,N_6338);
nand U6524 (N_6524,N_6363,N_6411);
or U6525 (N_6525,N_6423,N_6481);
xor U6526 (N_6526,N_6325,N_6274);
xor U6527 (N_6527,N_6473,N_6373);
or U6528 (N_6528,N_6441,N_6498);
xor U6529 (N_6529,N_6281,N_6254);
nor U6530 (N_6530,N_6302,N_6361);
nand U6531 (N_6531,N_6489,N_6276);
or U6532 (N_6532,N_6253,N_6493);
and U6533 (N_6533,N_6334,N_6353);
xnor U6534 (N_6534,N_6321,N_6465);
and U6535 (N_6535,N_6293,N_6391);
nor U6536 (N_6536,N_6356,N_6289);
nor U6537 (N_6537,N_6474,N_6284);
and U6538 (N_6538,N_6288,N_6349);
and U6539 (N_6539,N_6459,N_6399);
and U6540 (N_6540,N_6472,N_6311);
nand U6541 (N_6541,N_6394,N_6486);
xor U6542 (N_6542,N_6445,N_6331);
or U6543 (N_6543,N_6271,N_6345);
or U6544 (N_6544,N_6352,N_6393);
nand U6545 (N_6545,N_6336,N_6437);
xnor U6546 (N_6546,N_6357,N_6294);
nand U6547 (N_6547,N_6453,N_6419);
or U6548 (N_6548,N_6490,N_6269);
nor U6549 (N_6549,N_6450,N_6348);
nand U6550 (N_6550,N_6298,N_6263);
nand U6551 (N_6551,N_6327,N_6250);
nor U6552 (N_6552,N_6337,N_6438);
or U6553 (N_6553,N_6340,N_6312);
and U6554 (N_6554,N_6415,N_6301);
nor U6555 (N_6555,N_6480,N_6277);
and U6556 (N_6556,N_6444,N_6287);
nand U6557 (N_6557,N_6282,N_6479);
or U6558 (N_6558,N_6251,N_6280);
and U6559 (N_6559,N_6291,N_6461);
nor U6560 (N_6560,N_6292,N_6320);
or U6561 (N_6561,N_6330,N_6471);
or U6562 (N_6562,N_6272,N_6418);
nand U6563 (N_6563,N_6283,N_6428);
xnor U6564 (N_6564,N_6409,N_6378);
nor U6565 (N_6565,N_6463,N_6252);
xnor U6566 (N_6566,N_6257,N_6266);
or U6567 (N_6567,N_6279,N_6371);
nor U6568 (N_6568,N_6451,N_6341);
xnor U6569 (N_6569,N_6482,N_6468);
xnor U6570 (N_6570,N_6379,N_6420);
nor U6571 (N_6571,N_6499,N_6344);
nor U6572 (N_6572,N_6259,N_6300);
xnor U6573 (N_6573,N_6368,N_6412);
and U6574 (N_6574,N_6413,N_6261);
nor U6575 (N_6575,N_6256,N_6354);
and U6576 (N_6576,N_6492,N_6442);
nand U6577 (N_6577,N_6403,N_6475);
or U6578 (N_6578,N_6377,N_6314);
nand U6579 (N_6579,N_6395,N_6477);
nor U6580 (N_6580,N_6496,N_6365);
xor U6581 (N_6581,N_6404,N_6389);
and U6582 (N_6582,N_6390,N_6402);
and U6583 (N_6583,N_6408,N_6384);
and U6584 (N_6584,N_6483,N_6268);
xor U6585 (N_6585,N_6299,N_6421);
nor U6586 (N_6586,N_6359,N_6484);
and U6587 (N_6587,N_6439,N_6495);
nor U6588 (N_6588,N_6422,N_6426);
xor U6589 (N_6589,N_6458,N_6427);
xor U6590 (N_6590,N_6278,N_6306);
nand U6591 (N_6591,N_6469,N_6449);
or U6592 (N_6592,N_6313,N_6417);
and U6593 (N_6593,N_6262,N_6424);
nor U6594 (N_6594,N_6264,N_6386);
or U6595 (N_6595,N_6470,N_6443);
xor U6596 (N_6596,N_6462,N_6425);
xor U6597 (N_6597,N_6343,N_6303);
nand U6598 (N_6598,N_6355,N_6295);
xor U6599 (N_6599,N_6326,N_6317);
or U6600 (N_6600,N_6260,N_6375);
and U6601 (N_6601,N_6457,N_6360);
nand U6602 (N_6602,N_6335,N_6339);
xnor U6603 (N_6603,N_6382,N_6431);
or U6604 (N_6604,N_6362,N_6381);
or U6605 (N_6605,N_6296,N_6476);
xnor U6606 (N_6606,N_6346,N_6304);
or U6607 (N_6607,N_6396,N_6275);
and U6608 (N_6608,N_6328,N_6342);
nor U6609 (N_6609,N_6308,N_6385);
and U6610 (N_6610,N_6485,N_6405);
or U6611 (N_6611,N_6401,N_6369);
nand U6612 (N_6612,N_6487,N_6309);
xnor U6613 (N_6613,N_6270,N_6460);
nor U6614 (N_6614,N_6400,N_6491);
and U6615 (N_6615,N_6255,N_6433);
and U6616 (N_6616,N_6456,N_6316);
xnor U6617 (N_6617,N_6434,N_6478);
or U6618 (N_6618,N_6367,N_6374);
and U6619 (N_6619,N_6467,N_6350);
xor U6620 (N_6620,N_6380,N_6430);
xnor U6621 (N_6621,N_6464,N_6285);
and U6622 (N_6622,N_6323,N_6410);
nor U6623 (N_6623,N_6305,N_6397);
nand U6624 (N_6624,N_6307,N_6351);
xnor U6625 (N_6625,N_6281,N_6411);
nand U6626 (N_6626,N_6396,N_6408);
or U6627 (N_6627,N_6412,N_6250);
and U6628 (N_6628,N_6272,N_6298);
nand U6629 (N_6629,N_6362,N_6450);
or U6630 (N_6630,N_6490,N_6323);
nor U6631 (N_6631,N_6451,N_6470);
nand U6632 (N_6632,N_6436,N_6286);
nor U6633 (N_6633,N_6338,N_6408);
or U6634 (N_6634,N_6266,N_6408);
xor U6635 (N_6635,N_6380,N_6255);
nand U6636 (N_6636,N_6327,N_6252);
and U6637 (N_6637,N_6474,N_6341);
or U6638 (N_6638,N_6350,N_6439);
and U6639 (N_6639,N_6494,N_6262);
nand U6640 (N_6640,N_6342,N_6271);
nor U6641 (N_6641,N_6261,N_6391);
xnor U6642 (N_6642,N_6409,N_6341);
and U6643 (N_6643,N_6471,N_6454);
and U6644 (N_6644,N_6448,N_6375);
nand U6645 (N_6645,N_6381,N_6486);
and U6646 (N_6646,N_6455,N_6324);
and U6647 (N_6647,N_6477,N_6321);
xnor U6648 (N_6648,N_6360,N_6493);
or U6649 (N_6649,N_6318,N_6495);
nand U6650 (N_6650,N_6443,N_6429);
or U6651 (N_6651,N_6469,N_6274);
nor U6652 (N_6652,N_6311,N_6377);
and U6653 (N_6653,N_6480,N_6271);
or U6654 (N_6654,N_6441,N_6489);
and U6655 (N_6655,N_6333,N_6466);
and U6656 (N_6656,N_6397,N_6472);
nand U6657 (N_6657,N_6415,N_6352);
xnor U6658 (N_6658,N_6313,N_6349);
nand U6659 (N_6659,N_6415,N_6410);
and U6660 (N_6660,N_6257,N_6334);
xor U6661 (N_6661,N_6336,N_6455);
or U6662 (N_6662,N_6251,N_6265);
nand U6663 (N_6663,N_6490,N_6384);
nor U6664 (N_6664,N_6392,N_6441);
or U6665 (N_6665,N_6252,N_6269);
and U6666 (N_6666,N_6438,N_6484);
xor U6667 (N_6667,N_6336,N_6423);
xor U6668 (N_6668,N_6259,N_6253);
or U6669 (N_6669,N_6483,N_6480);
and U6670 (N_6670,N_6424,N_6358);
and U6671 (N_6671,N_6491,N_6383);
and U6672 (N_6672,N_6494,N_6497);
xor U6673 (N_6673,N_6359,N_6439);
xor U6674 (N_6674,N_6290,N_6270);
or U6675 (N_6675,N_6403,N_6414);
or U6676 (N_6676,N_6420,N_6342);
xnor U6677 (N_6677,N_6378,N_6490);
and U6678 (N_6678,N_6385,N_6319);
or U6679 (N_6679,N_6489,N_6499);
xnor U6680 (N_6680,N_6263,N_6300);
and U6681 (N_6681,N_6413,N_6355);
and U6682 (N_6682,N_6284,N_6368);
nor U6683 (N_6683,N_6305,N_6477);
xor U6684 (N_6684,N_6406,N_6437);
xor U6685 (N_6685,N_6498,N_6316);
nor U6686 (N_6686,N_6453,N_6478);
xnor U6687 (N_6687,N_6317,N_6340);
xor U6688 (N_6688,N_6317,N_6452);
and U6689 (N_6689,N_6320,N_6255);
and U6690 (N_6690,N_6489,N_6409);
xnor U6691 (N_6691,N_6446,N_6462);
or U6692 (N_6692,N_6329,N_6473);
or U6693 (N_6693,N_6392,N_6483);
nand U6694 (N_6694,N_6286,N_6498);
and U6695 (N_6695,N_6361,N_6457);
nand U6696 (N_6696,N_6450,N_6303);
nand U6697 (N_6697,N_6488,N_6484);
or U6698 (N_6698,N_6428,N_6261);
nand U6699 (N_6699,N_6300,N_6381);
nor U6700 (N_6700,N_6271,N_6386);
xnor U6701 (N_6701,N_6316,N_6409);
xnor U6702 (N_6702,N_6472,N_6283);
and U6703 (N_6703,N_6426,N_6493);
or U6704 (N_6704,N_6380,N_6328);
nand U6705 (N_6705,N_6468,N_6484);
or U6706 (N_6706,N_6469,N_6407);
and U6707 (N_6707,N_6287,N_6340);
or U6708 (N_6708,N_6293,N_6262);
and U6709 (N_6709,N_6335,N_6393);
nor U6710 (N_6710,N_6496,N_6338);
or U6711 (N_6711,N_6403,N_6291);
nor U6712 (N_6712,N_6448,N_6439);
nor U6713 (N_6713,N_6317,N_6450);
xor U6714 (N_6714,N_6272,N_6340);
or U6715 (N_6715,N_6496,N_6403);
and U6716 (N_6716,N_6321,N_6405);
and U6717 (N_6717,N_6473,N_6493);
nor U6718 (N_6718,N_6400,N_6365);
nor U6719 (N_6719,N_6308,N_6428);
nor U6720 (N_6720,N_6260,N_6439);
nor U6721 (N_6721,N_6355,N_6429);
nor U6722 (N_6722,N_6337,N_6275);
and U6723 (N_6723,N_6324,N_6453);
xor U6724 (N_6724,N_6338,N_6331);
and U6725 (N_6725,N_6488,N_6440);
or U6726 (N_6726,N_6365,N_6484);
xnor U6727 (N_6727,N_6415,N_6308);
nand U6728 (N_6728,N_6366,N_6468);
and U6729 (N_6729,N_6254,N_6322);
nor U6730 (N_6730,N_6363,N_6348);
xor U6731 (N_6731,N_6497,N_6440);
nor U6732 (N_6732,N_6328,N_6312);
and U6733 (N_6733,N_6489,N_6454);
nor U6734 (N_6734,N_6298,N_6350);
or U6735 (N_6735,N_6480,N_6387);
nor U6736 (N_6736,N_6497,N_6401);
or U6737 (N_6737,N_6352,N_6260);
and U6738 (N_6738,N_6339,N_6472);
nand U6739 (N_6739,N_6312,N_6301);
nand U6740 (N_6740,N_6360,N_6382);
xnor U6741 (N_6741,N_6372,N_6330);
xnor U6742 (N_6742,N_6270,N_6363);
xnor U6743 (N_6743,N_6347,N_6412);
nor U6744 (N_6744,N_6387,N_6499);
or U6745 (N_6745,N_6260,N_6373);
xor U6746 (N_6746,N_6388,N_6358);
xor U6747 (N_6747,N_6322,N_6333);
nand U6748 (N_6748,N_6263,N_6271);
xor U6749 (N_6749,N_6340,N_6327);
and U6750 (N_6750,N_6586,N_6693);
nor U6751 (N_6751,N_6574,N_6736);
and U6752 (N_6752,N_6580,N_6620);
xnor U6753 (N_6753,N_6566,N_6705);
nor U6754 (N_6754,N_6724,N_6717);
xor U6755 (N_6755,N_6641,N_6677);
nor U6756 (N_6756,N_6687,N_6697);
nand U6757 (N_6757,N_6730,N_6522);
xor U6758 (N_6758,N_6589,N_6619);
xor U6759 (N_6759,N_6639,N_6584);
and U6760 (N_6760,N_6531,N_6659);
nor U6761 (N_6761,N_6542,N_6636);
nand U6762 (N_6762,N_6595,N_6517);
and U6763 (N_6763,N_6640,N_6579);
or U6764 (N_6764,N_6544,N_6616);
xor U6765 (N_6765,N_6519,N_6568);
and U6766 (N_6766,N_6618,N_6582);
nor U6767 (N_6767,N_6699,N_6596);
nand U6768 (N_6768,N_6709,N_6622);
and U6769 (N_6769,N_6564,N_6602);
nor U6770 (N_6770,N_6534,N_6575);
or U6771 (N_6771,N_6681,N_6722);
or U6772 (N_6772,N_6538,N_6630);
nand U6773 (N_6773,N_6523,N_6704);
or U6774 (N_6774,N_6715,N_6621);
or U6775 (N_6775,N_6543,N_6701);
nand U6776 (N_6776,N_6707,N_6738);
and U6777 (N_6777,N_6652,N_6603);
or U6778 (N_6778,N_6708,N_6521);
nand U6779 (N_6779,N_6609,N_6626);
nand U6780 (N_6780,N_6668,N_6565);
xnor U6781 (N_6781,N_6550,N_6711);
xor U6782 (N_6782,N_6617,N_6578);
xor U6783 (N_6783,N_6663,N_6562);
nand U6784 (N_6784,N_6684,N_6665);
and U6785 (N_6785,N_6532,N_6552);
nor U6786 (N_6786,N_6624,N_6597);
and U6787 (N_6787,N_6694,N_6651);
nor U6788 (N_6788,N_6581,N_6655);
nor U6789 (N_6789,N_6572,N_6692);
nor U6790 (N_6790,N_6706,N_6607);
nor U6791 (N_6791,N_6653,N_6732);
nor U6792 (N_6792,N_6529,N_6551);
xnor U6793 (N_6793,N_6703,N_6537);
xnor U6794 (N_6794,N_6664,N_6669);
nor U6795 (N_6795,N_6646,N_6554);
and U6796 (N_6796,N_6576,N_6642);
or U6797 (N_6797,N_6737,N_6674);
or U6798 (N_6798,N_6747,N_6645);
and U6799 (N_6799,N_6745,N_6739);
and U6800 (N_6800,N_6726,N_6689);
nand U6801 (N_6801,N_6503,N_6506);
and U6802 (N_6802,N_6555,N_6556);
or U6803 (N_6803,N_6611,N_6656);
xnor U6804 (N_6804,N_6627,N_6673);
nand U6805 (N_6805,N_6746,N_6604);
xor U6806 (N_6806,N_6505,N_6593);
nand U6807 (N_6807,N_6546,N_6691);
and U6808 (N_6808,N_6508,N_6558);
xnor U6809 (N_6809,N_6649,N_6612);
and U6810 (N_6810,N_6741,N_6591);
or U6811 (N_6811,N_6535,N_6658);
or U6812 (N_6812,N_6567,N_6592);
xor U6813 (N_6813,N_6514,N_6749);
nand U6814 (N_6814,N_6650,N_6661);
and U6815 (N_6815,N_6524,N_6629);
or U6816 (N_6816,N_6507,N_6637);
xor U6817 (N_6817,N_6509,N_6520);
nor U6818 (N_6818,N_6539,N_6632);
and U6819 (N_6819,N_6504,N_6683);
nor U6820 (N_6820,N_6634,N_6744);
xnor U6821 (N_6821,N_6588,N_6710);
nor U6822 (N_6822,N_6561,N_6686);
nor U6823 (N_6823,N_6702,N_6608);
nand U6824 (N_6824,N_6599,N_6547);
or U6825 (N_6825,N_6571,N_6695);
and U6826 (N_6826,N_6671,N_6713);
and U6827 (N_6827,N_6500,N_6700);
nand U6828 (N_6828,N_6721,N_6698);
xnor U6829 (N_6829,N_6657,N_6635);
nand U6830 (N_6830,N_6676,N_6678);
xor U6831 (N_6831,N_6680,N_6728);
nor U6832 (N_6832,N_6557,N_6719);
xnor U6833 (N_6833,N_6569,N_6734);
nand U6834 (N_6834,N_6648,N_6615);
nor U6835 (N_6835,N_6605,N_6654);
and U6836 (N_6836,N_6696,N_6714);
nor U6837 (N_6837,N_6614,N_6525);
and U6838 (N_6838,N_6501,N_6563);
nor U6839 (N_6839,N_6553,N_6526);
nor U6840 (N_6840,N_6573,N_6548);
nand U6841 (N_6841,N_6590,N_6682);
xor U6842 (N_6842,N_6685,N_6540);
nor U6843 (N_6843,N_6512,N_6729);
nor U6844 (N_6844,N_6712,N_6577);
nand U6845 (N_6845,N_6670,N_6513);
xnor U6846 (N_6846,N_6583,N_6613);
and U6847 (N_6847,N_6533,N_6631);
or U6848 (N_6848,N_6528,N_6623);
or U6849 (N_6849,N_6672,N_6731);
xor U6850 (N_6850,N_6610,N_6587);
or U6851 (N_6851,N_6690,N_6725);
and U6852 (N_6852,N_6643,N_6723);
nand U6853 (N_6853,N_6510,N_6606);
xor U6854 (N_6854,N_6727,N_6600);
and U6855 (N_6855,N_6516,N_6735);
xor U6856 (N_6856,N_6570,N_6502);
nor U6857 (N_6857,N_6742,N_6559);
xnor U6858 (N_6858,N_6748,N_6718);
nor U6859 (N_6859,N_6625,N_6541);
nor U6860 (N_6860,N_6585,N_6515);
nor U6861 (N_6861,N_6511,N_6688);
or U6862 (N_6862,N_6660,N_6601);
nor U6863 (N_6863,N_6527,N_6667);
or U6864 (N_6864,N_6644,N_6679);
and U6865 (N_6865,N_6549,N_6666);
nand U6866 (N_6866,N_6518,N_6716);
nand U6867 (N_6867,N_6675,N_6740);
nand U6868 (N_6868,N_6560,N_6662);
or U6869 (N_6869,N_6598,N_6743);
nor U6870 (N_6870,N_6536,N_6530);
nor U6871 (N_6871,N_6647,N_6720);
or U6872 (N_6872,N_6628,N_6638);
nor U6873 (N_6873,N_6545,N_6733);
and U6874 (N_6874,N_6594,N_6633);
and U6875 (N_6875,N_6589,N_6597);
xnor U6876 (N_6876,N_6730,N_6601);
and U6877 (N_6877,N_6666,N_6714);
nand U6878 (N_6878,N_6555,N_6636);
or U6879 (N_6879,N_6537,N_6608);
nand U6880 (N_6880,N_6615,N_6724);
nand U6881 (N_6881,N_6658,N_6615);
or U6882 (N_6882,N_6660,N_6742);
nor U6883 (N_6883,N_6690,N_6634);
nand U6884 (N_6884,N_6527,N_6692);
nor U6885 (N_6885,N_6607,N_6743);
nor U6886 (N_6886,N_6507,N_6529);
and U6887 (N_6887,N_6742,N_6593);
or U6888 (N_6888,N_6624,N_6711);
or U6889 (N_6889,N_6743,N_6631);
nor U6890 (N_6890,N_6711,N_6710);
xnor U6891 (N_6891,N_6635,N_6532);
or U6892 (N_6892,N_6695,N_6598);
and U6893 (N_6893,N_6678,N_6574);
nand U6894 (N_6894,N_6650,N_6525);
xor U6895 (N_6895,N_6659,N_6642);
nor U6896 (N_6896,N_6727,N_6509);
xnor U6897 (N_6897,N_6578,N_6728);
xnor U6898 (N_6898,N_6519,N_6708);
xnor U6899 (N_6899,N_6527,N_6526);
nor U6900 (N_6900,N_6736,N_6718);
nand U6901 (N_6901,N_6693,N_6508);
nor U6902 (N_6902,N_6747,N_6740);
nor U6903 (N_6903,N_6559,N_6749);
xor U6904 (N_6904,N_6517,N_6501);
or U6905 (N_6905,N_6707,N_6713);
and U6906 (N_6906,N_6672,N_6704);
nor U6907 (N_6907,N_6661,N_6725);
or U6908 (N_6908,N_6639,N_6621);
nand U6909 (N_6909,N_6561,N_6707);
nand U6910 (N_6910,N_6573,N_6679);
nor U6911 (N_6911,N_6635,N_6699);
or U6912 (N_6912,N_6670,N_6501);
or U6913 (N_6913,N_6725,N_6572);
or U6914 (N_6914,N_6718,N_6521);
nor U6915 (N_6915,N_6678,N_6735);
or U6916 (N_6916,N_6518,N_6679);
or U6917 (N_6917,N_6504,N_6534);
nor U6918 (N_6918,N_6607,N_6521);
nor U6919 (N_6919,N_6701,N_6527);
and U6920 (N_6920,N_6500,N_6525);
xor U6921 (N_6921,N_6671,N_6589);
and U6922 (N_6922,N_6552,N_6568);
or U6923 (N_6923,N_6702,N_6698);
nand U6924 (N_6924,N_6719,N_6570);
xor U6925 (N_6925,N_6688,N_6615);
xor U6926 (N_6926,N_6508,N_6629);
or U6927 (N_6927,N_6615,N_6567);
nor U6928 (N_6928,N_6714,N_6531);
nand U6929 (N_6929,N_6582,N_6714);
and U6930 (N_6930,N_6680,N_6601);
nor U6931 (N_6931,N_6537,N_6734);
xor U6932 (N_6932,N_6623,N_6714);
or U6933 (N_6933,N_6676,N_6530);
and U6934 (N_6934,N_6690,N_6588);
xor U6935 (N_6935,N_6733,N_6569);
or U6936 (N_6936,N_6559,N_6727);
xnor U6937 (N_6937,N_6567,N_6706);
xor U6938 (N_6938,N_6745,N_6644);
and U6939 (N_6939,N_6535,N_6614);
or U6940 (N_6940,N_6603,N_6599);
nor U6941 (N_6941,N_6574,N_6676);
nand U6942 (N_6942,N_6540,N_6656);
and U6943 (N_6943,N_6551,N_6585);
or U6944 (N_6944,N_6505,N_6711);
nor U6945 (N_6945,N_6575,N_6621);
nor U6946 (N_6946,N_6685,N_6713);
nor U6947 (N_6947,N_6596,N_6535);
xor U6948 (N_6948,N_6658,N_6523);
and U6949 (N_6949,N_6573,N_6554);
and U6950 (N_6950,N_6670,N_6616);
and U6951 (N_6951,N_6582,N_6608);
xor U6952 (N_6952,N_6567,N_6590);
and U6953 (N_6953,N_6649,N_6590);
xnor U6954 (N_6954,N_6632,N_6692);
nor U6955 (N_6955,N_6534,N_6714);
nor U6956 (N_6956,N_6506,N_6573);
nor U6957 (N_6957,N_6749,N_6707);
or U6958 (N_6958,N_6637,N_6728);
and U6959 (N_6959,N_6731,N_6539);
or U6960 (N_6960,N_6747,N_6721);
xnor U6961 (N_6961,N_6521,N_6559);
nor U6962 (N_6962,N_6687,N_6620);
or U6963 (N_6963,N_6650,N_6585);
or U6964 (N_6964,N_6608,N_6737);
nor U6965 (N_6965,N_6641,N_6742);
nand U6966 (N_6966,N_6725,N_6711);
nor U6967 (N_6967,N_6574,N_6737);
nor U6968 (N_6968,N_6674,N_6700);
and U6969 (N_6969,N_6588,N_6528);
and U6970 (N_6970,N_6637,N_6658);
nor U6971 (N_6971,N_6671,N_6679);
nor U6972 (N_6972,N_6747,N_6596);
and U6973 (N_6973,N_6645,N_6679);
nand U6974 (N_6974,N_6653,N_6578);
nor U6975 (N_6975,N_6628,N_6510);
nand U6976 (N_6976,N_6561,N_6667);
xnor U6977 (N_6977,N_6654,N_6589);
nand U6978 (N_6978,N_6507,N_6677);
nand U6979 (N_6979,N_6669,N_6616);
nand U6980 (N_6980,N_6616,N_6511);
or U6981 (N_6981,N_6679,N_6681);
or U6982 (N_6982,N_6745,N_6538);
nor U6983 (N_6983,N_6736,N_6705);
or U6984 (N_6984,N_6742,N_6580);
xor U6985 (N_6985,N_6710,N_6530);
and U6986 (N_6986,N_6720,N_6523);
nand U6987 (N_6987,N_6702,N_6600);
or U6988 (N_6988,N_6533,N_6512);
and U6989 (N_6989,N_6704,N_6569);
xnor U6990 (N_6990,N_6691,N_6696);
or U6991 (N_6991,N_6719,N_6579);
and U6992 (N_6992,N_6560,N_6681);
and U6993 (N_6993,N_6607,N_6552);
xor U6994 (N_6994,N_6575,N_6696);
nor U6995 (N_6995,N_6568,N_6733);
or U6996 (N_6996,N_6616,N_6693);
nor U6997 (N_6997,N_6621,N_6544);
xor U6998 (N_6998,N_6613,N_6530);
nor U6999 (N_6999,N_6664,N_6714);
nor U7000 (N_7000,N_6990,N_6772);
and U7001 (N_7001,N_6947,N_6825);
nor U7002 (N_7002,N_6887,N_6890);
xor U7003 (N_7003,N_6861,N_6885);
nor U7004 (N_7004,N_6801,N_6935);
nand U7005 (N_7005,N_6831,N_6928);
nand U7006 (N_7006,N_6973,N_6921);
xor U7007 (N_7007,N_6770,N_6873);
or U7008 (N_7008,N_6846,N_6849);
or U7009 (N_7009,N_6858,N_6933);
and U7010 (N_7010,N_6970,N_6785);
nor U7011 (N_7011,N_6828,N_6917);
and U7012 (N_7012,N_6852,N_6905);
and U7013 (N_7013,N_6919,N_6775);
nor U7014 (N_7014,N_6945,N_6886);
xor U7015 (N_7015,N_6914,N_6755);
and U7016 (N_7016,N_6763,N_6868);
nand U7017 (N_7017,N_6881,N_6842);
xnor U7018 (N_7018,N_6994,N_6958);
xor U7019 (N_7019,N_6851,N_6844);
or U7020 (N_7020,N_6880,N_6957);
xor U7021 (N_7021,N_6894,N_6754);
xnor U7022 (N_7022,N_6901,N_6904);
nor U7023 (N_7023,N_6834,N_6789);
nand U7024 (N_7024,N_6984,N_6790);
nor U7025 (N_7025,N_6893,N_6792);
nor U7026 (N_7026,N_6767,N_6977);
nor U7027 (N_7027,N_6758,N_6929);
xnor U7028 (N_7028,N_6839,N_6757);
xnor U7029 (N_7029,N_6949,N_6938);
nor U7030 (N_7030,N_6830,N_6819);
and U7031 (N_7031,N_6814,N_6838);
and U7032 (N_7032,N_6804,N_6798);
nor U7033 (N_7033,N_6965,N_6840);
xnor U7034 (N_7034,N_6934,N_6907);
or U7035 (N_7035,N_6779,N_6912);
and U7036 (N_7036,N_6913,N_6824);
and U7037 (N_7037,N_6867,N_6930);
xor U7038 (N_7038,N_6948,N_6883);
xnor U7039 (N_7039,N_6997,N_6931);
xnor U7040 (N_7040,N_6972,N_6891);
or U7041 (N_7041,N_6897,N_6971);
or U7042 (N_7042,N_6769,N_6878);
and U7043 (N_7043,N_6969,N_6850);
nand U7044 (N_7044,N_6906,N_6916);
xnor U7045 (N_7045,N_6812,N_6974);
or U7046 (N_7046,N_6818,N_6955);
and U7047 (N_7047,N_6756,N_6799);
xor U7048 (N_7048,N_6855,N_6845);
or U7049 (N_7049,N_6899,N_6833);
and U7050 (N_7050,N_6927,N_6918);
or U7051 (N_7051,N_6988,N_6848);
or U7052 (N_7052,N_6764,N_6956);
xor U7053 (N_7053,N_6888,N_6787);
xor U7054 (N_7054,N_6778,N_6750);
or U7055 (N_7055,N_6966,N_6992);
xnor U7056 (N_7056,N_6832,N_6853);
and U7057 (N_7057,N_6835,N_6782);
xnor U7058 (N_7058,N_6946,N_6982);
nor U7059 (N_7059,N_6922,N_6866);
and U7060 (N_7060,N_6944,N_6978);
or U7061 (N_7061,N_6815,N_6877);
nand U7062 (N_7062,N_6869,N_6995);
nor U7063 (N_7063,N_6985,N_6963);
and U7064 (N_7064,N_6940,N_6797);
or U7065 (N_7065,N_6872,N_6765);
xnor U7066 (N_7066,N_6976,N_6937);
xnor U7067 (N_7067,N_6822,N_6908);
xor U7068 (N_7068,N_6968,N_6920);
nand U7069 (N_7069,N_6871,N_6820);
xnor U7070 (N_7070,N_6942,N_6816);
and U7071 (N_7071,N_6771,N_6943);
xor U7072 (N_7072,N_6898,N_6761);
nor U7073 (N_7073,N_6857,N_6788);
nand U7074 (N_7074,N_6903,N_6895);
xnor U7075 (N_7075,N_6875,N_6795);
xnor U7076 (N_7076,N_6776,N_6759);
xnor U7077 (N_7077,N_6975,N_6837);
or U7078 (N_7078,N_6941,N_6981);
xor U7079 (N_7079,N_6859,N_6962);
and U7080 (N_7080,N_6967,N_6959);
and U7081 (N_7081,N_6793,N_6987);
nand U7082 (N_7082,N_6915,N_6900);
or U7083 (N_7083,N_6829,N_6800);
nor U7084 (N_7084,N_6847,N_6999);
or U7085 (N_7085,N_6951,N_6989);
and U7086 (N_7086,N_6753,N_6760);
xnor U7087 (N_7087,N_6811,N_6983);
nand U7088 (N_7088,N_6932,N_6841);
xnor U7089 (N_7089,N_6817,N_6925);
and U7090 (N_7090,N_6993,N_6865);
and U7091 (N_7091,N_6784,N_6979);
nand U7092 (N_7092,N_6996,N_6980);
nand U7093 (N_7093,N_6860,N_6802);
nor U7094 (N_7094,N_6774,N_6936);
xor U7095 (N_7095,N_6773,N_6864);
or U7096 (N_7096,N_6964,N_6862);
xnor U7097 (N_7097,N_6889,N_6809);
xnor U7098 (N_7098,N_6808,N_6939);
nand U7099 (N_7099,N_6910,N_6896);
xor U7100 (N_7100,N_6783,N_6923);
nor U7101 (N_7101,N_6870,N_6892);
nand U7102 (N_7102,N_6836,N_6805);
and U7103 (N_7103,N_6777,N_6780);
nand U7104 (N_7104,N_6960,N_6879);
nor U7105 (N_7105,N_6986,N_6882);
nor U7106 (N_7106,N_6751,N_6961);
or U7107 (N_7107,N_6813,N_6926);
nor U7108 (N_7108,N_6781,N_6843);
nand U7109 (N_7109,N_6856,N_6794);
and U7110 (N_7110,N_6952,N_6806);
and U7111 (N_7111,N_6821,N_6924);
xor U7112 (N_7112,N_6766,N_6991);
xor U7113 (N_7113,N_6826,N_6854);
xnor U7114 (N_7114,N_6954,N_6909);
nor U7115 (N_7115,N_6998,N_6752);
and U7116 (N_7116,N_6807,N_6827);
xnor U7117 (N_7117,N_6874,N_6823);
nor U7118 (N_7118,N_6863,N_6768);
or U7119 (N_7119,N_6953,N_6876);
xnor U7120 (N_7120,N_6950,N_6791);
nor U7121 (N_7121,N_6810,N_6803);
and U7122 (N_7122,N_6911,N_6762);
nor U7123 (N_7123,N_6884,N_6902);
nand U7124 (N_7124,N_6786,N_6796);
nor U7125 (N_7125,N_6796,N_6887);
or U7126 (N_7126,N_6863,N_6988);
xor U7127 (N_7127,N_6912,N_6835);
and U7128 (N_7128,N_6824,N_6769);
or U7129 (N_7129,N_6895,N_6858);
or U7130 (N_7130,N_6960,N_6932);
nand U7131 (N_7131,N_6836,N_6812);
and U7132 (N_7132,N_6780,N_6903);
nor U7133 (N_7133,N_6990,N_6924);
nor U7134 (N_7134,N_6769,N_6935);
nand U7135 (N_7135,N_6851,N_6902);
or U7136 (N_7136,N_6877,N_6962);
nor U7137 (N_7137,N_6959,N_6955);
xnor U7138 (N_7138,N_6913,N_6906);
and U7139 (N_7139,N_6987,N_6976);
and U7140 (N_7140,N_6822,N_6877);
and U7141 (N_7141,N_6902,N_6785);
and U7142 (N_7142,N_6901,N_6949);
xor U7143 (N_7143,N_6889,N_6958);
nand U7144 (N_7144,N_6898,N_6909);
xnor U7145 (N_7145,N_6943,N_6942);
and U7146 (N_7146,N_6912,N_6951);
nand U7147 (N_7147,N_6820,N_6842);
xnor U7148 (N_7148,N_6991,N_6826);
and U7149 (N_7149,N_6879,N_6847);
nand U7150 (N_7150,N_6963,N_6872);
nor U7151 (N_7151,N_6855,N_6797);
and U7152 (N_7152,N_6968,N_6780);
or U7153 (N_7153,N_6759,N_6764);
and U7154 (N_7154,N_6822,N_6844);
xnor U7155 (N_7155,N_6999,N_6765);
or U7156 (N_7156,N_6783,N_6848);
or U7157 (N_7157,N_6823,N_6833);
nand U7158 (N_7158,N_6877,N_6927);
xnor U7159 (N_7159,N_6956,N_6988);
or U7160 (N_7160,N_6872,N_6981);
or U7161 (N_7161,N_6956,N_6762);
and U7162 (N_7162,N_6765,N_6783);
or U7163 (N_7163,N_6980,N_6750);
nand U7164 (N_7164,N_6964,N_6762);
or U7165 (N_7165,N_6847,N_6869);
and U7166 (N_7166,N_6910,N_6901);
nand U7167 (N_7167,N_6981,N_6973);
or U7168 (N_7168,N_6961,N_6773);
or U7169 (N_7169,N_6778,N_6861);
xor U7170 (N_7170,N_6921,N_6988);
and U7171 (N_7171,N_6784,N_6820);
or U7172 (N_7172,N_6930,N_6892);
nor U7173 (N_7173,N_6769,N_6944);
or U7174 (N_7174,N_6913,N_6893);
nor U7175 (N_7175,N_6897,N_6776);
nor U7176 (N_7176,N_6798,N_6764);
and U7177 (N_7177,N_6824,N_6823);
xnor U7178 (N_7178,N_6901,N_6853);
nand U7179 (N_7179,N_6844,N_6977);
nand U7180 (N_7180,N_6952,N_6893);
nor U7181 (N_7181,N_6865,N_6834);
xor U7182 (N_7182,N_6776,N_6981);
nand U7183 (N_7183,N_6836,N_6833);
nor U7184 (N_7184,N_6837,N_6910);
nand U7185 (N_7185,N_6754,N_6802);
nand U7186 (N_7186,N_6901,N_6959);
and U7187 (N_7187,N_6761,N_6878);
nor U7188 (N_7188,N_6979,N_6968);
nand U7189 (N_7189,N_6910,N_6766);
xnor U7190 (N_7190,N_6776,N_6843);
or U7191 (N_7191,N_6772,N_6885);
nand U7192 (N_7192,N_6831,N_6758);
nand U7193 (N_7193,N_6973,N_6859);
nor U7194 (N_7194,N_6910,N_6933);
and U7195 (N_7195,N_6923,N_6924);
nand U7196 (N_7196,N_6828,N_6820);
nand U7197 (N_7197,N_6913,N_6970);
nand U7198 (N_7198,N_6835,N_6925);
nor U7199 (N_7199,N_6889,N_6966);
or U7200 (N_7200,N_6904,N_6988);
and U7201 (N_7201,N_6870,N_6848);
or U7202 (N_7202,N_6862,N_6803);
nand U7203 (N_7203,N_6915,N_6771);
and U7204 (N_7204,N_6885,N_6830);
and U7205 (N_7205,N_6840,N_6948);
or U7206 (N_7206,N_6777,N_6805);
nor U7207 (N_7207,N_6893,N_6777);
nor U7208 (N_7208,N_6989,N_6820);
and U7209 (N_7209,N_6895,N_6865);
nor U7210 (N_7210,N_6896,N_6973);
or U7211 (N_7211,N_6832,N_6906);
nand U7212 (N_7212,N_6854,N_6828);
xor U7213 (N_7213,N_6805,N_6852);
or U7214 (N_7214,N_6925,N_6764);
and U7215 (N_7215,N_6810,N_6845);
nor U7216 (N_7216,N_6888,N_6977);
or U7217 (N_7217,N_6991,N_6760);
nand U7218 (N_7218,N_6917,N_6896);
or U7219 (N_7219,N_6954,N_6899);
nor U7220 (N_7220,N_6946,N_6887);
nor U7221 (N_7221,N_6839,N_6864);
nand U7222 (N_7222,N_6751,N_6836);
nor U7223 (N_7223,N_6794,N_6932);
nor U7224 (N_7224,N_6859,N_6984);
xor U7225 (N_7225,N_6942,N_6769);
nand U7226 (N_7226,N_6885,N_6766);
and U7227 (N_7227,N_6978,N_6823);
nand U7228 (N_7228,N_6827,N_6850);
or U7229 (N_7229,N_6913,N_6774);
or U7230 (N_7230,N_6947,N_6809);
nand U7231 (N_7231,N_6871,N_6910);
or U7232 (N_7232,N_6974,N_6797);
nor U7233 (N_7233,N_6873,N_6800);
and U7234 (N_7234,N_6926,N_6768);
xor U7235 (N_7235,N_6838,N_6840);
and U7236 (N_7236,N_6800,N_6847);
or U7237 (N_7237,N_6974,N_6977);
and U7238 (N_7238,N_6824,N_6847);
nor U7239 (N_7239,N_6967,N_6907);
nand U7240 (N_7240,N_6864,N_6888);
nor U7241 (N_7241,N_6789,N_6762);
xor U7242 (N_7242,N_6879,N_6873);
xnor U7243 (N_7243,N_6921,N_6908);
or U7244 (N_7244,N_6950,N_6989);
nor U7245 (N_7245,N_6986,N_6909);
and U7246 (N_7246,N_6939,N_6994);
xnor U7247 (N_7247,N_6894,N_6961);
xor U7248 (N_7248,N_6995,N_6808);
or U7249 (N_7249,N_6849,N_6786);
and U7250 (N_7250,N_7124,N_7221);
or U7251 (N_7251,N_7113,N_7181);
and U7252 (N_7252,N_7013,N_7174);
or U7253 (N_7253,N_7020,N_7232);
nand U7254 (N_7254,N_7139,N_7136);
nor U7255 (N_7255,N_7083,N_7141);
nand U7256 (N_7256,N_7234,N_7054);
nand U7257 (N_7257,N_7168,N_7241);
nor U7258 (N_7258,N_7009,N_7103);
or U7259 (N_7259,N_7215,N_7153);
nor U7260 (N_7260,N_7098,N_7143);
or U7261 (N_7261,N_7201,N_7178);
and U7262 (N_7262,N_7146,N_7203);
nor U7263 (N_7263,N_7014,N_7173);
nand U7264 (N_7264,N_7194,N_7188);
and U7265 (N_7265,N_7145,N_7017);
nand U7266 (N_7266,N_7069,N_7056);
xor U7267 (N_7267,N_7209,N_7092);
and U7268 (N_7268,N_7161,N_7055);
and U7269 (N_7269,N_7202,N_7175);
or U7270 (N_7270,N_7199,N_7224);
xor U7271 (N_7271,N_7245,N_7176);
xnor U7272 (N_7272,N_7072,N_7179);
or U7273 (N_7273,N_7063,N_7101);
nand U7274 (N_7274,N_7163,N_7147);
nand U7275 (N_7275,N_7090,N_7151);
xor U7276 (N_7276,N_7104,N_7213);
xor U7277 (N_7277,N_7105,N_7135);
nor U7278 (N_7278,N_7021,N_7002);
or U7279 (N_7279,N_7042,N_7015);
xnor U7280 (N_7280,N_7166,N_7027);
or U7281 (N_7281,N_7036,N_7067);
or U7282 (N_7282,N_7058,N_7133);
nor U7283 (N_7283,N_7074,N_7038);
nor U7284 (N_7284,N_7084,N_7210);
nand U7285 (N_7285,N_7010,N_7160);
or U7286 (N_7286,N_7087,N_7193);
and U7287 (N_7287,N_7190,N_7032);
nor U7288 (N_7288,N_7128,N_7080);
xnor U7289 (N_7289,N_7064,N_7100);
and U7290 (N_7290,N_7212,N_7137);
and U7291 (N_7291,N_7073,N_7066);
or U7292 (N_7292,N_7122,N_7220);
nand U7293 (N_7293,N_7109,N_7233);
or U7294 (N_7294,N_7004,N_7142);
xor U7295 (N_7295,N_7031,N_7205);
nand U7296 (N_7296,N_7140,N_7039);
and U7297 (N_7297,N_7244,N_7240);
nand U7298 (N_7298,N_7217,N_7247);
nor U7299 (N_7299,N_7115,N_7216);
nand U7300 (N_7300,N_7192,N_7119);
nand U7301 (N_7301,N_7062,N_7162);
and U7302 (N_7302,N_7195,N_7191);
nand U7303 (N_7303,N_7231,N_7048);
or U7304 (N_7304,N_7171,N_7030);
and U7305 (N_7305,N_7034,N_7094);
or U7306 (N_7306,N_7006,N_7189);
or U7307 (N_7307,N_7246,N_7249);
or U7308 (N_7308,N_7005,N_7076);
nor U7309 (N_7309,N_7184,N_7001);
nor U7310 (N_7310,N_7110,N_7214);
nand U7311 (N_7311,N_7060,N_7208);
nand U7312 (N_7312,N_7131,N_7125);
and U7313 (N_7313,N_7012,N_7235);
and U7314 (N_7314,N_7040,N_7126);
nand U7315 (N_7315,N_7046,N_7198);
nor U7316 (N_7316,N_7129,N_7047);
or U7317 (N_7317,N_7051,N_7061);
or U7318 (N_7318,N_7049,N_7117);
or U7319 (N_7319,N_7229,N_7230);
xor U7320 (N_7320,N_7099,N_7157);
xor U7321 (N_7321,N_7182,N_7070);
nor U7322 (N_7322,N_7077,N_7204);
or U7323 (N_7323,N_7223,N_7238);
xor U7324 (N_7324,N_7152,N_7120);
xnor U7325 (N_7325,N_7096,N_7127);
and U7326 (N_7326,N_7022,N_7035);
and U7327 (N_7327,N_7024,N_7025);
and U7328 (N_7328,N_7185,N_7097);
xnor U7329 (N_7329,N_7144,N_7075);
and U7330 (N_7330,N_7091,N_7052);
xnor U7331 (N_7331,N_7003,N_7134);
xnor U7332 (N_7332,N_7044,N_7148);
and U7333 (N_7333,N_7180,N_7078);
and U7334 (N_7334,N_7165,N_7079);
or U7335 (N_7335,N_7082,N_7023);
and U7336 (N_7336,N_7037,N_7007);
nor U7337 (N_7337,N_7222,N_7242);
and U7338 (N_7338,N_7111,N_7057);
or U7339 (N_7339,N_7239,N_7236);
or U7340 (N_7340,N_7130,N_7118);
and U7341 (N_7341,N_7237,N_7196);
and U7342 (N_7342,N_7187,N_7095);
nor U7343 (N_7343,N_7028,N_7200);
xnor U7344 (N_7344,N_7226,N_7041);
nand U7345 (N_7345,N_7159,N_7164);
and U7346 (N_7346,N_7207,N_7132);
xnor U7347 (N_7347,N_7008,N_7156);
nor U7348 (N_7348,N_7107,N_7116);
xor U7349 (N_7349,N_7065,N_7089);
xnor U7350 (N_7350,N_7154,N_7225);
xnor U7351 (N_7351,N_7093,N_7059);
nand U7352 (N_7352,N_7150,N_7088);
nand U7353 (N_7353,N_7243,N_7106);
nor U7354 (N_7354,N_7228,N_7011);
nand U7355 (N_7355,N_7050,N_7112);
or U7356 (N_7356,N_7000,N_7068);
xnor U7357 (N_7357,N_7033,N_7114);
nand U7358 (N_7358,N_7045,N_7071);
xnor U7359 (N_7359,N_7138,N_7197);
xor U7360 (N_7360,N_7206,N_7086);
nor U7361 (N_7361,N_7248,N_7155);
or U7362 (N_7362,N_7043,N_7121);
and U7363 (N_7363,N_7053,N_7016);
xor U7364 (N_7364,N_7183,N_7211);
xor U7365 (N_7365,N_7219,N_7123);
nand U7366 (N_7366,N_7029,N_7177);
or U7367 (N_7367,N_7158,N_7102);
or U7368 (N_7368,N_7186,N_7172);
nand U7369 (N_7369,N_7169,N_7227);
xnor U7370 (N_7370,N_7167,N_7108);
nor U7371 (N_7371,N_7149,N_7081);
and U7372 (N_7372,N_7019,N_7170);
nand U7373 (N_7373,N_7018,N_7218);
or U7374 (N_7374,N_7085,N_7026);
or U7375 (N_7375,N_7067,N_7095);
xnor U7376 (N_7376,N_7071,N_7199);
and U7377 (N_7377,N_7184,N_7221);
nor U7378 (N_7378,N_7194,N_7211);
and U7379 (N_7379,N_7141,N_7061);
nor U7380 (N_7380,N_7080,N_7068);
xnor U7381 (N_7381,N_7144,N_7231);
xor U7382 (N_7382,N_7189,N_7226);
xor U7383 (N_7383,N_7088,N_7160);
or U7384 (N_7384,N_7124,N_7110);
nor U7385 (N_7385,N_7204,N_7058);
or U7386 (N_7386,N_7138,N_7166);
xnor U7387 (N_7387,N_7088,N_7073);
xnor U7388 (N_7388,N_7161,N_7170);
xnor U7389 (N_7389,N_7248,N_7238);
or U7390 (N_7390,N_7182,N_7042);
xor U7391 (N_7391,N_7090,N_7087);
and U7392 (N_7392,N_7196,N_7144);
xor U7393 (N_7393,N_7147,N_7097);
and U7394 (N_7394,N_7075,N_7045);
nand U7395 (N_7395,N_7212,N_7073);
nor U7396 (N_7396,N_7132,N_7203);
nor U7397 (N_7397,N_7166,N_7120);
or U7398 (N_7398,N_7052,N_7067);
nor U7399 (N_7399,N_7074,N_7245);
nand U7400 (N_7400,N_7155,N_7013);
nand U7401 (N_7401,N_7062,N_7205);
xor U7402 (N_7402,N_7148,N_7211);
nor U7403 (N_7403,N_7072,N_7247);
nand U7404 (N_7404,N_7176,N_7139);
nor U7405 (N_7405,N_7180,N_7068);
xor U7406 (N_7406,N_7162,N_7087);
and U7407 (N_7407,N_7119,N_7003);
nand U7408 (N_7408,N_7169,N_7145);
xnor U7409 (N_7409,N_7193,N_7154);
nand U7410 (N_7410,N_7138,N_7064);
nand U7411 (N_7411,N_7098,N_7132);
and U7412 (N_7412,N_7057,N_7184);
xor U7413 (N_7413,N_7145,N_7007);
nor U7414 (N_7414,N_7238,N_7237);
nor U7415 (N_7415,N_7195,N_7245);
xnor U7416 (N_7416,N_7109,N_7060);
xnor U7417 (N_7417,N_7035,N_7217);
or U7418 (N_7418,N_7038,N_7201);
or U7419 (N_7419,N_7239,N_7243);
and U7420 (N_7420,N_7055,N_7076);
nand U7421 (N_7421,N_7072,N_7014);
nand U7422 (N_7422,N_7246,N_7179);
xnor U7423 (N_7423,N_7084,N_7093);
nand U7424 (N_7424,N_7085,N_7170);
nand U7425 (N_7425,N_7079,N_7124);
and U7426 (N_7426,N_7230,N_7123);
nand U7427 (N_7427,N_7098,N_7203);
xor U7428 (N_7428,N_7207,N_7086);
and U7429 (N_7429,N_7133,N_7197);
or U7430 (N_7430,N_7130,N_7246);
xor U7431 (N_7431,N_7139,N_7071);
and U7432 (N_7432,N_7115,N_7048);
or U7433 (N_7433,N_7020,N_7095);
nand U7434 (N_7434,N_7170,N_7191);
nor U7435 (N_7435,N_7027,N_7231);
nand U7436 (N_7436,N_7180,N_7130);
xor U7437 (N_7437,N_7007,N_7140);
and U7438 (N_7438,N_7198,N_7244);
nand U7439 (N_7439,N_7177,N_7240);
nand U7440 (N_7440,N_7116,N_7083);
or U7441 (N_7441,N_7141,N_7193);
and U7442 (N_7442,N_7027,N_7236);
and U7443 (N_7443,N_7120,N_7159);
nor U7444 (N_7444,N_7165,N_7141);
nor U7445 (N_7445,N_7163,N_7090);
and U7446 (N_7446,N_7146,N_7046);
xnor U7447 (N_7447,N_7230,N_7016);
nor U7448 (N_7448,N_7201,N_7213);
xor U7449 (N_7449,N_7156,N_7070);
or U7450 (N_7450,N_7058,N_7142);
and U7451 (N_7451,N_7142,N_7071);
or U7452 (N_7452,N_7145,N_7178);
or U7453 (N_7453,N_7249,N_7167);
and U7454 (N_7454,N_7123,N_7005);
nor U7455 (N_7455,N_7011,N_7007);
nor U7456 (N_7456,N_7054,N_7036);
nand U7457 (N_7457,N_7047,N_7234);
xnor U7458 (N_7458,N_7066,N_7136);
nor U7459 (N_7459,N_7008,N_7165);
nor U7460 (N_7460,N_7042,N_7121);
and U7461 (N_7461,N_7015,N_7152);
nand U7462 (N_7462,N_7205,N_7188);
nand U7463 (N_7463,N_7027,N_7063);
nor U7464 (N_7464,N_7156,N_7186);
xor U7465 (N_7465,N_7028,N_7226);
or U7466 (N_7466,N_7077,N_7070);
nor U7467 (N_7467,N_7163,N_7152);
or U7468 (N_7468,N_7195,N_7121);
nand U7469 (N_7469,N_7132,N_7126);
and U7470 (N_7470,N_7115,N_7108);
and U7471 (N_7471,N_7203,N_7110);
xnor U7472 (N_7472,N_7049,N_7085);
and U7473 (N_7473,N_7170,N_7240);
nand U7474 (N_7474,N_7015,N_7029);
or U7475 (N_7475,N_7243,N_7051);
xnor U7476 (N_7476,N_7145,N_7249);
xnor U7477 (N_7477,N_7209,N_7226);
xnor U7478 (N_7478,N_7153,N_7129);
nor U7479 (N_7479,N_7188,N_7028);
nor U7480 (N_7480,N_7000,N_7249);
or U7481 (N_7481,N_7139,N_7002);
xor U7482 (N_7482,N_7157,N_7082);
or U7483 (N_7483,N_7207,N_7243);
nor U7484 (N_7484,N_7065,N_7213);
and U7485 (N_7485,N_7120,N_7023);
nand U7486 (N_7486,N_7246,N_7117);
nor U7487 (N_7487,N_7027,N_7038);
nor U7488 (N_7488,N_7004,N_7236);
or U7489 (N_7489,N_7206,N_7103);
xnor U7490 (N_7490,N_7093,N_7120);
or U7491 (N_7491,N_7204,N_7136);
xor U7492 (N_7492,N_7062,N_7181);
and U7493 (N_7493,N_7152,N_7119);
xnor U7494 (N_7494,N_7133,N_7013);
and U7495 (N_7495,N_7191,N_7105);
nor U7496 (N_7496,N_7088,N_7051);
and U7497 (N_7497,N_7044,N_7171);
nand U7498 (N_7498,N_7152,N_7226);
nor U7499 (N_7499,N_7128,N_7005);
nor U7500 (N_7500,N_7492,N_7443);
and U7501 (N_7501,N_7439,N_7496);
xor U7502 (N_7502,N_7275,N_7335);
or U7503 (N_7503,N_7449,N_7351);
nor U7504 (N_7504,N_7280,N_7299);
xnor U7505 (N_7505,N_7352,N_7254);
nor U7506 (N_7506,N_7295,N_7377);
xnor U7507 (N_7507,N_7257,N_7328);
nor U7508 (N_7508,N_7376,N_7316);
or U7509 (N_7509,N_7445,N_7264);
and U7510 (N_7510,N_7251,N_7314);
and U7511 (N_7511,N_7262,N_7488);
nor U7512 (N_7512,N_7296,N_7321);
and U7513 (N_7513,N_7372,N_7491);
xor U7514 (N_7514,N_7386,N_7398);
nand U7515 (N_7515,N_7484,N_7287);
nand U7516 (N_7516,N_7320,N_7361);
or U7517 (N_7517,N_7409,N_7451);
nand U7518 (N_7518,N_7252,N_7349);
nor U7519 (N_7519,N_7271,N_7390);
or U7520 (N_7520,N_7489,N_7283);
or U7521 (N_7521,N_7428,N_7332);
nor U7522 (N_7522,N_7404,N_7456);
nand U7523 (N_7523,N_7460,N_7289);
and U7524 (N_7524,N_7303,N_7294);
nand U7525 (N_7525,N_7273,N_7269);
xor U7526 (N_7526,N_7437,N_7407);
and U7527 (N_7527,N_7319,N_7353);
xnor U7528 (N_7528,N_7309,N_7274);
nand U7529 (N_7529,N_7433,N_7356);
or U7530 (N_7530,N_7301,N_7438);
or U7531 (N_7531,N_7360,N_7440);
nand U7532 (N_7532,N_7276,N_7410);
and U7533 (N_7533,N_7324,N_7307);
nand U7534 (N_7534,N_7392,N_7461);
nor U7535 (N_7535,N_7282,N_7472);
xor U7536 (N_7536,N_7452,N_7260);
xor U7537 (N_7537,N_7476,N_7285);
xnor U7538 (N_7538,N_7483,N_7375);
nor U7539 (N_7539,N_7340,N_7418);
nor U7540 (N_7540,N_7434,N_7420);
xnor U7541 (N_7541,N_7290,N_7378);
nand U7542 (N_7542,N_7373,N_7387);
and U7543 (N_7543,N_7253,N_7325);
nor U7544 (N_7544,N_7308,N_7453);
xor U7545 (N_7545,N_7477,N_7468);
and U7546 (N_7546,N_7334,N_7388);
or U7547 (N_7547,N_7268,N_7494);
or U7548 (N_7548,N_7442,N_7481);
and U7549 (N_7549,N_7318,N_7354);
nor U7550 (N_7550,N_7322,N_7397);
nor U7551 (N_7551,N_7323,N_7256);
and U7552 (N_7552,N_7463,N_7329);
or U7553 (N_7553,N_7265,N_7368);
xnor U7554 (N_7554,N_7343,N_7408);
nand U7555 (N_7555,N_7411,N_7431);
or U7556 (N_7556,N_7374,N_7315);
nor U7557 (N_7557,N_7297,N_7311);
or U7558 (N_7558,N_7313,N_7288);
or U7559 (N_7559,N_7367,N_7339);
nor U7560 (N_7560,N_7281,N_7417);
or U7561 (N_7561,N_7458,N_7279);
and U7562 (N_7562,N_7277,N_7464);
nand U7563 (N_7563,N_7305,N_7263);
nand U7564 (N_7564,N_7389,N_7346);
and U7565 (N_7565,N_7424,N_7448);
xnor U7566 (N_7566,N_7363,N_7450);
and U7567 (N_7567,N_7487,N_7383);
or U7568 (N_7568,N_7402,N_7365);
and U7569 (N_7569,N_7446,N_7421);
nand U7570 (N_7570,N_7435,N_7401);
nor U7571 (N_7571,N_7490,N_7393);
or U7572 (N_7572,N_7459,N_7330);
or U7573 (N_7573,N_7406,N_7419);
xor U7574 (N_7574,N_7358,N_7357);
nor U7575 (N_7575,N_7344,N_7485);
nand U7576 (N_7576,N_7465,N_7403);
nor U7577 (N_7577,N_7486,N_7272);
nand U7578 (N_7578,N_7259,N_7342);
and U7579 (N_7579,N_7258,N_7336);
xor U7580 (N_7580,N_7391,N_7382);
nand U7581 (N_7581,N_7471,N_7326);
xor U7582 (N_7582,N_7345,N_7474);
and U7583 (N_7583,N_7454,N_7470);
and U7584 (N_7584,N_7473,N_7350);
and U7585 (N_7585,N_7466,N_7348);
or U7586 (N_7586,N_7480,N_7310);
nor U7587 (N_7587,N_7317,N_7385);
or U7588 (N_7588,N_7412,N_7298);
xor U7589 (N_7589,N_7455,N_7429);
nor U7590 (N_7590,N_7384,N_7413);
xnor U7591 (N_7591,N_7270,N_7284);
or U7592 (N_7592,N_7306,N_7359);
xor U7593 (N_7593,N_7379,N_7300);
or U7594 (N_7594,N_7366,N_7493);
and U7595 (N_7595,N_7278,N_7415);
xor U7596 (N_7596,N_7371,N_7399);
xor U7597 (N_7597,N_7400,N_7462);
or U7598 (N_7598,N_7497,N_7396);
xor U7599 (N_7599,N_7261,N_7355);
nor U7600 (N_7600,N_7302,N_7380);
xnor U7601 (N_7601,N_7250,N_7312);
nor U7602 (N_7602,N_7479,N_7495);
nand U7603 (N_7603,N_7416,N_7405);
or U7604 (N_7604,N_7347,N_7304);
and U7605 (N_7605,N_7364,N_7430);
xor U7606 (N_7606,N_7370,N_7291);
nand U7607 (N_7607,N_7436,N_7394);
and U7608 (N_7608,N_7498,N_7292);
and U7609 (N_7609,N_7381,N_7341);
nand U7610 (N_7610,N_7427,N_7255);
and U7611 (N_7611,N_7293,N_7432);
nor U7612 (N_7612,N_7457,N_7337);
nand U7613 (N_7613,N_7266,N_7362);
or U7614 (N_7614,N_7369,N_7478);
nand U7615 (N_7615,N_7441,N_7422);
and U7616 (N_7616,N_7327,N_7423);
nor U7617 (N_7617,N_7447,N_7444);
or U7618 (N_7618,N_7267,N_7425);
or U7619 (N_7619,N_7426,N_7414);
nor U7620 (N_7620,N_7395,N_7331);
nand U7621 (N_7621,N_7333,N_7469);
or U7622 (N_7622,N_7475,N_7499);
and U7623 (N_7623,N_7286,N_7482);
and U7624 (N_7624,N_7338,N_7467);
nor U7625 (N_7625,N_7498,N_7300);
and U7626 (N_7626,N_7334,N_7403);
xnor U7627 (N_7627,N_7257,N_7426);
nor U7628 (N_7628,N_7271,N_7292);
nand U7629 (N_7629,N_7317,N_7386);
and U7630 (N_7630,N_7451,N_7446);
and U7631 (N_7631,N_7334,N_7494);
and U7632 (N_7632,N_7458,N_7492);
nand U7633 (N_7633,N_7327,N_7364);
and U7634 (N_7634,N_7475,N_7440);
or U7635 (N_7635,N_7330,N_7416);
and U7636 (N_7636,N_7494,N_7276);
nand U7637 (N_7637,N_7393,N_7423);
or U7638 (N_7638,N_7313,N_7325);
and U7639 (N_7639,N_7288,N_7289);
nand U7640 (N_7640,N_7499,N_7366);
nand U7641 (N_7641,N_7274,N_7473);
or U7642 (N_7642,N_7378,N_7448);
xnor U7643 (N_7643,N_7325,N_7294);
and U7644 (N_7644,N_7319,N_7399);
nor U7645 (N_7645,N_7323,N_7250);
and U7646 (N_7646,N_7478,N_7362);
and U7647 (N_7647,N_7306,N_7282);
and U7648 (N_7648,N_7446,N_7274);
and U7649 (N_7649,N_7380,N_7315);
nand U7650 (N_7650,N_7367,N_7484);
and U7651 (N_7651,N_7485,N_7253);
or U7652 (N_7652,N_7254,N_7485);
and U7653 (N_7653,N_7443,N_7456);
or U7654 (N_7654,N_7485,N_7466);
nor U7655 (N_7655,N_7269,N_7474);
and U7656 (N_7656,N_7402,N_7358);
or U7657 (N_7657,N_7290,N_7491);
xor U7658 (N_7658,N_7349,N_7368);
xnor U7659 (N_7659,N_7370,N_7340);
or U7660 (N_7660,N_7397,N_7413);
and U7661 (N_7661,N_7431,N_7370);
xor U7662 (N_7662,N_7343,N_7288);
xnor U7663 (N_7663,N_7377,N_7252);
or U7664 (N_7664,N_7293,N_7263);
xnor U7665 (N_7665,N_7328,N_7426);
and U7666 (N_7666,N_7450,N_7485);
or U7667 (N_7667,N_7339,N_7490);
or U7668 (N_7668,N_7288,N_7279);
nor U7669 (N_7669,N_7499,N_7368);
xor U7670 (N_7670,N_7399,N_7481);
nand U7671 (N_7671,N_7261,N_7353);
or U7672 (N_7672,N_7465,N_7413);
xor U7673 (N_7673,N_7480,N_7264);
nand U7674 (N_7674,N_7390,N_7410);
xor U7675 (N_7675,N_7345,N_7435);
nand U7676 (N_7676,N_7468,N_7320);
and U7677 (N_7677,N_7427,N_7394);
nand U7678 (N_7678,N_7471,N_7295);
xor U7679 (N_7679,N_7468,N_7258);
xnor U7680 (N_7680,N_7421,N_7288);
or U7681 (N_7681,N_7464,N_7291);
nand U7682 (N_7682,N_7323,N_7308);
and U7683 (N_7683,N_7319,N_7437);
xnor U7684 (N_7684,N_7394,N_7345);
and U7685 (N_7685,N_7419,N_7269);
or U7686 (N_7686,N_7398,N_7448);
and U7687 (N_7687,N_7277,N_7431);
and U7688 (N_7688,N_7492,N_7394);
nor U7689 (N_7689,N_7279,N_7290);
nand U7690 (N_7690,N_7259,N_7447);
xnor U7691 (N_7691,N_7438,N_7360);
xor U7692 (N_7692,N_7430,N_7392);
nor U7693 (N_7693,N_7292,N_7463);
nor U7694 (N_7694,N_7266,N_7453);
and U7695 (N_7695,N_7364,N_7356);
xor U7696 (N_7696,N_7461,N_7252);
and U7697 (N_7697,N_7339,N_7434);
and U7698 (N_7698,N_7278,N_7353);
and U7699 (N_7699,N_7437,N_7395);
xnor U7700 (N_7700,N_7452,N_7303);
xor U7701 (N_7701,N_7277,N_7272);
and U7702 (N_7702,N_7453,N_7267);
nor U7703 (N_7703,N_7300,N_7389);
nor U7704 (N_7704,N_7408,N_7482);
nand U7705 (N_7705,N_7491,N_7292);
nor U7706 (N_7706,N_7403,N_7456);
or U7707 (N_7707,N_7362,N_7448);
and U7708 (N_7708,N_7333,N_7312);
xnor U7709 (N_7709,N_7350,N_7330);
and U7710 (N_7710,N_7336,N_7261);
nand U7711 (N_7711,N_7477,N_7275);
xnor U7712 (N_7712,N_7433,N_7393);
nor U7713 (N_7713,N_7308,N_7388);
nor U7714 (N_7714,N_7365,N_7288);
nor U7715 (N_7715,N_7372,N_7257);
nor U7716 (N_7716,N_7281,N_7283);
nor U7717 (N_7717,N_7402,N_7476);
nor U7718 (N_7718,N_7361,N_7403);
and U7719 (N_7719,N_7269,N_7342);
xnor U7720 (N_7720,N_7412,N_7492);
and U7721 (N_7721,N_7474,N_7372);
nor U7722 (N_7722,N_7262,N_7370);
or U7723 (N_7723,N_7487,N_7494);
nand U7724 (N_7724,N_7495,N_7427);
nor U7725 (N_7725,N_7418,N_7495);
xor U7726 (N_7726,N_7335,N_7263);
and U7727 (N_7727,N_7379,N_7465);
or U7728 (N_7728,N_7250,N_7342);
xnor U7729 (N_7729,N_7475,N_7409);
or U7730 (N_7730,N_7253,N_7270);
nand U7731 (N_7731,N_7395,N_7450);
xor U7732 (N_7732,N_7492,N_7280);
xnor U7733 (N_7733,N_7388,N_7303);
or U7734 (N_7734,N_7387,N_7287);
xor U7735 (N_7735,N_7453,N_7333);
nor U7736 (N_7736,N_7468,N_7481);
or U7737 (N_7737,N_7354,N_7277);
nand U7738 (N_7738,N_7297,N_7414);
xnor U7739 (N_7739,N_7344,N_7367);
xnor U7740 (N_7740,N_7366,N_7383);
xor U7741 (N_7741,N_7469,N_7402);
or U7742 (N_7742,N_7394,N_7499);
xnor U7743 (N_7743,N_7258,N_7420);
xor U7744 (N_7744,N_7317,N_7483);
or U7745 (N_7745,N_7371,N_7308);
and U7746 (N_7746,N_7490,N_7351);
nand U7747 (N_7747,N_7396,N_7329);
nor U7748 (N_7748,N_7431,N_7401);
nand U7749 (N_7749,N_7459,N_7390);
nor U7750 (N_7750,N_7508,N_7653);
or U7751 (N_7751,N_7741,N_7634);
xor U7752 (N_7752,N_7579,N_7600);
nor U7753 (N_7753,N_7660,N_7694);
or U7754 (N_7754,N_7528,N_7604);
nor U7755 (N_7755,N_7509,N_7716);
nor U7756 (N_7756,N_7587,N_7501);
or U7757 (N_7757,N_7519,N_7710);
or U7758 (N_7758,N_7621,N_7623);
xor U7759 (N_7759,N_7591,N_7713);
or U7760 (N_7760,N_7651,N_7636);
nand U7761 (N_7761,N_7675,N_7539);
xor U7762 (N_7762,N_7613,N_7569);
or U7763 (N_7763,N_7626,N_7719);
nand U7764 (N_7764,N_7622,N_7659);
nand U7765 (N_7765,N_7732,N_7730);
nor U7766 (N_7766,N_7693,N_7689);
and U7767 (N_7767,N_7520,N_7566);
or U7768 (N_7768,N_7684,N_7647);
nor U7769 (N_7769,N_7688,N_7642);
or U7770 (N_7770,N_7705,N_7568);
nand U7771 (N_7771,N_7500,N_7745);
nand U7772 (N_7772,N_7633,N_7582);
or U7773 (N_7773,N_7690,N_7644);
nor U7774 (N_7774,N_7707,N_7607);
nand U7775 (N_7775,N_7529,N_7665);
nor U7776 (N_7776,N_7672,N_7619);
or U7777 (N_7777,N_7699,N_7679);
xnor U7778 (N_7778,N_7525,N_7590);
nor U7779 (N_7779,N_7744,N_7532);
xor U7780 (N_7780,N_7577,N_7718);
and U7781 (N_7781,N_7656,N_7541);
nand U7782 (N_7782,N_7724,N_7668);
nor U7783 (N_7783,N_7740,N_7534);
and U7784 (N_7784,N_7543,N_7542);
and U7785 (N_7785,N_7637,N_7686);
nand U7786 (N_7786,N_7734,N_7558);
xor U7787 (N_7787,N_7666,N_7748);
or U7788 (N_7788,N_7583,N_7655);
and U7789 (N_7789,N_7547,N_7551);
or U7790 (N_7790,N_7669,N_7620);
and U7791 (N_7791,N_7511,N_7612);
nand U7792 (N_7792,N_7564,N_7595);
nand U7793 (N_7793,N_7517,N_7578);
or U7794 (N_7794,N_7737,N_7504);
or U7795 (N_7795,N_7720,N_7611);
and U7796 (N_7796,N_7625,N_7527);
nand U7797 (N_7797,N_7536,N_7585);
xor U7798 (N_7798,N_7738,N_7557);
nand U7799 (N_7799,N_7700,N_7503);
nor U7800 (N_7800,N_7550,N_7567);
nor U7801 (N_7801,N_7714,N_7616);
xnor U7802 (N_7802,N_7725,N_7721);
and U7803 (N_7803,N_7728,N_7681);
xor U7804 (N_7804,N_7584,N_7507);
xnor U7805 (N_7805,N_7592,N_7601);
nand U7806 (N_7806,N_7629,N_7606);
nor U7807 (N_7807,N_7524,N_7698);
nor U7808 (N_7808,N_7530,N_7513);
and U7809 (N_7809,N_7664,N_7514);
or U7810 (N_7810,N_7602,N_7533);
or U7811 (N_7811,N_7537,N_7657);
and U7812 (N_7812,N_7739,N_7512);
nor U7813 (N_7813,N_7749,N_7597);
xnor U7814 (N_7814,N_7617,N_7631);
nor U7815 (N_7815,N_7560,N_7711);
or U7816 (N_7816,N_7701,N_7522);
and U7817 (N_7817,N_7575,N_7561);
nor U7818 (N_7818,N_7593,N_7505);
xor U7819 (N_7819,N_7540,N_7704);
and U7820 (N_7820,N_7695,N_7735);
nand U7821 (N_7821,N_7717,N_7729);
xor U7822 (N_7822,N_7702,N_7731);
nand U7823 (N_7823,N_7652,N_7608);
and U7824 (N_7824,N_7639,N_7663);
xnor U7825 (N_7825,N_7538,N_7683);
xnor U7826 (N_7826,N_7654,N_7706);
or U7827 (N_7827,N_7521,N_7516);
xor U7828 (N_7828,N_7552,N_7649);
and U7829 (N_7829,N_7555,N_7630);
nand U7830 (N_7830,N_7742,N_7697);
nand U7831 (N_7831,N_7682,N_7571);
or U7832 (N_7832,N_7546,N_7615);
or U7833 (N_7833,N_7589,N_7596);
or U7834 (N_7834,N_7570,N_7641);
nor U7835 (N_7835,N_7722,N_7586);
or U7836 (N_7836,N_7662,N_7610);
nand U7837 (N_7837,N_7559,N_7609);
xnor U7838 (N_7838,N_7573,N_7526);
nand U7839 (N_7839,N_7632,N_7523);
nor U7840 (N_7840,N_7671,N_7554);
or U7841 (N_7841,N_7556,N_7650);
nor U7842 (N_7842,N_7549,N_7605);
xor U7843 (N_7843,N_7726,N_7747);
nand U7844 (N_7844,N_7618,N_7581);
or U7845 (N_7845,N_7628,N_7677);
nor U7846 (N_7846,N_7614,N_7598);
nor U7847 (N_7847,N_7658,N_7643);
xnor U7848 (N_7848,N_7680,N_7510);
or U7849 (N_7849,N_7535,N_7599);
xnor U7850 (N_7850,N_7574,N_7506);
xor U7851 (N_7851,N_7661,N_7580);
or U7852 (N_7852,N_7563,N_7723);
nor U7853 (N_7853,N_7667,N_7624);
nand U7854 (N_7854,N_7572,N_7708);
xnor U7855 (N_7855,N_7635,N_7638);
and U7856 (N_7856,N_7648,N_7545);
nand U7857 (N_7857,N_7548,N_7553);
or U7858 (N_7858,N_7692,N_7691);
nor U7859 (N_7859,N_7703,N_7727);
xor U7860 (N_7860,N_7544,N_7674);
xnor U7861 (N_7861,N_7646,N_7576);
and U7862 (N_7862,N_7670,N_7640);
nor U7863 (N_7863,N_7685,N_7594);
nand U7864 (N_7864,N_7518,N_7736);
xor U7865 (N_7865,N_7743,N_7645);
xor U7866 (N_7866,N_7603,N_7588);
nand U7867 (N_7867,N_7676,N_7565);
nand U7868 (N_7868,N_7696,N_7531);
nor U7869 (N_7869,N_7678,N_7709);
xnor U7870 (N_7870,N_7515,N_7502);
and U7871 (N_7871,N_7712,N_7746);
xor U7872 (N_7872,N_7733,N_7715);
or U7873 (N_7873,N_7562,N_7673);
nor U7874 (N_7874,N_7687,N_7627);
nand U7875 (N_7875,N_7730,N_7594);
nor U7876 (N_7876,N_7550,N_7658);
or U7877 (N_7877,N_7739,N_7647);
xor U7878 (N_7878,N_7565,N_7693);
or U7879 (N_7879,N_7549,N_7687);
nor U7880 (N_7880,N_7519,N_7559);
nor U7881 (N_7881,N_7557,N_7674);
and U7882 (N_7882,N_7540,N_7572);
xnor U7883 (N_7883,N_7602,N_7507);
xnor U7884 (N_7884,N_7735,N_7597);
nor U7885 (N_7885,N_7740,N_7552);
and U7886 (N_7886,N_7646,N_7681);
nand U7887 (N_7887,N_7699,N_7630);
nand U7888 (N_7888,N_7678,N_7667);
nor U7889 (N_7889,N_7523,N_7733);
and U7890 (N_7890,N_7620,N_7659);
or U7891 (N_7891,N_7609,N_7654);
xor U7892 (N_7892,N_7615,N_7541);
nand U7893 (N_7893,N_7674,N_7519);
xor U7894 (N_7894,N_7652,N_7659);
xnor U7895 (N_7895,N_7633,N_7730);
xor U7896 (N_7896,N_7704,N_7502);
xnor U7897 (N_7897,N_7685,N_7535);
and U7898 (N_7898,N_7653,N_7562);
and U7899 (N_7899,N_7634,N_7643);
xor U7900 (N_7900,N_7620,N_7513);
nand U7901 (N_7901,N_7617,N_7719);
nor U7902 (N_7902,N_7694,N_7662);
or U7903 (N_7903,N_7679,N_7693);
nand U7904 (N_7904,N_7729,N_7633);
nand U7905 (N_7905,N_7520,N_7584);
nand U7906 (N_7906,N_7728,N_7517);
xnor U7907 (N_7907,N_7607,N_7718);
xnor U7908 (N_7908,N_7746,N_7593);
and U7909 (N_7909,N_7654,N_7748);
or U7910 (N_7910,N_7748,N_7527);
and U7911 (N_7911,N_7612,N_7518);
nor U7912 (N_7912,N_7664,N_7571);
xnor U7913 (N_7913,N_7594,N_7508);
or U7914 (N_7914,N_7714,N_7565);
and U7915 (N_7915,N_7662,N_7586);
nand U7916 (N_7916,N_7645,N_7735);
nand U7917 (N_7917,N_7510,N_7595);
or U7918 (N_7918,N_7552,N_7671);
or U7919 (N_7919,N_7614,N_7721);
and U7920 (N_7920,N_7742,N_7653);
or U7921 (N_7921,N_7579,N_7737);
nor U7922 (N_7922,N_7696,N_7592);
and U7923 (N_7923,N_7508,N_7718);
nand U7924 (N_7924,N_7559,N_7641);
and U7925 (N_7925,N_7669,N_7626);
or U7926 (N_7926,N_7611,N_7710);
xor U7927 (N_7927,N_7565,N_7709);
xor U7928 (N_7928,N_7567,N_7686);
nor U7929 (N_7929,N_7715,N_7554);
nor U7930 (N_7930,N_7731,N_7501);
and U7931 (N_7931,N_7641,N_7530);
xor U7932 (N_7932,N_7580,N_7639);
nand U7933 (N_7933,N_7686,N_7526);
or U7934 (N_7934,N_7502,N_7604);
xor U7935 (N_7935,N_7678,N_7613);
nor U7936 (N_7936,N_7645,N_7572);
xor U7937 (N_7937,N_7723,N_7661);
xor U7938 (N_7938,N_7515,N_7660);
and U7939 (N_7939,N_7644,N_7620);
or U7940 (N_7940,N_7562,N_7511);
xnor U7941 (N_7941,N_7624,N_7512);
nor U7942 (N_7942,N_7555,N_7536);
nor U7943 (N_7943,N_7635,N_7664);
xnor U7944 (N_7944,N_7709,N_7520);
xor U7945 (N_7945,N_7668,N_7543);
nor U7946 (N_7946,N_7730,N_7576);
nor U7947 (N_7947,N_7503,N_7720);
and U7948 (N_7948,N_7592,N_7726);
nand U7949 (N_7949,N_7684,N_7539);
or U7950 (N_7950,N_7511,N_7729);
nand U7951 (N_7951,N_7591,N_7553);
nor U7952 (N_7952,N_7667,N_7708);
or U7953 (N_7953,N_7729,N_7708);
nand U7954 (N_7954,N_7602,N_7582);
xor U7955 (N_7955,N_7500,N_7681);
and U7956 (N_7956,N_7724,N_7721);
xnor U7957 (N_7957,N_7730,N_7703);
and U7958 (N_7958,N_7678,N_7532);
or U7959 (N_7959,N_7548,N_7720);
or U7960 (N_7960,N_7660,N_7564);
and U7961 (N_7961,N_7683,N_7511);
nor U7962 (N_7962,N_7500,N_7525);
xnor U7963 (N_7963,N_7683,N_7728);
nor U7964 (N_7964,N_7694,N_7565);
nor U7965 (N_7965,N_7644,N_7694);
xor U7966 (N_7966,N_7743,N_7615);
and U7967 (N_7967,N_7600,N_7667);
nand U7968 (N_7968,N_7513,N_7517);
or U7969 (N_7969,N_7708,N_7589);
nand U7970 (N_7970,N_7508,N_7714);
and U7971 (N_7971,N_7717,N_7593);
or U7972 (N_7972,N_7727,N_7505);
nand U7973 (N_7973,N_7569,N_7608);
and U7974 (N_7974,N_7601,N_7556);
or U7975 (N_7975,N_7593,N_7736);
xor U7976 (N_7976,N_7721,N_7531);
and U7977 (N_7977,N_7703,N_7624);
or U7978 (N_7978,N_7676,N_7516);
xnor U7979 (N_7979,N_7520,N_7646);
nand U7980 (N_7980,N_7669,N_7681);
xor U7981 (N_7981,N_7513,N_7648);
nor U7982 (N_7982,N_7573,N_7664);
or U7983 (N_7983,N_7572,N_7672);
nor U7984 (N_7984,N_7673,N_7629);
xor U7985 (N_7985,N_7719,N_7502);
nand U7986 (N_7986,N_7534,N_7525);
xnor U7987 (N_7987,N_7748,N_7736);
nor U7988 (N_7988,N_7699,N_7733);
xnor U7989 (N_7989,N_7732,N_7724);
nor U7990 (N_7990,N_7509,N_7682);
nand U7991 (N_7991,N_7659,N_7514);
xnor U7992 (N_7992,N_7683,N_7589);
nand U7993 (N_7993,N_7646,N_7599);
nor U7994 (N_7994,N_7700,N_7623);
and U7995 (N_7995,N_7625,N_7600);
and U7996 (N_7996,N_7654,N_7731);
or U7997 (N_7997,N_7553,N_7682);
or U7998 (N_7998,N_7636,N_7580);
or U7999 (N_7999,N_7658,N_7739);
or U8000 (N_8000,N_7843,N_7867);
and U8001 (N_8001,N_7979,N_7857);
xnor U8002 (N_8002,N_7800,N_7769);
or U8003 (N_8003,N_7931,N_7865);
and U8004 (N_8004,N_7901,N_7791);
and U8005 (N_8005,N_7951,N_7798);
nor U8006 (N_8006,N_7909,N_7773);
nand U8007 (N_8007,N_7897,N_7835);
nor U8008 (N_8008,N_7993,N_7795);
or U8009 (N_8009,N_7772,N_7997);
xor U8010 (N_8010,N_7853,N_7977);
and U8011 (N_8011,N_7988,N_7986);
nand U8012 (N_8012,N_7811,N_7994);
or U8013 (N_8013,N_7809,N_7814);
and U8014 (N_8014,N_7796,N_7849);
or U8015 (N_8015,N_7904,N_7771);
xor U8016 (N_8016,N_7870,N_7875);
and U8017 (N_8017,N_7783,N_7834);
and U8018 (N_8018,N_7836,N_7964);
and U8019 (N_8019,N_7837,N_7912);
and U8020 (N_8020,N_7876,N_7813);
nor U8021 (N_8021,N_7871,N_7942);
or U8022 (N_8022,N_7840,N_7957);
and U8023 (N_8023,N_7845,N_7943);
nor U8024 (N_8024,N_7950,N_7919);
and U8025 (N_8025,N_7763,N_7767);
and U8026 (N_8026,N_7802,N_7799);
and U8027 (N_8027,N_7898,N_7778);
nand U8028 (N_8028,N_7818,N_7883);
and U8029 (N_8029,N_7900,N_7775);
and U8030 (N_8030,N_7996,N_7765);
and U8031 (N_8031,N_7963,N_7753);
and U8032 (N_8032,N_7970,N_7754);
or U8033 (N_8033,N_7862,N_7922);
and U8034 (N_8034,N_7838,N_7820);
nor U8035 (N_8035,N_7945,N_7929);
nor U8036 (N_8036,N_7946,N_7873);
nand U8037 (N_8037,N_7864,N_7866);
xnor U8038 (N_8038,N_7930,N_7887);
nand U8039 (N_8039,N_7882,N_7751);
xnor U8040 (N_8040,N_7955,N_7804);
nor U8041 (N_8041,N_7832,N_7850);
or U8042 (N_8042,N_7868,N_7932);
nor U8043 (N_8043,N_7907,N_7856);
and U8044 (N_8044,N_7768,N_7935);
nand U8045 (N_8045,N_7911,N_7817);
xor U8046 (N_8046,N_7992,N_7842);
xnor U8047 (N_8047,N_7894,N_7939);
and U8048 (N_8048,N_7784,N_7891);
nor U8049 (N_8049,N_7937,N_7782);
xor U8050 (N_8050,N_7831,N_7859);
xnor U8051 (N_8051,N_7833,N_7756);
or U8052 (N_8052,N_7969,N_7777);
and U8053 (N_8053,N_7889,N_7913);
nor U8054 (N_8054,N_7830,N_7899);
nor U8055 (N_8055,N_7967,N_7790);
or U8056 (N_8056,N_7801,N_7954);
nor U8057 (N_8057,N_7948,N_7910);
nand U8058 (N_8058,N_7826,N_7956);
or U8059 (N_8059,N_7808,N_7982);
and U8060 (N_8060,N_7884,N_7947);
and U8061 (N_8061,N_7863,N_7774);
nand U8062 (N_8062,N_7750,N_7781);
nor U8063 (N_8063,N_7881,N_7788);
xnor U8064 (N_8064,N_7908,N_7807);
or U8065 (N_8065,N_7819,N_7823);
nand U8066 (N_8066,N_7987,N_7878);
and U8067 (N_8067,N_7825,N_7880);
and U8068 (N_8068,N_7905,N_7933);
or U8069 (N_8069,N_7760,N_7961);
and U8070 (N_8070,N_7812,N_7851);
or U8071 (N_8071,N_7816,N_7789);
and U8072 (N_8072,N_7803,N_7786);
and U8073 (N_8073,N_7938,N_7787);
and U8074 (N_8074,N_7861,N_7949);
nand U8075 (N_8075,N_7779,N_7770);
xnor U8076 (N_8076,N_7995,N_7761);
nand U8077 (N_8077,N_7903,N_7920);
and U8078 (N_8078,N_7879,N_7810);
nor U8079 (N_8079,N_7981,N_7978);
nor U8080 (N_8080,N_7959,N_7998);
nand U8081 (N_8081,N_7855,N_7915);
xor U8082 (N_8082,N_7968,N_7973);
xnor U8083 (N_8083,N_7766,N_7828);
nor U8084 (N_8084,N_7827,N_7764);
nor U8085 (N_8085,N_7852,N_7794);
xnor U8086 (N_8086,N_7877,N_7983);
xor U8087 (N_8087,N_7759,N_7934);
and U8088 (N_8088,N_7928,N_7846);
nor U8089 (N_8089,N_7966,N_7960);
nor U8090 (N_8090,N_7940,N_7829);
nor U8091 (N_8091,N_7985,N_7841);
nand U8092 (N_8092,N_7780,N_7971);
nor U8093 (N_8093,N_7989,N_7975);
nand U8094 (N_8094,N_7902,N_7785);
nand U8095 (N_8095,N_7792,N_7872);
and U8096 (N_8096,N_7848,N_7762);
nor U8097 (N_8097,N_7874,N_7923);
and U8098 (N_8098,N_7847,N_7793);
nor U8099 (N_8099,N_7944,N_7974);
and U8100 (N_8100,N_7844,N_7917);
or U8101 (N_8101,N_7805,N_7984);
and U8102 (N_8102,N_7888,N_7755);
nand U8103 (N_8103,N_7965,N_7927);
and U8104 (N_8104,N_7918,N_7962);
nand U8105 (N_8105,N_7952,N_7980);
and U8106 (N_8106,N_7924,N_7886);
and U8107 (N_8107,N_7941,N_7892);
or U8108 (N_8108,N_7869,N_7776);
and U8109 (N_8109,N_7916,N_7953);
or U8110 (N_8110,N_7958,N_7921);
nor U8111 (N_8111,N_7914,N_7821);
and U8112 (N_8112,N_7893,N_7815);
xnor U8113 (N_8113,N_7895,N_7824);
or U8114 (N_8114,N_7752,N_7822);
nand U8115 (N_8115,N_7925,N_7860);
and U8116 (N_8116,N_7896,N_7890);
xor U8117 (N_8117,N_7854,N_7976);
nor U8118 (N_8118,N_7757,N_7999);
xnor U8119 (N_8119,N_7797,N_7972);
and U8120 (N_8120,N_7926,N_7990);
nor U8121 (N_8121,N_7936,N_7758);
xor U8122 (N_8122,N_7858,N_7991);
or U8123 (N_8123,N_7885,N_7806);
nor U8124 (N_8124,N_7906,N_7839);
xnor U8125 (N_8125,N_7936,N_7968);
nor U8126 (N_8126,N_7988,N_7915);
nand U8127 (N_8127,N_7780,N_7762);
nand U8128 (N_8128,N_7826,N_7908);
or U8129 (N_8129,N_7950,N_7841);
nand U8130 (N_8130,N_7973,N_7775);
nor U8131 (N_8131,N_7968,N_7920);
nor U8132 (N_8132,N_7822,N_7764);
and U8133 (N_8133,N_7774,N_7880);
and U8134 (N_8134,N_7909,N_7906);
and U8135 (N_8135,N_7790,N_7753);
xnor U8136 (N_8136,N_7860,N_7974);
or U8137 (N_8137,N_7828,N_7790);
xor U8138 (N_8138,N_7784,N_7948);
nor U8139 (N_8139,N_7949,N_7862);
nor U8140 (N_8140,N_7809,N_7980);
nor U8141 (N_8141,N_7927,N_7948);
and U8142 (N_8142,N_7993,N_7983);
or U8143 (N_8143,N_7933,N_7836);
and U8144 (N_8144,N_7854,N_7933);
and U8145 (N_8145,N_7790,N_7806);
and U8146 (N_8146,N_7872,N_7921);
nor U8147 (N_8147,N_7802,N_7830);
or U8148 (N_8148,N_7944,N_7916);
nand U8149 (N_8149,N_7768,N_7939);
nor U8150 (N_8150,N_7813,N_7858);
nand U8151 (N_8151,N_7967,N_7784);
and U8152 (N_8152,N_7849,N_7981);
xor U8153 (N_8153,N_7882,N_7963);
nand U8154 (N_8154,N_7883,N_7853);
and U8155 (N_8155,N_7771,N_7768);
or U8156 (N_8156,N_7768,N_7928);
xor U8157 (N_8157,N_7926,N_7988);
xor U8158 (N_8158,N_7909,N_7943);
or U8159 (N_8159,N_7750,N_7987);
xnor U8160 (N_8160,N_7906,N_7900);
and U8161 (N_8161,N_7955,N_7794);
nand U8162 (N_8162,N_7910,N_7853);
xor U8163 (N_8163,N_7792,N_7827);
or U8164 (N_8164,N_7891,N_7908);
or U8165 (N_8165,N_7895,N_7876);
or U8166 (N_8166,N_7794,N_7944);
and U8167 (N_8167,N_7870,N_7834);
nand U8168 (N_8168,N_7791,N_7815);
nor U8169 (N_8169,N_7848,N_7948);
xor U8170 (N_8170,N_7826,N_7988);
or U8171 (N_8171,N_7874,N_7917);
xor U8172 (N_8172,N_7764,N_7909);
nor U8173 (N_8173,N_7994,N_7842);
or U8174 (N_8174,N_7956,N_7946);
and U8175 (N_8175,N_7982,N_7889);
and U8176 (N_8176,N_7888,N_7826);
and U8177 (N_8177,N_7809,N_7841);
xor U8178 (N_8178,N_7905,N_7951);
xnor U8179 (N_8179,N_7919,N_7773);
and U8180 (N_8180,N_7779,N_7784);
and U8181 (N_8181,N_7760,N_7777);
nand U8182 (N_8182,N_7972,N_7955);
or U8183 (N_8183,N_7758,N_7850);
or U8184 (N_8184,N_7871,N_7995);
xor U8185 (N_8185,N_7891,N_7758);
and U8186 (N_8186,N_7985,N_7919);
xor U8187 (N_8187,N_7987,N_7849);
nand U8188 (N_8188,N_7967,N_7950);
or U8189 (N_8189,N_7910,N_7806);
xnor U8190 (N_8190,N_7758,N_7837);
xor U8191 (N_8191,N_7783,N_7898);
and U8192 (N_8192,N_7910,N_7846);
xor U8193 (N_8193,N_7780,N_7995);
and U8194 (N_8194,N_7819,N_7906);
or U8195 (N_8195,N_7994,N_7978);
and U8196 (N_8196,N_7828,N_7928);
or U8197 (N_8197,N_7881,N_7822);
nor U8198 (N_8198,N_7897,N_7762);
nand U8199 (N_8199,N_7813,N_7896);
nand U8200 (N_8200,N_7905,N_7949);
nor U8201 (N_8201,N_7761,N_7752);
nand U8202 (N_8202,N_7905,N_7831);
nor U8203 (N_8203,N_7918,N_7932);
nor U8204 (N_8204,N_7774,N_7759);
nor U8205 (N_8205,N_7836,N_7816);
or U8206 (N_8206,N_7851,N_7791);
nor U8207 (N_8207,N_7811,N_7833);
and U8208 (N_8208,N_7808,N_7912);
and U8209 (N_8209,N_7810,N_7987);
and U8210 (N_8210,N_7889,N_7891);
nand U8211 (N_8211,N_7789,N_7882);
nand U8212 (N_8212,N_7772,N_7978);
nor U8213 (N_8213,N_7817,N_7753);
nor U8214 (N_8214,N_7982,N_7937);
nand U8215 (N_8215,N_7849,N_7917);
and U8216 (N_8216,N_7784,N_7780);
nand U8217 (N_8217,N_7824,N_7929);
or U8218 (N_8218,N_7946,N_7829);
and U8219 (N_8219,N_7923,N_7768);
or U8220 (N_8220,N_7933,N_7778);
nor U8221 (N_8221,N_7867,N_7971);
nand U8222 (N_8222,N_7998,N_7904);
nand U8223 (N_8223,N_7889,N_7856);
and U8224 (N_8224,N_7892,N_7911);
nor U8225 (N_8225,N_7805,N_7966);
or U8226 (N_8226,N_7762,N_7784);
nor U8227 (N_8227,N_7771,N_7772);
xor U8228 (N_8228,N_7882,N_7934);
nand U8229 (N_8229,N_7978,N_7790);
xor U8230 (N_8230,N_7997,N_7845);
nand U8231 (N_8231,N_7871,N_7802);
nand U8232 (N_8232,N_7901,N_7786);
and U8233 (N_8233,N_7971,N_7759);
or U8234 (N_8234,N_7979,N_7837);
nand U8235 (N_8235,N_7948,N_7888);
nand U8236 (N_8236,N_7799,N_7916);
or U8237 (N_8237,N_7993,N_7917);
nand U8238 (N_8238,N_7927,N_7895);
nand U8239 (N_8239,N_7839,N_7967);
nor U8240 (N_8240,N_7931,N_7819);
xor U8241 (N_8241,N_7875,N_7857);
or U8242 (N_8242,N_7855,N_7981);
or U8243 (N_8243,N_7839,N_7963);
or U8244 (N_8244,N_7768,N_7927);
nand U8245 (N_8245,N_7872,N_7869);
or U8246 (N_8246,N_7922,N_7850);
xor U8247 (N_8247,N_7994,N_7766);
or U8248 (N_8248,N_7809,N_7959);
or U8249 (N_8249,N_7924,N_7791);
and U8250 (N_8250,N_8206,N_8120);
nand U8251 (N_8251,N_8221,N_8012);
and U8252 (N_8252,N_8238,N_8212);
or U8253 (N_8253,N_8237,N_8224);
nor U8254 (N_8254,N_8200,N_8075);
nor U8255 (N_8255,N_8061,N_8193);
xor U8256 (N_8256,N_8234,N_8108);
nor U8257 (N_8257,N_8197,N_8124);
and U8258 (N_8258,N_8078,N_8008);
and U8259 (N_8259,N_8134,N_8015);
nor U8260 (N_8260,N_8016,N_8140);
xor U8261 (N_8261,N_8100,N_8165);
xnor U8262 (N_8262,N_8035,N_8005);
nor U8263 (N_8263,N_8211,N_8004);
and U8264 (N_8264,N_8045,N_8202);
nor U8265 (N_8265,N_8065,N_8222);
xor U8266 (N_8266,N_8157,N_8204);
or U8267 (N_8267,N_8219,N_8069);
nor U8268 (N_8268,N_8137,N_8166);
and U8269 (N_8269,N_8168,N_8205);
xor U8270 (N_8270,N_8225,N_8087);
nor U8271 (N_8271,N_8125,N_8163);
or U8272 (N_8272,N_8044,N_8024);
nand U8273 (N_8273,N_8018,N_8091);
nand U8274 (N_8274,N_8171,N_8214);
and U8275 (N_8275,N_8092,N_8080);
nand U8276 (N_8276,N_8002,N_8175);
or U8277 (N_8277,N_8119,N_8076);
nand U8278 (N_8278,N_8043,N_8066);
nand U8279 (N_8279,N_8198,N_8046);
or U8280 (N_8280,N_8097,N_8117);
and U8281 (N_8281,N_8006,N_8195);
xnor U8282 (N_8282,N_8031,N_8241);
nand U8283 (N_8283,N_8128,N_8239);
nand U8284 (N_8284,N_8083,N_8235);
nor U8285 (N_8285,N_8010,N_8199);
xor U8286 (N_8286,N_8118,N_8164);
and U8287 (N_8287,N_8074,N_8247);
xnor U8288 (N_8288,N_8077,N_8126);
nand U8289 (N_8289,N_8033,N_8215);
nand U8290 (N_8290,N_8057,N_8052);
and U8291 (N_8291,N_8217,N_8232);
and U8292 (N_8292,N_8155,N_8153);
or U8293 (N_8293,N_8228,N_8220);
nand U8294 (N_8294,N_8019,N_8090);
nor U8295 (N_8295,N_8230,N_8013);
nor U8296 (N_8296,N_8032,N_8151);
or U8297 (N_8297,N_8072,N_8014);
nor U8298 (N_8298,N_8192,N_8114);
xor U8299 (N_8299,N_8067,N_8139);
or U8300 (N_8300,N_8194,N_8007);
and U8301 (N_8301,N_8187,N_8161);
nor U8302 (N_8302,N_8009,N_8079);
or U8303 (N_8303,N_8056,N_8203);
nor U8304 (N_8304,N_8226,N_8047);
nor U8305 (N_8305,N_8174,N_8093);
nand U8306 (N_8306,N_8158,N_8081);
nand U8307 (N_8307,N_8185,N_8243);
or U8308 (N_8308,N_8152,N_8244);
nand U8309 (N_8309,N_8156,N_8180);
xnor U8310 (N_8310,N_8130,N_8233);
or U8311 (N_8311,N_8104,N_8173);
or U8312 (N_8312,N_8089,N_8162);
nand U8313 (N_8313,N_8053,N_8001);
nand U8314 (N_8314,N_8223,N_8142);
nand U8315 (N_8315,N_8169,N_8184);
nand U8316 (N_8316,N_8102,N_8229);
and U8317 (N_8317,N_8101,N_8148);
and U8318 (N_8318,N_8034,N_8105);
and U8319 (N_8319,N_8003,N_8021);
nand U8320 (N_8320,N_8154,N_8096);
xnor U8321 (N_8321,N_8115,N_8048);
nor U8322 (N_8322,N_8133,N_8064);
or U8323 (N_8323,N_8107,N_8136);
or U8324 (N_8324,N_8022,N_8094);
and U8325 (N_8325,N_8240,N_8160);
or U8326 (N_8326,N_8071,N_8138);
and U8327 (N_8327,N_8172,N_8179);
or U8328 (N_8328,N_8000,N_8141);
xor U8329 (N_8329,N_8216,N_8149);
nor U8330 (N_8330,N_8088,N_8189);
and U8331 (N_8331,N_8131,N_8025);
or U8332 (N_8332,N_8054,N_8038);
and U8333 (N_8333,N_8082,N_8248);
and U8334 (N_8334,N_8062,N_8040);
or U8335 (N_8335,N_8042,N_8182);
nor U8336 (N_8336,N_8188,N_8178);
and U8337 (N_8337,N_8030,N_8208);
and U8338 (N_8338,N_8111,N_8236);
or U8339 (N_8339,N_8084,N_8086);
nand U8340 (N_8340,N_8210,N_8041);
nor U8341 (N_8341,N_8143,N_8186);
nor U8342 (N_8342,N_8181,N_8207);
or U8343 (N_8343,N_8249,N_8058);
xnor U8344 (N_8344,N_8113,N_8049);
xnor U8345 (N_8345,N_8196,N_8099);
or U8346 (N_8346,N_8085,N_8147);
nand U8347 (N_8347,N_8146,N_8055);
nand U8348 (N_8348,N_8068,N_8098);
nor U8349 (N_8349,N_8135,N_8170);
nand U8350 (N_8350,N_8011,N_8017);
nand U8351 (N_8351,N_8059,N_8073);
xor U8352 (N_8352,N_8070,N_8027);
xor U8353 (N_8353,N_8121,N_8127);
xnor U8354 (N_8354,N_8109,N_8150);
xnor U8355 (N_8355,N_8218,N_8122);
xnor U8356 (N_8356,N_8242,N_8029);
and U8357 (N_8357,N_8190,N_8132);
or U8358 (N_8358,N_8039,N_8110);
xnor U8359 (N_8359,N_8051,N_8103);
nand U8360 (N_8360,N_8028,N_8063);
and U8361 (N_8361,N_8209,N_8176);
nor U8362 (N_8362,N_8116,N_8112);
or U8363 (N_8363,N_8201,N_8095);
nand U8364 (N_8364,N_8023,N_8145);
or U8365 (N_8365,N_8231,N_8246);
nor U8366 (N_8366,N_8213,N_8177);
nor U8367 (N_8367,N_8060,N_8129);
or U8368 (N_8368,N_8191,N_8144);
or U8369 (N_8369,N_8167,N_8159);
nand U8370 (N_8370,N_8020,N_8183);
xnor U8371 (N_8371,N_8106,N_8227);
or U8372 (N_8372,N_8026,N_8036);
nor U8373 (N_8373,N_8037,N_8245);
xor U8374 (N_8374,N_8123,N_8050);
or U8375 (N_8375,N_8006,N_8220);
xnor U8376 (N_8376,N_8045,N_8210);
nand U8377 (N_8377,N_8007,N_8072);
nor U8378 (N_8378,N_8172,N_8092);
nand U8379 (N_8379,N_8031,N_8128);
or U8380 (N_8380,N_8016,N_8105);
or U8381 (N_8381,N_8087,N_8067);
xor U8382 (N_8382,N_8179,N_8214);
xnor U8383 (N_8383,N_8118,N_8082);
nand U8384 (N_8384,N_8046,N_8078);
nand U8385 (N_8385,N_8244,N_8009);
nand U8386 (N_8386,N_8170,N_8142);
or U8387 (N_8387,N_8192,N_8113);
or U8388 (N_8388,N_8186,N_8155);
or U8389 (N_8389,N_8173,N_8190);
nand U8390 (N_8390,N_8232,N_8184);
or U8391 (N_8391,N_8070,N_8235);
and U8392 (N_8392,N_8166,N_8004);
xor U8393 (N_8393,N_8232,N_8091);
nand U8394 (N_8394,N_8148,N_8001);
or U8395 (N_8395,N_8244,N_8113);
xnor U8396 (N_8396,N_8181,N_8081);
nand U8397 (N_8397,N_8192,N_8240);
nor U8398 (N_8398,N_8227,N_8065);
or U8399 (N_8399,N_8186,N_8079);
nand U8400 (N_8400,N_8082,N_8169);
or U8401 (N_8401,N_8235,N_8146);
xnor U8402 (N_8402,N_8235,N_8194);
nor U8403 (N_8403,N_8193,N_8024);
xor U8404 (N_8404,N_8094,N_8163);
xnor U8405 (N_8405,N_8225,N_8125);
nand U8406 (N_8406,N_8230,N_8112);
xor U8407 (N_8407,N_8087,N_8050);
nor U8408 (N_8408,N_8076,N_8244);
xnor U8409 (N_8409,N_8140,N_8178);
and U8410 (N_8410,N_8099,N_8249);
nor U8411 (N_8411,N_8054,N_8089);
and U8412 (N_8412,N_8105,N_8204);
nor U8413 (N_8413,N_8104,N_8137);
xnor U8414 (N_8414,N_8127,N_8237);
or U8415 (N_8415,N_8143,N_8032);
xnor U8416 (N_8416,N_8143,N_8220);
nor U8417 (N_8417,N_8115,N_8166);
and U8418 (N_8418,N_8232,N_8233);
xnor U8419 (N_8419,N_8185,N_8179);
nand U8420 (N_8420,N_8006,N_8080);
and U8421 (N_8421,N_8064,N_8249);
nand U8422 (N_8422,N_8040,N_8137);
or U8423 (N_8423,N_8124,N_8076);
nor U8424 (N_8424,N_8213,N_8083);
nor U8425 (N_8425,N_8024,N_8186);
or U8426 (N_8426,N_8045,N_8244);
xor U8427 (N_8427,N_8137,N_8060);
nor U8428 (N_8428,N_8024,N_8228);
nor U8429 (N_8429,N_8053,N_8077);
nor U8430 (N_8430,N_8182,N_8088);
or U8431 (N_8431,N_8177,N_8026);
xnor U8432 (N_8432,N_8027,N_8127);
or U8433 (N_8433,N_8086,N_8146);
or U8434 (N_8434,N_8181,N_8169);
nor U8435 (N_8435,N_8134,N_8144);
nand U8436 (N_8436,N_8186,N_8135);
and U8437 (N_8437,N_8238,N_8202);
and U8438 (N_8438,N_8011,N_8224);
nor U8439 (N_8439,N_8184,N_8193);
xnor U8440 (N_8440,N_8032,N_8229);
xnor U8441 (N_8441,N_8011,N_8095);
and U8442 (N_8442,N_8140,N_8108);
nor U8443 (N_8443,N_8029,N_8192);
and U8444 (N_8444,N_8222,N_8175);
nor U8445 (N_8445,N_8056,N_8076);
xnor U8446 (N_8446,N_8162,N_8060);
xor U8447 (N_8447,N_8215,N_8176);
nand U8448 (N_8448,N_8086,N_8097);
and U8449 (N_8449,N_8207,N_8205);
nor U8450 (N_8450,N_8035,N_8032);
or U8451 (N_8451,N_8063,N_8181);
and U8452 (N_8452,N_8089,N_8233);
xor U8453 (N_8453,N_8064,N_8075);
and U8454 (N_8454,N_8198,N_8065);
nand U8455 (N_8455,N_8139,N_8246);
xnor U8456 (N_8456,N_8158,N_8228);
xor U8457 (N_8457,N_8161,N_8240);
or U8458 (N_8458,N_8065,N_8100);
nor U8459 (N_8459,N_8099,N_8015);
and U8460 (N_8460,N_8119,N_8087);
and U8461 (N_8461,N_8069,N_8220);
xor U8462 (N_8462,N_8173,N_8077);
xnor U8463 (N_8463,N_8100,N_8142);
nor U8464 (N_8464,N_8160,N_8110);
or U8465 (N_8465,N_8228,N_8106);
nor U8466 (N_8466,N_8194,N_8245);
and U8467 (N_8467,N_8218,N_8082);
xnor U8468 (N_8468,N_8148,N_8025);
and U8469 (N_8469,N_8070,N_8066);
xnor U8470 (N_8470,N_8227,N_8104);
xnor U8471 (N_8471,N_8038,N_8200);
nor U8472 (N_8472,N_8022,N_8144);
nor U8473 (N_8473,N_8211,N_8049);
nand U8474 (N_8474,N_8067,N_8112);
and U8475 (N_8475,N_8164,N_8018);
and U8476 (N_8476,N_8195,N_8000);
nor U8477 (N_8477,N_8219,N_8109);
xor U8478 (N_8478,N_8141,N_8133);
nor U8479 (N_8479,N_8207,N_8224);
nor U8480 (N_8480,N_8062,N_8048);
xor U8481 (N_8481,N_8044,N_8246);
nand U8482 (N_8482,N_8096,N_8061);
xnor U8483 (N_8483,N_8094,N_8186);
and U8484 (N_8484,N_8026,N_8029);
or U8485 (N_8485,N_8183,N_8235);
xnor U8486 (N_8486,N_8019,N_8096);
and U8487 (N_8487,N_8017,N_8164);
xor U8488 (N_8488,N_8106,N_8091);
nor U8489 (N_8489,N_8105,N_8227);
nand U8490 (N_8490,N_8052,N_8037);
or U8491 (N_8491,N_8070,N_8077);
nand U8492 (N_8492,N_8198,N_8013);
or U8493 (N_8493,N_8124,N_8224);
and U8494 (N_8494,N_8237,N_8110);
nand U8495 (N_8495,N_8191,N_8183);
or U8496 (N_8496,N_8034,N_8168);
or U8497 (N_8497,N_8203,N_8100);
and U8498 (N_8498,N_8228,N_8055);
nand U8499 (N_8499,N_8073,N_8035);
or U8500 (N_8500,N_8477,N_8406);
nor U8501 (N_8501,N_8493,N_8367);
xnor U8502 (N_8502,N_8482,N_8463);
nand U8503 (N_8503,N_8468,N_8464);
and U8504 (N_8504,N_8473,N_8401);
xnor U8505 (N_8505,N_8404,N_8390);
nor U8506 (N_8506,N_8480,N_8460);
xnor U8507 (N_8507,N_8489,N_8283);
nor U8508 (N_8508,N_8313,N_8327);
xor U8509 (N_8509,N_8474,N_8402);
nand U8510 (N_8510,N_8415,N_8341);
nand U8511 (N_8511,N_8369,N_8353);
and U8512 (N_8512,N_8487,N_8368);
nand U8513 (N_8513,N_8403,N_8481);
and U8514 (N_8514,N_8329,N_8488);
and U8515 (N_8515,N_8413,N_8393);
nand U8516 (N_8516,N_8264,N_8301);
xor U8517 (N_8517,N_8395,N_8285);
nor U8518 (N_8518,N_8490,N_8436);
nor U8519 (N_8519,N_8443,N_8337);
and U8520 (N_8520,N_8437,N_8491);
or U8521 (N_8521,N_8499,N_8262);
nor U8522 (N_8522,N_8304,N_8438);
and U8523 (N_8523,N_8323,N_8379);
and U8524 (N_8524,N_8457,N_8392);
nor U8525 (N_8525,N_8391,N_8287);
xnor U8526 (N_8526,N_8296,N_8378);
xnor U8527 (N_8527,N_8260,N_8440);
xnor U8528 (N_8528,N_8351,N_8326);
and U8529 (N_8529,N_8373,N_8309);
and U8530 (N_8530,N_8299,N_8428);
xnor U8531 (N_8531,N_8348,N_8498);
nor U8532 (N_8532,N_8282,N_8427);
and U8533 (N_8533,N_8270,N_8442);
nand U8534 (N_8534,N_8412,N_8332);
and U8535 (N_8535,N_8446,N_8445);
or U8536 (N_8536,N_8462,N_8444);
xor U8537 (N_8537,N_8383,N_8279);
nor U8538 (N_8538,N_8343,N_8385);
or U8539 (N_8539,N_8336,N_8452);
and U8540 (N_8540,N_8324,N_8448);
nand U8541 (N_8541,N_8382,N_8459);
or U8542 (N_8542,N_8286,N_8295);
nor U8543 (N_8543,N_8338,N_8265);
nor U8544 (N_8544,N_8478,N_8257);
xor U8545 (N_8545,N_8307,N_8424);
nor U8546 (N_8546,N_8451,N_8453);
and U8547 (N_8547,N_8356,N_8305);
nand U8548 (N_8548,N_8435,N_8409);
nor U8549 (N_8549,N_8273,N_8398);
nand U8550 (N_8550,N_8430,N_8416);
nor U8551 (N_8551,N_8303,N_8344);
nand U8552 (N_8552,N_8253,N_8274);
xnor U8553 (N_8553,N_8342,N_8288);
nor U8554 (N_8554,N_8420,N_8358);
and U8555 (N_8555,N_8476,N_8399);
nor U8556 (N_8556,N_8370,N_8330);
or U8557 (N_8557,N_8300,N_8492);
or U8558 (N_8558,N_8471,N_8458);
or U8559 (N_8559,N_8456,N_8362);
or U8560 (N_8560,N_8429,N_8466);
nor U8561 (N_8561,N_8447,N_8345);
and U8562 (N_8562,N_8278,N_8423);
and U8563 (N_8563,N_8350,N_8387);
nand U8564 (N_8564,N_8419,N_8479);
nor U8565 (N_8565,N_8414,N_8467);
xor U8566 (N_8566,N_8441,N_8418);
and U8567 (N_8567,N_8255,N_8352);
and U8568 (N_8568,N_8258,N_8365);
nand U8569 (N_8569,N_8312,N_8455);
or U8570 (N_8570,N_8410,N_8340);
nand U8571 (N_8571,N_8417,N_8461);
and U8572 (N_8572,N_8310,N_8267);
nand U8573 (N_8573,N_8268,N_8275);
and U8574 (N_8574,N_8334,N_8497);
nand U8575 (N_8575,N_8449,N_8389);
nor U8576 (N_8576,N_8317,N_8355);
or U8577 (N_8577,N_8266,N_8276);
nor U8578 (N_8578,N_8363,N_8291);
xor U8579 (N_8579,N_8251,N_8431);
and U8580 (N_8580,N_8306,N_8290);
nand U8581 (N_8581,N_8421,N_8360);
or U8582 (N_8582,N_8321,N_8281);
and U8583 (N_8583,N_8354,N_8347);
nand U8584 (N_8584,N_8375,N_8320);
nor U8585 (N_8585,N_8472,N_8366);
nor U8586 (N_8586,N_8484,N_8261);
nor U8587 (N_8587,N_8280,N_8361);
nand U8588 (N_8588,N_8432,N_8494);
and U8589 (N_8589,N_8434,N_8465);
or U8590 (N_8590,N_8376,N_8394);
xor U8591 (N_8591,N_8397,N_8349);
nand U8592 (N_8592,N_8311,N_8308);
nor U8593 (N_8593,N_8318,N_8316);
nor U8594 (N_8594,N_8293,N_8495);
xor U8595 (N_8595,N_8314,N_8439);
and U8596 (N_8596,N_8298,N_8377);
nor U8597 (N_8597,N_8372,N_8277);
nor U8598 (N_8598,N_8289,N_8256);
xor U8599 (N_8599,N_8259,N_8322);
nand U8600 (N_8600,N_8380,N_8388);
and U8601 (N_8601,N_8405,N_8359);
nor U8602 (N_8602,N_8292,N_8450);
nor U8603 (N_8603,N_8483,N_8319);
nor U8604 (N_8604,N_8271,N_8470);
and U8605 (N_8605,N_8400,N_8254);
xnor U8606 (N_8606,N_8374,N_8315);
or U8607 (N_8607,N_8284,N_8485);
nor U8608 (N_8608,N_8486,N_8294);
or U8609 (N_8609,N_8331,N_8263);
xor U8610 (N_8610,N_8335,N_8346);
nand U8611 (N_8611,N_8433,N_8422);
or U8612 (N_8612,N_8339,N_8364);
nand U8613 (N_8613,N_8328,N_8469);
xor U8614 (N_8614,N_8297,N_8408);
nor U8615 (N_8615,N_8386,N_8302);
xnor U8616 (N_8616,N_8371,N_8496);
xnor U8617 (N_8617,N_8357,N_8252);
and U8618 (N_8618,N_8411,N_8454);
xnor U8619 (N_8619,N_8407,N_8426);
nand U8620 (N_8620,N_8269,N_8425);
nor U8621 (N_8621,N_8381,N_8333);
and U8622 (N_8622,N_8384,N_8396);
and U8623 (N_8623,N_8325,N_8272);
nor U8624 (N_8624,N_8250,N_8475);
nand U8625 (N_8625,N_8321,N_8373);
nand U8626 (N_8626,N_8378,N_8453);
and U8627 (N_8627,N_8335,N_8474);
and U8628 (N_8628,N_8374,N_8255);
nor U8629 (N_8629,N_8475,N_8412);
nand U8630 (N_8630,N_8415,N_8367);
and U8631 (N_8631,N_8461,N_8472);
xor U8632 (N_8632,N_8473,N_8361);
nand U8633 (N_8633,N_8443,N_8393);
nand U8634 (N_8634,N_8418,N_8308);
nor U8635 (N_8635,N_8331,N_8410);
and U8636 (N_8636,N_8308,N_8490);
and U8637 (N_8637,N_8467,N_8416);
nor U8638 (N_8638,N_8344,N_8274);
or U8639 (N_8639,N_8315,N_8360);
nor U8640 (N_8640,N_8388,N_8279);
nor U8641 (N_8641,N_8309,N_8464);
and U8642 (N_8642,N_8278,N_8332);
nand U8643 (N_8643,N_8389,N_8455);
or U8644 (N_8644,N_8390,N_8453);
and U8645 (N_8645,N_8379,N_8391);
nor U8646 (N_8646,N_8260,N_8436);
nand U8647 (N_8647,N_8300,N_8277);
nor U8648 (N_8648,N_8314,N_8474);
nor U8649 (N_8649,N_8416,N_8425);
and U8650 (N_8650,N_8344,N_8470);
or U8651 (N_8651,N_8351,N_8481);
nand U8652 (N_8652,N_8499,N_8288);
or U8653 (N_8653,N_8392,N_8270);
or U8654 (N_8654,N_8339,N_8340);
and U8655 (N_8655,N_8308,N_8382);
nand U8656 (N_8656,N_8437,N_8300);
and U8657 (N_8657,N_8433,N_8397);
and U8658 (N_8658,N_8469,N_8394);
nand U8659 (N_8659,N_8375,N_8459);
nand U8660 (N_8660,N_8475,N_8435);
nand U8661 (N_8661,N_8458,N_8431);
or U8662 (N_8662,N_8374,N_8300);
and U8663 (N_8663,N_8387,N_8432);
and U8664 (N_8664,N_8287,N_8250);
or U8665 (N_8665,N_8388,N_8291);
nor U8666 (N_8666,N_8261,N_8442);
and U8667 (N_8667,N_8363,N_8399);
and U8668 (N_8668,N_8268,N_8369);
nand U8669 (N_8669,N_8283,N_8475);
nor U8670 (N_8670,N_8425,N_8353);
and U8671 (N_8671,N_8294,N_8390);
and U8672 (N_8672,N_8335,N_8338);
nand U8673 (N_8673,N_8260,N_8398);
xnor U8674 (N_8674,N_8310,N_8442);
nand U8675 (N_8675,N_8258,N_8353);
or U8676 (N_8676,N_8285,N_8411);
nor U8677 (N_8677,N_8285,N_8364);
nor U8678 (N_8678,N_8377,N_8491);
or U8679 (N_8679,N_8392,N_8258);
xor U8680 (N_8680,N_8431,N_8250);
nand U8681 (N_8681,N_8388,N_8370);
nand U8682 (N_8682,N_8345,N_8419);
nor U8683 (N_8683,N_8332,N_8474);
xor U8684 (N_8684,N_8414,N_8308);
xor U8685 (N_8685,N_8374,N_8351);
nor U8686 (N_8686,N_8282,N_8357);
or U8687 (N_8687,N_8319,N_8366);
and U8688 (N_8688,N_8444,N_8452);
and U8689 (N_8689,N_8422,N_8336);
or U8690 (N_8690,N_8275,N_8484);
nand U8691 (N_8691,N_8314,N_8352);
nand U8692 (N_8692,N_8475,N_8384);
xnor U8693 (N_8693,N_8480,N_8281);
and U8694 (N_8694,N_8409,N_8285);
and U8695 (N_8695,N_8299,N_8345);
nand U8696 (N_8696,N_8350,N_8493);
and U8697 (N_8697,N_8359,N_8458);
or U8698 (N_8698,N_8300,N_8319);
nor U8699 (N_8699,N_8372,N_8340);
and U8700 (N_8700,N_8316,N_8295);
or U8701 (N_8701,N_8279,N_8267);
nor U8702 (N_8702,N_8419,N_8451);
nor U8703 (N_8703,N_8495,N_8371);
nor U8704 (N_8704,N_8282,N_8466);
xnor U8705 (N_8705,N_8257,N_8407);
xnor U8706 (N_8706,N_8439,N_8431);
and U8707 (N_8707,N_8355,N_8251);
and U8708 (N_8708,N_8480,N_8458);
and U8709 (N_8709,N_8383,N_8387);
nor U8710 (N_8710,N_8258,N_8295);
nor U8711 (N_8711,N_8367,N_8320);
nand U8712 (N_8712,N_8483,N_8261);
or U8713 (N_8713,N_8298,N_8494);
or U8714 (N_8714,N_8326,N_8407);
nor U8715 (N_8715,N_8315,N_8420);
or U8716 (N_8716,N_8424,N_8431);
nand U8717 (N_8717,N_8479,N_8347);
and U8718 (N_8718,N_8305,N_8290);
nand U8719 (N_8719,N_8282,N_8474);
and U8720 (N_8720,N_8480,N_8253);
nand U8721 (N_8721,N_8421,N_8260);
nor U8722 (N_8722,N_8375,N_8352);
or U8723 (N_8723,N_8359,N_8390);
and U8724 (N_8724,N_8493,N_8449);
nand U8725 (N_8725,N_8374,N_8466);
and U8726 (N_8726,N_8472,N_8309);
nor U8727 (N_8727,N_8470,N_8320);
xnor U8728 (N_8728,N_8388,N_8438);
nor U8729 (N_8729,N_8473,N_8257);
nand U8730 (N_8730,N_8346,N_8441);
or U8731 (N_8731,N_8276,N_8411);
and U8732 (N_8732,N_8405,N_8265);
nand U8733 (N_8733,N_8437,N_8267);
nand U8734 (N_8734,N_8405,N_8424);
xnor U8735 (N_8735,N_8332,N_8468);
or U8736 (N_8736,N_8448,N_8315);
nand U8737 (N_8737,N_8496,N_8470);
nor U8738 (N_8738,N_8488,N_8270);
or U8739 (N_8739,N_8297,N_8321);
nor U8740 (N_8740,N_8373,N_8438);
nand U8741 (N_8741,N_8405,N_8355);
and U8742 (N_8742,N_8401,N_8254);
xnor U8743 (N_8743,N_8413,N_8430);
xnor U8744 (N_8744,N_8312,N_8321);
and U8745 (N_8745,N_8292,N_8330);
xnor U8746 (N_8746,N_8309,N_8337);
and U8747 (N_8747,N_8453,N_8322);
nand U8748 (N_8748,N_8441,N_8359);
nor U8749 (N_8749,N_8296,N_8346);
nor U8750 (N_8750,N_8656,N_8731);
xnor U8751 (N_8751,N_8566,N_8554);
nand U8752 (N_8752,N_8721,N_8599);
nor U8753 (N_8753,N_8693,N_8629);
or U8754 (N_8754,N_8519,N_8606);
nand U8755 (N_8755,N_8543,N_8607);
xnor U8756 (N_8756,N_8655,N_8735);
and U8757 (N_8757,N_8512,N_8671);
nand U8758 (N_8758,N_8501,N_8712);
nand U8759 (N_8759,N_8636,N_8610);
xnor U8760 (N_8760,N_8609,N_8649);
or U8761 (N_8761,N_8570,N_8624);
nand U8762 (N_8762,N_8746,N_8654);
nor U8763 (N_8763,N_8679,N_8627);
nand U8764 (N_8764,N_8640,N_8520);
nor U8765 (N_8765,N_8727,N_8544);
nor U8766 (N_8766,N_8711,N_8601);
nand U8767 (N_8767,N_8719,N_8515);
xor U8768 (N_8768,N_8676,N_8552);
or U8769 (N_8769,N_8533,N_8733);
and U8770 (N_8770,N_8696,N_8685);
nand U8771 (N_8771,N_8535,N_8739);
and U8772 (N_8772,N_8562,N_8557);
and U8773 (N_8773,N_8532,N_8509);
nor U8774 (N_8774,N_8677,N_8621);
nor U8775 (N_8775,N_8556,N_8672);
nand U8776 (N_8776,N_8738,N_8540);
and U8777 (N_8777,N_8652,N_8615);
and U8778 (N_8778,N_8580,N_8740);
nand U8779 (N_8779,N_8527,N_8588);
and U8780 (N_8780,N_8747,N_8567);
nor U8781 (N_8781,N_8718,N_8593);
or U8782 (N_8782,N_8638,N_8653);
or U8783 (N_8783,N_8635,N_8691);
nand U8784 (N_8784,N_8591,N_8600);
nor U8785 (N_8785,N_8542,N_8732);
or U8786 (N_8786,N_8612,N_8553);
nor U8787 (N_8787,N_8661,N_8651);
xnor U8788 (N_8788,N_8680,N_8716);
nor U8789 (N_8789,N_8645,N_8689);
nand U8790 (N_8790,N_8604,N_8673);
nor U8791 (N_8791,N_8648,N_8717);
or U8792 (N_8792,N_8703,N_8521);
nand U8793 (N_8793,N_8575,N_8741);
nor U8794 (N_8794,N_8634,N_8724);
nor U8795 (N_8795,N_8614,N_8547);
nor U8796 (N_8796,N_8744,N_8524);
xnor U8797 (N_8797,N_8686,N_8569);
nor U8798 (N_8798,N_8626,N_8688);
or U8799 (N_8799,N_8595,N_8608);
nor U8800 (N_8800,N_8734,N_8526);
xor U8801 (N_8801,N_8537,N_8590);
xor U8802 (N_8802,N_8522,N_8517);
nor U8803 (N_8803,N_8650,N_8674);
xnor U8804 (N_8804,N_8505,N_8538);
xnor U8805 (N_8805,N_8572,N_8563);
nand U8806 (N_8806,N_8558,N_8713);
or U8807 (N_8807,N_8702,N_8597);
xor U8808 (N_8808,N_8578,N_8619);
xnor U8809 (N_8809,N_8613,N_8571);
nor U8810 (N_8810,N_8545,N_8700);
xor U8811 (N_8811,N_8715,N_8698);
or U8812 (N_8812,N_8546,N_8748);
and U8813 (N_8813,N_8589,N_8549);
xor U8814 (N_8814,N_8514,N_8692);
or U8815 (N_8815,N_8705,N_8617);
nand U8816 (N_8816,N_8723,N_8564);
or U8817 (N_8817,N_8534,N_8602);
or U8818 (N_8818,N_8667,N_8637);
and U8819 (N_8819,N_8603,N_8631);
nand U8820 (N_8820,N_8706,N_8525);
xor U8821 (N_8821,N_8592,N_8523);
or U8822 (N_8822,N_8632,N_8539);
or U8823 (N_8823,N_8708,N_8678);
or U8824 (N_8824,N_8611,N_8681);
and U8825 (N_8825,N_8647,N_8714);
nand U8826 (N_8826,N_8630,N_8669);
nor U8827 (N_8827,N_8749,N_8694);
nor U8828 (N_8828,N_8555,N_8577);
and U8829 (N_8829,N_8559,N_8502);
xor U8830 (N_8830,N_8548,N_8729);
and U8831 (N_8831,N_8664,N_8642);
and U8832 (N_8832,N_8507,N_8684);
and U8833 (N_8833,N_8536,N_8516);
nor U8834 (N_8834,N_8662,N_8551);
nor U8835 (N_8835,N_8581,N_8699);
and U8836 (N_8836,N_8665,N_8720);
xor U8837 (N_8837,N_8568,N_8529);
xor U8838 (N_8838,N_8618,N_8683);
nand U8839 (N_8839,N_8510,N_8710);
and U8840 (N_8840,N_8709,N_8730);
xor U8841 (N_8841,N_8528,N_8668);
or U8842 (N_8842,N_8639,N_8643);
nor U8843 (N_8843,N_8701,N_8728);
nor U8844 (N_8844,N_8736,N_8646);
and U8845 (N_8845,N_8531,N_8504);
and U8846 (N_8846,N_8541,N_8579);
nand U8847 (N_8847,N_8625,N_8726);
nor U8848 (N_8848,N_8508,N_8573);
and U8849 (N_8849,N_8560,N_8704);
xnor U8850 (N_8850,N_8585,N_8513);
and U8851 (N_8851,N_8687,N_8628);
nor U8852 (N_8852,N_8596,N_8722);
and U8853 (N_8853,N_8666,N_8743);
or U8854 (N_8854,N_8574,N_8511);
or U8855 (N_8855,N_8745,N_8695);
or U8856 (N_8856,N_8565,N_8576);
nand U8857 (N_8857,N_8658,N_8616);
or U8858 (N_8858,N_8605,N_8657);
or U8859 (N_8859,N_8550,N_8584);
nand U8860 (N_8860,N_8518,N_8622);
nand U8861 (N_8861,N_8682,N_8697);
nor U8862 (N_8862,N_8623,N_8500);
nand U8863 (N_8863,N_8503,N_8663);
or U8864 (N_8864,N_8587,N_8506);
nand U8865 (N_8865,N_8530,N_8620);
and U8866 (N_8866,N_8670,N_8675);
or U8867 (N_8867,N_8598,N_8641);
and U8868 (N_8868,N_8660,N_8707);
nand U8869 (N_8869,N_8586,N_8742);
and U8870 (N_8870,N_8583,N_8582);
or U8871 (N_8871,N_8594,N_8633);
or U8872 (N_8872,N_8659,N_8690);
or U8873 (N_8873,N_8737,N_8561);
and U8874 (N_8874,N_8725,N_8644);
and U8875 (N_8875,N_8667,N_8741);
nor U8876 (N_8876,N_8694,N_8608);
and U8877 (N_8877,N_8503,N_8536);
nand U8878 (N_8878,N_8510,N_8614);
nand U8879 (N_8879,N_8560,N_8631);
xnor U8880 (N_8880,N_8669,N_8500);
nand U8881 (N_8881,N_8564,N_8500);
nand U8882 (N_8882,N_8578,N_8505);
or U8883 (N_8883,N_8581,N_8692);
nor U8884 (N_8884,N_8542,N_8520);
xnor U8885 (N_8885,N_8722,N_8708);
nor U8886 (N_8886,N_8657,N_8506);
xor U8887 (N_8887,N_8695,N_8532);
nor U8888 (N_8888,N_8693,N_8577);
xnor U8889 (N_8889,N_8745,N_8683);
xnor U8890 (N_8890,N_8561,N_8593);
nor U8891 (N_8891,N_8533,N_8702);
xor U8892 (N_8892,N_8596,N_8733);
or U8893 (N_8893,N_8733,N_8682);
or U8894 (N_8894,N_8715,N_8533);
nor U8895 (N_8895,N_8522,N_8642);
nor U8896 (N_8896,N_8638,N_8697);
nand U8897 (N_8897,N_8639,N_8710);
nand U8898 (N_8898,N_8549,N_8615);
nand U8899 (N_8899,N_8538,N_8700);
nor U8900 (N_8900,N_8602,N_8674);
and U8901 (N_8901,N_8626,N_8619);
or U8902 (N_8902,N_8532,N_8607);
and U8903 (N_8903,N_8713,N_8637);
xor U8904 (N_8904,N_8572,N_8621);
nand U8905 (N_8905,N_8613,N_8603);
and U8906 (N_8906,N_8558,N_8644);
nand U8907 (N_8907,N_8717,N_8708);
xnor U8908 (N_8908,N_8654,N_8626);
nand U8909 (N_8909,N_8697,N_8657);
and U8910 (N_8910,N_8601,N_8568);
xor U8911 (N_8911,N_8726,N_8658);
xor U8912 (N_8912,N_8686,N_8724);
and U8913 (N_8913,N_8527,N_8535);
nand U8914 (N_8914,N_8618,N_8713);
or U8915 (N_8915,N_8557,N_8504);
or U8916 (N_8916,N_8730,N_8638);
or U8917 (N_8917,N_8600,N_8720);
or U8918 (N_8918,N_8640,N_8707);
xor U8919 (N_8919,N_8506,N_8626);
nand U8920 (N_8920,N_8659,N_8632);
or U8921 (N_8921,N_8695,N_8632);
or U8922 (N_8922,N_8741,N_8526);
xor U8923 (N_8923,N_8598,N_8584);
nor U8924 (N_8924,N_8714,N_8742);
nand U8925 (N_8925,N_8723,N_8553);
nor U8926 (N_8926,N_8722,N_8665);
or U8927 (N_8927,N_8740,N_8506);
nor U8928 (N_8928,N_8605,N_8516);
xor U8929 (N_8929,N_8587,N_8593);
xnor U8930 (N_8930,N_8627,N_8749);
and U8931 (N_8931,N_8529,N_8632);
xnor U8932 (N_8932,N_8744,N_8540);
or U8933 (N_8933,N_8603,N_8667);
or U8934 (N_8934,N_8599,N_8552);
nand U8935 (N_8935,N_8517,N_8585);
nor U8936 (N_8936,N_8649,N_8544);
nor U8937 (N_8937,N_8550,N_8576);
xnor U8938 (N_8938,N_8541,N_8632);
nor U8939 (N_8939,N_8513,N_8549);
nor U8940 (N_8940,N_8707,N_8739);
or U8941 (N_8941,N_8601,N_8634);
nor U8942 (N_8942,N_8743,N_8545);
xor U8943 (N_8943,N_8612,N_8661);
and U8944 (N_8944,N_8692,N_8567);
and U8945 (N_8945,N_8634,N_8607);
xor U8946 (N_8946,N_8581,N_8510);
xor U8947 (N_8947,N_8679,N_8500);
or U8948 (N_8948,N_8588,N_8739);
nand U8949 (N_8949,N_8618,N_8541);
nand U8950 (N_8950,N_8655,N_8715);
nand U8951 (N_8951,N_8555,N_8710);
and U8952 (N_8952,N_8682,N_8640);
xnor U8953 (N_8953,N_8717,N_8638);
and U8954 (N_8954,N_8697,N_8710);
nor U8955 (N_8955,N_8696,N_8637);
nand U8956 (N_8956,N_8691,N_8572);
and U8957 (N_8957,N_8563,N_8630);
nor U8958 (N_8958,N_8591,N_8603);
xor U8959 (N_8959,N_8524,N_8509);
nand U8960 (N_8960,N_8622,N_8621);
and U8961 (N_8961,N_8533,N_8647);
nor U8962 (N_8962,N_8500,N_8739);
xor U8963 (N_8963,N_8602,N_8710);
xor U8964 (N_8964,N_8551,N_8694);
nand U8965 (N_8965,N_8648,N_8678);
nor U8966 (N_8966,N_8676,N_8524);
nor U8967 (N_8967,N_8549,N_8579);
and U8968 (N_8968,N_8670,N_8612);
and U8969 (N_8969,N_8675,N_8740);
and U8970 (N_8970,N_8589,N_8550);
nand U8971 (N_8971,N_8749,N_8504);
nor U8972 (N_8972,N_8518,N_8566);
nand U8973 (N_8973,N_8605,N_8529);
and U8974 (N_8974,N_8577,N_8717);
nor U8975 (N_8975,N_8705,N_8535);
and U8976 (N_8976,N_8696,N_8705);
nor U8977 (N_8977,N_8523,N_8665);
or U8978 (N_8978,N_8700,N_8637);
nor U8979 (N_8979,N_8524,N_8656);
xnor U8980 (N_8980,N_8599,N_8722);
or U8981 (N_8981,N_8583,N_8578);
nand U8982 (N_8982,N_8693,N_8578);
and U8983 (N_8983,N_8694,N_8668);
or U8984 (N_8984,N_8527,N_8639);
nor U8985 (N_8985,N_8729,N_8694);
nor U8986 (N_8986,N_8594,N_8567);
and U8987 (N_8987,N_8540,N_8613);
xor U8988 (N_8988,N_8700,N_8573);
or U8989 (N_8989,N_8539,N_8529);
or U8990 (N_8990,N_8573,N_8600);
nand U8991 (N_8991,N_8568,N_8523);
and U8992 (N_8992,N_8696,N_8673);
nand U8993 (N_8993,N_8527,N_8713);
nand U8994 (N_8994,N_8740,N_8546);
and U8995 (N_8995,N_8546,N_8744);
nor U8996 (N_8996,N_8526,N_8748);
nor U8997 (N_8997,N_8534,N_8544);
nor U8998 (N_8998,N_8653,N_8566);
nand U8999 (N_8999,N_8663,N_8671);
or U9000 (N_9000,N_8827,N_8850);
nor U9001 (N_9001,N_8764,N_8923);
and U9002 (N_9002,N_8924,N_8918);
xnor U9003 (N_9003,N_8871,N_8881);
nand U9004 (N_9004,N_8932,N_8831);
and U9005 (N_9005,N_8919,N_8822);
nor U9006 (N_9006,N_8814,N_8756);
nor U9007 (N_9007,N_8848,N_8864);
nand U9008 (N_9008,N_8970,N_8836);
and U9009 (N_9009,N_8821,N_8784);
and U9010 (N_9010,N_8948,N_8809);
and U9011 (N_9011,N_8907,N_8761);
nand U9012 (N_9012,N_8963,N_8802);
xnor U9013 (N_9013,N_8755,N_8812);
xnor U9014 (N_9014,N_8771,N_8837);
xor U9015 (N_9015,N_8853,N_8886);
nand U9016 (N_9016,N_8928,N_8855);
nor U9017 (N_9017,N_8934,N_8898);
nor U9018 (N_9018,N_8752,N_8950);
and U9019 (N_9019,N_8843,N_8975);
nand U9020 (N_9020,N_8854,N_8753);
nand U9021 (N_9021,N_8816,N_8922);
xnor U9022 (N_9022,N_8800,N_8778);
nor U9023 (N_9023,N_8791,N_8883);
or U9024 (N_9024,N_8862,N_8940);
xor U9025 (N_9025,N_8914,N_8960);
xor U9026 (N_9026,N_8949,N_8786);
nand U9027 (N_9027,N_8795,N_8751);
and U9028 (N_9028,N_8829,N_8895);
xnor U9029 (N_9029,N_8917,N_8890);
nand U9030 (N_9030,N_8893,N_8964);
nor U9031 (N_9031,N_8952,N_8787);
nor U9032 (N_9032,N_8840,N_8776);
or U9033 (N_9033,N_8842,N_8900);
xnor U9034 (N_9034,N_8982,N_8988);
and U9035 (N_9035,N_8887,N_8997);
and U9036 (N_9036,N_8773,N_8845);
nor U9037 (N_9037,N_8983,N_8971);
nor U9038 (N_9038,N_8911,N_8832);
xor U9039 (N_9039,N_8856,N_8966);
and U9040 (N_9040,N_8878,N_8985);
and U9041 (N_9041,N_8852,N_8959);
nor U9042 (N_9042,N_8772,N_8980);
nand U9043 (N_9043,N_8847,N_8808);
or U9044 (N_9044,N_8750,N_8879);
or U9045 (N_9045,N_8978,N_8910);
nand U9046 (N_9046,N_8803,N_8921);
nor U9047 (N_9047,N_8873,N_8758);
and U9048 (N_9048,N_8861,N_8799);
and U9049 (N_9049,N_8989,N_8986);
xor U9050 (N_9050,N_8781,N_8830);
or U9051 (N_9051,N_8849,N_8815);
and U9052 (N_9052,N_8884,N_8951);
or U9053 (N_9053,N_8869,N_8782);
nor U9054 (N_9054,N_8927,N_8860);
xor U9055 (N_9055,N_8806,N_8838);
nand U9056 (N_9056,N_8942,N_8996);
or U9057 (N_9057,N_8903,N_8759);
xor U9058 (N_9058,N_8793,N_8954);
nor U9059 (N_9059,N_8804,N_8851);
xnor U9060 (N_9060,N_8790,N_8930);
nand U9061 (N_9061,N_8823,N_8828);
xnor U9062 (N_9062,N_8945,N_8969);
nand U9063 (N_9063,N_8768,N_8817);
and U9064 (N_9064,N_8767,N_8925);
xor U9065 (N_9065,N_8798,N_8866);
xor U9066 (N_9066,N_8833,N_8763);
nor U9067 (N_9067,N_8901,N_8953);
and U9068 (N_9068,N_8859,N_8888);
or U9069 (N_9069,N_8944,N_8825);
nor U9070 (N_9070,N_8984,N_8958);
nor U9071 (N_9071,N_8957,N_8788);
or U9072 (N_9072,N_8754,N_8991);
and U9073 (N_9073,N_8874,N_8968);
and U9074 (N_9074,N_8870,N_8813);
and U9075 (N_9075,N_8766,N_8857);
or U9076 (N_9076,N_8899,N_8805);
xor U9077 (N_9077,N_8769,N_8965);
or U9078 (N_9078,N_8834,N_8913);
nor U9079 (N_9079,N_8777,N_8933);
nor U9080 (N_9080,N_8894,N_8915);
xor U9081 (N_9081,N_8955,N_8939);
nor U9082 (N_9082,N_8889,N_8877);
and U9083 (N_9083,N_8908,N_8875);
xnor U9084 (N_9084,N_8844,N_8826);
or U9085 (N_9085,N_8868,N_8990);
xor U9086 (N_9086,N_8938,N_8946);
nand U9087 (N_9087,N_8937,N_8780);
nor U9088 (N_9088,N_8882,N_8792);
and U9089 (N_9089,N_8762,N_8858);
nand U9090 (N_9090,N_8846,N_8775);
or U9091 (N_9091,N_8824,N_8962);
or U9092 (N_9092,N_8811,N_8891);
nor U9093 (N_9093,N_8906,N_8797);
or U9094 (N_9094,N_8794,N_8789);
nor U9095 (N_9095,N_8785,N_8912);
xnor U9096 (N_9096,N_8979,N_8757);
xor U9097 (N_9097,N_8760,N_8920);
and U9098 (N_9098,N_8936,N_8976);
nor U9099 (N_9099,N_8972,N_8981);
nand U9100 (N_9100,N_8892,N_8876);
nor U9101 (N_9101,N_8841,N_8867);
or U9102 (N_9102,N_8896,N_8779);
nand U9103 (N_9103,N_8941,N_8796);
nor U9104 (N_9104,N_8992,N_8905);
nor U9105 (N_9105,N_8943,N_8931);
nand U9106 (N_9106,N_8774,N_8902);
nand U9107 (N_9107,N_8765,N_8999);
and U9108 (N_9108,N_8807,N_8977);
and U9109 (N_9109,N_8885,N_8929);
nand U9110 (N_9110,N_8935,N_8926);
and U9111 (N_9111,N_8904,N_8947);
or U9112 (N_9112,N_8916,N_8993);
xnor U9113 (N_9113,N_8897,N_8994);
nand U9114 (N_9114,N_8801,N_8819);
nand U9115 (N_9115,N_8995,N_8810);
xor U9116 (N_9116,N_8820,N_8872);
and U9117 (N_9117,N_8835,N_8961);
nand U9118 (N_9118,N_8987,N_8973);
xor U9119 (N_9119,N_8998,N_8865);
or U9120 (N_9120,N_8770,N_8783);
xnor U9121 (N_9121,N_8967,N_8909);
or U9122 (N_9122,N_8880,N_8956);
nor U9123 (N_9123,N_8974,N_8818);
xor U9124 (N_9124,N_8839,N_8863);
nor U9125 (N_9125,N_8778,N_8866);
nand U9126 (N_9126,N_8814,N_8879);
xor U9127 (N_9127,N_8801,N_8972);
and U9128 (N_9128,N_8783,N_8865);
and U9129 (N_9129,N_8966,N_8798);
or U9130 (N_9130,N_8940,N_8951);
xor U9131 (N_9131,N_8832,N_8921);
or U9132 (N_9132,N_8986,N_8979);
xnor U9133 (N_9133,N_8798,N_8842);
xnor U9134 (N_9134,N_8912,N_8977);
xor U9135 (N_9135,N_8791,N_8937);
and U9136 (N_9136,N_8910,N_8918);
nor U9137 (N_9137,N_8805,N_8971);
nand U9138 (N_9138,N_8939,N_8891);
and U9139 (N_9139,N_8786,N_8845);
nor U9140 (N_9140,N_8824,N_8806);
nor U9141 (N_9141,N_8943,N_8984);
xor U9142 (N_9142,N_8771,N_8977);
or U9143 (N_9143,N_8865,N_8948);
nor U9144 (N_9144,N_8871,N_8994);
nor U9145 (N_9145,N_8788,N_8834);
nor U9146 (N_9146,N_8916,N_8909);
and U9147 (N_9147,N_8830,N_8765);
xor U9148 (N_9148,N_8869,N_8985);
nor U9149 (N_9149,N_8773,N_8778);
or U9150 (N_9150,N_8904,N_8942);
or U9151 (N_9151,N_8858,N_8776);
xnor U9152 (N_9152,N_8997,N_8969);
nand U9153 (N_9153,N_8894,N_8839);
xnor U9154 (N_9154,N_8849,N_8969);
nor U9155 (N_9155,N_8859,N_8928);
nand U9156 (N_9156,N_8973,N_8845);
nor U9157 (N_9157,N_8798,N_8816);
nand U9158 (N_9158,N_8864,N_8967);
or U9159 (N_9159,N_8885,N_8971);
xor U9160 (N_9160,N_8822,N_8817);
xor U9161 (N_9161,N_8822,N_8767);
and U9162 (N_9162,N_8965,N_8825);
nor U9163 (N_9163,N_8930,N_8763);
xnor U9164 (N_9164,N_8765,N_8998);
xnor U9165 (N_9165,N_8911,N_8962);
and U9166 (N_9166,N_8882,N_8808);
and U9167 (N_9167,N_8761,N_8990);
nand U9168 (N_9168,N_8912,N_8790);
or U9169 (N_9169,N_8812,N_8967);
or U9170 (N_9170,N_8932,N_8964);
xor U9171 (N_9171,N_8975,N_8844);
and U9172 (N_9172,N_8882,N_8816);
xnor U9173 (N_9173,N_8788,N_8862);
nand U9174 (N_9174,N_8950,N_8964);
or U9175 (N_9175,N_8894,N_8842);
and U9176 (N_9176,N_8817,N_8789);
nor U9177 (N_9177,N_8940,N_8860);
xor U9178 (N_9178,N_8878,N_8955);
nor U9179 (N_9179,N_8769,N_8885);
and U9180 (N_9180,N_8754,N_8777);
nand U9181 (N_9181,N_8889,N_8995);
nand U9182 (N_9182,N_8830,N_8887);
xnor U9183 (N_9183,N_8863,N_8882);
and U9184 (N_9184,N_8973,N_8920);
nor U9185 (N_9185,N_8766,N_8927);
nor U9186 (N_9186,N_8867,N_8953);
nand U9187 (N_9187,N_8775,N_8770);
nand U9188 (N_9188,N_8840,N_8824);
nand U9189 (N_9189,N_8947,N_8857);
nand U9190 (N_9190,N_8982,N_8769);
nand U9191 (N_9191,N_8774,N_8835);
xor U9192 (N_9192,N_8775,N_8904);
and U9193 (N_9193,N_8766,N_8878);
and U9194 (N_9194,N_8856,N_8953);
nand U9195 (N_9195,N_8915,N_8863);
xor U9196 (N_9196,N_8778,N_8977);
nand U9197 (N_9197,N_8936,N_8914);
and U9198 (N_9198,N_8918,N_8936);
or U9199 (N_9199,N_8835,N_8930);
or U9200 (N_9200,N_8906,N_8951);
and U9201 (N_9201,N_8799,N_8848);
or U9202 (N_9202,N_8855,N_8874);
or U9203 (N_9203,N_8794,N_8887);
nor U9204 (N_9204,N_8935,N_8915);
or U9205 (N_9205,N_8880,N_8782);
and U9206 (N_9206,N_8959,N_8776);
nor U9207 (N_9207,N_8759,N_8914);
nand U9208 (N_9208,N_8762,N_8933);
or U9209 (N_9209,N_8761,N_8915);
xor U9210 (N_9210,N_8781,N_8760);
or U9211 (N_9211,N_8841,N_8997);
and U9212 (N_9212,N_8832,N_8929);
and U9213 (N_9213,N_8784,N_8977);
nand U9214 (N_9214,N_8828,N_8881);
or U9215 (N_9215,N_8799,N_8884);
or U9216 (N_9216,N_8767,N_8880);
or U9217 (N_9217,N_8757,N_8893);
nor U9218 (N_9218,N_8940,N_8892);
and U9219 (N_9219,N_8999,N_8952);
xnor U9220 (N_9220,N_8932,N_8772);
or U9221 (N_9221,N_8926,N_8906);
xnor U9222 (N_9222,N_8764,N_8860);
or U9223 (N_9223,N_8897,N_8824);
nor U9224 (N_9224,N_8813,N_8890);
xor U9225 (N_9225,N_8898,N_8770);
nand U9226 (N_9226,N_8802,N_8806);
nor U9227 (N_9227,N_8766,N_8818);
nand U9228 (N_9228,N_8898,N_8831);
xor U9229 (N_9229,N_8753,N_8771);
or U9230 (N_9230,N_8942,N_8938);
xor U9231 (N_9231,N_8941,N_8856);
xor U9232 (N_9232,N_8953,N_8962);
nand U9233 (N_9233,N_8805,N_8918);
nand U9234 (N_9234,N_8755,N_8823);
or U9235 (N_9235,N_8901,N_8899);
and U9236 (N_9236,N_8913,N_8787);
xor U9237 (N_9237,N_8830,N_8951);
xnor U9238 (N_9238,N_8852,N_8840);
xor U9239 (N_9239,N_8835,N_8773);
xor U9240 (N_9240,N_8885,N_8977);
xor U9241 (N_9241,N_8981,N_8778);
nor U9242 (N_9242,N_8967,N_8896);
or U9243 (N_9243,N_8769,N_8926);
nand U9244 (N_9244,N_8786,N_8986);
and U9245 (N_9245,N_8893,N_8945);
nor U9246 (N_9246,N_8893,N_8954);
or U9247 (N_9247,N_8757,N_8980);
xnor U9248 (N_9248,N_8826,N_8869);
and U9249 (N_9249,N_8774,N_8827);
nand U9250 (N_9250,N_9163,N_9098);
and U9251 (N_9251,N_9090,N_9201);
or U9252 (N_9252,N_9030,N_9192);
or U9253 (N_9253,N_9121,N_9248);
nor U9254 (N_9254,N_9020,N_9158);
and U9255 (N_9255,N_9213,N_9058);
nand U9256 (N_9256,N_9203,N_9228);
xor U9257 (N_9257,N_9231,N_9091);
nor U9258 (N_9258,N_9145,N_9195);
nor U9259 (N_9259,N_9147,N_9205);
nor U9260 (N_9260,N_9156,N_9002);
and U9261 (N_9261,N_9193,N_9104);
and U9262 (N_9262,N_9016,N_9120);
or U9263 (N_9263,N_9107,N_9161);
nor U9264 (N_9264,N_9187,N_9202);
xnor U9265 (N_9265,N_9131,N_9073);
nand U9266 (N_9266,N_9071,N_9190);
xnor U9267 (N_9267,N_9197,N_9103);
xnor U9268 (N_9268,N_9003,N_9047);
or U9269 (N_9269,N_9166,N_9046);
nand U9270 (N_9270,N_9083,N_9208);
or U9271 (N_9271,N_9061,N_9008);
and U9272 (N_9272,N_9137,N_9175);
and U9273 (N_9273,N_9100,N_9066);
or U9274 (N_9274,N_9031,N_9136);
nand U9275 (N_9275,N_9113,N_9233);
or U9276 (N_9276,N_9128,N_9212);
or U9277 (N_9277,N_9246,N_9057);
and U9278 (N_9278,N_9139,N_9112);
nand U9279 (N_9279,N_9168,N_9235);
nor U9280 (N_9280,N_9155,N_9093);
xnor U9281 (N_9281,N_9078,N_9127);
nand U9282 (N_9282,N_9040,N_9005);
nor U9283 (N_9283,N_9063,N_9075);
nor U9284 (N_9284,N_9105,N_9179);
nor U9285 (N_9285,N_9207,N_9159);
and U9286 (N_9286,N_9010,N_9176);
xnor U9287 (N_9287,N_9004,N_9000);
nor U9288 (N_9288,N_9189,N_9217);
nand U9289 (N_9289,N_9056,N_9037);
nor U9290 (N_9290,N_9026,N_9064);
or U9291 (N_9291,N_9108,N_9196);
nor U9292 (N_9292,N_9021,N_9164);
nor U9293 (N_9293,N_9007,N_9157);
xor U9294 (N_9294,N_9178,N_9094);
nand U9295 (N_9295,N_9132,N_9012);
nand U9296 (N_9296,N_9124,N_9150);
nand U9297 (N_9297,N_9223,N_9059);
nor U9298 (N_9298,N_9028,N_9045);
nor U9299 (N_9299,N_9013,N_9060);
or U9300 (N_9300,N_9216,N_9015);
and U9301 (N_9301,N_9034,N_9019);
xor U9302 (N_9302,N_9162,N_9080);
and U9303 (N_9303,N_9067,N_9238);
or U9304 (N_9304,N_9226,N_9215);
or U9305 (N_9305,N_9109,N_9169);
nor U9306 (N_9306,N_9022,N_9143);
and U9307 (N_9307,N_9245,N_9204);
and U9308 (N_9308,N_9017,N_9036);
nor U9309 (N_9309,N_9018,N_9119);
nand U9310 (N_9310,N_9134,N_9088);
nor U9311 (N_9311,N_9247,N_9129);
and U9312 (N_9312,N_9051,N_9011);
nand U9313 (N_9313,N_9009,N_9234);
nand U9314 (N_9314,N_9240,N_9133);
xor U9315 (N_9315,N_9032,N_9230);
xor U9316 (N_9316,N_9210,N_9183);
and U9317 (N_9317,N_9111,N_9182);
nand U9318 (N_9318,N_9087,N_9221);
and U9319 (N_9319,N_9086,N_9116);
nor U9320 (N_9320,N_9224,N_9077);
nor U9321 (N_9321,N_9001,N_9149);
nor U9322 (N_9322,N_9138,N_9023);
and U9323 (N_9323,N_9106,N_9052);
or U9324 (N_9324,N_9042,N_9101);
or U9325 (N_9325,N_9171,N_9033);
nand U9326 (N_9326,N_9135,N_9027);
or U9327 (N_9327,N_9154,N_9229);
nand U9328 (N_9328,N_9095,N_9014);
and U9329 (N_9329,N_9099,N_9110);
nor U9330 (N_9330,N_9082,N_9118);
and U9331 (N_9331,N_9089,N_9214);
xor U9332 (N_9332,N_9170,N_9173);
or U9333 (N_9333,N_9115,N_9122);
xor U9334 (N_9334,N_9041,N_9184);
nand U9335 (N_9335,N_9102,N_9079);
and U9336 (N_9336,N_9249,N_9172);
and U9337 (N_9337,N_9244,N_9242);
nor U9338 (N_9338,N_9188,N_9084);
nand U9339 (N_9339,N_9243,N_9029);
nand U9340 (N_9340,N_9220,N_9125);
and U9341 (N_9341,N_9048,N_9072);
nor U9342 (N_9342,N_9076,N_9055);
nand U9343 (N_9343,N_9241,N_9069);
or U9344 (N_9344,N_9024,N_9236);
nand U9345 (N_9345,N_9123,N_9081);
and U9346 (N_9346,N_9160,N_9092);
or U9347 (N_9347,N_9209,N_9065);
nor U9348 (N_9348,N_9074,N_9181);
and U9349 (N_9349,N_9146,N_9219);
and U9350 (N_9350,N_9044,N_9237);
and U9351 (N_9351,N_9211,N_9227);
nor U9352 (N_9352,N_9025,N_9177);
and U9353 (N_9353,N_9199,N_9232);
xor U9354 (N_9354,N_9126,N_9039);
nand U9355 (N_9355,N_9054,N_9097);
and U9356 (N_9356,N_9148,N_9006);
and U9357 (N_9357,N_9239,N_9165);
xnor U9358 (N_9358,N_9141,N_9218);
nand U9359 (N_9359,N_9186,N_9152);
and U9360 (N_9360,N_9043,N_9050);
nor U9361 (N_9361,N_9153,N_9198);
nor U9362 (N_9362,N_9140,N_9035);
or U9363 (N_9363,N_9062,N_9151);
nor U9364 (N_9364,N_9167,N_9053);
or U9365 (N_9365,N_9185,N_9191);
xor U9366 (N_9366,N_9096,N_9222);
nor U9367 (N_9367,N_9180,N_9194);
nand U9368 (N_9368,N_9117,N_9070);
and U9369 (N_9369,N_9142,N_9049);
nor U9370 (N_9370,N_9206,N_9144);
nand U9371 (N_9371,N_9130,N_9200);
nand U9372 (N_9372,N_9225,N_9114);
nand U9373 (N_9373,N_9085,N_9068);
nand U9374 (N_9374,N_9038,N_9174);
nand U9375 (N_9375,N_9070,N_9247);
or U9376 (N_9376,N_9063,N_9237);
xor U9377 (N_9377,N_9125,N_9086);
nor U9378 (N_9378,N_9131,N_9234);
nand U9379 (N_9379,N_9043,N_9072);
nor U9380 (N_9380,N_9006,N_9127);
and U9381 (N_9381,N_9125,N_9153);
and U9382 (N_9382,N_9152,N_9004);
xnor U9383 (N_9383,N_9087,N_9053);
or U9384 (N_9384,N_9120,N_9024);
xor U9385 (N_9385,N_9232,N_9210);
and U9386 (N_9386,N_9112,N_9118);
nand U9387 (N_9387,N_9075,N_9180);
nor U9388 (N_9388,N_9072,N_9178);
and U9389 (N_9389,N_9185,N_9092);
and U9390 (N_9390,N_9116,N_9180);
or U9391 (N_9391,N_9173,N_9180);
nor U9392 (N_9392,N_9046,N_9093);
xnor U9393 (N_9393,N_9049,N_9008);
and U9394 (N_9394,N_9109,N_9086);
nand U9395 (N_9395,N_9064,N_9222);
nor U9396 (N_9396,N_9081,N_9066);
xor U9397 (N_9397,N_9121,N_9048);
or U9398 (N_9398,N_9242,N_9206);
nor U9399 (N_9399,N_9149,N_9047);
and U9400 (N_9400,N_9219,N_9181);
nand U9401 (N_9401,N_9097,N_9125);
and U9402 (N_9402,N_9126,N_9213);
xor U9403 (N_9403,N_9193,N_9124);
or U9404 (N_9404,N_9036,N_9183);
nand U9405 (N_9405,N_9022,N_9190);
xor U9406 (N_9406,N_9225,N_9044);
or U9407 (N_9407,N_9097,N_9175);
or U9408 (N_9408,N_9043,N_9197);
xor U9409 (N_9409,N_9100,N_9246);
and U9410 (N_9410,N_9198,N_9050);
and U9411 (N_9411,N_9248,N_9118);
or U9412 (N_9412,N_9043,N_9144);
nor U9413 (N_9413,N_9066,N_9204);
or U9414 (N_9414,N_9051,N_9016);
nand U9415 (N_9415,N_9235,N_9248);
and U9416 (N_9416,N_9044,N_9024);
or U9417 (N_9417,N_9060,N_9131);
xor U9418 (N_9418,N_9183,N_9122);
nor U9419 (N_9419,N_9007,N_9191);
xor U9420 (N_9420,N_9145,N_9110);
nor U9421 (N_9421,N_9044,N_9052);
or U9422 (N_9422,N_9178,N_9040);
and U9423 (N_9423,N_9017,N_9038);
and U9424 (N_9424,N_9229,N_9060);
or U9425 (N_9425,N_9124,N_9231);
xnor U9426 (N_9426,N_9201,N_9156);
and U9427 (N_9427,N_9123,N_9125);
xor U9428 (N_9428,N_9000,N_9064);
or U9429 (N_9429,N_9132,N_9076);
or U9430 (N_9430,N_9027,N_9099);
xor U9431 (N_9431,N_9094,N_9063);
nand U9432 (N_9432,N_9212,N_9231);
nand U9433 (N_9433,N_9007,N_9248);
nand U9434 (N_9434,N_9084,N_9080);
xor U9435 (N_9435,N_9088,N_9068);
xor U9436 (N_9436,N_9231,N_9102);
or U9437 (N_9437,N_9150,N_9033);
and U9438 (N_9438,N_9068,N_9195);
or U9439 (N_9439,N_9114,N_9158);
nor U9440 (N_9440,N_9176,N_9063);
nand U9441 (N_9441,N_9103,N_9155);
or U9442 (N_9442,N_9033,N_9160);
nor U9443 (N_9443,N_9177,N_9004);
nand U9444 (N_9444,N_9232,N_9167);
xor U9445 (N_9445,N_9059,N_9014);
and U9446 (N_9446,N_9129,N_9188);
or U9447 (N_9447,N_9214,N_9142);
xor U9448 (N_9448,N_9215,N_9232);
and U9449 (N_9449,N_9120,N_9125);
nor U9450 (N_9450,N_9174,N_9142);
nand U9451 (N_9451,N_9074,N_9152);
and U9452 (N_9452,N_9165,N_9033);
xnor U9453 (N_9453,N_9248,N_9003);
and U9454 (N_9454,N_9000,N_9115);
nand U9455 (N_9455,N_9159,N_9180);
nor U9456 (N_9456,N_9010,N_9167);
or U9457 (N_9457,N_9232,N_9233);
nor U9458 (N_9458,N_9099,N_9015);
xnor U9459 (N_9459,N_9233,N_9168);
nand U9460 (N_9460,N_9097,N_9196);
and U9461 (N_9461,N_9065,N_9088);
nand U9462 (N_9462,N_9241,N_9095);
or U9463 (N_9463,N_9005,N_9212);
or U9464 (N_9464,N_9118,N_9005);
nand U9465 (N_9465,N_9203,N_9242);
or U9466 (N_9466,N_9128,N_9024);
nor U9467 (N_9467,N_9208,N_9089);
or U9468 (N_9468,N_9091,N_9217);
or U9469 (N_9469,N_9200,N_9102);
xnor U9470 (N_9470,N_9237,N_9124);
xnor U9471 (N_9471,N_9144,N_9182);
nand U9472 (N_9472,N_9002,N_9208);
nor U9473 (N_9473,N_9233,N_9000);
xor U9474 (N_9474,N_9175,N_9245);
or U9475 (N_9475,N_9143,N_9012);
xor U9476 (N_9476,N_9137,N_9041);
or U9477 (N_9477,N_9214,N_9139);
nor U9478 (N_9478,N_9241,N_9072);
or U9479 (N_9479,N_9200,N_9146);
and U9480 (N_9480,N_9178,N_9200);
and U9481 (N_9481,N_9226,N_9090);
nand U9482 (N_9482,N_9214,N_9105);
nand U9483 (N_9483,N_9198,N_9214);
nand U9484 (N_9484,N_9203,N_9207);
or U9485 (N_9485,N_9150,N_9039);
xor U9486 (N_9486,N_9143,N_9211);
xnor U9487 (N_9487,N_9018,N_9059);
and U9488 (N_9488,N_9047,N_9134);
and U9489 (N_9489,N_9039,N_9241);
nand U9490 (N_9490,N_9095,N_9194);
xnor U9491 (N_9491,N_9047,N_9233);
nor U9492 (N_9492,N_9248,N_9021);
and U9493 (N_9493,N_9129,N_9139);
nor U9494 (N_9494,N_9097,N_9112);
nor U9495 (N_9495,N_9098,N_9193);
nand U9496 (N_9496,N_9213,N_9128);
or U9497 (N_9497,N_9030,N_9066);
or U9498 (N_9498,N_9194,N_9128);
xnor U9499 (N_9499,N_9085,N_9047);
nor U9500 (N_9500,N_9424,N_9255);
or U9501 (N_9501,N_9263,N_9326);
xnor U9502 (N_9502,N_9496,N_9342);
nand U9503 (N_9503,N_9406,N_9468);
nand U9504 (N_9504,N_9315,N_9266);
or U9505 (N_9505,N_9412,N_9321);
or U9506 (N_9506,N_9498,N_9331);
nor U9507 (N_9507,N_9335,N_9323);
xor U9508 (N_9508,N_9257,N_9332);
and U9509 (N_9509,N_9491,N_9402);
xor U9510 (N_9510,N_9314,N_9298);
and U9511 (N_9511,N_9436,N_9419);
or U9512 (N_9512,N_9297,N_9482);
and U9513 (N_9513,N_9432,N_9348);
nand U9514 (N_9514,N_9413,N_9281);
nor U9515 (N_9515,N_9429,N_9327);
nand U9516 (N_9516,N_9428,N_9350);
nand U9517 (N_9517,N_9441,N_9273);
xnor U9518 (N_9518,N_9489,N_9380);
xnor U9519 (N_9519,N_9279,N_9269);
or U9520 (N_9520,N_9365,N_9361);
nand U9521 (N_9521,N_9336,N_9448);
and U9522 (N_9522,N_9345,N_9346);
xnor U9523 (N_9523,N_9292,N_9253);
or U9524 (N_9524,N_9392,N_9294);
and U9525 (N_9525,N_9304,N_9311);
nand U9526 (N_9526,N_9407,N_9290);
nor U9527 (N_9527,N_9264,N_9289);
xnor U9528 (N_9528,N_9453,N_9283);
xnor U9529 (N_9529,N_9459,N_9357);
nand U9530 (N_9530,N_9285,N_9438);
xnor U9531 (N_9531,N_9486,N_9389);
nor U9532 (N_9532,N_9379,N_9494);
nand U9533 (N_9533,N_9296,N_9262);
nand U9534 (N_9534,N_9464,N_9352);
and U9535 (N_9535,N_9261,N_9347);
nor U9536 (N_9536,N_9369,N_9287);
nand U9537 (N_9537,N_9470,N_9268);
xnor U9538 (N_9538,N_9394,N_9386);
or U9539 (N_9539,N_9343,N_9322);
nand U9540 (N_9540,N_9473,N_9267);
nor U9541 (N_9541,N_9434,N_9404);
or U9542 (N_9542,N_9420,N_9320);
nand U9543 (N_9543,N_9480,N_9403);
xor U9544 (N_9544,N_9272,N_9339);
nor U9545 (N_9545,N_9445,N_9463);
xnor U9546 (N_9546,N_9430,N_9373);
xor U9547 (N_9547,N_9274,N_9426);
and U9548 (N_9548,N_9368,N_9443);
or U9549 (N_9549,N_9446,N_9461);
nand U9550 (N_9550,N_9308,N_9467);
and U9551 (N_9551,N_9252,N_9431);
nor U9552 (N_9552,N_9395,N_9447);
or U9553 (N_9553,N_9405,N_9258);
xor U9554 (N_9554,N_9301,N_9425);
nand U9555 (N_9555,N_9449,N_9318);
and U9556 (N_9556,N_9276,N_9417);
nor U9557 (N_9557,N_9465,N_9495);
and U9558 (N_9558,N_9400,N_9251);
and U9559 (N_9559,N_9398,N_9329);
nand U9560 (N_9560,N_9487,N_9362);
or U9561 (N_9561,N_9344,N_9370);
or U9562 (N_9562,N_9367,N_9377);
and U9563 (N_9563,N_9390,N_9401);
nor U9564 (N_9564,N_9422,N_9359);
nand U9565 (N_9565,N_9456,N_9440);
and U9566 (N_9566,N_9260,N_9375);
or U9567 (N_9567,N_9391,N_9305);
and U9568 (N_9568,N_9397,N_9310);
nand U9569 (N_9569,N_9475,N_9421);
nand U9570 (N_9570,N_9499,N_9372);
and U9571 (N_9571,N_9270,N_9312);
nor U9572 (N_9572,N_9313,N_9460);
nand U9573 (N_9573,N_9490,N_9277);
xnor U9574 (N_9574,N_9280,N_9250);
or U9575 (N_9575,N_9358,N_9484);
nor U9576 (N_9576,N_9286,N_9493);
or U9577 (N_9577,N_9488,N_9408);
xor U9578 (N_9578,N_9334,N_9317);
and U9579 (N_9579,N_9471,N_9374);
or U9580 (N_9580,N_9256,N_9437);
and U9581 (N_9581,N_9457,N_9485);
or U9582 (N_9582,N_9450,N_9384);
xor U9583 (N_9583,N_9462,N_9416);
or U9584 (N_9584,N_9415,N_9492);
nand U9585 (N_9585,N_9458,N_9309);
or U9586 (N_9586,N_9444,N_9481);
or U9587 (N_9587,N_9371,N_9385);
and U9588 (N_9588,N_9483,N_9288);
or U9589 (N_9589,N_9338,N_9469);
nor U9590 (N_9590,N_9254,N_9410);
or U9591 (N_9591,N_9376,N_9478);
nor U9592 (N_9592,N_9455,N_9306);
nor U9593 (N_9593,N_9423,N_9300);
xnor U9594 (N_9594,N_9466,N_9328);
nand U9595 (N_9595,N_9452,N_9497);
nand U9596 (N_9596,N_9387,N_9340);
and U9597 (N_9597,N_9477,N_9325);
and U9598 (N_9598,N_9479,N_9442);
or U9599 (N_9599,N_9299,N_9472);
nor U9600 (N_9600,N_9378,N_9454);
nor U9601 (N_9601,N_9265,N_9364);
xor U9602 (N_9602,N_9316,N_9302);
nor U9603 (N_9603,N_9259,N_9330);
or U9604 (N_9604,N_9381,N_9319);
xor U9605 (N_9605,N_9293,N_9278);
and U9606 (N_9606,N_9476,N_9356);
and U9607 (N_9607,N_9303,N_9282);
nand U9608 (N_9608,N_9399,N_9353);
nand U9609 (N_9609,N_9355,N_9409);
nor U9610 (N_9610,N_9324,N_9451);
and U9611 (N_9611,N_9435,N_9351);
or U9612 (N_9612,N_9284,N_9393);
and U9613 (N_9613,N_9349,N_9414);
nand U9614 (N_9614,N_9333,N_9360);
xor U9615 (N_9615,N_9427,N_9271);
or U9616 (N_9616,N_9396,N_9337);
or U9617 (N_9617,N_9341,N_9433);
and U9618 (N_9618,N_9291,N_9295);
nor U9619 (N_9619,N_9388,N_9382);
nor U9620 (N_9620,N_9411,N_9363);
nand U9621 (N_9621,N_9366,N_9383);
nor U9622 (N_9622,N_9307,N_9474);
xnor U9623 (N_9623,N_9418,N_9275);
xnor U9624 (N_9624,N_9439,N_9354);
nand U9625 (N_9625,N_9356,N_9421);
nand U9626 (N_9626,N_9252,N_9380);
and U9627 (N_9627,N_9287,N_9496);
xor U9628 (N_9628,N_9264,N_9344);
and U9629 (N_9629,N_9357,N_9476);
xnor U9630 (N_9630,N_9276,N_9361);
xor U9631 (N_9631,N_9454,N_9305);
and U9632 (N_9632,N_9350,N_9412);
and U9633 (N_9633,N_9280,N_9440);
nand U9634 (N_9634,N_9407,N_9346);
and U9635 (N_9635,N_9354,N_9272);
nor U9636 (N_9636,N_9488,N_9298);
nand U9637 (N_9637,N_9318,N_9386);
xor U9638 (N_9638,N_9492,N_9263);
nand U9639 (N_9639,N_9262,N_9450);
or U9640 (N_9640,N_9477,N_9395);
nand U9641 (N_9641,N_9429,N_9273);
nor U9642 (N_9642,N_9386,N_9350);
or U9643 (N_9643,N_9310,N_9416);
and U9644 (N_9644,N_9414,N_9291);
xor U9645 (N_9645,N_9277,N_9473);
xnor U9646 (N_9646,N_9401,N_9385);
nor U9647 (N_9647,N_9288,N_9332);
or U9648 (N_9648,N_9283,N_9388);
and U9649 (N_9649,N_9351,N_9279);
nor U9650 (N_9650,N_9293,N_9373);
or U9651 (N_9651,N_9301,N_9376);
nand U9652 (N_9652,N_9368,N_9317);
xnor U9653 (N_9653,N_9428,N_9395);
xnor U9654 (N_9654,N_9289,N_9273);
or U9655 (N_9655,N_9252,N_9433);
nand U9656 (N_9656,N_9496,N_9373);
nand U9657 (N_9657,N_9359,N_9480);
xor U9658 (N_9658,N_9437,N_9376);
or U9659 (N_9659,N_9443,N_9285);
nand U9660 (N_9660,N_9361,N_9291);
nand U9661 (N_9661,N_9393,N_9422);
nor U9662 (N_9662,N_9369,N_9417);
nor U9663 (N_9663,N_9303,N_9338);
nand U9664 (N_9664,N_9472,N_9470);
nand U9665 (N_9665,N_9309,N_9359);
or U9666 (N_9666,N_9259,N_9262);
nand U9667 (N_9667,N_9351,N_9363);
nand U9668 (N_9668,N_9343,N_9288);
nor U9669 (N_9669,N_9273,N_9496);
and U9670 (N_9670,N_9498,N_9333);
nand U9671 (N_9671,N_9489,N_9278);
or U9672 (N_9672,N_9325,N_9287);
xnor U9673 (N_9673,N_9468,N_9347);
or U9674 (N_9674,N_9342,N_9283);
or U9675 (N_9675,N_9421,N_9287);
or U9676 (N_9676,N_9414,N_9496);
or U9677 (N_9677,N_9285,N_9429);
xor U9678 (N_9678,N_9334,N_9493);
xor U9679 (N_9679,N_9350,N_9298);
and U9680 (N_9680,N_9376,N_9461);
or U9681 (N_9681,N_9396,N_9493);
nor U9682 (N_9682,N_9386,N_9450);
xnor U9683 (N_9683,N_9291,N_9370);
and U9684 (N_9684,N_9334,N_9288);
xnor U9685 (N_9685,N_9454,N_9370);
nand U9686 (N_9686,N_9485,N_9423);
and U9687 (N_9687,N_9309,N_9417);
and U9688 (N_9688,N_9398,N_9445);
xnor U9689 (N_9689,N_9276,N_9314);
xor U9690 (N_9690,N_9443,N_9301);
and U9691 (N_9691,N_9306,N_9385);
or U9692 (N_9692,N_9346,N_9425);
nor U9693 (N_9693,N_9354,N_9468);
xor U9694 (N_9694,N_9496,N_9408);
or U9695 (N_9695,N_9257,N_9442);
xnor U9696 (N_9696,N_9369,N_9472);
xnor U9697 (N_9697,N_9305,N_9465);
and U9698 (N_9698,N_9420,N_9378);
nor U9699 (N_9699,N_9297,N_9465);
xnor U9700 (N_9700,N_9428,N_9275);
or U9701 (N_9701,N_9338,N_9257);
nor U9702 (N_9702,N_9387,N_9426);
and U9703 (N_9703,N_9425,N_9370);
nand U9704 (N_9704,N_9308,N_9337);
and U9705 (N_9705,N_9439,N_9343);
and U9706 (N_9706,N_9390,N_9452);
nor U9707 (N_9707,N_9389,N_9418);
or U9708 (N_9708,N_9367,N_9279);
and U9709 (N_9709,N_9357,N_9350);
and U9710 (N_9710,N_9314,N_9426);
or U9711 (N_9711,N_9444,N_9294);
nand U9712 (N_9712,N_9458,N_9456);
and U9713 (N_9713,N_9417,N_9404);
and U9714 (N_9714,N_9454,N_9436);
or U9715 (N_9715,N_9430,N_9476);
or U9716 (N_9716,N_9348,N_9315);
nor U9717 (N_9717,N_9407,N_9374);
nor U9718 (N_9718,N_9366,N_9392);
nand U9719 (N_9719,N_9395,N_9361);
and U9720 (N_9720,N_9359,N_9299);
xor U9721 (N_9721,N_9466,N_9346);
nor U9722 (N_9722,N_9346,N_9421);
nor U9723 (N_9723,N_9453,N_9357);
xnor U9724 (N_9724,N_9420,N_9333);
nand U9725 (N_9725,N_9352,N_9469);
nand U9726 (N_9726,N_9292,N_9430);
nor U9727 (N_9727,N_9458,N_9433);
xnor U9728 (N_9728,N_9278,N_9442);
xor U9729 (N_9729,N_9433,N_9393);
nand U9730 (N_9730,N_9460,N_9396);
and U9731 (N_9731,N_9292,N_9296);
xnor U9732 (N_9732,N_9478,N_9445);
nand U9733 (N_9733,N_9389,N_9448);
and U9734 (N_9734,N_9328,N_9388);
and U9735 (N_9735,N_9432,N_9381);
nand U9736 (N_9736,N_9468,N_9319);
or U9737 (N_9737,N_9379,N_9260);
nor U9738 (N_9738,N_9358,N_9493);
nor U9739 (N_9739,N_9491,N_9393);
and U9740 (N_9740,N_9371,N_9389);
xor U9741 (N_9741,N_9268,N_9389);
nand U9742 (N_9742,N_9467,N_9273);
xor U9743 (N_9743,N_9444,N_9418);
nand U9744 (N_9744,N_9259,N_9294);
nand U9745 (N_9745,N_9285,N_9474);
or U9746 (N_9746,N_9461,N_9454);
or U9747 (N_9747,N_9499,N_9426);
nor U9748 (N_9748,N_9482,N_9290);
or U9749 (N_9749,N_9367,N_9337);
or U9750 (N_9750,N_9500,N_9745);
nand U9751 (N_9751,N_9697,N_9569);
xor U9752 (N_9752,N_9547,N_9715);
nand U9753 (N_9753,N_9650,N_9657);
nor U9754 (N_9754,N_9574,N_9624);
nand U9755 (N_9755,N_9572,N_9519);
nand U9756 (N_9756,N_9638,N_9730);
xor U9757 (N_9757,N_9501,N_9557);
xnor U9758 (N_9758,N_9734,N_9568);
nand U9759 (N_9759,N_9582,N_9630);
nand U9760 (N_9760,N_9720,N_9728);
xor U9761 (N_9761,N_9552,N_9513);
xor U9762 (N_9762,N_9604,N_9558);
and U9763 (N_9763,N_9725,N_9690);
nor U9764 (N_9764,N_9625,N_9525);
or U9765 (N_9765,N_9660,N_9607);
or U9766 (N_9766,N_9692,N_9649);
and U9767 (N_9767,N_9531,N_9546);
nor U9768 (N_9768,N_9696,N_9590);
nor U9769 (N_9769,N_9645,N_9623);
nor U9770 (N_9770,N_9526,N_9654);
nor U9771 (N_9771,N_9632,N_9661);
nand U9772 (N_9772,N_9567,N_9549);
nor U9773 (N_9773,N_9676,N_9640);
and U9774 (N_9774,N_9586,N_9608);
and U9775 (N_9775,N_9707,N_9641);
nand U9776 (N_9776,N_9562,N_9612);
nand U9777 (N_9777,N_9556,N_9721);
xor U9778 (N_9778,N_9711,N_9603);
nand U9779 (N_9779,N_9701,N_9744);
or U9780 (N_9780,N_9722,N_9702);
or U9781 (N_9781,N_9663,N_9600);
nand U9782 (N_9782,N_9714,N_9679);
nand U9783 (N_9783,N_9597,N_9550);
nor U9784 (N_9784,N_9735,N_9646);
nand U9785 (N_9785,N_9621,N_9723);
nor U9786 (N_9786,N_9553,N_9512);
and U9787 (N_9787,N_9741,N_9508);
xor U9788 (N_9788,N_9626,N_9566);
nor U9789 (N_9789,N_9554,N_9509);
nand U9790 (N_9790,N_9505,N_9511);
xnor U9791 (N_9791,N_9693,N_9529);
xnor U9792 (N_9792,N_9743,N_9565);
and U9793 (N_9793,N_9610,N_9524);
nor U9794 (N_9794,N_9631,N_9680);
nand U9795 (N_9795,N_9536,N_9606);
and U9796 (N_9796,N_9635,N_9618);
nor U9797 (N_9797,N_9732,N_9539);
xor U9798 (N_9798,N_9592,N_9644);
and U9799 (N_9799,N_9619,N_9677);
or U9800 (N_9800,N_9598,N_9520);
nor U9801 (N_9801,N_9543,N_9545);
xnor U9802 (N_9802,N_9541,N_9736);
or U9803 (N_9803,N_9538,N_9577);
xnor U9804 (N_9804,N_9749,N_9727);
nand U9805 (N_9805,N_9652,N_9616);
nor U9806 (N_9806,N_9533,N_9578);
and U9807 (N_9807,N_9601,N_9561);
nor U9808 (N_9808,N_9563,N_9564);
and U9809 (N_9809,N_9684,N_9651);
xor U9810 (N_9810,N_9605,N_9587);
xor U9811 (N_9811,N_9589,N_9689);
and U9812 (N_9812,N_9682,N_9705);
and U9813 (N_9813,N_9602,N_9738);
nor U9814 (N_9814,N_9609,N_9615);
and U9815 (N_9815,N_9585,N_9662);
nor U9816 (N_9816,N_9570,N_9724);
xnor U9817 (N_9817,N_9523,N_9530);
nand U9818 (N_9818,N_9614,N_9559);
or U9819 (N_9819,N_9656,N_9670);
xnor U9820 (N_9820,N_9703,N_9528);
xor U9821 (N_9821,N_9726,N_9532);
xor U9822 (N_9822,N_9731,N_9594);
nor U9823 (N_9823,N_9622,N_9687);
or U9824 (N_9824,N_9571,N_9573);
nand U9825 (N_9825,N_9713,N_9746);
nand U9826 (N_9826,N_9542,N_9580);
or U9827 (N_9827,N_9748,N_9637);
nand U9828 (N_9828,N_9686,N_9504);
xnor U9829 (N_9829,N_9659,N_9584);
and U9830 (N_9830,N_9678,N_9716);
nor U9831 (N_9831,N_9629,N_9555);
nor U9832 (N_9832,N_9611,N_9522);
xor U9833 (N_9833,N_9515,N_9516);
or U9834 (N_9834,N_9503,N_9648);
or U9835 (N_9835,N_9636,N_9737);
xnor U9836 (N_9836,N_9643,N_9665);
nor U9837 (N_9837,N_9583,N_9627);
xor U9838 (N_9838,N_9642,N_9708);
nand U9839 (N_9839,N_9514,N_9639);
and U9840 (N_9840,N_9595,N_9667);
and U9841 (N_9841,N_9706,N_9634);
nor U9842 (N_9842,N_9633,N_9694);
nor U9843 (N_9843,N_9695,N_9527);
xnor U9844 (N_9844,N_9506,N_9588);
or U9845 (N_9845,N_9698,N_9647);
xnor U9846 (N_9846,N_9709,N_9719);
xor U9847 (N_9847,N_9540,N_9518);
and U9848 (N_9848,N_9733,N_9718);
xnor U9849 (N_9849,N_9537,N_9658);
xor U9850 (N_9850,N_9674,N_9683);
and U9851 (N_9851,N_9510,N_9628);
or U9852 (N_9852,N_9613,N_9681);
nor U9853 (N_9853,N_9581,N_9653);
nor U9854 (N_9854,N_9669,N_9675);
nand U9855 (N_9855,N_9579,N_9699);
xnor U9856 (N_9856,N_9671,N_9544);
nand U9857 (N_9857,N_9535,N_9666);
nand U9858 (N_9858,N_9691,N_9502);
nand U9859 (N_9859,N_9576,N_9688);
or U9860 (N_9860,N_9710,N_9620);
xnor U9861 (N_9861,N_9717,N_9596);
nand U9862 (N_9862,N_9593,N_9617);
xnor U9863 (N_9863,N_9704,N_9672);
or U9864 (N_9864,N_9712,N_9521);
xor U9865 (N_9865,N_9517,N_9685);
xor U9866 (N_9866,N_9655,N_9560);
or U9867 (N_9867,N_9747,N_9700);
xnor U9868 (N_9868,N_9534,N_9739);
nand U9869 (N_9869,N_9673,N_9599);
nor U9870 (N_9870,N_9729,N_9664);
nor U9871 (N_9871,N_9740,N_9742);
nand U9872 (N_9872,N_9551,N_9575);
or U9873 (N_9873,N_9548,N_9591);
nand U9874 (N_9874,N_9507,N_9668);
and U9875 (N_9875,N_9624,N_9733);
or U9876 (N_9876,N_9701,N_9523);
nand U9877 (N_9877,N_9706,N_9557);
or U9878 (N_9878,N_9695,N_9743);
or U9879 (N_9879,N_9507,N_9707);
nand U9880 (N_9880,N_9738,N_9619);
xnor U9881 (N_9881,N_9721,N_9679);
and U9882 (N_9882,N_9682,N_9577);
xnor U9883 (N_9883,N_9730,N_9526);
or U9884 (N_9884,N_9514,N_9678);
or U9885 (N_9885,N_9613,N_9556);
or U9886 (N_9886,N_9678,N_9695);
xor U9887 (N_9887,N_9662,N_9710);
nor U9888 (N_9888,N_9624,N_9712);
or U9889 (N_9889,N_9556,N_9515);
and U9890 (N_9890,N_9601,N_9588);
xor U9891 (N_9891,N_9610,N_9679);
xnor U9892 (N_9892,N_9626,N_9744);
or U9893 (N_9893,N_9655,N_9721);
nor U9894 (N_9894,N_9583,N_9590);
nor U9895 (N_9895,N_9629,N_9571);
nor U9896 (N_9896,N_9742,N_9744);
xnor U9897 (N_9897,N_9688,N_9556);
nand U9898 (N_9898,N_9659,N_9594);
xnor U9899 (N_9899,N_9652,N_9598);
xnor U9900 (N_9900,N_9609,N_9664);
nand U9901 (N_9901,N_9559,N_9530);
or U9902 (N_9902,N_9720,N_9624);
xor U9903 (N_9903,N_9545,N_9748);
nor U9904 (N_9904,N_9729,N_9500);
nor U9905 (N_9905,N_9599,N_9693);
nor U9906 (N_9906,N_9580,N_9512);
nand U9907 (N_9907,N_9735,N_9526);
and U9908 (N_9908,N_9658,N_9732);
nand U9909 (N_9909,N_9553,N_9640);
nand U9910 (N_9910,N_9665,N_9636);
nor U9911 (N_9911,N_9578,N_9598);
or U9912 (N_9912,N_9736,N_9545);
nand U9913 (N_9913,N_9566,N_9661);
or U9914 (N_9914,N_9738,N_9546);
or U9915 (N_9915,N_9716,N_9535);
and U9916 (N_9916,N_9530,N_9544);
or U9917 (N_9917,N_9537,N_9711);
or U9918 (N_9918,N_9578,N_9713);
nand U9919 (N_9919,N_9719,N_9689);
and U9920 (N_9920,N_9609,N_9559);
xnor U9921 (N_9921,N_9733,N_9615);
xnor U9922 (N_9922,N_9597,N_9731);
xor U9923 (N_9923,N_9707,N_9653);
and U9924 (N_9924,N_9643,N_9545);
or U9925 (N_9925,N_9517,N_9600);
and U9926 (N_9926,N_9519,N_9723);
xnor U9927 (N_9927,N_9668,N_9581);
xnor U9928 (N_9928,N_9714,N_9600);
nand U9929 (N_9929,N_9704,N_9639);
nor U9930 (N_9930,N_9555,N_9594);
or U9931 (N_9931,N_9559,N_9687);
nand U9932 (N_9932,N_9731,N_9632);
nand U9933 (N_9933,N_9708,N_9600);
xnor U9934 (N_9934,N_9657,N_9726);
or U9935 (N_9935,N_9567,N_9640);
and U9936 (N_9936,N_9615,N_9585);
nor U9937 (N_9937,N_9504,N_9680);
xor U9938 (N_9938,N_9506,N_9580);
nor U9939 (N_9939,N_9676,N_9573);
and U9940 (N_9940,N_9716,N_9608);
nor U9941 (N_9941,N_9522,N_9605);
and U9942 (N_9942,N_9719,N_9582);
nand U9943 (N_9943,N_9532,N_9574);
xnor U9944 (N_9944,N_9561,N_9648);
or U9945 (N_9945,N_9661,N_9616);
nor U9946 (N_9946,N_9715,N_9575);
nor U9947 (N_9947,N_9708,N_9587);
nand U9948 (N_9948,N_9722,N_9644);
or U9949 (N_9949,N_9701,N_9541);
nand U9950 (N_9950,N_9580,N_9725);
xor U9951 (N_9951,N_9688,N_9587);
nor U9952 (N_9952,N_9611,N_9588);
xnor U9953 (N_9953,N_9693,N_9612);
nand U9954 (N_9954,N_9655,N_9533);
xor U9955 (N_9955,N_9679,N_9727);
nor U9956 (N_9956,N_9548,N_9574);
or U9957 (N_9957,N_9648,N_9714);
and U9958 (N_9958,N_9613,N_9540);
or U9959 (N_9959,N_9708,N_9537);
nand U9960 (N_9960,N_9716,N_9573);
xnor U9961 (N_9961,N_9686,N_9748);
xor U9962 (N_9962,N_9600,N_9622);
xnor U9963 (N_9963,N_9655,N_9608);
nand U9964 (N_9964,N_9542,N_9604);
nor U9965 (N_9965,N_9653,N_9622);
and U9966 (N_9966,N_9563,N_9704);
or U9967 (N_9967,N_9678,N_9594);
or U9968 (N_9968,N_9550,N_9667);
or U9969 (N_9969,N_9612,N_9626);
and U9970 (N_9970,N_9749,N_9581);
or U9971 (N_9971,N_9660,N_9669);
or U9972 (N_9972,N_9537,N_9531);
nand U9973 (N_9973,N_9574,N_9520);
or U9974 (N_9974,N_9576,N_9625);
and U9975 (N_9975,N_9711,N_9674);
nor U9976 (N_9976,N_9703,N_9633);
nor U9977 (N_9977,N_9700,N_9508);
or U9978 (N_9978,N_9634,N_9681);
xor U9979 (N_9979,N_9638,N_9532);
and U9980 (N_9980,N_9739,N_9702);
or U9981 (N_9981,N_9695,N_9579);
or U9982 (N_9982,N_9545,N_9632);
and U9983 (N_9983,N_9715,N_9525);
nor U9984 (N_9984,N_9564,N_9742);
nand U9985 (N_9985,N_9719,N_9516);
and U9986 (N_9986,N_9710,N_9626);
nand U9987 (N_9987,N_9716,N_9655);
and U9988 (N_9988,N_9712,N_9529);
nand U9989 (N_9989,N_9577,N_9681);
and U9990 (N_9990,N_9682,N_9721);
or U9991 (N_9991,N_9670,N_9638);
and U9992 (N_9992,N_9592,N_9706);
nand U9993 (N_9993,N_9559,N_9721);
xor U9994 (N_9994,N_9709,N_9570);
and U9995 (N_9995,N_9634,N_9631);
or U9996 (N_9996,N_9608,N_9587);
or U9997 (N_9997,N_9739,N_9743);
and U9998 (N_9998,N_9530,N_9502);
nor U9999 (N_9999,N_9574,N_9610);
xnor U10000 (N_10000,N_9928,N_9886);
nor U10001 (N_10001,N_9781,N_9973);
xor U10002 (N_10002,N_9846,N_9937);
or U10003 (N_10003,N_9757,N_9858);
nor U10004 (N_10004,N_9870,N_9956);
and U10005 (N_10005,N_9777,N_9950);
xnor U10006 (N_10006,N_9823,N_9821);
or U10007 (N_10007,N_9959,N_9774);
nand U10008 (N_10008,N_9915,N_9944);
or U10009 (N_10009,N_9907,N_9824);
nand U10010 (N_10010,N_9993,N_9790);
nor U10011 (N_10011,N_9912,N_9980);
nand U10012 (N_10012,N_9841,N_9802);
xor U10013 (N_10013,N_9866,N_9987);
nand U10014 (N_10014,N_9854,N_9796);
or U10015 (N_10015,N_9772,N_9815);
xor U10016 (N_10016,N_9831,N_9754);
and U10017 (N_10017,N_9755,N_9779);
xnor U10018 (N_10018,N_9999,N_9951);
and U10019 (N_10019,N_9767,N_9964);
nand U10020 (N_10020,N_9998,N_9863);
and U10021 (N_10021,N_9989,N_9817);
and U10022 (N_10022,N_9942,N_9752);
nor U10023 (N_10023,N_9996,N_9933);
xor U10024 (N_10024,N_9906,N_9893);
nand U10025 (N_10025,N_9939,N_9760);
nand U10026 (N_10026,N_9862,N_9877);
nand U10027 (N_10027,N_9921,N_9968);
and U10028 (N_10028,N_9842,N_9806);
nor U10029 (N_10029,N_9764,N_9927);
nor U10030 (N_10030,N_9851,N_9897);
nor U10031 (N_10031,N_9931,N_9936);
xor U10032 (N_10032,N_9967,N_9888);
xnor U10033 (N_10033,N_9822,N_9799);
and U10034 (N_10034,N_9955,N_9938);
xnor U10035 (N_10035,N_9788,N_9972);
or U10036 (N_10036,N_9830,N_9759);
xnor U10037 (N_10037,N_9920,N_9995);
and U10038 (N_10038,N_9975,N_9868);
xnor U10039 (N_10039,N_9916,N_9768);
xor U10040 (N_10040,N_9874,N_9826);
nand U10041 (N_10041,N_9839,N_9780);
nor U10042 (N_10042,N_9794,N_9840);
nand U10043 (N_10043,N_9895,N_9911);
or U10044 (N_10044,N_9930,N_9843);
nor U10045 (N_10045,N_9983,N_9929);
xnor U10046 (N_10046,N_9940,N_9856);
nand U10047 (N_10047,N_9766,N_9871);
xor U10048 (N_10048,N_9900,N_9855);
or U10049 (N_10049,N_9885,N_9773);
nand U10050 (N_10050,N_9953,N_9905);
or U10051 (N_10051,N_9859,N_9988);
nand U10052 (N_10052,N_9803,N_9876);
and U10053 (N_10053,N_9827,N_9816);
nand U10054 (N_10054,N_9976,N_9879);
nand U10055 (N_10055,N_9808,N_9832);
xnor U10056 (N_10056,N_9994,N_9904);
nor U10057 (N_10057,N_9836,N_9919);
nand U10058 (N_10058,N_9926,N_9801);
and U10059 (N_10059,N_9889,N_9984);
nand U10060 (N_10060,N_9800,N_9834);
nor U10061 (N_10061,N_9902,N_9852);
and U10062 (N_10062,N_9786,N_9974);
nand U10063 (N_10063,N_9761,N_9848);
and U10064 (N_10064,N_9878,N_9835);
or U10065 (N_10065,N_9756,N_9820);
xor U10066 (N_10066,N_9981,N_9966);
nor U10067 (N_10067,N_9833,N_9943);
or U10068 (N_10068,N_9914,N_9785);
and U10069 (N_10069,N_9861,N_9782);
nor U10070 (N_10070,N_9963,N_9997);
and U10071 (N_10071,N_9853,N_9962);
nor U10072 (N_10072,N_9978,N_9810);
or U10073 (N_10073,N_9991,N_9961);
nand U10074 (N_10074,N_9797,N_9946);
nand U10075 (N_10075,N_9908,N_9941);
or U10076 (N_10076,N_9825,N_9947);
nor U10077 (N_10077,N_9898,N_9935);
and U10078 (N_10078,N_9872,N_9882);
and U10079 (N_10079,N_9762,N_9867);
or U10080 (N_10080,N_9804,N_9828);
nor U10081 (N_10081,N_9892,N_9844);
nor U10082 (N_10082,N_9925,N_9857);
xor U10083 (N_10083,N_9783,N_9753);
nor U10084 (N_10084,N_9850,N_9869);
xnor U10085 (N_10085,N_9977,N_9784);
xor U10086 (N_10086,N_9901,N_9865);
nand U10087 (N_10087,N_9812,N_9899);
or U10088 (N_10088,N_9965,N_9880);
xnor U10089 (N_10089,N_9934,N_9917);
nor U10090 (N_10090,N_9918,N_9805);
nand U10091 (N_10091,N_9873,N_9979);
and U10092 (N_10092,N_9948,N_9903);
xor U10093 (N_10093,N_9849,N_9818);
nor U10094 (N_10094,N_9949,N_9985);
or U10095 (N_10095,N_9791,N_9894);
nand U10096 (N_10096,N_9957,N_9798);
and U10097 (N_10097,N_9838,N_9758);
or U10098 (N_10098,N_9795,N_9982);
and U10099 (N_10099,N_9971,N_9891);
and U10100 (N_10100,N_9778,N_9945);
xnor U10101 (N_10101,N_9771,N_9775);
nor U10102 (N_10102,N_9881,N_9884);
or U10103 (N_10103,N_9992,N_9763);
and U10104 (N_10104,N_9807,N_9913);
or U10105 (N_10105,N_9909,N_9932);
nor U10106 (N_10106,N_9793,N_9792);
xor U10107 (N_10107,N_9837,N_9864);
nand U10108 (N_10108,N_9890,N_9910);
or U10109 (N_10109,N_9789,N_9970);
nand U10110 (N_10110,N_9787,N_9960);
xor U10111 (N_10111,N_9952,N_9896);
nand U10112 (N_10112,N_9954,N_9922);
xnor U10113 (N_10113,N_9860,N_9887);
and U10114 (N_10114,N_9819,N_9776);
nand U10115 (N_10115,N_9769,N_9770);
xor U10116 (N_10116,N_9969,N_9845);
and U10117 (N_10117,N_9765,N_9813);
or U10118 (N_10118,N_9958,N_9875);
and U10119 (N_10119,N_9814,N_9811);
nor U10120 (N_10120,N_9923,N_9847);
and U10121 (N_10121,N_9924,N_9990);
nor U10122 (N_10122,N_9750,N_9829);
or U10123 (N_10123,N_9751,N_9986);
xor U10124 (N_10124,N_9809,N_9883);
and U10125 (N_10125,N_9957,N_9993);
nand U10126 (N_10126,N_9843,N_9848);
and U10127 (N_10127,N_9986,N_9850);
or U10128 (N_10128,N_9963,N_9938);
and U10129 (N_10129,N_9779,N_9893);
and U10130 (N_10130,N_9979,N_9832);
nand U10131 (N_10131,N_9836,N_9966);
nand U10132 (N_10132,N_9994,N_9871);
nor U10133 (N_10133,N_9872,N_9970);
or U10134 (N_10134,N_9867,N_9994);
or U10135 (N_10135,N_9907,N_9931);
nand U10136 (N_10136,N_9816,N_9867);
xor U10137 (N_10137,N_9986,N_9908);
xnor U10138 (N_10138,N_9769,N_9879);
nor U10139 (N_10139,N_9998,N_9975);
and U10140 (N_10140,N_9851,N_9959);
or U10141 (N_10141,N_9935,N_9906);
and U10142 (N_10142,N_9761,N_9783);
or U10143 (N_10143,N_9833,N_9791);
xor U10144 (N_10144,N_9952,N_9898);
or U10145 (N_10145,N_9852,N_9954);
and U10146 (N_10146,N_9851,N_9816);
and U10147 (N_10147,N_9954,N_9887);
nand U10148 (N_10148,N_9872,N_9823);
nor U10149 (N_10149,N_9751,N_9797);
nor U10150 (N_10150,N_9936,N_9873);
or U10151 (N_10151,N_9831,N_9758);
nand U10152 (N_10152,N_9772,N_9952);
xnor U10153 (N_10153,N_9775,N_9875);
or U10154 (N_10154,N_9986,N_9911);
nor U10155 (N_10155,N_9930,N_9989);
nand U10156 (N_10156,N_9904,N_9788);
nand U10157 (N_10157,N_9766,N_9910);
or U10158 (N_10158,N_9882,N_9927);
nand U10159 (N_10159,N_9939,N_9940);
nor U10160 (N_10160,N_9882,N_9777);
nand U10161 (N_10161,N_9992,N_9860);
or U10162 (N_10162,N_9955,N_9810);
or U10163 (N_10163,N_9957,N_9845);
and U10164 (N_10164,N_9797,N_9963);
xor U10165 (N_10165,N_9791,N_9785);
and U10166 (N_10166,N_9956,N_9753);
nor U10167 (N_10167,N_9755,N_9762);
and U10168 (N_10168,N_9857,N_9952);
xnor U10169 (N_10169,N_9751,N_9972);
or U10170 (N_10170,N_9762,N_9896);
nand U10171 (N_10171,N_9867,N_9837);
nor U10172 (N_10172,N_9793,N_9759);
nor U10173 (N_10173,N_9802,N_9896);
nor U10174 (N_10174,N_9785,N_9864);
or U10175 (N_10175,N_9839,N_9830);
and U10176 (N_10176,N_9955,N_9948);
xor U10177 (N_10177,N_9799,N_9886);
nand U10178 (N_10178,N_9791,N_9773);
xnor U10179 (N_10179,N_9788,N_9980);
xor U10180 (N_10180,N_9970,N_9845);
nand U10181 (N_10181,N_9751,N_9800);
nor U10182 (N_10182,N_9885,N_9979);
xor U10183 (N_10183,N_9815,N_9944);
nand U10184 (N_10184,N_9843,N_9822);
nand U10185 (N_10185,N_9978,N_9812);
and U10186 (N_10186,N_9959,N_9926);
xor U10187 (N_10187,N_9957,N_9787);
nor U10188 (N_10188,N_9827,N_9757);
xnor U10189 (N_10189,N_9890,N_9780);
or U10190 (N_10190,N_9760,N_9776);
xor U10191 (N_10191,N_9824,N_9761);
nand U10192 (N_10192,N_9769,N_9763);
nand U10193 (N_10193,N_9808,N_9785);
xnor U10194 (N_10194,N_9837,N_9847);
nor U10195 (N_10195,N_9921,N_9868);
xor U10196 (N_10196,N_9984,N_9981);
and U10197 (N_10197,N_9775,N_9925);
and U10198 (N_10198,N_9886,N_9916);
or U10199 (N_10199,N_9912,N_9890);
nor U10200 (N_10200,N_9837,N_9869);
xnor U10201 (N_10201,N_9849,N_9954);
or U10202 (N_10202,N_9897,N_9817);
xnor U10203 (N_10203,N_9952,N_9757);
nor U10204 (N_10204,N_9787,N_9951);
or U10205 (N_10205,N_9793,N_9972);
nor U10206 (N_10206,N_9752,N_9784);
nor U10207 (N_10207,N_9919,N_9759);
nor U10208 (N_10208,N_9889,N_9883);
or U10209 (N_10209,N_9966,N_9806);
or U10210 (N_10210,N_9893,N_9869);
and U10211 (N_10211,N_9886,N_9948);
nor U10212 (N_10212,N_9970,N_9823);
nand U10213 (N_10213,N_9852,N_9811);
nor U10214 (N_10214,N_9985,N_9866);
xor U10215 (N_10215,N_9862,N_9756);
and U10216 (N_10216,N_9782,N_9875);
xnor U10217 (N_10217,N_9764,N_9777);
and U10218 (N_10218,N_9841,N_9756);
or U10219 (N_10219,N_9864,N_9929);
and U10220 (N_10220,N_9855,N_9793);
nand U10221 (N_10221,N_9894,N_9756);
and U10222 (N_10222,N_9924,N_9995);
and U10223 (N_10223,N_9789,N_9928);
nor U10224 (N_10224,N_9819,N_9985);
nor U10225 (N_10225,N_9829,N_9943);
or U10226 (N_10226,N_9931,N_9781);
xnor U10227 (N_10227,N_9813,N_9864);
xor U10228 (N_10228,N_9883,N_9901);
and U10229 (N_10229,N_9757,N_9842);
and U10230 (N_10230,N_9806,N_9950);
and U10231 (N_10231,N_9755,N_9952);
and U10232 (N_10232,N_9879,N_9917);
xnor U10233 (N_10233,N_9902,N_9758);
or U10234 (N_10234,N_9785,N_9783);
or U10235 (N_10235,N_9942,N_9915);
nor U10236 (N_10236,N_9845,N_9777);
nor U10237 (N_10237,N_9809,N_9968);
or U10238 (N_10238,N_9778,N_9912);
nor U10239 (N_10239,N_9929,N_9972);
xor U10240 (N_10240,N_9889,N_9820);
nand U10241 (N_10241,N_9901,N_9910);
xor U10242 (N_10242,N_9842,N_9868);
nand U10243 (N_10243,N_9773,N_9946);
xnor U10244 (N_10244,N_9935,N_9995);
and U10245 (N_10245,N_9921,N_9821);
xor U10246 (N_10246,N_9963,N_9783);
or U10247 (N_10247,N_9955,N_9836);
nand U10248 (N_10248,N_9826,N_9988);
nand U10249 (N_10249,N_9757,N_9885);
nand U10250 (N_10250,N_10187,N_10141);
nand U10251 (N_10251,N_10172,N_10221);
or U10252 (N_10252,N_10129,N_10211);
nor U10253 (N_10253,N_10117,N_10003);
or U10254 (N_10254,N_10208,N_10166);
xnor U10255 (N_10255,N_10138,N_10159);
nor U10256 (N_10256,N_10157,N_10025);
or U10257 (N_10257,N_10073,N_10043);
and U10258 (N_10258,N_10072,N_10191);
and U10259 (N_10259,N_10074,N_10107);
nand U10260 (N_10260,N_10127,N_10203);
nand U10261 (N_10261,N_10177,N_10120);
or U10262 (N_10262,N_10088,N_10012);
nand U10263 (N_10263,N_10122,N_10022);
or U10264 (N_10264,N_10000,N_10091);
xnor U10265 (N_10265,N_10198,N_10086);
xor U10266 (N_10266,N_10100,N_10053);
nand U10267 (N_10267,N_10149,N_10011);
xnor U10268 (N_10268,N_10069,N_10031);
nand U10269 (N_10269,N_10087,N_10225);
or U10270 (N_10270,N_10179,N_10034);
or U10271 (N_10271,N_10089,N_10081);
and U10272 (N_10272,N_10229,N_10170);
xnor U10273 (N_10273,N_10192,N_10212);
nor U10274 (N_10274,N_10215,N_10099);
nand U10275 (N_10275,N_10226,N_10005);
xnor U10276 (N_10276,N_10112,N_10189);
and U10277 (N_10277,N_10180,N_10158);
and U10278 (N_10278,N_10119,N_10249);
or U10279 (N_10279,N_10206,N_10142);
and U10280 (N_10280,N_10101,N_10028);
or U10281 (N_10281,N_10001,N_10181);
xor U10282 (N_10282,N_10106,N_10083);
nand U10283 (N_10283,N_10194,N_10143);
xor U10284 (N_10284,N_10241,N_10248);
nor U10285 (N_10285,N_10111,N_10125);
xnor U10286 (N_10286,N_10118,N_10245);
and U10287 (N_10287,N_10210,N_10048);
or U10288 (N_10288,N_10196,N_10124);
xor U10289 (N_10289,N_10044,N_10244);
or U10290 (N_10290,N_10024,N_10155);
xnor U10291 (N_10291,N_10169,N_10137);
nand U10292 (N_10292,N_10015,N_10193);
xnor U10293 (N_10293,N_10236,N_10200);
or U10294 (N_10294,N_10145,N_10134);
nor U10295 (N_10295,N_10114,N_10183);
or U10296 (N_10296,N_10017,N_10049);
nor U10297 (N_10297,N_10230,N_10063);
nor U10298 (N_10298,N_10080,N_10161);
and U10299 (N_10299,N_10160,N_10057);
or U10300 (N_10300,N_10219,N_10102);
or U10301 (N_10301,N_10110,N_10010);
or U10302 (N_10302,N_10037,N_10235);
nand U10303 (N_10303,N_10078,N_10128);
and U10304 (N_10304,N_10204,N_10123);
nor U10305 (N_10305,N_10202,N_10121);
nor U10306 (N_10306,N_10064,N_10108);
nand U10307 (N_10307,N_10103,N_10041);
and U10308 (N_10308,N_10071,N_10054);
and U10309 (N_10309,N_10116,N_10199);
or U10310 (N_10310,N_10097,N_10197);
xnor U10311 (N_10311,N_10126,N_10239);
nor U10312 (N_10312,N_10154,N_10171);
or U10313 (N_10313,N_10029,N_10018);
and U10314 (N_10314,N_10032,N_10213);
or U10315 (N_10315,N_10228,N_10033);
or U10316 (N_10316,N_10217,N_10077);
or U10317 (N_10317,N_10209,N_10163);
and U10318 (N_10318,N_10195,N_10201);
nand U10319 (N_10319,N_10184,N_10051);
nor U10320 (N_10320,N_10168,N_10045);
nand U10321 (N_10321,N_10167,N_10014);
or U10322 (N_10322,N_10223,N_10079);
nand U10323 (N_10323,N_10098,N_10020);
nand U10324 (N_10324,N_10084,N_10094);
or U10325 (N_10325,N_10027,N_10113);
xnor U10326 (N_10326,N_10040,N_10013);
and U10327 (N_10327,N_10095,N_10038);
nand U10328 (N_10328,N_10058,N_10153);
nand U10329 (N_10329,N_10006,N_10065);
nand U10330 (N_10330,N_10062,N_10021);
nand U10331 (N_10331,N_10234,N_10085);
xnor U10332 (N_10332,N_10061,N_10056);
nor U10333 (N_10333,N_10220,N_10055);
xor U10334 (N_10334,N_10035,N_10232);
nand U10335 (N_10335,N_10009,N_10246);
xnor U10336 (N_10336,N_10115,N_10036);
nor U10337 (N_10337,N_10165,N_10139);
or U10338 (N_10338,N_10075,N_10176);
xnor U10339 (N_10339,N_10218,N_10185);
and U10340 (N_10340,N_10247,N_10136);
nand U10341 (N_10341,N_10090,N_10147);
nor U10342 (N_10342,N_10224,N_10093);
or U10343 (N_10343,N_10214,N_10151);
nor U10344 (N_10344,N_10207,N_10042);
nand U10345 (N_10345,N_10076,N_10131);
nor U10346 (N_10346,N_10070,N_10162);
nand U10347 (N_10347,N_10156,N_10144);
and U10348 (N_10348,N_10233,N_10240);
and U10349 (N_10349,N_10060,N_10109);
and U10350 (N_10350,N_10178,N_10135);
or U10351 (N_10351,N_10002,N_10205);
nor U10352 (N_10352,N_10148,N_10004);
or U10353 (N_10353,N_10243,N_10007);
nand U10354 (N_10354,N_10237,N_10188);
or U10355 (N_10355,N_10146,N_10105);
or U10356 (N_10356,N_10186,N_10238);
or U10357 (N_10357,N_10059,N_10132);
nand U10358 (N_10358,N_10173,N_10133);
and U10359 (N_10359,N_10066,N_10050);
or U10360 (N_10360,N_10222,N_10052);
or U10361 (N_10361,N_10190,N_10216);
and U10362 (N_10362,N_10026,N_10130);
xnor U10363 (N_10363,N_10092,N_10182);
xnor U10364 (N_10364,N_10030,N_10242);
nor U10365 (N_10365,N_10164,N_10175);
xnor U10366 (N_10366,N_10019,N_10152);
xnor U10367 (N_10367,N_10227,N_10067);
xnor U10368 (N_10368,N_10068,N_10096);
or U10369 (N_10369,N_10082,N_10104);
or U10370 (N_10370,N_10023,N_10008);
xnor U10371 (N_10371,N_10150,N_10047);
nor U10372 (N_10372,N_10016,N_10174);
xnor U10373 (N_10373,N_10039,N_10046);
or U10374 (N_10374,N_10140,N_10231);
xor U10375 (N_10375,N_10084,N_10210);
and U10376 (N_10376,N_10076,N_10054);
nor U10377 (N_10377,N_10189,N_10237);
and U10378 (N_10378,N_10085,N_10022);
nor U10379 (N_10379,N_10214,N_10164);
nor U10380 (N_10380,N_10082,N_10080);
nand U10381 (N_10381,N_10077,N_10242);
and U10382 (N_10382,N_10248,N_10003);
or U10383 (N_10383,N_10162,N_10151);
nand U10384 (N_10384,N_10020,N_10022);
or U10385 (N_10385,N_10127,N_10081);
nor U10386 (N_10386,N_10070,N_10186);
nor U10387 (N_10387,N_10164,N_10145);
nor U10388 (N_10388,N_10193,N_10051);
and U10389 (N_10389,N_10006,N_10082);
nor U10390 (N_10390,N_10165,N_10007);
nor U10391 (N_10391,N_10113,N_10233);
nor U10392 (N_10392,N_10195,N_10176);
nand U10393 (N_10393,N_10248,N_10130);
xor U10394 (N_10394,N_10022,N_10100);
or U10395 (N_10395,N_10180,N_10088);
or U10396 (N_10396,N_10182,N_10112);
nor U10397 (N_10397,N_10049,N_10235);
nand U10398 (N_10398,N_10163,N_10036);
nand U10399 (N_10399,N_10135,N_10110);
nor U10400 (N_10400,N_10199,N_10060);
and U10401 (N_10401,N_10196,N_10032);
xor U10402 (N_10402,N_10107,N_10089);
nand U10403 (N_10403,N_10010,N_10219);
nor U10404 (N_10404,N_10113,N_10176);
nor U10405 (N_10405,N_10150,N_10176);
nor U10406 (N_10406,N_10033,N_10145);
nand U10407 (N_10407,N_10191,N_10230);
or U10408 (N_10408,N_10115,N_10035);
or U10409 (N_10409,N_10240,N_10199);
nor U10410 (N_10410,N_10137,N_10009);
or U10411 (N_10411,N_10037,N_10167);
and U10412 (N_10412,N_10036,N_10123);
or U10413 (N_10413,N_10166,N_10145);
nor U10414 (N_10414,N_10148,N_10168);
nand U10415 (N_10415,N_10092,N_10173);
and U10416 (N_10416,N_10085,N_10152);
xor U10417 (N_10417,N_10086,N_10042);
xnor U10418 (N_10418,N_10110,N_10186);
or U10419 (N_10419,N_10103,N_10233);
nor U10420 (N_10420,N_10031,N_10172);
and U10421 (N_10421,N_10222,N_10012);
or U10422 (N_10422,N_10029,N_10013);
or U10423 (N_10423,N_10008,N_10248);
xnor U10424 (N_10424,N_10221,N_10167);
nand U10425 (N_10425,N_10034,N_10150);
xnor U10426 (N_10426,N_10191,N_10149);
nand U10427 (N_10427,N_10222,N_10170);
and U10428 (N_10428,N_10245,N_10013);
and U10429 (N_10429,N_10092,N_10022);
or U10430 (N_10430,N_10051,N_10077);
and U10431 (N_10431,N_10015,N_10200);
and U10432 (N_10432,N_10212,N_10119);
nor U10433 (N_10433,N_10217,N_10111);
xnor U10434 (N_10434,N_10166,N_10211);
or U10435 (N_10435,N_10165,N_10021);
or U10436 (N_10436,N_10248,N_10196);
and U10437 (N_10437,N_10011,N_10118);
and U10438 (N_10438,N_10047,N_10161);
nand U10439 (N_10439,N_10084,N_10169);
or U10440 (N_10440,N_10228,N_10100);
xnor U10441 (N_10441,N_10098,N_10221);
nor U10442 (N_10442,N_10198,N_10080);
or U10443 (N_10443,N_10106,N_10214);
xnor U10444 (N_10444,N_10093,N_10181);
xor U10445 (N_10445,N_10073,N_10047);
nand U10446 (N_10446,N_10204,N_10202);
xnor U10447 (N_10447,N_10165,N_10231);
and U10448 (N_10448,N_10168,N_10070);
xor U10449 (N_10449,N_10116,N_10230);
xnor U10450 (N_10450,N_10072,N_10056);
xnor U10451 (N_10451,N_10115,N_10144);
xor U10452 (N_10452,N_10131,N_10040);
and U10453 (N_10453,N_10111,N_10016);
nand U10454 (N_10454,N_10245,N_10030);
nor U10455 (N_10455,N_10119,N_10208);
and U10456 (N_10456,N_10072,N_10244);
or U10457 (N_10457,N_10144,N_10069);
xor U10458 (N_10458,N_10235,N_10004);
or U10459 (N_10459,N_10226,N_10010);
nor U10460 (N_10460,N_10230,N_10000);
nor U10461 (N_10461,N_10131,N_10003);
nand U10462 (N_10462,N_10035,N_10209);
nand U10463 (N_10463,N_10211,N_10032);
nor U10464 (N_10464,N_10098,N_10161);
or U10465 (N_10465,N_10100,N_10126);
or U10466 (N_10466,N_10054,N_10221);
or U10467 (N_10467,N_10223,N_10067);
and U10468 (N_10468,N_10146,N_10211);
nand U10469 (N_10469,N_10225,N_10035);
nor U10470 (N_10470,N_10017,N_10052);
nand U10471 (N_10471,N_10087,N_10219);
xnor U10472 (N_10472,N_10222,N_10163);
or U10473 (N_10473,N_10087,N_10053);
xnor U10474 (N_10474,N_10179,N_10190);
nor U10475 (N_10475,N_10197,N_10236);
nand U10476 (N_10476,N_10024,N_10171);
xnor U10477 (N_10477,N_10247,N_10142);
xnor U10478 (N_10478,N_10249,N_10145);
or U10479 (N_10479,N_10211,N_10064);
nand U10480 (N_10480,N_10187,N_10209);
nand U10481 (N_10481,N_10036,N_10113);
nor U10482 (N_10482,N_10216,N_10243);
xor U10483 (N_10483,N_10164,N_10070);
nand U10484 (N_10484,N_10155,N_10217);
xor U10485 (N_10485,N_10095,N_10101);
xnor U10486 (N_10486,N_10071,N_10079);
xor U10487 (N_10487,N_10197,N_10093);
nand U10488 (N_10488,N_10215,N_10240);
xnor U10489 (N_10489,N_10059,N_10221);
or U10490 (N_10490,N_10046,N_10117);
and U10491 (N_10491,N_10185,N_10137);
and U10492 (N_10492,N_10025,N_10127);
or U10493 (N_10493,N_10093,N_10129);
and U10494 (N_10494,N_10208,N_10207);
nand U10495 (N_10495,N_10164,N_10012);
xnor U10496 (N_10496,N_10071,N_10126);
xor U10497 (N_10497,N_10112,N_10224);
or U10498 (N_10498,N_10192,N_10029);
or U10499 (N_10499,N_10227,N_10242);
or U10500 (N_10500,N_10451,N_10375);
xor U10501 (N_10501,N_10377,N_10479);
nor U10502 (N_10502,N_10268,N_10405);
nor U10503 (N_10503,N_10373,N_10411);
or U10504 (N_10504,N_10335,N_10454);
xor U10505 (N_10505,N_10472,N_10303);
and U10506 (N_10506,N_10499,N_10402);
nand U10507 (N_10507,N_10280,N_10469);
nor U10508 (N_10508,N_10354,N_10302);
or U10509 (N_10509,N_10367,N_10274);
nand U10510 (N_10510,N_10407,N_10379);
xnor U10511 (N_10511,N_10344,N_10482);
xor U10512 (N_10512,N_10273,N_10259);
nor U10513 (N_10513,N_10319,N_10459);
and U10514 (N_10514,N_10348,N_10265);
nor U10515 (N_10515,N_10384,N_10279);
xnor U10516 (N_10516,N_10276,N_10342);
nand U10517 (N_10517,N_10463,N_10301);
nor U10518 (N_10518,N_10250,N_10368);
or U10519 (N_10519,N_10448,N_10272);
xor U10520 (N_10520,N_10455,N_10423);
and U10521 (N_10521,N_10307,N_10442);
or U10522 (N_10522,N_10270,N_10325);
nor U10523 (N_10523,N_10324,N_10452);
nor U10524 (N_10524,N_10326,N_10471);
nor U10525 (N_10525,N_10428,N_10410);
nand U10526 (N_10526,N_10358,N_10421);
nand U10527 (N_10527,N_10416,N_10441);
nor U10528 (N_10528,N_10362,N_10450);
nor U10529 (N_10529,N_10356,N_10341);
nor U10530 (N_10530,N_10371,N_10460);
and U10531 (N_10531,N_10339,N_10308);
nand U10532 (N_10532,N_10281,N_10269);
and U10533 (N_10533,N_10489,N_10266);
xor U10534 (N_10534,N_10298,N_10425);
nand U10535 (N_10535,N_10386,N_10412);
or U10536 (N_10536,N_10256,N_10284);
and U10537 (N_10537,N_10456,N_10444);
xnor U10538 (N_10538,N_10312,N_10398);
and U10539 (N_10539,N_10262,N_10491);
xor U10540 (N_10540,N_10419,N_10283);
nor U10541 (N_10541,N_10253,N_10395);
xnor U10542 (N_10542,N_10457,N_10490);
xnor U10543 (N_10543,N_10409,N_10327);
nand U10544 (N_10544,N_10349,N_10493);
nor U10545 (N_10545,N_10294,N_10372);
or U10546 (N_10546,N_10436,N_10288);
nand U10547 (N_10547,N_10278,N_10285);
nor U10548 (N_10548,N_10484,N_10264);
nand U10549 (N_10549,N_10275,N_10439);
nor U10550 (N_10550,N_10314,N_10487);
nand U10551 (N_10551,N_10435,N_10306);
and U10552 (N_10552,N_10400,N_10477);
nand U10553 (N_10553,N_10364,N_10385);
or U10554 (N_10554,N_10432,N_10346);
nand U10555 (N_10555,N_10474,N_10426);
nand U10556 (N_10556,N_10404,N_10378);
or U10557 (N_10557,N_10347,N_10486);
or U10558 (N_10558,N_10461,N_10291);
nor U10559 (N_10559,N_10252,N_10406);
or U10560 (N_10560,N_10429,N_10470);
or U10561 (N_10561,N_10260,N_10458);
and U10562 (N_10562,N_10392,N_10462);
or U10563 (N_10563,N_10351,N_10271);
or U10564 (N_10564,N_10257,N_10258);
nor U10565 (N_10565,N_10391,N_10465);
nand U10566 (N_10566,N_10464,N_10343);
xnor U10567 (N_10567,N_10267,N_10316);
nand U10568 (N_10568,N_10445,N_10337);
and U10569 (N_10569,N_10295,N_10481);
or U10570 (N_10570,N_10360,N_10417);
and U10571 (N_10571,N_10315,N_10413);
xnor U10572 (N_10572,N_10488,N_10447);
nand U10573 (N_10573,N_10390,N_10374);
xnor U10574 (N_10574,N_10443,N_10311);
nor U10575 (N_10575,N_10383,N_10415);
and U10576 (N_10576,N_10387,N_10330);
xor U10577 (N_10577,N_10446,N_10338);
nand U10578 (N_10578,N_10332,N_10287);
xnor U10579 (N_10579,N_10366,N_10399);
nor U10580 (N_10580,N_10345,N_10309);
xnor U10581 (N_10581,N_10261,N_10478);
nor U10582 (N_10582,N_10318,N_10313);
nor U10583 (N_10583,N_10480,N_10468);
nand U10584 (N_10584,N_10473,N_10427);
nand U10585 (N_10585,N_10255,N_10297);
xor U10586 (N_10586,N_10369,N_10299);
xor U10587 (N_10587,N_10476,N_10485);
xnor U10588 (N_10588,N_10393,N_10431);
nand U10589 (N_10589,N_10289,N_10420);
or U10590 (N_10590,N_10370,N_10494);
nand U10591 (N_10591,N_10353,N_10251);
or U10592 (N_10592,N_10430,N_10437);
nor U10593 (N_10593,N_10336,N_10483);
nand U10594 (N_10594,N_10440,N_10350);
nor U10595 (N_10595,N_10422,N_10263);
and U10596 (N_10596,N_10290,N_10414);
and U10597 (N_10597,N_10389,N_10492);
xnor U10598 (N_10598,N_10333,N_10453);
nor U10599 (N_10599,N_10334,N_10282);
xor U10600 (N_10600,N_10498,N_10331);
nor U10601 (N_10601,N_10495,N_10467);
and U10602 (N_10602,N_10449,N_10359);
or U10603 (N_10603,N_10363,N_10380);
nor U10604 (N_10604,N_10296,N_10376);
or U10605 (N_10605,N_10394,N_10497);
and U10606 (N_10606,N_10310,N_10475);
nand U10607 (N_10607,N_10286,N_10434);
nand U10608 (N_10608,N_10305,N_10300);
nor U10609 (N_10609,N_10340,N_10397);
and U10610 (N_10610,N_10317,N_10424);
or U10611 (N_10611,N_10293,N_10381);
or U10612 (N_10612,N_10355,N_10328);
nand U10613 (N_10613,N_10357,N_10396);
nand U10614 (N_10614,N_10254,N_10321);
xor U10615 (N_10615,N_10403,N_10433);
nand U10616 (N_10616,N_10408,N_10304);
or U10617 (N_10617,N_10361,N_10388);
nand U10618 (N_10618,N_10292,N_10401);
and U10619 (N_10619,N_10365,N_10277);
or U10620 (N_10620,N_10352,N_10329);
nand U10621 (N_10621,N_10466,N_10418);
nor U10622 (N_10622,N_10438,N_10496);
xor U10623 (N_10623,N_10323,N_10320);
xor U10624 (N_10624,N_10322,N_10382);
xor U10625 (N_10625,N_10402,N_10362);
and U10626 (N_10626,N_10423,N_10280);
xnor U10627 (N_10627,N_10297,N_10374);
and U10628 (N_10628,N_10453,N_10416);
nand U10629 (N_10629,N_10319,N_10469);
xor U10630 (N_10630,N_10336,N_10467);
or U10631 (N_10631,N_10467,N_10494);
xor U10632 (N_10632,N_10452,N_10456);
nand U10633 (N_10633,N_10337,N_10457);
or U10634 (N_10634,N_10279,N_10428);
or U10635 (N_10635,N_10277,N_10315);
nand U10636 (N_10636,N_10360,N_10477);
nand U10637 (N_10637,N_10361,N_10336);
or U10638 (N_10638,N_10486,N_10456);
xnor U10639 (N_10639,N_10277,N_10377);
nand U10640 (N_10640,N_10308,N_10306);
nor U10641 (N_10641,N_10422,N_10437);
or U10642 (N_10642,N_10435,N_10453);
nand U10643 (N_10643,N_10331,N_10304);
nor U10644 (N_10644,N_10431,N_10483);
nor U10645 (N_10645,N_10320,N_10365);
nor U10646 (N_10646,N_10349,N_10277);
and U10647 (N_10647,N_10293,N_10441);
or U10648 (N_10648,N_10280,N_10397);
nor U10649 (N_10649,N_10442,N_10488);
or U10650 (N_10650,N_10303,N_10413);
and U10651 (N_10651,N_10277,N_10412);
or U10652 (N_10652,N_10462,N_10474);
xnor U10653 (N_10653,N_10480,N_10384);
xnor U10654 (N_10654,N_10337,N_10493);
or U10655 (N_10655,N_10346,N_10423);
or U10656 (N_10656,N_10497,N_10285);
xnor U10657 (N_10657,N_10286,N_10420);
nand U10658 (N_10658,N_10318,N_10330);
nor U10659 (N_10659,N_10371,N_10450);
nand U10660 (N_10660,N_10403,N_10349);
nor U10661 (N_10661,N_10384,N_10449);
nor U10662 (N_10662,N_10389,N_10274);
and U10663 (N_10663,N_10417,N_10453);
nand U10664 (N_10664,N_10319,N_10456);
or U10665 (N_10665,N_10416,N_10263);
nand U10666 (N_10666,N_10319,N_10301);
xnor U10667 (N_10667,N_10436,N_10396);
nor U10668 (N_10668,N_10493,N_10298);
nand U10669 (N_10669,N_10406,N_10432);
xor U10670 (N_10670,N_10451,N_10258);
nor U10671 (N_10671,N_10305,N_10406);
nor U10672 (N_10672,N_10268,N_10406);
nor U10673 (N_10673,N_10437,N_10433);
or U10674 (N_10674,N_10259,N_10399);
and U10675 (N_10675,N_10496,N_10331);
or U10676 (N_10676,N_10289,N_10293);
nor U10677 (N_10677,N_10344,N_10481);
xor U10678 (N_10678,N_10397,N_10461);
nand U10679 (N_10679,N_10409,N_10256);
nor U10680 (N_10680,N_10445,N_10370);
xor U10681 (N_10681,N_10472,N_10435);
nor U10682 (N_10682,N_10267,N_10471);
nor U10683 (N_10683,N_10294,N_10293);
xnor U10684 (N_10684,N_10477,N_10356);
nand U10685 (N_10685,N_10378,N_10442);
and U10686 (N_10686,N_10397,N_10302);
or U10687 (N_10687,N_10439,N_10414);
nand U10688 (N_10688,N_10254,N_10275);
and U10689 (N_10689,N_10477,N_10307);
or U10690 (N_10690,N_10412,N_10314);
nor U10691 (N_10691,N_10344,N_10318);
xnor U10692 (N_10692,N_10488,N_10324);
or U10693 (N_10693,N_10389,N_10348);
nand U10694 (N_10694,N_10446,N_10453);
or U10695 (N_10695,N_10269,N_10440);
and U10696 (N_10696,N_10417,N_10299);
and U10697 (N_10697,N_10482,N_10288);
or U10698 (N_10698,N_10429,N_10445);
nand U10699 (N_10699,N_10287,N_10410);
or U10700 (N_10700,N_10409,N_10368);
xor U10701 (N_10701,N_10422,N_10285);
or U10702 (N_10702,N_10315,N_10274);
nor U10703 (N_10703,N_10474,N_10422);
and U10704 (N_10704,N_10373,N_10455);
and U10705 (N_10705,N_10348,N_10309);
xor U10706 (N_10706,N_10293,N_10262);
xnor U10707 (N_10707,N_10474,N_10352);
xnor U10708 (N_10708,N_10422,N_10253);
and U10709 (N_10709,N_10345,N_10394);
and U10710 (N_10710,N_10402,N_10406);
nor U10711 (N_10711,N_10327,N_10347);
and U10712 (N_10712,N_10258,N_10456);
or U10713 (N_10713,N_10363,N_10448);
nor U10714 (N_10714,N_10470,N_10419);
nand U10715 (N_10715,N_10452,N_10397);
nor U10716 (N_10716,N_10293,N_10323);
nor U10717 (N_10717,N_10438,N_10260);
or U10718 (N_10718,N_10266,N_10311);
or U10719 (N_10719,N_10258,N_10263);
or U10720 (N_10720,N_10450,N_10490);
and U10721 (N_10721,N_10465,N_10432);
and U10722 (N_10722,N_10389,N_10345);
and U10723 (N_10723,N_10306,N_10457);
nand U10724 (N_10724,N_10289,N_10380);
nor U10725 (N_10725,N_10333,N_10365);
xor U10726 (N_10726,N_10369,N_10353);
and U10727 (N_10727,N_10274,N_10455);
or U10728 (N_10728,N_10356,N_10363);
and U10729 (N_10729,N_10485,N_10449);
and U10730 (N_10730,N_10293,N_10400);
or U10731 (N_10731,N_10359,N_10343);
nor U10732 (N_10732,N_10355,N_10378);
nand U10733 (N_10733,N_10277,N_10306);
xnor U10734 (N_10734,N_10393,N_10325);
nor U10735 (N_10735,N_10347,N_10462);
xor U10736 (N_10736,N_10435,N_10321);
nand U10737 (N_10737,N_10404,N_10455);
xor U10738 (N_10738,N_10252,N_10318);
or U10739 (N_10739,N_10340,N_10331);
nand U10740 (N_10740,N_10467,N_10323);
xnor U10741 (N_10741,N_10395,N_10361);
nand U10742 (N_10742,N_10411,N_10334);
nor U10743 (N_10743,N_10329,N_10395);
nand U10744 (N_10744,N_10427,N_10448);
nor U10745 (N_10745,N_10328,N_10261);
and U10746 (N_10746,N_10343,N_10250);
and U10747 (N_10747,N_10293,N_10461);
xnor U10748 (N_10748,N_10284,N_10352);
xor U10749 (N_10749,N_10460,N_10490);
and U10750 (N_10750,N_10573,N_10726);
and U10751 (N_10751,N_10574,N_10519);
xnor U10752 (N_10752,N_10630,N_10559);
or U10753 (N_10753,N_10557,N_10718);
or U10754 (N_10754,N_10662,N_10571);
xor U10755 (N_10755,N_10595,N_10584);
nand U10756 (N_10756,N_10683,N_10547);
nand U10757 (N_10757,N_10748,N_10535);
nand U10758 (N_10758,N_10621,N_10694);
or U10759 (N_10759,N_10672,N_10505);
xor U10760 (N_10760,N_10551,N_10667);
nor U10761 (N_10761,N_10615,N_10616);
or U10762 (N_10762,N_10634,N_10742);
nand U10763 (N_10763,N_10706,N_10578);
or U10764 (N_10764,N_10632,N_10503);
nor U10765 (N_10765,N_10721,N_10597);
xnor U10766 (N_10766,N_10717,N_10545);
and U10767 (N_10767,N_10715,N_10564);
nor U10768 (N_10768,N_10534,N_10620);
nor U10769 (N_10769,N_10655,N_10511);
and U10770 (N_10770,N_10522,N_10506);
or U10771 (N_10771,N_10515,N_10661);
xor U10772 (N_10772,N_10541,N_10539);
and U10773 (N_10773,N_10657,N_10603);
or U10774 (N_10774,N_10733,N_10724);
xnor U10775 (N_10775,N_10658,N_10692);
xor U10776 (N_10776,N_10599,N_10647);
and U10777 (N_10777,N_10636,N_10668);
or U10778 (N_10778,N_10702,N_10690);
or U10779 (N_10779,N_10542,N_10622);
and U10780 (N_10780,N_10691,N_10625);
xnor U10781 (N_10781,N_10654,N_10745);
or U10782 (N_10782,N_10725,N_10653);
and U10783 (N_10783,N_10652,N_10612);
nor U10784 (N_10784,N_10558,N_10619);
nand U10785 (N_10785,N_10642,N_10592);
or U10786 (N_10786,N_10714,N_10637);
xor U10787 (N_10787,N_10671,N_10749);
xnor U10788 (N_10788,N_10656,N_10582);
xnor U10789 (N_10789,N_10727,N_10530);
and U10790 (N_10790,N_10593,N_10518);
nand U10791 (N_10791,N_10602,N_10645);
nand U10792 (N_10792,N_10739,N_10605);
or U10793 (N_10793,N_10737,N_10532);
nor U10794 (N_10794,N_10586,N_10549);
xnor U10795 (N_10795,N_10588,N_10626);
xor U10796 (N_10796,N_10562,N_10705);
and U10797 (N_10797,N_10719,N_10546);
nor U10798 (N_10798,N_10536,N_10666);
xor U10799 (N_10799,N_10650,N_10569);
nor U10800 (N_10800,N_10713,N_10531);
nand U10801 (N_10801,N_10644,N_10677);
and U10802 (N_10802,N_10663,N_10529);
nand U10803 (N_10803,N_10501,N_10675);
xnor U10804 (N_10804,N_10591,N_10512);
xor U10805 (N_10805,N_10608,N_10516);
or U10806 (N_10806,N_10553,N_10500);
and U10807 (N_10807,N_10638,N_10684);
nand U10808 (N_10808,N_10579,N_10596);
nor U10809 (N_10809,N_10716,N_10627);
or U10810 (N_10810,N_10740,N_10681);
and U10811 (N_10811,N_10635,N_10695);
nand U10812 (N_10812,N_10561,N_10728);
or U10813 (N_10813,N_10746,N_10665);
and U10814 (N_10814,N_10700,N_10701);
or U10815 (N_10815,N_10686,N_10523);
nor U10816 (N_10816,N_10707,N_10651);
and U10817 (N_10817,N_10673,N_10628);
and U10818 (N_10818,N_10556,N_10618);
nand U10819 (N_10819,N_10720,N_10570);
or U10820 (N_10820,N_10659,N_10576);
and U10821 (N_10821,N_10696,N_10687);
and U10822 (N_10822,N_10572,N_10709);
xnor U10823 (N_10823,N_10682,N_10697);
xnor U10824 (N_10824,N_10712,N_10688);
or U10825 (N_10825,N_10544,N_10533);
xor U10826 (N_10826,N_10566,N_10670);
and U10827 (N_10827,N_10587,N_10722);
and U10828 (N_10828,N_10540,N_10736);
xnor U10829 (N_10829,N_10674,N_10604);
or U10830 (N_10830,N_10509,N_10743);
nor U10831 (N_10831,N_10563,N_10669);
xnor U10832 (N_10832,N_10548,N_10575);
xor U10833 (N_10833,N_10565,N_10710);
or U10834 (N_10834,N_10679,N_10731);
nand U10835 (N_10835,N_10648,N_10611);
nor U10836 (N_10836,N_10585,N_10598);
nor U10837 (N_10837,N_10521,N_10730);
nor U10838 (N_10838,N_10744,N_10610);
and U10839 (N_10839,N_10525,N_10560);
xnor U10840 (N_10840,N_10685,N_10550);
nand U10841 (N_10841,N_10704,N_10617);
xnor U10842 (N_10842,N_10678,N_10711);
nor U10843 (N_10843,N_10643,N_10580);
and U10844 (N_10844,N_10732,N_10528);
and U10845 (N_10845,N_10640,N_10581);
or U10846 (N_10846,N_10641,N_10689);
and U10847 (N_10847,N_10624,N_10589);
and U10848 (N_10848,N_10676,N_10504);
and U10849 (N_10849,N_10698,N_10514);
xnor U10850 (N_10850,N_10583,N_10601);
nor U10851 (N_10851,N_10507,N_10554);
nor U10852 (N_10852,N_10664,N_10524);
and U10853 (N_10853,N_10629,N_10510);
nand U10854 (N_10854,N_10508,N_10609);
xor U10855 (N_10855,N_10741,N_10623);
and U10856 (N_10856,N_10708,N_10607);
xor U10857 (N_10857,N_10649,N_10680);
or U10858 (N_10858,N_10552,N_10555);
nand U10859 (N_10859,N_10568,N_10590);
nand U10860 (N_10860,N_10633,N_10537);
xor U10861 (N_10861,N_10660,N_10520);
or U10862 (N_10862,N_10594,N_10738);
nor U10863 (N_10863,N_10543,N_10639);
and U10864 (N_10864,N_10747,N_10729);
and U10865 (N_10865,N_10735,N_10577);
or U10866 (N_10866,N_10693,N_10606);
xnor U10867 (N_10867,N_10502,N_10723);
or U10868 (N_10868,N_10513,N_10646);
xor U10869 (N_10869,N_10631,N_10734);
and U10870 (N_10870,N_10538,N_10614);
and U10871 (N_10871,N_10703,N_10699);
xnor U10872 (N_10872,N_10527,N_10600);
or U10873 (N_10873,N_10613,N_10567);
or U10874 (N_10874,N_10517,N_10526);
or U10875 (N_10875,N_10528,N_10551);
nor U10876 (N_10876,N_10665,N_10642);
nand U10877 (N_10877,N_10720,N_10564);
nand U10878 (N_10878,N_10749,N_10701);
and U10879 (N_10879,N_10566,N_10664);
and U10880 (N_10880,N_10557,N_10611);
and U10881 (N_10881,N_10684,N_10729);
or U10882 (N_10882,N_10698,N_10602);
xnor U10883 (N_10883,N_10544,N_10604);
nor U10884 (N_10884,N_10545,N_10724);
nor U10885 (N_10885,N_10646,N_10625);
and U10886 (N_10886,N_10664,N_10647);
or U10887 (N_10887,N_10591,N_10720);
or U10888 (N_10888,N_10660,N_10528);
or U10889 (N_10889,N_10712,N_10594);
nor U10890 (N_10890,N_10660,N_10561);
nand U10891 (N_10891,N_10545,N_10728);
nand U10892 (N_10892,N_10670,N_10691);
nand U10893 (N_10893,N_10513,N_10704);
nand U10894 (N_10894,N_10598,N_10550);
nand U10895 (N_10895,N_10681,N_10626);
xor U10896 (N_10896,N_10508,N_10600);
nor U10897 (N_10897,N_10600,N_10574);
nor U10898 (N_10898,N_10614,N_10728);
nor U10899 (N_10899,N_10524,N_10523);
nand U10900 (N_10900,N_10538,N_10600);
and U10901 (N_10901,N_10565,N_10547);
xor U10902 (N_10902,N_10598,N_10577);
xnor U10903 (N_10903,N_10555,N_10564);
xnor U10904 (N_10904,N_10675,N_10523);
xnor U10905 (N_10905,N_10541,N_10722);
or U10906 (N_10906,N_10700,N_10634);
and U10907 (N_10907,N_10621,N_10605);
xor U10908 (N_10908,N_10542,N_10589);
nand U10909 (N_10909,N_10565,N_10665);
nand U10910 (N_10910,N_10618,N_10562);
nand U10911 (N_10911,N_10596,N_10685);
or U10912 (N_10912,N_10673,N_10597);
nor U10913 (N_10913,N_10610,N_10532);
or U10914 (N_10914,N_10540,N_10713);
and U10915 (N_10915,N_10570,N_10545);
and U10916 (N_10916,N_10664,N_10571);
nand U10917 (N_10917,N_10683,N_10681);
or U10918 (N_10918,N_10668,N_10565);
nand U10919 (N_10919,N_10572,N_10616);
and U10920 (N_10920,N_10540,N_10718);
xnor U10921 (N_10921,N_10506,N_10703);
or U10922 (N_10922,N_10739,N_10737);
and U10923 (N_10923,N_10578,N_10542);
or U10924 (N_10924,N_10609,N_10504);
and U10925 (N_10925,N_10676,N_10641);
xnor U10926 (N_10926,N_10601,N_10691);
nor U10927 (N_10927,N_10716,N_10576);
and U10928 (N_10928,N_10568,N_10579);
nand U10929 (N_10929,N_10604,N_10726);
xor U10930 (N_10930,N_10533,N_10574);
nand U10931 (N_10931,N_10526,N_10658);
xnor U10932 (N_10932,N_10511,N_10652);
xor U10933 (N_10933,N_10622,N_10646);
nand U10934 (N_10934,N_10610,N_10596);
or U10935 (N_10935,N_10681,N_10667);
or U10936 (N_10936,N_10654,N_10671);
nor U10937 (N_10937,N_10736,N_10589);
xor U10938 (N_10938,N_10706,N_10679);
nor U10939 (N_10939,N_10660,N_10665);
and U10940 (N_10940,N_10666,N_10574);
and U10941 (N_10941,N_10540,N_10560);
xor U10942 (N_10942,N_10682,N_10718);
nor U10943 (N_10943,N_10628,N_10535);
or U10944 (N_10944,N_10604,N_10517);
xor U10945 (N_10945,N_10574,N_10749);
or U10946 (N_10946,N_10549,N_10657);
xor U10947 (N_10947,N_10597,N_10682);
xnor U10948 (N_10948,N_10530,N_10636);
nor U10949 (N_10949,N_10728,N_10619);
and U10950 (N_10950,N_10677,N_10735);
nand U10951 (N_10951,N_10721,N_10677);
xor U10952 (N_10952,N_10638,N_10703);
and U10953 (N_10953,N_10594,N_10581);
nor U10954 (N_10954,N_10743,N_10615);
nand U10955 (N_10955,N_10526,N_10701);
nor U10956 (N_10956,N_10607,N_10536);
xor U10957 (N_10957,N_10581,N_10559);
or U10958 (N_10958,N_10747,N_10716);
nand U10959 (N_10959,N_10699,N_10505);
or U10960 (N_10960,N_10672,N_10700);
xor U10961 (N_10961,N_10516,N_10639);
nand U10962 (N_10962,N_10646,N_10577);
xor U10963 (N_10963,N_10676,N_10534);
nand U10964 (N_10964,N_10609,N_10601);
or U10965 (N_10965,N_10544,N_10521);
or U10966 (N_10966,N_10745,N_10691);
and U10967 (N_10967,N_10624,N_10675);
xor U10968 (N_10968,N_10575,N_10738);
xor U10969 (N_10969,N_10564,N_10695);
nor U10970 (N_10970,N_10722,N_10617);
nand U10971 (N_10971,N_10728,N_10684);
xnor U10972 (N_10972,N_10501,N_10689);
xor U10973 (N_10973,N_10551,N_10711);
xnor U10974 (N_10974,N_10568,N_10550);
xor U10975 (N_10975,N_10519,N_10715);
xor U10976 (N_10976,N_10741,N_10603);
or U10977 (N_10977,N_10569,N_10548);
or U10978 (N_10978,N_10647,N_10644);
nand U10979 (N_10979,N_10697,N_10641);
and U10980 (N_10980,N_10709,N_10720);
or U10981 (N_10981,N_10617,N_10711);
nor U10982 (N_10982,N_10692,N_10728);
nand U10983 (N_10983,N_10665,N_10695);
nor U10984 (N_10984,N_10736,N_10516);
xor U10985 (N_10985,N_10625,N_10708);
or U10986 (N_10986,N_10545,N_10689);
nor U10987 (N_10987,N_10596,N_10605);
or U10988 (N_10988,N_10517,N_10567);
and U10989 (N_10989,N_10521,N_10714);
nor U10990 (N_10990,N_10672,N_10613);
and U10991 (N_10991,N_10588,N_10691);
or U10992 (N_10992,N_10511,N_10589);
or U10993 (N_10993,N_10687,N_10727);
and U10994 (N_10994,N_10501,N_10648);
or U10995 (N_10995,N_10601,N_10737);
or U10996 (N_10996,N_10745,N_10520);
and U10997 (N_10997,N_10683,N_10625);
and U10998 (N_10998,N_10641,N_10660);
and U10999 (N_10999,N_10639,N_10576);
or U11000 (N_11000,N_10992,N_10790);
xor U11001 (N_11001,N_10989,N_10924);
or U11002 (N_11002,N_10791,N_10877);
and U11003 (N_11003,N_10847,N_10946);
xnor U11004 (N_11004,N_10975,N_10968);
nor U11005 (N_11005,N_10866,N_10917);
and U11006 (N_11006,N_10762,N_10773);
xor U11007 (N_11007,N_10965,N_10853);
and U11008 (N_11008,N_10950,N_10964);
xnor U11009 (N_11009,N_10770,N_10991);
nor U11010 (N_11010,N_10801,N_10810);
nand U11011 (N_11011,N_10829,N_10761);
xor U11012 (N_11012,N_10880,N_10831);
nor U11013 (N_11013,N_10833,N_10851);
or U11014 (N_11014,N_10916,N_10875);
and U11015 (N_11015,N_10813,N_10784);
nand U11016 (N_11016,N_10912,N_10905);
xnor U11017 (N_11017,N_10815,N_10857);
nor U11018 (N_11018,N_10915,N_10780);
xor U11019 (N_11019,N_10963,N_10892);
and U11020 (N_11020,N_10842,N_10838);
xor U11021 (N_11021,N_10942,N_10819);
or U11022 (N_11022,N_10993,N_10805);
nor U11023 (N_11023,N_10800,N_10835);
xnor U11024 (N_11024,N_10961,N_10795);
nor U11025 (N_11025,N_10903,N_10985);
nand U11026 (N_11026,N_10919,N_10854);
nand U11027 (N_11027,N_10870,N_10824);
nand U11028 (N_11028,N_10941,N_10890);
nand U11029 (N_11029,N_10914,N_10765);
xor U11030 (N_11030,N_10803,N_10883);
and U11031 (N_11031,N_10966,N_10797);
and U11032 (N_11032,N_10984,N_10774);
or U11033 (N_11033,N_10972,N_10856);
nor U11034 (N_11034,N_10879,N_10977);
nor U11035 (N_11035,N_10830,N_10889);
and U11036 (N_11036,N_10812,N_10758);
or U11037 (N_11037,N_10982,N_10816);
nand U11038 (N_11038,N_10909,N_10954);
xnor U11039 (N_11039,N_10911,N_10873);
nand U11040 (N_11040,N_10988,N_10973);
xor U11041 (N_11041,N_10969,N_10848);
xor U11042 (N_11042,N_10974,N_10841);
nor U11043 (N_11043,N_10760,N_10771);
and U11044 (N_11044,N_10979,N_10840);
and U11045 (N_11045,N_10769,N_10821);
nor U11046 (N_11046,N_10750,N_10827);
and U11047 (N_11047,N_10957,N_10926);
nor U11048 (N_11048,N_10996,N_10887);
and U11049 (N_11049,N_10976,N_10978);
or U11050 (N_11050,N_10757,N_10898);
nand U11051 (N_11051,N_10987,N_10896);
or U11052 (N_11052,N_10967,N_10958);
nor U11053 (N_11053,N_10846,N_10931);
and U11054 (N_11054,N_10820,N_10882);
nor U11055 (N_11055,N_10995,N_10871);
and U11056 (N_11056,N_10955,N_10849);
nand U11057 (N_11057,N_10834,N_10939);
xnor U11058 (N_11058,N_10895,N_10763);
xnor U11059 (N_11059,N_10861,N_10855);
nand U11060 (N_11060,N_10913,N_10802);
xnor U11061 (N_11061,N_10822,N_10766);
nand U11062 (N_11062,N_10845,N_10990);
nor U11063 (N_11063,N_10865,N_10920);
xor U11064 (N_11064,N_10867,N_10893);
and U11065 (N_11065,N_10899,N_10828);
nor U11066 (N_11066,N_10789,N_10778);
xnor U11067 (N_11067,N_10852,N_10863);
and U11068 (N_11068,N_10804,N_10793);
nor U11069 (N_11069,N_10811,N_10951);
nor U11070 (N_11070,N_10809,N_10994);
nand U11071 (N_11071,N_10962,N_10904);
nor U11072 (N_11072,N_10799,N_10874);
and U11073 (N_11073,N_10936,N_10885);
nand U11074 (N_11074,N_10859,N_10807);
nand U11075 (N_11075,N_10923,N_10754);
nand U11076 (N_11076,N_10823,N_10782);
nand U11077 (N_11077,N_10953,N_10886);
or U11078 (N_11078,N_10792,N_10935);
xor U11079 (N_11079,N_10970,N_10876);
and U11080 (N_11080,N_10925,N_10943);
or U11081 (N_11081,N_10844,N_10868);
and U11082 (N_11082,N_10928,N_10759);
and U11083 (N_11083,N_10858,N_10999);
and U11084 (N_11084,N_10772,N_10971);
nand U11085 (N_11085,N_10836,N_10767);
nor U11086 (N_11086,N_10775,N_10983);
nor U11087 (N_11087,N_10753,N_10927);
nand U11088 (N_11088,N_10755,N_10832);
or U11089 (N_11089,N_10952,N_10947);
nor U11090 (N_11090,N_10897,N_10768);
nor U11091 (N_11091,N_10907,N_10906);
and U11092 (N_11092,N_10940,N_10843);
nor U11093 (N_11093,N_10945,N_10788);
nor U11094 (N_11094,N_10937,N_10756);
and U11095 (N_11095,N_10959,N_10888);
xor U11096 (N_11096,N_10938,N_10948);
xnor U11097 (N_11097,N_10817,N_10839);
nor U11098 (N_11098,N_10777,N_10826);
nand U11099 (N_11099,N_10918,N_10956);
xnor U11100 (N_11100,N_10864,N_10900);
or U11101 (N_11101,N_10910,N_10881);
xnor U11102 (N_11102,N_10860,N_10781);
or U11103 (N_11103,N_10798,N_10901);
and U11104 (N_11104,N_10776,N_10808);
and U11105 (N_11105,N_10997,N_10869);
and U11106 (N_11106,N_10894,N_10785);
nor U11107 (N_11107,N_10752,N_10986);
nor U11108 (N_11108,N_10908,N_10786);
or U11109 (N_11109,N_10932,N_10751);
nand U11110 (N_11110,N_10764,N_10825);
and U11111 (N_11111,N_10960,N_10998);
and U11112 (N_11112,N_10934,N_10806);
or U11113 (N_11113,N_10814,N_10922);
nand U11114 (N_11114,N_10884,N_10862);
and U11115 (N_11115,N_10944,N_10818);
and U11116 (N_11116,N_10850,N_10929);
and U11117 (N_11117,N_10878,N_10933);
and U11118 (N_11118,N_10796,N_10837);
or U11119 (N_11119,N_10981,N_10902);
nor U11120 (N_11120,N_10872,N_10949);
xnor U11121 (N_11121,N_10930,N_10891);
and U11122 (N_11122,N_10787,N_10783);
xor U11123 (N_11123,N_10921,N_10794);
nand U11124 (N_11124,N_10980,N_10779);
nand U11125 (N_11125,N_10877,N_10943);
and U11126 (N_11126,N_10824,N_10809);
nand U11127 (N_11127,N_10954,N_10800);
and U11128 (N_11128,N_10991,N_10825);
and U11129 (N_11129,N_10834,N_10931);
and U11130 (N_11130,N_10774,N_10786);
xnor U11131 (N_11131,N_10928,N_10965);
nor U11132 (N_11132,N_10957,N_10820);
and U11133 (N_11133,N_10934,N_10901);
or U11134 (N_11134,N_10925,N_10854);
nand U11135 (N_11135,N_10882,N_10781);
xnor U11136 (N_11136,N_10838,N_10876);
or U11137 (N_11137,N_10931,N_10761);
and U11138 (N_11138,N_10945,N_10931);
or U11139 (N_11139,N_10808,N_10789);
and U11140 (N_11140,N_10950,N_10840);
xor U11141 (N_11141,N_10925,N_10771);
nor U11142 (N_11142,N_10833,N_10933);
or U11143 (N_11143,N_10828,N_10923);
and U11144 (N_11144,N_10874,N_10980);
xor U11145 (N_11145,N_10813,N_10882);
or U11146 (N_11146,N_10771,N_10947);
xnor U11147 (N_11147,N_10802,N_10809);
nor U11148 (N_11148,N_10862,N_10903);
or U11149 (N_11149,N_10937,N_10994);
xnor U11150 (N_11150,N_10857,N_10914);
nand U11151 (N_11151,N_10792,N_10787);
nor U11152 (N_11152,N_10952,N_10804);
xor U11153 (N_11153,N_10804,N_10774);
xor U11154 (N_11154,N_10862,N_10944);
nand U11155 (N_11155,N_10867,N_10817);
nand U11156 (N_11156,N_10874,N_10806);
xor U11157 (N_11157,N_10853,N_10953);
nand U11158 (N_11158,N_10797,N_10919);
and U11159 (N_11159,N_10917,N_10957);
or U11160 (N_11160,N_10978,N_10968);
or U11161 (N_11161,N_10812,N_10829);
nand U11162 (N_11162,N_10870,N_10774);
and U11163 (N_11163,N_10787,N_10973);
and U11164 (N_11164,N_10895,N_10881);
or U11165 (N_11165,N_10977,N_10968);
nand U11166 (N_11166,N_10933,N_10967);
xor U11167 (N_11167,N_10756,N_10797);
xnor U11168 (N_11168,N_10771,N_10990);
nor U11169 (N_11169,N_10933,N_10759);
xor U11170 (N_11170,N_10946,N_10930);
nand U11171 (N_11171,N_10776,N_10990);
nand U11172 (N_11172,N_10901,N_10872);
or U11173 (N_11173,N_10932,N_10837);
nand U11174 (N_11174,N_10910,N_10790);
or U11175 (N_11175,N_10846,N_10872);
nand U11176 (N_11176,N_10787,N_10938);
nor U11177 (N_11177,N_10825,N_10781);
and U11178 (N_11178,N_10770,N_10994);
nand U11179 (N_11179,N_10997,N_10891);
nand U11180 (N_11180,N_10905,N_10931);
nor U11181 (N_11181,N_10898,N_10857);
or U11182 (N_11182,N_10901,N_10850);
or U11183 (N_11183,N_10892,N_10843);
and U11184 (N_11184,N_10811,N_10756);
nor U11185 (N_11185,N_10949,N_10859);
nor U11186 (N_11186,N_10847,N_10931);
or U11187 (N_11187,N_10841,N_10925);
and U11188 (N_11188,N_10851,N_10829);
or U11189 (N_11189,N_10770,N_10929);
or U11190 (N_11190,N_10918,N_10941);
xor U11191 (N_11191,N_10972,N_10761);
xnor U11192 (N_11192,N_10833,N_10912);
nand U11193 (N_11193,N_10900,N_10835);
and U11194 (N_11194,N_10756,N_10940);
nor U11195 (N_11195,N_10952,N_10833);
or U11196 (N_11196,N_10887,N_10808);
or U11197 (N_11197,N_10767,N_10948);
and U11198 (N_11198,N_10873,N_10972);
or U11199 (N_11199,N_10831,N_10790);
or U11200 (N_11200,N_10982,N_10766);
xnor U11201 (N_11201,N_10786,N_10776);
nand U11202 (N_11202,N_10753,N_10830);
or U11203 (N_11203,N_10829,N_10918);
xor U11204 (N_11204,N_10950,N_10944);
and U11205 (N_11205,N_10958,N_10915);
or U11206 (N_11206,N_10991,N_10767);
or U11207 (N_11207,N_10756,N_10959);
nor U11208 (N_11208,N_10848,N_10831);
xor U11209 (N_11209,N_10982,N_10964);
or U11210 (N_11210,N_10818,N_10974);
nor U11211 (N_11211,N_10819,N_10947);
xnor U11212 (N_11212,N_10924,N_10905);
nand U11213 (N_11213,N_10848,N_10923);
and U11214 (N_11214,N_10984,N_10772);
or U11215 (N_11215,N_10807,N_10806);
nand U11216 (N_11216,N_10814,N_10908);
nand U11217 (N_11217,N_10983,N_10944);
xnor U11218 (N_11218,N_10940,N_10798);
xor U11219 (N_11219,N_10816,N_10862);
nor U11220 (N_11220,N_10812,N_10760);
xnor U11221 (N_11221,N_10938,N_10817);
and U11222 (N_11222,N_10840,N_10774);
or U11223 (N_11223,N_10928,N_10921);
and U11224 (N_11224,N_10790,N_10846);
xor U11225 (N_11225,N_10901,N_10810);
or U11226 (N_11226,N_10930,N_10820);
nand U11227 (N_11227,N_10776,N_10985);
nor U11228 (N_11228,N_10787,N_10891);
and U11229 (N_11229,N_10891,N_10803);
xnor U11230 (N_11230,N_10982,N_10776);
or U11231 (N_11231,N_10861,N_10752);
or U11232 (N_11232,N_10984,N_10891);
xor U11233 (N_11233,N_10949,N_10908);
and U11234 (N_11234,N_10874,N_10791);
xor U11235 (N_11235,N_10891,N_10969);
or U11236 (N_11236,N_10824,N_10813);
nor U11237 (N_11237,N_10895,N_10918);
nand U11238 (N_11238,N_10833,N_10895);
or U11239 (N_11239,N_10846,N_10794);
or U11240 (N_11240,N_10831,N_10855);
or U11241 (N_11241,N_10808,N_10937);
nand U11242 (N_11242,N_10842,N_10888);
or U11243 (N_11243,N_10965,N_10976);
or U11244 (N_11244,N_10895,N_10916);
and U11245 (N_11245,N_10966,N_10798);
or U11246 (N_11246,N_10988,N_10881);
or U11247 (N_11247,N_10785,N_10821);
nand U11248 (N_11248,N_10914,N_10828);
and U11249 (N_11249,N_10881,N_10838);
nor U11250 (N_11250,N_11002,N_11149);
or U11251 (N_11251,N_11192,N_11176);
xor U11252 (N_11252,N_11233,N_11068);
nor U11253 (N_11253,N_11171,N_11000);
xor U11254 (N_11254,N_11051,N_11064);
nand U11255 (N_11255,N_11090,N_11080);
nor U11256 (N_11256,N_11032,N_11052);
nor U11257 (N_11257,N_11040,N_11054);
and U11258 (N_11258,N_11129,N_11136);
and U11259 (N_11259,N_11004,N_11109);
nand U11260 (N_11260,N_11062,N_11173);
xnor U11261 (N_11261,N_11200,N_11238);
and U11262 (N_11262,N_11013,N_11063);
and U11263 (N_11263,N_11222,N_11061);
and U11264 (N_11264,N_11150,N_11164);
nand U11265 (N_11265,N_11014,N_11157);
xnor U11266 (N_11266,N_11087,N_11199);
or U11267 (N_11267,N_11135,N_11028);
nand U11268 (N_11268,N_11158,N_11193);
nand U11269 (N_11269,N_11147,N_11019);
xnor U11270 (N_11270,N_11196,N_11152);
nor U11271 (N_11271,N_11031,N_11160);
nand U11272 (N_11272,N_11228,N_11181);
nor U11273 (N_11273,N_11104,N_11183);
nor U11274 (N_11274,N_11131,N_11094);
nand U11275 (N_11275,N_11122,N_11232);
nand U11276 (N_11276,N_11174,N_11120);
nand U11277 (N_11277,N_11175,N_11026);
xor U11278 (N_11278,N_11075,N_11249);
nor U11279 (N_11279,N_11151,N_11029);
and U11280 (N_11280,N_11037,N_11108);
nor U11281 (N_11281,N_11177,N_11143);
or U11282 (N_11282,N_11214,N_11021);
nor U11283 (N_11283,N_11246,N_11025);
or U11284 (N_11284,N_11016,N_11146);
nor U11285 (N_11285,N_11206,N_11119);
xnor U11286 (N_11286,N_11057,N_11117);
nand U11287 (N_11287,N_11212,N_11209);
nand U11288 (N_11288,N_11207,N_11053);
and U11289 (N_11289,N_11069,N_11163);
nand U11290 (N_11290,N_11186,N_11070);
nor U11291 (N_11291,N_11015,N_11046);
and U11292 (N_11292,N_11034,N_11114);
xnor U11293 (N_11293,N_11167,N_11049);
nor U11294 (N_11294,N_11097,N_11170);
nor U11295 (N_11295,N_11127,N_11191);
or U11296 (N_11296,N_11009,N_11010);
nor U11297 (N_11297,N_11126,N_11165);
nand U11298 (N_11298,N_11081,N_11133);
nor U11299 (N_11299,N_11156,N_11103);
xor U11300 (N_11300,N_11239,N_11017);
or U11301 (N_11301,N_11182,N_11084);
nor U11302 (N_11302,N_11138,N_11036);
xnor U11303 (N_11303,N_11216,N_11027);
or U11304 (N_11304,N_11047,N_11226);
and U11305 (N_11305,N_11142,N_11022);
xnor U11306 (N_11306,N_11244,N_11240);
xnor U11307 (N_11307,N_11130,N_11153);
nand U11308 (N_11308,N_11248,N_11145);
nor U11309 (N_11309,N_11106,N_11030);
nor U11310 (N_11310,N_11161,N_11189);
and U11311 (N_11311,N_11201,N_11033);
nand U11312 (N_11312,N_11217,N_11243);
xor U11313 (N_11313,N_11166,N_11237);
nor U11314 (N_11314,N_11071,N_11005);
or U11315 (N_11315,N_11065,N_11188);
or U11316 (N_11316,N_11213,N_11059);
or U11317 (N_11317,N_11091,N_11221);
nor U11318 (N_11318,N_11204,N_11007);
xnor U11319 (N_11319,N_11086,N_11154);
nand U11320 (N_11320,N_11144,N_11008);
or U11321 (N_11321,N_11044,N_11045);
or U11322 (N_11322,N_11218,N_11234);
and U11323 (N_11323,N_11236,N_11098);
nand U11324 (N_11324,N_11134,N_11224);
nand U11325 (N_11325,N_11060,N_11208);
nand U11326 (N_11326,N_11185,N_11024);
nand U11327 (N_11327,N_11194,N_11159);
nor U11328 (N_11328,N_11168,N_11006);
or U11329 (N_11329,N_11125,N_11211);
nand U11330 (N_11330,N_11227,N_11123);
nor U11331 (N_11331,N_11105,N_11078);
nand U11332 (N_11332,N_11148,N_11231);
xnor U11333 (N_11333,N_11111,N_11110);
nor U11334 (N_11334,N_11179,N_11095);
xnor U11335 (N_11335,N_11116,N_11018);
or U11336 (N_11336,N_11203,N_11137);
nor U11337 (N_11337,N_11077,N_11225);
xnor U11338 (N_11338,N_11169,N_11083);
and U11339 (N_11339,N_11139,N_11118);
and U11340 (N_11340,N_11195,N_11223);
nand U11341 (N_11341,N_11241,N_11011);
nand U11342 (N_11342,N_11082,N_11162);
and U11343 (N_11343,N_11210,N_11205);
nor U11344 (N_11344,N_11102,N_11190);
and U11345 (N_11345,N_11041,N_11115);
or U11346 (N_11346,N_11215,N_11020);
xor U11347 (N_11347,N_11229,N_11132);
nand U11348 (N_11348,N_11187,N_11178);
nor U11349 (N_11349,N_11112,N_11067);
nand U11350 (N_11350,N_11073,N_11124);
nand U11351 (N_11351,N_11096,N_11058);
nand U11352 (N_11352,N_11001,N_11056);
or U11353 (N_11353,N_11089,N_11072);
or U11354 (N_11354,N_11085,N_11055);
and U11355 (N_11355,N_11100,N_11099);
or U11356 (N_11356,N_11092,N_11235);
or U11357 (N_11357,N_11113,N_11039);
nand U11358 (N_11358,N_11074,N_11140);
nor U11359 (N_11359,N_11184,N_11180);
xor U11360 (N_11360,N_11066,N_11141);
xnor U11361 (N_11361,N_11198,N_11012);
xnor U11362 (N_11362,N_11023,N_11242);
nand U11363 (N_11363,N_11202,N_11035);
nor U11364 (N_11364,N_11043,N_11245);
and U11365 (N_11365,N_11128,N_11042);
xnor U11366 (N_11366,N_11121,N_11155);
and U11367 (N_11367,N_11003,N_11172);
xor U11368 (N_11368,N_11101,N_11050);
and U11369 (N_11369,N_11247,N_11048);
nand U11370 (N_11370,N_11079,N_11107);
or U11371 (N_11371,N_11038,N_11197);
nor U11372 (N_11372,N_11088,N_11219);
nand U11373 (N_11373,N_11220,N_11076);
xor U11374 (N_11374,N_11230,N_11093);
or U11375 (N_11375,N_11023,N_11071);
and U11376 (N_11376,N_11141,N_11006);
or U11377 (N_11377,N_11038,N_11032);
and U11378 (N_11378,N_11248,N_11227);
nor U11379 (N_11379,N_11220,N_11147);
nor U11380 (N_11380,N_11159,N_11192);
and U11381 (N_11381,N_11159,N_11061);
xnor U11382 (N_11382,N_11155,N_11098);
and U11383 (N_11383,N_11020,N_11216);
and U11384 (N_11384,N_11186,N_11128);
xor U11385 (N_11385,N_11163,N_11131);
or U11386 (N_11386,N_11213,N_11029);
or U11387 (N_11387,N_11202,N_11073);
nor U11388 (N_11388,N_11181,N_11185);
xnor U11389 (N_11389,N_11163,N_11128);
nor U11390 (N_11390,N_11218,N_11055);
nand U11391 (N_11391,N_11115,N_11000);
xnor U11392 (N_11392,N_11027,N_11147);
or U11393 (N_11393,N_11070,N_11146);
nor U11394 (N_11394,N_11214,N_11058);
and U11395 (N_11395,N_11074,N_11223);
nor U11396 (N_11396,N_11241,N_11128);
nand U11397 (N_11397,N_11109,N_11100);
nor U11398 (N_11398,N_11138,N_11040);
and U11399 (N_11399,N_11042,N_11124);
xor U11400 (N_11400,N_11013,N_11192);
xor U11401 (N_11401,N_11020,N_11212);
and U11402 (N_11402,N_11032,N_11129);
or U11403 (N_11403,N_11121,N_11073);
nor U11404 (N_11404,N_11081,N_11229);
xnor U11405 (N_11405,N_11089,N_11222);
and U11406 (N_11406,N_11101,N_11148);
and U11407 (N_11407,N_11043,N_11103);
and U11408 (N_11408,N_11182,N_11119);
and U11409 (N_11409,N_11084,N_11009);
and U11410 (N_11410,N_11009,N_11146);
xnor U11411 (N_11411,N_11030,N_11174);
and U11412 (N_11412,N_11036,N_11106);
nor U11413 (N_11413,N_11039,N_11169);
and U11414 (N_11414,N_11247,N_11099);
and U11415 (N_11415,N_11141,N_11009);
xnor U11416 (N_11416,N_11103,N_11206);
xor U11417 (N_11417,N_11142,N_11077);
nand U11418 (N_11418,N_11091,N_11242);
or U11419 (N_11419,N_11143,N_11088);
xnor U11420 (N_11420,N_11064,N_11163);
nand U11421 (N_11421,N_11179,N_11193);
xor U11422 (N_11422,N_11183,N_11182);
nand U11423 (N_11423,N_11145,N_11037);
or U11424 (N_11424,N_11046,N_11188);
nand U11425 (N_11425,N_11196,N_11089);
or U11426 (N_11426,N_11144,N_11031);
or U11427 (N_11427,N_11200,N_11129);
or U11428 (N_11428,N_11247,N_11102);
and U11429 (N_11429,N_11046,N_11138);
and U11430 (N_11430,N_11210,N_11229);
nor U11431 (N_11431,N_11123,N_11166);
nand U11432 (N_11432,N_11129,N_11139);
xnor U11433 (N_11433,N_11053,N_11096);
nand U11434 (N_11434,N_11158,N_11145);
nor U11435 (N_11435,N_11080,N_11070);
or U11436 (N_11436,N_11001,N_11234);
nand U11437 (N_11437,N_11132,N_11160);
xor U11438 (N_11438,N_11034,N_11083);
xor U11439 (N_11439,N_11203,N_11195);
nand U11440 (N_11440,N_11049,N_11150);
xor U11441 (N_11441,N_11064,N_11158);
and U11442 (N_11442,N_11248,N_11141);
xor U11443 (N_11443,N_11090,N_11010);
or U11444 (N_11444,N_11172,N_11002);
nor U11445 (N_11445,N_11090,N_11099);
nor U11446 (N_11446,N_11119,N_11092);
xor U11447 (N_11447,N_11242,N_11232);
nor U11448 (N_11448,N_11122,N_11132);
and U11449 (N_11449,N_11075,N_11118);
and U11450 (N_11450,N_11242,N_11046);
and U11451 (N_11451,N_11038,N_11128);
and U11452 (N_11452,N_11021,N_11130);
xor U11453 (N_11453,N_11049,N_11001);
xor U11454 (N_11454,N_11118,N_11115);
nor U11455 (N_11455,N_11222,N_11039);
xor U11456 (N_11456,N_11029,N_11019);
nand U11457 (N_11457,N_11183,N_11087);
xnor U11458 (N_11458,N_11136,N_11068);
xnor U11459 (N_11459,N_11110,N_11016);
or U11460 (N_11460,N_11206,N_11074);
or U11461 (N_11461,N_11236,N_11174);
or U11462 (N_11462,N_11009,N_11030);
nor U11463 (N_11463,N_11015,N_11202);
nand U11464 (N_11464,N_11119,N_11088);
nor U11465 (N_11465,N_11011,N_11175);
nor U11466 (N_11466,N_11092,N_11087);
xnor U11467 (N_11467,N_11066,N_11022);
nor U11468 (N_11468,N_11245,N_11063);
and U11469 (N_11469,N_11179,N_11241);
or U11470 (N_11470,N_11064,N_11132);
or U11471 (N_11471,N_11037,N_11159);
nand U11472 (N_11472,N_11093,N_11218);
nor U11473 (N_11473,N_11084,N_11015);
nand U11474 (N_11474,N_11123,N_11014);
xor U11475 (N_11475,N_11149,N_11162);
nor U11476 (N_11476,N_11173,N_11023);
nor U11477 (N_11477,N_11218,N_11132);
or U11478 (N_11478,N_11186,N_11155);
nor U11479 (N_11479,N_11058,N_11209);
and U11480 (N_11480,N_11088,N_11170);
or U11481 (N_11481,N_11209,N_11124);
and U11482 (N_11482,N_11056,N_11090);
nor U11483 (N_11483,N_11170,N_11108);
nand U11484 (N_11484,N_11038,N_11122);
xor U11485 (N_11485,N_11236,N_11064);
nor U11486 (N_11486,N_11105,N_11198);
or U11487 (N_11487,N_11124,N_11134);
or U11488 (N_11488,N_11042,N_11112);
and U11489 (N_11489,N_11140,N_11024);
nand U11490 (N_11490,N_11102,N_11038);
or U11491 (N_11491,N_11237,N_11024);
xor U11492 (N_11492,N_11085,N_11067);
or U11493 (N_11493,N_11184,N_11089);
and U11494 (N_11494,N_11070,N_11099);
nand U11495 (N_11495,N_11041,N_11087);
and U11496 (N_11496,N_11013,N_11225);
nand U11497 (N_11497,N_11061,N_11143);
xnor U11498 (N_11498,N_11028,N_11140);
xor U11499 (N_11499,N_11132,N_11172);
nor U11500 (N_11500,N_11251,N_11471);
nor U11501 (N_11501,N_11398,N_11314);
and U11502 (N_11502,N_11412,N_11420);
nor U11503 (N_11503,N_11435,N_11271);
xnor U11504 (N_11504,N_11369,N_11440);
and U11505 (N_11505,N_11282,N_11352);
nor U11506 (N_11506,N_11430,N_11351);
or U11507 (N_11507,N_11274,N_11312);
nor U11508 (N_11508,N_11275,N_11496);
nor U11509 (N_11509,N_11475,N_11405);
and U11510 (N_11510,N_11468,N_11480);
nand U11511 (N_11511,N_11451,N_11493);
nand U11512 (N_11512,N_11368,N_11490);
xor U11513 (N_11513,N_11346,N_11392);
nor U11514 (N_11514,N_11305,N_11456);
or U11515 (N_11515,N_11260,N_11444);
and U11516 (N_11516,N_11272,N_11299);
nand U11517 (N_11517,N_11259,N_11486);
or U11518 (N_11518,N_11296,N_11457);
and U11519 (N_11519,N_11337,N_11421);
and U11520 (N_11520,N_11443,N_11488);
or U11521 (N_11521,N_11393,N_11336);
and U11522 (N_11522,N_11283,N_11495);
or U11523 (N_11523,N_11466,N_11441);
xnor U11524 (N_11524,N_11343,N_11463);
or U11525 (N_11525,N_11257,N_11325);
nor U11526 (N_11526,N_11404,N_11384);
nor U11527 (N_11527,N_11254,N_11383);
nand U11528 (N_11528,N_11400,N_11303);
and U11529 (N_11529,N_11419,N_11379);
and U11530 (N_11530,N_11386,N_11367);
nand U11531 (N_11531,N_11285,N_11313);
and U11532 (N_11532,N_11366,N_11357);
xnor U11533 (N_11533,N_11338,N_11418);
or U11534 (N_11534,N_11479,N_11464);
xnor U11535 (N_11535,N_11447,N_11465);
xor U11536 (N_11536,N_11494,N_11356);
nand U11537 (N_11537,N_11327,N_11453);
nor U11538 (N_11538,N_11316,N_11281);
nor U11539 (N_11539,N_11310,N_11334);
nand U11540 (N_11540,N_11446,N_11333);
nor U11541 (N_11541,N_11395,N_11317);
and U11542 (N_11542,N_11311,N_11360);
nand U11543 (N_11543,N_11270,N_11458);
or U11544 (N_11544,N_11492,N_11345);
xnor U11545 (N_11545,N_11497,N_11349);
or U11546 (N_11546,N_11477,N_11280);
nor U11547 (N_11547,N_11445,N_11476);
nand U11548 (N_11548,N_11307,N_11295);
nor U11549 (N_11549,N_11264,N_11429);
and U11550 (N_11550,N_11373,N_11265);
and U11551 (N_11551,N_11425,N_11415);
and U11552 (N_11552,N_11442,N_11321);
nor U11553 (N_11553,N_11335,N_11365);
xnor U11554 (N_11554,N_11481,N_11407);
nor U11555 (N_11555,N_11328,N_11382);
nand U11556 (N_11556,N_11426,N_11250);
xnor U11557 (N_11557,N_11266,N_11460);
and U11558 (N_11558,N_11252,N_11498);
nand U11559 (N_11559,N_11402,N_11487);
and U11560 (N_11560,N_11406,N_11473);
nor U11561 (N_11561,N_11306,N_11290);
and U11562 (N_11562,N_11267,N_11399);
nor U11563 (N_11563,N_11339,N_11376);
nand U11564 (N_11564,N_11436,N_11347);
nor U11565 (N_11565,N_11273,N_11268);
nand U11566 (N_11566,N_11315,N_11432);
nand U11567 (N_11567,N_11291,N_11454);
nor U11568 (N_11568,N_11455,N_11323);
xor U11569 (N_11569,N_11380,N_11298);
nand U11570 (N_11570,N_11396,N_11439);
or U11571 (N_11571,N_11474,N_11324);
and U11572 (N_11572,N_11340,N_11363);
nor U11573 (N_11573,N_11362,N_11284);
xor U11574 (N_11574,N_11329,N_11433);
and U11575 (N_11575,N_11297,N_11422);
nor U11576 (N_11576,N_11279,N_11469);
xnor U11577 (N_11577,N_11423,N_11342);
and U11578 (N_11578,N_11318,N_11322);
and U11579 (N_11579,N_11332,N_11377);
nand U11580 (N_11580,N_11350,N_11277);
nor U11581 (N_11581,N_11408,N_11416);
and U11582 (N_11582,N_11253,N_11262);
nor U11583 (N_11583,N_11459,N_11410);
nor U11584 (N_11584,N_11258,N_11438);
xnor U11585 (N_11585,N_11427,N_11448);
nand U11586 (N_11586,N_11403,N_11478);
xor U11587 (N_11587,N_11491,N_11301);
nor U11588 (N_11588,N_11302,N_11385);
or U11589 (N_11589,N_11292,N_11359);
or U11590 (N_11590,N_11355,N_11326);
nand U11591 (N_11591,N_11387,N_11483);
nor U11592 (N_11592,N_11358,N_11341);
xor U11593 (N_11593,N_11289,N_11391);
nor U11594 (N_11594,N_11381,N_11348);
xnor U11595 (N_11595,N_11411,N_11278);
xor U11596 (N_11596,N_11388,N_11294);
or U11597 (N_11597,N_11320,N_11309);
nor U11598 (N_11598,N_11417,N_11390);
and U11599 (N_11599,N_11344,N_11485);
and U11600 (N_11600,N_11434,N_11304);
xnor U11601 (N_11601,N_11462,N_11397);
or U11602 (N_11602,N_11300,N_11261);
xnor U11603 (N_11603,N_11353,N_11375);
nor U11604 (N_11604,N_11293,N_11489);
nand U11605 (N_11605,N_11437,N_11389);
and U11606 (N_11606,N_11330,N_11431);
nand U11607 (N_11607,N_11374,N_11482);
nand U11608 (N_11608,N_11409,N_11499);
xor U11609 (N_11609,N_11461,N_11286);
nor U11610 (N_11610,N_11450,N_11287);
and U11611 (N_11611,N_11256,N_11401);
nand U11612 (N_11612,N_11276,N_11472);
nor U11613 (N_11613,N_11414,N_11370);
or U11614 (N_11614,N_11452,N_11378);
or U11615 (N_11615,N_11394,N_11319);
or U11616 (N_11616,N_11428,N_11467);
and U11617 (N_11617,N_11354,N_11255);
nand U11618 (N_11618,N_11424,N_11449);
and U11619 (N_11619,N_11331,N_11308);
nand U11620 (N_11620,N_11372,N_11484);
nor U11621 (N_11621,N_11413,N_11263);
or U11622 (N_11622,N_11364,N_11470);
or U11623 (N_11623,N_11288,N_11269);
xnor U11624 (N_11624,N_11361,N_11371);
and U11625 (N_11625,N_11407,N_11258);
and U11626 (N_11626,N_11439,N_11357);
nand U11627 (N_11627,N_11469,N_11410);
nor U11628 (N_11628,N_11489,N_11423);
xnor U11629 (N_11629,N_11460,N_11477);
and U11630 (N_11630,N_11303,N_11480);
xnor U11631 (N_11631,N_11317,N_11342);
nor U11632 (N_11632,N_11458,N_11272);
or U11633 (N_11633,N_11420,N_11458);
nor U11634 (N_11634,N_11417,N_11358);
nand U11635 (N_11635,N_11272,N_11416);
xor U11636 (N_11636,N_11295,N_11302);
nand U11637 (N_11637,N_11312,N_11390);
nor U11638 (N_11638,N_11311,N_11332);
nor U11639 (N_11639,N_11470,N_11371);
nor U11640 (N_11640,N_11349,N_11316);
xnor U11641 (N_11641,N_11274,N_11372);
or U11642 (N_11642,N_11352,N_11267);
xor U11643 (N_11643,N_11358,N_11340);
nor U11644 (N_11644,N_11421,N_11345);
or U11645 (N_11645,N_11431,N_11465);
nand U11646 (N_11646,N_11359,N_11462);
xnor U11647 (N_11647,N_11440,N_11329);
or U11648 (N_11648,N_11264,N_11317);
and U11649 (N_11649,N_11418,N_11278);
and U11650 (N_11650,N_11282,N_11414);
and U11651 (N_11651,N_11359,N_11420);
xnor U11652 (N_11652,N_11281,N_11420);
nor U11653 (N_11653,N_11401,N_11285);
or U11654 (N_11654,N_11250,N_11323);
or U11655 (N_11655,N_11395,N_11324);
and U11656 (N_11656,N_11418,N_11463);
nor U11657 (N_11657,N_11347,N_11443);
and U11658 (N_11658,N_11478,N_11370);
nand U11659 (N_11659,N_11419,N_11360);
nand U11660 (N_11660,N_11447,N_11402);
xor U11661 (N_11661,N_11415,N_11295);
and U11662 (N_11662,N_11315,N_11442);
xor U11663 (N_11663,N_11401,N_11309);
nor U11664 (N_11664,N_11493,N_11316);
xor U11665 (N_11665,N_11427,N_11442);
and U11666 (N_11666,N_11485,N_11315);
nand U11667 (N_11667,N_11285,N_11470);
or U11668 (N_11668,N_11265,N_11499);
nor U11669 (N_11669,N_11269,N_11437);
xor U11670 (N_11670,N_11288,N_11302);
xnor U11671 (N_11671,N_11495,N_11463);
nor U11672 (N_11672,N_11451,N_11360);
xor U11673 (N_11673,N_11385,N_11421);
and U11674 (N_11674,N_11341,N_11254);
nor U11675 (N_11675,N_11361,N_11484);
nand U11676 (N_11676,N_11322,N_11276);
nand U11677 (N_11677,N_11296,N_11345);
xnor U11678 (N_11678,N_11323,N_11267);
nor U11679 (N_11679,N_11390,N_11349);
and U11680 (N_11680,N_11267,N_11438);
xor U11681 (N_11681,N_11487,N_11340);
and U11682 (N_11682,N_11357,N_11259);
nand U11683 (N_11683,N_11343,N_11301);
xor U11684 (N_11684,N_11341,N_11481);
xor U11685 (N_11685,N_11350,N_11424);
or U11686 (N_11686,N_11379,N_11411);
nor U11687 (N_11687,N_11422,N_11307);
nor U11688 (N_11688,N_11478,N_11469);
or U11689 (N_11689,N_11440,N_11293);
and U11690 (N_11690,N_11388,N_11300);
nand U11691 (N_11691,N_11331,N_11416);
nand U11692 (N_11692,N_11281,N_11499);
or U11693 (N_11693,N_11332,N_11470);
nor U11694 (N_11694,N_11266,N_11273);
xnor U11695 (N_11695,N_11470,N_11453);
nor U11696 (N_11696,N_11447,N_11350);
nand U11697 (N_11697,N_11294,N_11261);
nor U11698 (N_11698,N_11269,N_11337);
nor U11699 (N_11699,N_11392,N_11453);
and U11700 (N_11700,N_11405,N_11385);
and U11701 (N_11701,N_11386,N_11328);
nor U11702 (N_11702,N_11338,N_11275);
and U11703 (N_11703,N_11428,N_11477);
xor U11704 (N_11704,N_11291,N_11282);
or U11705 (N_11705,N_11269,N_11379);
xnor U11706 (N_11706,N_11406,N_11426);
and U11707 (N_11707,N_11496,N_11440);
xnor U11708 (N_11708,N_11326,N_11493);
or U11709 (N_11709,N_11463,N_11496);
and U11710 (N_11710,N_11343,N_11376);
xnor U11711 (N_11711,N_11290,N_11254);
xnor U11712 (N_11712,N_11357,N_11271);
xor U11713 (N_11713,N_11466,N_11250);
nand U11714 (N_11714,N_11457,N_11489);
nor U11715 (N_11715,N_11360,N_11347);
nor U11716 (N_11716,N_11444,N_11447);
and U11717 (N_11717,N_11393,N_11433);
xor U11718 (N_11718,N_11303,N_11319);
and U11719 (N_11719,N_11263,N_11422);
and U11720 (N_11720,N_11445,N_11257);
nor U11721 (N_11721,N_11312,N_11293);
nand U11722 (N_11722,N_11322,N_11449);
nand U11723 (N_11723,N_11415,N_11354);
and U11724 (N_11724,N_11327,N_11325);
xnor U11725 (N_11725,N_11420,N_11452);
nand U11726 (N_11726,N_11382,N_11413);
or U11727 (N_11727,N_11381,N_11382);
xor U11728 (N_11728,N_11267,N_11372);
nand U11729 (N_11729,N_11460,N_11260);
xor U11730 (N_11730,N_11388,N_11260);
or U11731 (N_11731,N_11498,N_11304);
xnor U11732 (N_11732,N_11341,N_11416);
xnor U11733 (N_11733,N_11409,N_11352);
nor U11734 (N_11734,N_11415,N_11370);
or U11735 (N_11735,N_11478,N_11367);
and U11736 (N_11736,N_11296,N_11342);
xnor U11737 (N_11737,N_11271,N_11252);
xnor U11738 (N_11738,N_11473,N_11480);
or U11739 (N_11739,N_11399,N_11467);
nand U11740 (N_11740,N_11417,N_11447);
nor U11741 (N_11741,N_11255,N_11318);
nor U11742 (N_11742,N_11252,N_11291);
or U11743 (N_11743,N_11359,N_11430);
xnor U11744 (N_11744,N_11454,N_11448);
xor U11745 (N_11745,N_11436,N_11419);
nor U11746 (N_11746,N_11252,N_11440);
xor U11747 (N_11747,N_11494,N_11295);
nor U11748 (N_11748,N_11358,N_11395);
and U11749 (N_11749,N_11375,N_11401);
xnor U11750 (N_11750,N_11719,N_11699);
nand U11751 (N_11751,N_11731,N_11655);
nand U11752 (N_11752,N_11665,N_11529);
nor U11753 (N_11753,N_11684,N_11634);
xor U11754 (N_11754,N_11696,N_11693);
nand U11755 (N_11755,N_11686,N_11552);
nor U11756 (N_11756,N_11536,N_11593);
and U11757 (N_11757,N_11578,N_11538);
xor U11758 (N_11758,N_11666,N_11690);
xor U11759 (N_11759,N_11742,N_11676);
or U11760 (N_11760,N_11592,N_11501);
xor U11761 (N_11761,N_11576,N_11632);
xor U11762 (N_11762,N_11747,N_11626);
xor U11763 (N_11763,N_11688,N_11566);
nand U11764 (N_11764,N_11553,N_11681);
nor U11765 (N_11765,N_11711,N_11638);
xnor U11766 (N_11766,N_11737,N_11509);
nand U11767 (N_11767,N_11672,N_11537);
and U11768 (N_11768,N_11570,N_11730);
or U11769 (N_11769,N_11703,N_11528);
xnor U11770 (N_11770,N_11544,N_11519);
xor U11771 (N_11771,N_11667,N_11645);
xor U11772 (N_11772,N_11517,N_11649);
and U11773 (N_11773,N_11714,N_11694);
xor U11774 (N_11774,N_11644,N_11643);
nor U11775 (N_11775,N_11627,N_11591);
and U11776 (N_11776,N_11506,N_11505);
and U11777 (N_11777,N_11508,N_11654);
nand U11778 (N_11778,N_11700,N_11746);
or U11779 (N_11779,N_11616,N_11574);
or U11780 (N_11780,N_11594,N_11522);
xnor U11781 (N_11781,N_11656,N_11702);
and U11782 (N_11782,N_11743,N_11585);
xnor U11783 (N_11783,N_11558,N_11604);
xnor U11784 (N_11784,N_11733,N_11586);
xor U11785 (N_11785,N_11587,N_11677);
xor U11786 (N_11786,N_11512,N_11521);
xnor U11787 (N_11787,N_11556,N_11560);
or U11788 (N_11788,N_11642,N_11657);
or U11789 (N_11789,N_11662,N_11663);
nor U11790 (N_11790,N_11562,N_11597);
xnor U11791 (N_11791,N_11631,N_11674);
and U11792 (N_11792,N_11748,N_11708);
or U11793 (N_11793,N_11736,N_11550);
xnor U11794 (N_11794,N_11596,N_11551);
and U11795 (N_11795,N_11607,N_11671);
nor U11796 (N_11796,N_11510,N_11739);
and U11797 (N_11797,N_11548,N_11695);
and U11798 (N_11798,N_11727,N_11575);
or U11799 (N_11799,N_11641,N_11682);
nand U11800 (N_11800,N_11543,N_11534);
or U11801 (N_11801,N_11650,N_11615);
or U11802 (N_11802,N_11706,N_11533);
nor U11803 (N_11803,N_11687,N_11721);
and U11804 (N_11804,N_11648,N_11569);
xor U11805 (N_11805,N_11541,N_11523);
or U11806 (N_11806,N_11633,N_11602);
nand U11807 (N_11807,N_11680,N_11659);
nor U11808 (N_11808,N_11514,N_11526);
xnor U11809 (N_11809,N_11718,N_11564);
nor U11810 (N_11810,N_11668,N_11625);
and U11811 (N_11811,N_11571,N_11636);
or U11812 (N_11812,N_11545,N_11673);
or U11813 (N_11813,N_11549,N_11669);
nor U11814 (N_11814,N_11697,N_11664);
or U11815 (N_11815,N_11606,N_11608);
or U11816 (N_11816,N_11647,N_11722);
and U11817 (N_11817,N_11715,N_11609);
nand U11818 (N_11818,N_11502,N_11621);
or U11819 (N_11819,N_11653,N_11559);
and U11820 (N_11820,N_11723,N_11651);
xor U11821 (N_11821,N_11590,N_11527);
or U11822 (N_11822,N_11554,N_11623);
and U11823 (N_11823,N_11745,N_11735);
and U11824 (N_11824,N_11709,N_11704);
or U11825 (N_11825,N_11573,N_11613);
nor U11826 (N_11826,N_11741,N_11691);
nor U11827 (N_11827,N_11614,N_11732);
and U11828 (N_11828,N_11675,N_11525);
xor U11829 (N_11829,N_11532,N_11720);
xor U11830 (N_11830,N_11535,N_11520);
nand U11831 (N_11831,N_11629,N_11503);
xnor U11832 (N_11832,N_11725,N_11622);
or U11833 (N_11833,N_11581,N_11580);
or U11834 (N_11834,N_11524,N_11716);
and U11835 (N_11835,N_11572,N_11692);
and U11836 (N_11836,N_11628,N_11710);
or U11837 (N_11837,N_11530,N_11579);
xnor U11838 (N_11838,N_11712,N_11547);
nor U11839 (N_11839,N_11707,N_11515);
or U11840 (N_11840,N_11583,N_11611);
and U11841 (N_11841,N_11740,N_11661);
nor U11842 (N_11842,N_11504,N_11595);
xor U11843 (N_11843,N_11635,N_11652);
and U11844 (N_11844,N_11539,N_11640);
xor U11845 (N_11845,N_11749,N_11679);
and U11846 (N_11846,N_11738,N_11546);
xor U11847 (N_11847,N_11705,N_11624);
nand U11848 (N_11848,N_11701,N_11620);
or U11849 (N_11849,N_11658,N_11513);
nand U11850 (N_11850,N_11577,N_11518);
nor U11851 (N_11851,N_11588,N_11612);
xnor U11852 (N_11852,N_11600,N_11683);
or U11853 (N_11853,N_11542,N_11555);
nor U11854 (N_11854,N_11557,N_11582);
nor U11855 (N_11855,N_11726,N_11610);
nor U11856 (N_11856,N_11617,N_11618);
and U11857 (N_11857,N_11729,N_11744);
or U11858 (N_11858,N_11531,N_11717);
nor U11859 (N_11859,N_11678,N_11619);
and U11860 (N_11860,N_11601,N_11698);
nor U11861 (N_11861,N_11637,N_11670);
nor U11862 (N_11862,N_11646,N_11728);
nand U11863 (N_11863,N_11507,N_11685);
and U11864 (N_11864,N_11540,N_11598);
nand U11865 (N_11865,N_11713,N_11511);
and U11866 (N_11866,N_11516,N_11724);
and U11867 (N_11867,N_11605,N_11689);
xnor U11868 (N_11868,N_11603,N_11565);
nor U11869 (N_11869,N_11630,N_11639);
and U11870 (N_11870,N_11563,N_11734);
nand U11871 (N_11871,N_11568,N_11584);
and U11872 (N_11872,N_11567,N_11561);
or U11873 (N_11873,N_11500,N_11589);
xnor U11874 (N_11874,N_11599,N_11660);
xor U11875 (N_11875,N_11607,N_11595);
xnor U11876 (N_11876,N_11680,N_11586);
nor U11877 (N_11877,N_11639,N_11660);
or U11878 (N_11878,N_11718,N_11652);
and U11879 (N_11879,N_11734,N_11510);
nor U11880 (N_11880,N_11585,N_11522);
nor U11881 (N_11881,N_11656,N_11522);
or U11882 (N_11882,N_11704,N_11646);
nand U11883 (N_11883,N_11669,N_11595);
nand U11884 (N_11884,N_11506,N_11598);
and U11885 (N_11885,N_11686,N_11688);
and U11886 (N_11886,N_11616,N_11690);
nand U11887 (N_11887,N_11578,N_11609);
or U11888 (N_11888,N_11672,N_11614);
and U11889 (N_11889,N_11694,N_11623);
xnor U11890 (N_11890,N_11573,N_11611);
xor U11891 (N_11891,N_11510,N_11530);
and U11892 (N_11892,N_11569,N_11566);
or U11893 (N_11893,N_11714,N_11730);
nand U11894 (N_11894,N_11669,N_11691);
nand U11895 (N_11895,N_11613,N_11683);
nand U11896 (N_11896,N_11610,N_11570);
nor U11897 (N_11897,N_11731,N_11738);
and U11898 (N_11898,N_11551,N_11520);
nor U11899 (N_11899,N_11533,N_11532);
nor U11900 (N_11900,N_11522,N_11706);
nor U11901 (N_11901,N_11707,N_11639);
xor U11902 (N_11902,N_11631,N_11546);
xor U11903 (N_11903,N_11713,N_11577);
and U11904 (N_11904,N_11675,N_11631);
nand U11905 (N_11905,N_11565,N_11729);
and U11906 (N_11906,N_11689,N_11663);
xor U11907 (N_11907,N_11552,N_11523);
nand U11908 (N_11908,N_11597,N_11696);
xnor U11909 (N_11909,N_11630,N_11656);
nand U11910 (N_11910,N_11583,N_11524);
or U11911 (N_11911,N_11719,N_11516);
and U11912 (N_11912,N_11612,N_11593);
nor U11913 (N_11913,N_11531,N_11616);
xnor U11914 (N_11914,N_11522,N_11602);
and U11915 (N_11915,N_11553,N_11500);
xnor U11916 (N_11916,N_11565,N_11526);
and U11917 (N_11917,N_11718,N_11568);
and U11918 (N_11918,N_11637,N_11602);
xor U11919 (N_11919,N_11626,N_11664);
or U11920 (N_11920,N_11517,N_11689);
or U11921 (N_11921,N_11612,N_11651);
nand U11922 (N_11922,N_11514,N_11727);
or U11923 (N_11923,N_11629,N_11606);
or U11924 (N_11924,N_11552,N_11724);
or U11925 (N_11925,N_11713,N_11582);
nand U11926 (N_11926,N_11526,N_11530);
or U11927 (N_11927,N_11585,N_11613);
nor U11928 (N_11928,N_11530,N_11695);
nor U11929 (N_11929,N_11645,N_11627);
and U11930 (N_11930,N_11567,N_11525);
and U11931 (N_11931,N_11554,N_11704);
nor U11932 (N_11932,N_11717,N_11657);
nand U11933 (N_11933,N_11725,N_11670);
or U11934 (N_11934,N_11571,N_11742);
xnor U11935 (N_11935,N_11700,N_11669);
or U11936 (N_11936,N_11597,N_11583);
nand U11937 (N_11937,N_11580,N_11537);
nand U11938 (N_11938,N_11701,N_11561);
and U11939 (N_11939,N_11701,N_11662);
nor U11940 (N_11940,N_11700,N_11656);
and U11941 (N_11941,N_11701,N_11698);
xnor U11942 (N_11942,N_11540,N_11664);
nor U11943 (N_11943,N_11667,N_11599);
or U11944 (N_11944,N_11561,N_11603);
nand U11945 (N_11945,N_11706,N_11710);
and U11946 (N_11946,N_11517,N_11663);
xnor U11947 (N_11947,N_11682,N_11634);
and U11948 (N_11948,N_11704,N_11597);
or U11949 (N_11949,N_11728,N_11736);
nand U11950 (N_11950,N_11700,N_11689);
nor U11951 (N_11951,N_11521,N_11607);
nor U11952 (N_11952,N_11580,N_11583);
xnor U11953 (N_11953,N_11685,N_11603);
and U11954 (N_11954,N_11614,N_11722);
nand U11955 (N_11955,N_11541,N_11670);
nand U11956 (N_11956,N_11576,N_11564);
nor U11957 (N_11957,N_11738,N_11558);
nor U11958 (N_11958,N_11547,N_11597);
nand U11959 (N_11959,N_11630,N_11734);
or U11960 (N_11960,N_11663,N_11697);
nand U11961 (N_11961,N_11747,N_11631);
nor U11962 (N_11962,N_11677,N_11648);
nor U11963 (N_11963,N_11607,N_11672);
and U11964 (N_11964,N_11660,N_11686);
and U11965 (N_11965,N_11665,N_11500);
nand U11966 (N_11966,N_11558,N_11695);
xor U11967 (N_11967,N_11608,N_11577);
xor U11968 (N_11968,N_11502,N_11598);
and U11969 (N_11969,N_11616,N_11706);
xor U11970 (N_11970,N_11581,N_11717);
xor U11971 (N_11971,N_11665,N_11690);
and U11972 (N_11972,N_11662,N_11575);
and U11973 (N_11973,N_11698,N_11538);
and U11974 (N_11974,N_11559,N_11580);
or U11975 (N_11975,N_11704,N_11640);
nor U11976 (N_11976,N_11691,N_11564);
nor U11977 (N_11977,N_11646,N_11584);
and U11978 (N_11978,N_11727,N_11649);
or U11979 (N_11979,N_11658,N_11682);
or U11980 (N_11980,N_11578,N_11540);
nor U11981 (N_11981,N_11749,N_11552);
xnor U11982 (N_11982,N_11531,N_11691);
nand U11983 (N_11983,N_11720,N_11596);
nor U11984 (N_11984,N_11619,N_11667);
nor U11985 (N_11985,N_11673,N_11520);
xnor U11986 (N_11986,N_11515,N_11663);
xnor U11987 (N_11987,N_11667,N_11618);
nand U11988 (N_11988,N_11638,N_11665);
nor U11989 (N_11989,N_11747,N_11546);
or U11990 (N_11990,N_11707,N_11636);
nand U11991 (N_11991,N_11666,N_11713);
and U11992 (N_11992,N_11508,N_11638);
nor U11993 (N_11993,N_11608,N_11689);
or U11994 (N_11994,N_11688,N_11637);
xnor U11995 (N_11995,N_11693,N_11701);
and U11996 (N_11996,N_11616,N_11660);
nand U11997 (N_11997,N_11554,N_11691);
or U11998 (N_11998,N_11634,N_11648);
nand U11999 (N_11999,N_11508,N_11533);
or U12000 (N_12000,N_11941,N_11880);
and U12001 (N_12001,N_11799,N_11981);
nand U12002 (N_12002,N_11842,N_11985);
nand U12003 (N_12003,N_11840,N_11751);
or U12004 (N_12004,N_11939,N_11844);
or U12005 (N_12005,N_11806,N_11934);
and U12006 (N_12006,N_11925,N_11963);
nor U12007 (N_12007,N_11801,N_11750);
nand U12008 (N_12008,N_11815,N_11976);
nor U12009 (N_12009,N_11940,N_11950);
xnor U12010 (N_12010,N_11933,N_11878);
nor U12011 (N_12011,N_11891,N_11920);
or U12012 (N_12012,N_11886,N_11958);
xnor U12013 (N_12013,N_11970,N_11856);
xnor U12014 (N_12014,N_11947,N_11851);
nor U12015 (N_12015,N_11854,N_11987);
nand U12016 (N_12016,N_11811,N_11752);
nor U12017 (N_12017,N_11902,N_11757);
nor U12018 (N_12018,N_11841,N_11991);
nand U12019 (N_12019,N_11767,N_11901);
nor U12020 (N_12020,N_11848,N_11897);
nand U12021 (N_12021,N_11870,N_11833);
and U12022 (N_12022,N_11805,N_11969);
nand U12023 (N_12023,N_11988,N_11974);
nand U12024 (N_12024,N_11753,N_11913);
nor U12025 (N_12025,N_11930,N_11966);
or U12026 (N_12026,N_11849,N_11781);
or U12027 (N_12027,N_11834,N_11879);
nand U12028 (N_12028,N_11760,N_11826);
or U12029 (N_12029,N_11807,N_11926);
or U12030 (N_12030,N_11876,N_11894);
nand U12031 (N_12031,N_11911,N_11997);
or U12032 (N_12032,N_11973,N_11838);
nor U12033 (N_12033,N_11924,N_11756);
nand U12034 (N_12034,N_11775,N_11980);
and U12035 (N_12035,N_11899,N_11915);
nor U12036 (N_12036,N_11783,N_11818);
nand U12037 (N_12037,N_11758,N_11754);
and U12038 (N_12038,N_11786,N_11763);
xnor U12039 (N_12039,N_11782,N_11852);
xnor U12040 (N_12040,N_11889,N_11813);
nand U12041 (N_12041,N_11916,N_11983);
nor U12042 (N_12042,N_11762,N_11964);
and U12043 (N_12043,N_11793,N_11855);
xnor U12044 (N_12044,N_11797,N_11817);
or U12045 (N_12045,N_11798,N_11977);
xor U12046 (N_12046,N_11837,N_11955);
xor U12047 (N_12047,N_11984,N_11904);
nor U12048 (N_12048,N_11875,N_11839);
nand U12049 (N_12049,N_11772,N_11954);
xnor U12050 (N_12050,N_11895,N_11887);
or U12051 (N_12051,N_11867,N_11907);
and U12052 (N_12052,N_11770,N_11943);
xor U12053 (N_12053,N_11912,N_11814);
and U12054 (N_12054,N_11975,N_11996);
nor U12055 (N_12055,N_11932,N_11951);
or U12056 (N_12056,N_11865,N_11860);
xnor U12057 (N_12057,N_11909,N_11810);
nor U12058 (N_12058,N_11905,N_11803);
xnor U12059 (N_12059,N_11847,N_11900);
nor U12060 (N_12060,N_11968,N_11960);
or U12061 (N_12061,N_11885,N_11931);
or U12062 (N_12062,N_11825,N_11824);
xor U12063 (N_12063,N_11993,N_11859);
xor U12064 (N_12064,N_11937,N_11771);
xnor U12065 (N_12065,N_11881,N_11888);
nand U12066 (N_12066,N_11890,N_11938);
nor U12067 (N_12067,N_11828,N_11942);
nor U12068 (N_12068,N_11967,N_11787);
xnor U12069 (N_12069,N_11928,N_11918);
and U12070 (N_12070,N_11866,N_11784);
xor U12071 (N_12071,N_11795,N_11831);
nand U12072 (N_12072,N_11830,N_11789);
nand U12073 (N_12073,N_11884,N_11995);
xor U12074 (N_12074,N_11906,N_11769);
xnor U12075 (N_12075,N_11800,N_11998);
nor U12076 (N_12076,N_11919,N_11858);
nor U12077 (N_12077,N_11823,N_11898);
nor U12078 (N_12078,N_11883,N_11764);
nor U12079 (N_12079,N_11990,N_11761);
xnor U12080 (N_12080,N_11843,N_11863);
nor U12081 (N_12081,N_11896,N_11779);
nor U12082 (N_12082,N_11809,N_11873);
nor U12083 (N_12083,N_11829,N_11804);
nand U12084 (N_12084,N_11796,N_11978);
or U12085 (N_12085,N_11945,N_11949);
nor U12086 (N_12086,N_11872,N_11908);
xor U12087 (N_12087,N_11965,N_11929);
nand U12088 (N_12088,N_11808,N_11759);
and U12089 (N_12089,N_11982,N_11952);
nand U12090 (N_12090,N_11862,N_11816);
nor U12091 (N_12091,N_11836,N_11790);
nor U12092 (N_12092,N_11874,N_11944);
and U12093 (N_12093,N_11845,N_11868);
nand U12094 (N_12094,N_11877,N_11893);
and U12095 (N_12095,N_11802,N_11927);
and U12096 (N_12096,N_11794,N_11882);
nor U12097 (N_12097,N_11853,N_11957);
nor U12098 (N_12098,N_11979,N_11791);
and U12099 (N_12099,N_11785,N_11936);
or U12100 (N_12100,N_11864,N_11972);
or U12101 (N_12101,N_11755,N_11788);
and U12102 (N_12102,N_11821,N_11910);
nand U12103 (N_12103,N_11792,N_11959);
xor U12104 (N_12104,N_11871,N_11846);
nor U12105 (N_12105,N_11953,N_11903);
nor U12106 (N_12106,N_11948,N_11780);
or U12107 (N_12107,N_11922,N_11819);
or U12108 (N_12108,N_11776,N_11914);
nand U12109 (N_12109,N_11777,N_11861);
nand U12110 (N_12110,N_11835,N_11989);
nand U12111 (N_12111,N_11961,N_11857);
and U12112 (N_12112,N_11935,N_11869);
xor U12113 (N_12113,N_11820,N_11923);
and U12114 (N_12114,N_11765,N_11768);
nand U12115 (N_12115,N_11994,N_11827);
and U12116 (N_12116,N_11992,N_11892);
and U12117 (N_12117,N_11986,N_11999);
xnor U12118 (N_12118,N_11773,N_11774);
xnor U12119 (N_12119,N_11778,N_11850);
and U12120 (N_12120,N_11822,N_11946);
and U12121 (N_12121,N_11962,N_11971);
nor U12122 (N_12122,N_11832,N_11956);
xor U12123 (N_12123,N_11766,N_11917);
nand U12124 (N_12124,N_11921,N_11812);
and U12125 (N_12125,N_11756,N_11935);
nor U12126 (N_12126,N_11925,N_11820);
nor U12127 (N_12127,N_11828,N_11950);
and U12128 (N_12128,N_11910,N_11993);
or U12129 (N_12129,N_11967,N_11821);
xnor U12130 (N_12130,N_11951,N_11778);
and U12131 (N_12131,N_11880,N_11863);
and U12132 (N_12132,N_11945,N_11786);
xor U12133 (N_12133,N_11931,N_11902);
and U12134 (N_12134,N_11805,N_11912);
or U12135 (N_12135,N_11957,N_11868);
nor U12136 (N_12136,N_11928,N_11804);
nand U12137 (N_12137,N_11837,N_11957);
and U12138 (N_12138,N_11900,N_11933);
and U12139 (N_12139,N_11807,N_11826);
nand U12140 (N_12140,N_11794,N_11819);
nor U12141 (N_12141,N_11834,N_11829);
nand U12142 (N_12142,N_11985,N_11892);
or U12143 (N_12143,N_11773,N_11978);
xor U12144 (N_12144,N_11814,N_11832);
nor U12145 (N_12145,N_11982,N_11942);
nor U12146 (N_12146,N_11895,N_11964);
nor U12147 (N_12147,N_11865,N_11936);
nor U12148 (N_12148,N_11830,N_11907);
or U12149 (N_12149,N_11932,N_11953);
or U12150 (N_12150,N_11824,N_11833);
and U12151 (N_12151,N_11767,N_11945);
and U12152 (N_12152,N_11873,N_11786);
or U12153 (N_12153,N_11984,N_11828);
nand U12154 (N_12154,N_11980,N_11861);
xnor U12155 (N_12155,N_11844,N_11914);
nand U12156 (N_12156,N_11914,N_11796);
or U12157 (N_12157,N_11761,N_11904);
xnor U12158 (N_12158,N_11783,N_11899);
and U12159 (N_12159,N_11980,N_11766);
xnor U12160 (N_12160,N_11762,N_11882);
or U12161 (N_12161,N_11823,N_11870);
xnor U12162 (N_12162,N_11878,N_11905);
xor U12163 (N_12163,N_11970,N_11822);
and U12164 (N_12164,N_11968,N_11827);
and U12165 (N_12165,N_11845,N_11797);
or U12166 (N_12166,N_11820,N_11971);
nand U12167 (N_12167,N_11941,N_11758);
xor U12168 (N_12168,N_11838,N_11814);
xor U12169 (N_12169,N_11954,N_11771);
and U12170 (N_12170,N_11993,N_11863);
nor U12171 (N_12171,N_11909,N_11890);
or U12172 (N_12172,N_11928,N_11945);
nor U12173 (N_12173,N_11860,N_11763);
nor U12174 (N_12174,N_11975,N_11943);
nand U12175 (N_12175,N_11881,N_11905);
and U12176 (N_12176,N_11888,N_11872);
nand U12177 (N_12177,N_11779,N_11841);
or U12178 (N_12178,N_11970,N_11755);
nor U12179 (N_12179,N_11807,N_11828);
nor U12180 (N_12180,N_11928,N_11911);
xnor U12181 (N_12181,N_11905,N_11956);
nor U12182 (N_12182,N_11946,N_11783);
or U12183 (N_12183,N_11980,N_11801);
or U12184 (N_12184,N_11818,N_11892);
xor U12185 (N_12185,N_11974,N_11920);
xnor U12186 (N_12186,N_11845,N_11863);
nor U12187 (N_12187,N_11761,N_11824);
nor U12188 (N_12188,N_11918,N_11779);
xnor U12189 (N_12189,N_11877,N_11836);
xor U12190 (N_12190,N_11762,N_11758);
nor U12191 (N_12191,N_11856,N_11911);
nand U12192 (N_12192,N_11788,N_11770);
nor U12193 (N_12193,N_11791,N_11893);
nor U12194 (N_12194,N_11911,N_11763);
nor U12195 (N_12195,N_11815,N_11937);
nor U12196 (N_12196,N_11804,N_11883);
nand U12197 (N_12197,N_11938,N_11931);
nand U12198 (N_12198,N_11892,N_11829);
nor U12199 (N_12199,N_11752,N_11767);
or U12200 (N_12200,N_11915,N_11862);
xnor U12201 (N_12201,N_11920,N_11904);
xor U12202 (N_12202,N_11887,N_11778);
nor U12203 (N_12203,N_11986,N_11805);
xor U12204 (N_12204,N_11766,N_11758);
nor U12205 (N_12205,N_11995,N_11896);
xnor U12206 (N_12206,N_11933,N_11771);
nor U12207 (N_12207,N_11854,N_11828);
nand U12208 (N_12208,N_11831,N_11889);
or U12209 (N_12209,N_11792,N_11828);
nor U12210 (N_12210,N_11934,N_11989);
nor U12211 (N_12211,N_11907,N_11858);
nor U12212 (N_12212,N_11852,N_11769);
nand U12213 (N_12213,N_11763,N_11875);
or U12214 (N_12214,N_11939,N_11976);
nand U12215 (N_12215,N_11883,N_11867);
xor U12216 (N_12216,N_11800,N_11889);
nand U12217 (N_12217,N_11874,N_11792);
xor U12218 (N_12218,N_11933,N_11853);
nor U12219 (N_12219,N_11935,N_11937);
nor U12220 (N_12220,N_11980,N_11925);
nand U12221 (N_12221,N_11893,N_11940);
nand U12222 (N_12222,N_11825,N_11795);
nand U12223 (N_12223,N_11783,N_11924);
and U12224 (N_12224,N_11971,N_11783);
and U12225 (N_12225,N_11838,N_11972);
nand U12226 (N_12226,N_11879,N_11904);
and U12227 (N_12227,N_11969,N_11917);
and U12228 (N_12228,N_11871,N_11955);
or U12229 (N_12229,N_11806,N_11836);
xor U12230 (N_12230,N_11806,N_11880);
nand U12231 (N_12231,N_11886,N_11836);
and U12232 (N_12232,N_11822,N_11987);
or U12233 (N_12233,N_11907,N_11811);
and U12234 (N_12234,N_11860,N_11786);
or U12235 (N_12235,N_11805,N_11860);
and U12236 (N_12236,N_11942,N_11875);
nand U12237 (N_12237,N_11777,N_11909);
and U12238 (N_12238,N_11800,N_11881);
or U12239 (N_12239,N_11903,N_11873);
or U12240 (N_12240,N_11799,N_11894);
nor U12241 (N_12241,N_11999,N_11979);
nor U12242 (N_12242,N_11754,N_11952);
or U12243 (N_12243,N_11881,N_11868);
and U12244 (N_12244,N_11922,N_11800);
and U12245 (N_12245,N_11965,N_11857);
xor U12246 (N_12246,N_11886,N_11755);
or U12247 (N_12247,N_11788,N_11913);
nor U12248 (N_12248,N_11966,N_11816);
nor U12249 (N_12249,N_11897,N_11822);
nor U12250 (N_12250,N_12082,N_12035);
or U12251 (N_12251,N_12216,N_12225);
and U12252 (N_12252,N_12073,N_12143);
or U12253 (N_12253,N_12162,N_12196);
and U12254 (N_12254,N_12034,N_12069);
xor U12255 (N_12255,N_12207,N_12235);
xnor U12256 (N_12256,N_12201,N_12057);
and U12257 (N_12257,N_12134,N_12240);
and U12258 (N_12258,N_12155,N_12222);
and U12259 (N_12259,N_12019,N_12077);
and U12260 (N_12260,N_12211,N_12189);
nand U12261 (N_12261,N_12132,N_12109);
and U12262 (N_12262,N_12098,N_12040);
nor U12263 (N_12263,N_12179,N_12228);
xor U12264 (N_12264,N_12099,N_12024);
or U12265 (N_12265,N_12011,N_12091);
and U12266 (N_12266,N_12059,N_12202);
nor U12267 (N_12267,N_12242,N_12088);
xnor U12268 (N_12268,N_12171,N_12147);
nor U12269 (N_12269,N_12145,N_12041);
xor U12270 (N_12270,N_12137,N_12039);
xnor U12271 (N_12271,N_12043,N_12022);
nand U12272 (N_12272,N_12151,N_12053);
nand U12273 (N_12273,N_12241,N_12046);
nand U12274 (N_12274,N_12094,N_12093);
or U12275 (N_12275,N_12101,N_12133);
nand U12276 (N_12276,N_12020,N_12018);
xnor U12277 (N_12277,N_12186,N_12025);
or U12278 (N_12278,N_12033,N_12215);
and U12279 (N_12279,N_12183,N_12135);
or U12280 (N_12280,N_12173,N_12191);
and U12281 (N_12281,N_12006,N_12097);
nor U12282 (N_12282,N_12014,N_12037);
nor U12283 (N_12283,N_12070,N_12227);
and U12284 (N_12284,N_12122,N_12166);
xnor U12285 (N_12285,N_12214,N_12128);
or U12286 (N_12286,N_12075,N_12004);
nor U12287 (N_12287,N_12198,N_12238);
xnor U12288 (N_12288,N_12218,N_12068);
xor U12289 (N_12289,N_12000,N_12009);
or U12290 (N_12290,N_12148,N_12178);
nand U12291 (N_12291,N_12114,N_12078);
nor U12292 (N_12292,N_12095,N_12153);
nand U12293 (N_12293,N_12203,N_12003);
xnor U12294 (N_12294,N_12029,N_12038);
and U12295 (N_12295,N_12236,N_12175);
nand U12296 (N_12296,N_12209,N_12237);
nor U12297 (N_12297,N_12158,N_12194);
nand U12298 (N_12298,N_12146,N_12027);
and U12299 (N_12299,N_12219,N_12013);
or U12300 (N_12300,N_12234,N_12050);
nor U12301 (N_12301,N_12061,N_12233);
or U12302 (N_12302,N_12051,N_12052);
nor U12303 (N_12303,N_12049,N_12100);
or U12304 (N_12304,N_12089,N_12054);
or U12305 (N_12305,N_12205,N_12048);
xnor U12306 (N_12306,N_12200,N_12032);
xnor U12307 (N_12307,N_12181,N_12017);
nor U12308 (N_12308,N_12249,N_12079);
and U12309 (N_12309,N_12152,N_12110);
nor U12310 (N_12310,N_12087,N_12223);
xnor U12311 (N_12311,N_12138,N_12107);
nor U12312 (N_12312,N_12012,N_12174);
nor U12313 (N_12313,N_12026,N_12168);
nand U12314 (N_12314,N_12023,N_12065);
nor U12315 (N_12315,N_12170,N_12131);
nand U12316 (N_12316,N_12090,N_12117);
or U12317 (N_12317,N_12144,N_12184);
xnor U12318 (N_12318,N_12142,N_12103);
xnor U12319 (N_12319,N_12112,N_12185);
nor U12320 (N_12320,N_12229,N_12149);
or U12321 (N_12321,N_12115,N_12028);
nand U12322 (N_12322,N_12047,N_12129);
nor U12323 (N_12323,N_12120,N_12244);
nor U12324 (N_12324,N_12096,N_12002);
or U12325 (N_12325,N_12139,N_12164);
nor U12326 (N_12326,N_12126,N_12212);
and U12327 (N_12327,N_12187,N_12169);
xor U12328 (N_12328,N_12001,N_12167);
nand U12329 (N_12329,N_12010,N_12058);
nand U12330 (N_12330,N_12230,N_12072);
and U12331 (N_12331,N_12016,N_12124);
or U12332 (N_12332,N_12177,N_12176);
xnor U12333 (N_12333,N_12042,N_12182);
xnor U12334 (N_12334,N_12030,N_12193);
nor U12335 (N_12335,N_12118,N_12157);
or U12336 (N_12336,N_12005,N_12031);
and U12337 (N_12337,N_12188,N_12141);
nand U12338 (N_12338,N_12159,N_12081);
and U12339 (N_12339,N_12217,N_12080);
xor U12340 (N_12340,N_12245,N_12106);
nand U12341 (N_12341,N_12232,N_12130);
nor U12342 (N_12342,N_12021,N_12192);
and U12343 (N_12343,N_12161,N_12045);
or U12344 (N_12344,N_12111,N_12008);
or U12345 (N_12345,N_12204,N_12160);
or U12346 (N_12346,N_12062,N_12190);
or U12347 (N_12347,N_12246,N_12197);
nand U12348 (N_12348,N_12067,N_12066);
and U12349 (N_12349,N_12056,N_12116);
and U12350 (N_12350,N_12156,N_12210);
or U12351 (N_12351,N_12199,N_12221);
or U12352 (N_12352,N_12123,N_12108);
xnor U12353 (N_12353,N_12247,N_12074);
or U12354 (N_12354,N_12076,N_12136);
xor U12355 (N_12355,N_12113,N_12195);
or U12356 (N_12356,N_12083,N_12150);
nand U12357 (N_12357,N_12044,N_12243);
nand U12358 (N_12358,N_12248,N_12121);
nand U12359 (N_12359,N_12085,N_12206);
xnor U12360 (N_12360,N_12154,N_12226);
nand U12361 (N_12361,N_12208,N_12060);
or U12362 (N_12362,N_12036,N_12119);
and U12363 (N_12363,N_12127,N_12172);
nand U12364 (N_12364,N_12007,N_12140);
nand U12365 (N_12365,N_12084,N_12105);
nand U12366 (N_12366,N_12071,N_12092);
nor U12367 (N_12367,N_12213,N_12220);
xor U12368 (N_12368,N_12055,N_12102);
xor U12369 (N_12369,N_12163,N_12165);
nand U12370 (N_12370,N_12104,N_12224);
nand U12371 (N_12371,N_12015,N_12063);
nand U12372 (N_12372,N_12064,N_12086);
and U12373 (N_12373,N_12125,N_12239);
nand U12374 (N_12374,N_12180,N_12231);
xnor U12375 (N_12375,N_12007,N_12109);
nor U12376 (N_12376,N_12181,N_12111);
and U12377 (N_12377,N_12237,N_12163);
xor U12378 (N_12378,N_12104,N_12119);
and U12379 (N_12379,N_12204,N_12216);
and U12380 (N_12380,N_12026,N_12196);
and U12381 (N_12381,N_12035,N_12210);
nor U12382 (N_12382,N_12120,N_12086);
and U12383 (N_12383,N_12060,N_12140);
xor U12384 (N_12384,N_12090,N_12190);
nand U12385 (N_12385,N_12034,N_12087);
xnor U12386 (N_12386,N_12197,N_12104);
xnor U12387 (N_12387,N_12016,N_12073);
or U12388 (N_12388,N_12143,N_12047);
xnor U12389 (N_12389,N_12223,N_12165);
nand U12390 (N_12390,N_12227,N_12222);
nand U12391 (N_12391,N_12210,N_12183);
or U12392 (N_12392,N_12014,N_12052);
or U12393 (N_12393,N_12199,N_12071);
xor U12394 (N_12394,N_12175,N_12140);
and U12395 (N_12395,N_12170,N_12068);
xnor U12396 (N_12396,N_12178,N_12137);
or U12397 (N_12397,N_12243,N_12157);
and U12398 (N_12398,N_12023,N_12163);
nand U12399 (N_12399,N_12176,N_12126);
nor U12400 (N_12400,N_12208,N_12148);
xnor U12401 (N_12401,N_12022,N_12082);
xor U12402 (N_12402,N_12190,N_12113);
xnor U12403 (N_12403,N_12137,N_12082);
or U12404 (N_12404,N_12061,N_12249);
or U12405 (N_12405,N_12141,N_12128);
or U12406 (N_12406,N_12122,N_12062);
xnor U12407 (N_12407,N_12169,N_12214);
xor U12408 (N_12408,N_12050,N_12091);
and U12409 (N_12409,N_12030,N_12104);
nand U12410 (N_12410,N_12131,N_12243);
xor U12411 (N_12411,N_12135,N_12004);
xnor U12412 (N_12412,N_12039,N_12145);
nand U12413 (N_12413,N_12039,N_12187);
or U12414 (N_12414,N_12097,N_12119);
nand U12415 (N_12415,N_12247,N_12136);
xor U12416 (N_12416,N_12054,N_12120);
xor U12417 (N_12417,N_12079,N_12142);
xor U12418 (N_12418,N_12125,N_12238);
or U12419 (N_12419,N_12023,N_12155);
xnor U12420 (N_12420,N_12038,N_12115);
nor U12421 (N_12421,N_12203,N_12048);
xnor U12422 (N_12422,N_12098,N_12079);
nand U12423 (N_12423,N_12171,N_12194);
nand U12424 (N_12424,N_12002,N_12123);
or U12425 (N_12425,N_12158,N_12131);
or U12426 (N_12426,N_12234,N_12113);
and U12427 (N_12427,N_12114,N_12229);
or U12428 (N_12428,N_12184,N_12215);
and U12429 (N_12429,N_12112,N_12105);
xnor U12430 (N_12430,N_12233,N_12160);
or U12431 (N_12431,N_12008,N_12234);
and U12432 (N_12432,N_12218,N_12089);
and U12433 (N_12433,N_12110,N_12224);
xnor U12434 (N_12434,N_12227,N_12061);
nand U12435 (N_12435,N_12079,N_12202);
or U12436 (N_12436,N_12130,N_12131);
xnor U12437 (N_12437,N_12057,N_12077);
xnor U12438 (N_12438,N_12025,N_12205);
nand U12439 (N_12439,N_12053,N_12224);
and U12440 (N_12440,N_12184,N_12175);
nand U12441 (N_12441,N_12160,N_12031);
and U12442 (N_12442,N_12235,N_12154);
xnor U12443 (N_12443,N_12244,N_12208);
nor U12444 (N_12444,N_12154,N_12072);
nand U12445 (N_12445,N_12046,N_12130);
or U12446 (N_12446,N_12100,N_12065);
xnor U12447 (N_12447,N_12171,N_12107);
xnor U12448 (N_12448,N_12185,N_12139);
or U12449 (N_12449,N_12091,N_12016);
nor U12450 (N_12450,N_12086,N_12167);
or U12451 (N_12451,N_12066,N_12038);
nor U12452 (N_12452,N_12194,N_12232);
and U12453 (N_12453,N_12138,N_12195);
and U12454 (N_12454,N_12008,N_12086);
nor U12455 (N_12455,N_12058,N_12113);
xor U12456 (N_12456,N_12208,N_12091);
xnor U12457 (N_12457,N_12085,N_12150);
or U12458 (N_12458,N_12118,N_12082);
nor U12459 (N_12459,N_12219,N_12182);
nor U12460 (N_12460,N_12236,N_12243);
xor U12461 (N_12461,N_12048,N_12248);
and U12462 (N_12462,N_12217,N_12043);
or U12463 (N_12463,N_12060,N_12172);
nor U12464 (N_12464,N_12177,N_12226);
xor U12465 (N_12465,N_12028,N_12094);
or U12466 (N_12466,N_12186,N_12013);
nand U12467 (N_12467,N_12218,N_12232);
or U12468 (N_12468,N_12102,N_12146);
nand U12469 (N_12469,N_12212,N_12172);
or U12470 (N_12470,N_12026,N_12030);
or U12471 (N_12471,N_12061,N_12012);
nand U12472 (N_12472,N_12003,N_12081);
nor U12473 (N_12473,N_12145,N_12192);
nand U12474 (N_12474,N_12182,N_12132);
nand U12475 (N_12475,N_12192,N_12089);
xor U12476 (N_12476,N_12082,N_12181);
nand U12477 (N_12477,N_12206,N_12029);
or U12478 (N_12478,N_12013,N_12131);
and U12479 (N_12479,N_12030,N_12220);
xor U12480 (N_12480,N_12123,N_12195);
nand U12481 (N_12481,N_12137,N_12217);
nand U12482 (N_12482,N_12046,N_12106);
or U12483 (N_12483,N_12075,N_12148);
or U12484 (N_12484,N_12081,N_12036);
xnor U12485 (N_12485,N_12064,N_12184);
nand U12486 (N_12486,N_12249,N_12038);
nand U12487 (N_12487,N_12186,N_12135);
or U12488 (N_12488,N_12241,N_12063);
nand U12489 (N_12489,N_12196,N_12080);
nand U12490 (N_12490,N_12199,N_12107);
nor U12491 (N_12491,N_12102,N_12243);
xor U12492 (N_12492,N_12115,N_12079);
nor U12493 (N_12493,N_12137,N_12165);
xnor U12494 (N_12494,N_12132,N_12038);
nand U12495 (N_12495,N_12022,N_12196);
and U12496 (N_12496,N_12201,N_12073);
nor U12497 (N_12497,N_12077,N_12106);
and U12498 (N_12498,N_12114,N_12028);
or U12499 (N_12499,N_12212,N_12229);
nand U12500 (N_12500,N_12268,N_12342);
and U12501 (N_12501,N_12396,N_12479);
or U12502 (N_12502,N_12443,N_12339);
nand U12503 (N_12503,N_12420,N_12252);
and U12504 (N_12504,N_12429,N_12474);
nand U12505 (N_12505,N_12343,N_12300);
nand U12506 (N_12506,N_12451,N_12325);
nand U12507 (N_12507,N_12489,N_12494);
and U12508 (N_12508,N_12311,N_12280);
xor U12509 (N_12509,N_12402,N_12266);
xnor U12510 (N_12510,N_12362,N_12336);
nor U12511 (N_12511,N_12285,N_12434);
nor U12512 (N_12512,N_12265,N_12351);
nand U12513 (N_12513,N_12259,N_12347);
nor U12514 (N_12514,N_12377,N_12477);
and U12515 (N_12515,N_12297,N_12334);
nor U12516 (N_12516,N_12427,N_12462);
and U12517 (N_12517,N_12312,N_12296);
xor U12518 (N_12518,N_12263,N_12290);
and U12519 (N_12519,N_12452,N_12492);
nor U12520 (N_12520,N_12475,N_12305);
nand U12521 (N_12521,N_12272,N_12408);
xnor U12522 (N_12522,N_12433,N_12391);
xnor U12523 (N_12523,N_12275,N_12364);
nor U12524 (N_12524,N_12359,N_12431);
and U12525 (N_12525,N_12306,N_12409);
xnor U12526 (N_12526,N_12289,N_12395);
nand U12527 (N_12527,N_12470,N_12419);
xnor U12528 (N_12528,N_12307,N_12301);
nand U12529 (N_12529,N_12484,N_12276);
or U12530 (N_12530,N_12495,N_12374);
or U12531 (N_12531,N_12369,N_12398);
nand U12532 (N_12532,N_12328,N_12264);
nor U12533 (N_12533,N_12424,N_12482);
xnor U12534 (N_12534,N_12304,N_12318);
nor U12535 (N_12535,N_12386,N_12426);
xor U12536 (N_12536,N_12279,N_12379);
xnor U12537 (N_12537,N_12271,N_12250);
xnor U12538 (N_12538,N_12321,N_12308);
nor U12539 (N_12539,N_12381,N_12358);
xnor U12540 (N_12540,N_12410,N_12341);
or U12541 (N_12541,N_12442,N_12473);
xnor U12542 (N_12542,N_12335,N_12380);
nor U12543 (N_12543,N_12357,N_12338);
nor U12544 (N_12544,N_12422,N_12363);
or U12545 (N_12545,N_12367,N_12417);
and U12546 (N_12546,N_12303,N_12487);
nand U12547 (N_12547,N_12385,N_12388);
and U12548 (N_12548,N_12444,N_12485);
xnor U12549 (N_12549,N_12319,N_12387);
nand U12550 (N_12550,N_12413,N_12498);
nor U12551 (N_12551,N_12293,N_12428);
nor U12552 (N_12552,N_12288,N_12486);
and U12553 (N_12553,N_12267,N_12382);
or U12554 (N_12554,N_12361,N_12394);
nor U12555 (N_12555,N_12436,N_12281);
nand U12556 (N_12556,N_12283,N_12468);
xnor U12557 (N_12557,N_12414,N_12471);
xnor U12558 (N_12558,N_12375,N_12399);
and U12559 (N_12559,N_12320,N_12491);
nor U12560 (N_12560,N_12469,N_12286);
xnor U12561 (N_12561,N_12333,N_12432);
and U12562 (N_12562,N_12340,N_12449);
nand U12563 (N_12563,N_12316,N_12284);
xnor U12564 (N_12564,N_12454,N_12464);
or U12565 (N_12565,N_12353,N_12365);
or U12566 (N_12566,N_12423,N_12314);
nand U12567 (N_12567,N_12329,N_12287);
xnor U12568 (N_12568,N_12448,N_12256);
nand U12569 (N_12569,N_12425,N_12261);
and U12570 (N_12570,N_12371,N_12488);
or U12571 (N_12571,N_12463,N_12456);
nor U12572 (N_12572,N_12352,N_12404);
nor U12573 (N_12573,N_12258,N_12348);
or U12574 (N_12574,N_12274,N_12481);
nor U12575 (N_12575,N_12439,N_12445);
nor U12576 (N_12576,N_12373,N_12277);
or U12577 (N_12577,N_12360,N_12397);
xnor U12578 (N_12578,N_12400,N_12356);
nor U12579 (N_12579,N_12326,N_12383);
or U12580 (N_12580,N_12384,N_12295);
xnor U12581 (N_12581,N_12490,N_12302);
nand U12582 (N_12582,N_12415,N_12337);
nor U12583 (N_12583,N_12298,N_12330);
nor U12584 (N_12584,N_12313,N_12260);
or U12585 (N_12585,N_12331,N_12344);
nand U12586 (N_12586,N_12376,N_12472);
nand U12587 (N_12587,N_12401,N_12406);
nor U12588 (N_12588,N_12255,N_12346);
nand U12589 (N_12589,N_12253,N_12478);
nor U12590 (N_12590,N_12291,N_12476);
or U12591 (N_12591,N_12269,N_12412);
xor U12592 (N_12592,N_12349,N_12350);
or U12593 (N_12593,N_12372,N_12262);
and U12594 (N_12594,N_12254,N_12332);
and U12595 (N_12595,N_12446,N_12460);
xor U12596 (N_12596,N_12389,N_12309);
xor U12597 (N_12597,N_12458,N_12496);
nand U12598 (N_12598,N_12497,N_12323);
nand U12599 (N_12599,N_12317,N_12392);
xor U12600 (N_12600,N_12294,N_12273);
nor U12601 (N_12601,N_12324,N_12459);
xor U12602 (N_12602,N_12270,N_12453);
xor U12603 (N_12603,N_12430,N_12345);
nor U12604 (N_12604,N_12299,N_12390);
xor U12605 (N_12605,N_12315,N_12407);
or U12606 (N_12606,N_12292,N_12354);
xor U12607 (N_12607,N_12405,N_12322);
and U12608 (N_12608,N_12282,N_12447);
nand U12609 (N_12609,N_12368,N_12355);
or U12610 (N_12610,N_12440,N_12378);
or U12611 (N_12611,N_12437,N_12327);
nor U12612 (N_12612,N_12421,N_12251);
nor U12613 (N_12613,N_12310,N_12416);
nand U12614 (N_12614,N_12499,N_12403);
and U12615 (N_12615,N_12366,N_12450);
nor U12616 (N_12616,N_12441,N_12438);
or U12617 (N_12617,N_12493,N_12370);
nand U12618 (N_12618,N_12467,N_12435);
or U12619 (N_12619,N_12457,N_12411);
nand U12620 (N_12620,N_12466,N_12393);
and U12621 (N_12621,N_12461,N_12480);
nand U12622 (N_12622,N_12465,N_12483);
xor U12623 (N_12623,N_12278,N_12455);
nor U12624 (N_12624,N_12418,N_12257);
nor U12625 (N_12625,N_12336,N_12250);
and U12626 (N_12626,N_12487,N_12423);
and U12627 (N_12627,N_12441,N_12403);
and U12628 (N_12628,N_12293,N_12254);
and U12629 (N_12629,N_12326,N_12380);
nor U12630 (N_12630,N_12432,N_12281);
nand U12631 (N_12631,N_12449,N_12330);
nor U12632 (N_12632,N_12318,N_12295);
or U12633 (N_12633,N_12390,N_12378);
nand U12634 (N_12634,N_12284,N_12330);
or U12635 (N_12635,N_12392,N_12451);
nand U12636 (N_12636,N_12455,N_12491);
or U12637 (N_12637,N_12363,N_12448);
and U12638 (N_12638,N_12365,N_12482);
nor U12639 (N_12639,N_12432,N_12334);
and U12640 (N_12640,N_12267,N_12358);
or U12641 (N_12641,N_12280,N_12493);
or U12642 (N_12642,N_12361,N_12281);
and U12643 (N_12643,N_12352,N_12264);
and U12644 (N_12644,N_12440,N_12439);
nor U12645 (N_12645,N_12279,N_12323);
xnor U12646 (N_12646,N_12370,N_12286);
and U12647 (N_12647,N_12266,N_12483);
nand U12648 (N_12648,N_12292,N_12443);
or U12649 (N_12649,N_12295,N_12274);
xnor U12650 (N_12650,N_12417,N_12389);
xor U12651 (N_12651,N_12258,N_12302);
or U12652 (N_12652,N_12405,N_12323);
nor U12653 (N_12653,N_12327,N_12403);
or U12654 (N_12654,N_12423,N_12307);
and U12655 (N_12655,N_12276,N_12426);
or U12656 (N_12656,N_12353,N_12412);
nor U12657 (N_12657,N_12301,N_12324);
xnor U12658 (N_12658,N_12326,N_12335);
nand U12659 (N_12659,N_12413,N_12390);
nand U12660 (N_12660,N_12412,N_12436);
nor U12661 (N_12661,N_12487,N_12427);
and U12662 (N_12662,N_12363,N_12486);
nand U12663 (N_12663,N_12332,N_12458);
or U12664 (N_12664,N_12411,N_12357);
nor U12665 (N_12665,N_12445,N_12327);
nor U12666 (N_12666,N_12363,N_12444);
nand U12667 (N_12667,N_12265,N_12403);
or U12668 (N_12668,N_12478,N_12372);
xnor U12669 (N_12669,N_12351,N_12266);
and U12670 (N_12670,N_12311,N_12326);
nand U12671 (N_12671,N_12336,N_12288);
nor U12672 (N_12672,N_12257,N_12407);
nor U12673 (N_12673,N_12404,N_12496);
xor U12674 (N_12674,N_12386,N_12272);
xor U12675 (N_12675,N_12490,N_12334);
xnor U12676 (N_12676,N_12291,N_12414);
nand U12677 (N_12677,N_12281,N_12369);
and U12678 (N_12678,N_12382,N_12377);
or U12679 (N_12679,N_12378,N_12493);
or U12680 (N_12680,N_12463,N_12346);
nor U12681 (N_12681,N_12302,N_12482);
and U12682 (N_12682,N_12419,N_12319);
nor U12683 (N_12683,N_12436,N_12470);
nand U12684 (N_12684,N_12452,N_12349);
nor U12685 (N_12685,N_12338,N_12475);
xnor U12686 (N_12686,N_12302,N_12422);
and U12687 (N_12687,N_12366,N_12390);
and U12688 (N_12688,N_12281,N_12452);
or U12689 (N_12689,N_12355,N_12274);
nand U12690 (N_12690,N_12468,N_12352);
nor U12691 (N_12691,N_12424,N_12425);
or U12692 (N_12692,N_12432,N_12496);
xor U12693 (N_12693,N_12383,N_12398);
or U12694 (N_12694,N_12452,N_12464);
nand U12695 (N_12695,N_12457,N_12280);
or U12696 (N_12696,N_12453,N_12433);
or U12697 (N_12697,N_12357,N_12478);
nor U12698 (N_12698,N_12260,N_12443);
xor U12699 (N_12699,N_12451,N_12351);
xnor U12700 (N_12700,N_12294,N_12490);
nand U12701 (N_12701,N_12499,N_12419);
nor U12702 (N_12702,N_12429,N_12371);
nand U12703 (N_12703,N_12465,N_12439);
and U12704 (N_12704,N_12411,N_12374);
nand U12705 (N_12705,N_12486,N_12252);
nand U12706 (N_12706,N_12417,N_12259);
nand U12707 (N_12707,N_12350,N_12436);
and U12708 (N_12708,N_12259,N_12402);
nor U12709 (N_12709,N_12268,N_12433);
or U12710 (N_12710,N_12489,N_12284);
and U12711 (N_12711,N_12325,N_12411);
and U12712 (N_12712,N_12462,N_12444);
and U12713 (N_12713,N_12404,N_12429);
nand U12714 (N_12714,N_12259,N_12405);
xor U12715 (N_12715,N_12384,N_12380);
nor U12716 (N_12716,N_12369,N_12447);
and U12717 (N_12717,N_12486,N_12294);
nor U12718 (N_12718,N_12327,N_12376);
nand U12719 (N_12719,N_12346,N_12294);
and U12720 (N_12720,N_12372,N_12295);
and U12721 (N_12721,N_12416,N_12480);
nand U12722 (N_12722,N_12426,N_12365);
or U12723 (N_12723,N_12355,N_12374);
nand U12724 (N_12724,N_12263,N_12344);
nor U12725 (N_12725,N_12253,N_12388);
and U12726 (N_12726,N_12450,N_12497);
nor U12727 (N_12727,N_12368,N_12370);
nand U12728 (N_12728,N_12330,N_12365);
nand U12729 (N_12729,N_12296,N_12261);
nand U12730 (N_12730,N_12400,N_12265);
or U12731 (N_12731,N_12382,N_12282);
and U12732 (N_12732,N_12413,N_12323);
nor U12733 (N_12733,N_12409,N_12265);
and U12734 (N_12734,N_12404,N_12382);
and U12735 (N_12735,N_12453,N_12397);
nor U12736 (N_12736,N_12440,N_12326);
and U12737 (N_12737,N_12367,N_12425);
nor U12738 (N_12738,N_12347,N_12452);
nand U12739 (N_12739,N_12336,N_12476);
or U12740 (N_12740,N_12277,N_12414);
or U12741 (N_12741,N_12418,N_12474);
xnor U12742 (N_12742,N_12335,N_12430);
or U12743 (N_12743,N_12473,N_12260);
nor U12744 (N_12744,N_12461,N_12382);
nand U12745 (N_12745,N_12491,N_12267);
xnor U12746 (N_12746,N_12318,N_12444);
nand U12747 (N_12747,N_12492,N_12448);
nand U12748 (N_12748,N_12259,N_12340);
and U12749 (N_12749,N_12253,N_12281);
nor U12750 (N_12750,N_12520,N_12742);
or U12751 (N_12751,N_12688,N_12718);
nand U12752 (N_12752,N_12734,N_12673);
xnor U12753 (N_12753,N_12512,N_12537);
nor U12754 (N_12754,N_12651,N_12642);
nand U12755 (N_12755,N_12725,N_12635);
nand U12756 (N_12756,N_12667,N_12561);
nand U12757 (N_12757,N_12653,N_12728);
and U12758 (N_12758,N_12613,N_12618);
nand U12759 (N_12759,N_12549,N_12680);
or U12760 (N_12760,N_12581,N_12571);
or U12761 (N_12761,N_12593,N_12659);
or U12762 (N_12762,N_12647,N_12568);
xor U12763 (N_12763,N_12749,N_12553);
xor U12764 (N_12764,N_12617,N_12677);
xnor U12765 (N_12765,N_12563,N_12615);
nand U12766 (N_12766,N_12598,N_12574);
nand U12767 (N_12767,N_12610,N_12648);
xor U12768 (N_12768,N_12585,N_12560);
or U12769 (N_12769,N_12596,N_12562);
xor U12770 (N_12770,N_12518,N_12609);
nor U12771 (N_12771,N_12631,N_12645);
xnor U12772 (N_12772,N_12606,N_12692);
nand U12773 (N_12773,N_12736,N_12602);
nand U12774 (N_12774,N_12539,N_12729);
xor U12775 (N_12775,N_12541,N_12664);
xnor U12776 (N_12776,N_12723,N_12510);
or U12777 (N_12777,N_12592,N_12694);
or U12778 (N_12778,N_12545,N_12714);
and U12779 (N_12779,N_12501,N_12671);
nor U12780 (N_12780,N_12698,N_12589);
nand U12781 (N_12781,N_12579,N_12612);
xor U12782 (N_12782,N_12740,N_12731);
or U12783 (N_12783,N_12707,N_12614);
nor U12784 (N_12784,N_12576,N_12712);
nor U12785 (N_12785,N_12565,N_12661);
nor U12786 (N_12786,N_12535,N_12605);
and U12787 (N_12787,N_12687,N_12705);
nand U12788 (N_12788,N_12720,N_12670);
nor U12789 (N_12789,N_12538,N_12746);
and U12790 (N_12790,N_12646,N_12672);
xor U12791 (N_12791,N_12590,N_12511);
and U12792 (N_12792,N_12657,N_12516);
or U12793 (N_12793,N_12665,N_12638);
and U12794 (N_12794,N_12699,N_12679);
or U12795 (N_12795,N_12704,N_12587);
or U12796 (N_12796,N_12509,N_12675);
nor U12797 (N_12797,N_12683,N_12676);
nand U12798 (N_12798,N_12559,N_12633);
nor U12799 (N_12799,N_12662,N_12604);
nor U12800 (N_12800,N_12732,N_12548);
nand U12801 (N_12801,N_12722,N_12643);
and U12802 (N_12802,N_12697,N_12570);
nand U12803 (N_12803,N_12578,N_12564);
nor U12804 (N_12804,N_12626,N_12542);
and U12805 (N_12805,N_12678,N_12504);
or U12806 (N_12806,N_12572,N_12619);
and U12807 (N_12807,N_12706,N_12627);
nor U12808 (N_12808,N_12721,N_12715);
xor U12809 (N_12809,N_12573,N_12554);
nand U12810 (N_12810,N_12689,N_12555);
nor U12811 (N_12811,N_12621,N_12690);
and U12812 (N_12812,N_12650,N_12575);
or U12813 (N_12813,N_12517,N_12629);
nand U12814 (N_12814,N_12744,N_12558);
nor U12815 (N_12815,N_12603,N_12521);
and U12816 (N_12816,N_12727,N_12640);
nor U12817 (N_12817,N_12543,N_12547);
nand U12818 (N_12818,N_12591,N_12582);
nand U12819 (N_12819,N_12726,N_12717);
xor U12820 (N_12820,N_12616,N_12700);
or U12821 (N_12821,N_12710,N_12595);
nor U12822 (N_12822,N_12523,N_12551);
nand U12823 (N_12823,N_12569,N_12637);
or U12824 (N_12824,N_12533,N_12522);
nand U12825 (N_12825,N_12685,N_12524);
nor U12826 (N_12826,N_12682,N_12641);
nor U12827 (N_12827,N_12649,N_12703);
or U12828 (N_12828,N_12567,N_12748);
xor U12829 (N_12829,N_12654,N_12702);
and U12830 (N_12830,N_12639,N_12644);
nand U12831 (N_12831,N_12503,N_12634);
or U12832 (N_12832,N_12730,N_12508);
nor U12833 (N_12833,N_12527,N_12719);
nor U12834 (N_12834,N_12536,N_12530);
xnor U12835 (N_12835,N_12711,N_12599);
nor U12836 (N_12836,N_12684,N_12552);
nand U12837 (N_12837,N_12506,N_12745);
nor U12838 (N_12838,N_12695,N_12505);
or U12839 (N_12839,N_12630,N_12625);
or U12840 (N_12840,N_12611,N_12724);
nor U12841 (N_12841,N_12652,N_12566);
and U12842 (N_12842,N_12656,N_12636);
and U12843 (N_12843,N_12601,N_12747);
nand U12844 (N_12844,N_12507,N_12534);
nor U12845 (N_12845,N_12733,N_12686);
or U12846 (N_12846,N_12691,N_12577);
xor U12847 (N_12847,N_12738,N_12529);
nand U12848 (N_12848,N_12693,N_12655);
xnor U12849 (N_12849,N_12743,N_12594);
or U12850 (N_12850,N_12739,N_12531);
nor U12851 (N_12851,N_12584,N_12622);
xnor U12852 (N_12852,N_12623,N_12526);
nand U12853 (N_12853,N_12658,N_12546);
nand U12854 (N_12854,N_12586,N_12709);
and U12855 (N_12855,N_12532,N_12600);
and U12856 (N_12856,N_12624,N_12620);
xnor U12857 (N_12857,N_12663,N_12588);
nor U12858 (N_12858,N_12500,N_12701);
nor U12859 (N_12859,N_12525,N_12660);
or U12860 (N_12860,N_12674,N_12666);
nand U12861 (N_12861,N_12557,N_12607);
or U12862 (N_12862,N_12597,N_12540);
nor U12863 (N_12863,N_12556,N_12519);
and U12864 (N_12864,N_12696,N_12580);
or U12865 (N_12865,N_12583,N_12528);
or U12866 (N_12866,N_12669,N_12502);
nor U12867 (N_12867,N_12544,N_12708);
nor U12868 (N_12868,N_12737,N_12735);
xnor U12869 (N_12869,N_12632,N_12515);
nor U12870 (N_12870,N_12741,N_12513);
and U12871 (N_12871,N_12628,N_12713);
nand U12872 (N_12872,N_12514,N_12550);
nand U12873 (N_12873,N_12608,N_12681);
and U12874 (N_12874,N_12716,N_12668);
and U12875 (N_12875,N_12742,N_12748);
xnor U12876 (N_12876,N_12652,N_12704);
xnor U12877 (N_12877,N_12698,N_12531);
nor U12878 (N_12878,N_12646,N_12684);
xnor U12879 (N_12879,N_12624,N_12554);
and U12880 (N_12880,N_12560,N_12719);
or U12881 (N_12881,N_12713,N_12684);
nor U12882 (N_12882,N_12627,N_12660);
nor U12883 (N_12883,N_12550,N_12690);
or U12884 (N_12884,N_12572,N_12723);
or U12885 (N_12885,N_12531,N_12646);
nand U12886 (N_12886,N_12540,N_12501);
or U12887 (N_12887,N_12584,N_12559);
and U12888 (N_12888,N_12731,N_12644);
or U12889 (N_12889,N_12575,N_12742);
nand U12890 (N_12890,N_12557,N_12504);
nor U12891 (N_12891,N_12654,N_12679);
or U12892 (N_12892,N_12513,N_12694);
or U12893 (N_12893,N_12710,N_12732);
nor U12894 (N_12894,N_12608,N_12656);
and U12895 (N_12895,N_12591,N_12611);
and U12896 (N_12896,N_12539,N_12511);
and U12897 (N_12897,N_12709,N_12571);
nor U12898 (N_12898,N_12692,N_12639);
or U12899 (N_12899,N_12591,N_12643);
or U12900 (N_12900,N_12527,N_12537);
nor U12901 (N_12901,N_12597,N_12654);
xor U12902 (N_12902,N_12579,N_12608);
nor U12903 (N_12903,N_12565,N_12569);
nand U12904 (N_12904,N_12538,N_12695);
nor U12905 (N_12905,N_12615,N_12576);
and U12906 (N_12906,N_12525,N_12736);
or U12907 (N_12907,N_12507,N_12641);
nand U12908 (N_12908,N_12695,N_12526);
nand U12909 (N_12909,N_12580,N_12508);
nand U12910 (N_12910,N_12612,N_12657);
and U12911 (N_12911,N_12623,N_12716);
and U12912 (N_12912,N_12707,N_12746);
and U12913 (N_12913,N_12623,N_12525);
or U12914 (N_12914,N_12739,N_12659);
or U12915 (N_12915,N_12518,N_12743);
and U12916 (N_12916,N_12650,N_12545);
and U12917 (N_12917,N_12687,N_12542);
nand U12918 (N_12918,N_12522,N_12571);
and U12919 (N_12919,N_12622,N_12544);
nand U12920 (N_12920,N_12724,N_12648);
and U12921 (N_12921,N_12554,N_12716);
nand U12922 (N_12922,N_12627,N_12652);
nand U12923 (N_12923,N_12587,N_12575);
xor U12924 (N_12924,N_12592,N_12681);
xor U12925 (N_12925,N_12749,N_12724);
and U12926 (N_12926,N_12659,N_12707);
and U12927 (N_12927,N_12589,N_12576);
xor U12928 (N_12928,N_12635,N_12667);
or U12929 (N_12929,N_12520,N_12733);
or U12930 (N_12930,N_12658,N_12597);
nor U12931 (N_12931,N_12528,N_12551);
xor U12932 (N_12932,N_12598,N_12673);
or U12933 (N_12933,N_12582,N_12561);
nor U12934 (N_12934,N_12503,N_12729);
nand U12935 (N_12935,N_12540,N_12729);
nor U12936 (N_12936,N_12654,N_12621);
xor U12937 (N_12937,N_12609,N_12643);
and U12938 (N_12938,N_12669,N_12592);
xor U12939 (N_12939,N_12556,N_12590);
and U12940 (N_12940,N_12597,N_12659);
and U12941 (N_12941,N_12718,N_12597);
or U12942 (N_12942,N_12734,N_12516);
or U12943 (N_12943,N_12595,N_12508);
xor U12944 (N_12944,N_12745,N_12510);
nand U12945 (N_12945,N_12525,N_12697);
nor U12946 (N_12946,N_12653,N_12623);
and U12947 (N_12947,N_12708,N_12507);
nand U12948 (N_12948,N_12642,N_12521);
nand U12949 (N_12949,N_12688,N_12721);
nand U12950 (N_12950,N_12598,N_12576);
or U12951 (N_12951,N_12710,N_12612);
or U12952 (N_12952,N_12672,N_12560);
or U12953 (N_12953,N_12729,N_12506);
nand U12954 (N_12954,N_12691,N_12694);
nor U12955 (N_12955,N_12694,N_12714);
nand U12956 (N_12956,N_12606,N_12685);
nor U12957 (N_12957,N_12533,N_12580);
nor U12958 (N_12958,N_12596,N_12650);
xor U12959 (N_12959,N_12505,N_12575);
and U12960 (N_12960,N_12678,N_12568);
and U12961 (N_12961,N_12725,N_12664);
and U12962 (N_12962,N_12720,N_12710);
xnor U12963 (N_12963,N_12673,N_12540);
nand U12964 (N_12964,N_12672,N_12509);
nand U12965 (N_12965,N_12620,N_12724);
and U12966 (N_12966,N_12675,N_12731);
xor U12967 (N_12967,N_12582,N_12664);
nand U12968 (N_12968,N_12548,N_12674);
nor U12969 (N_12969,N_12535,N_12630);
nand U12970 (N_12970,N_12715,N_12696);
or U12971 (N_12971,N_12552,N_12691);
and U12972 (N_12972,N_12553,N_12557);
and U12973 (N_12973,N_12512,N_12661);
or U12974 (N_12974,N_12709,N_12597);
and U12975 (N_12975,N_12681,N_12734);
or U12976 (N_12976,N_12678,N_12632);
or U12977 (N_12977,N_12684,N_12553);
xnor U12978 (N_12978,N_12726,N_12685);
or U12979 (N_12979,N_12537,N_12690);
nor U12980 (N_12980,N_12540,N_12713);
xnor U12981 (N_12981,N_12748,N_12696);
xnor U12982 (N_12982,N_12527,N_12514);
and U12983 (N_12983,N_12684,N_12500);
nand U12984 (N_12984,N_12520,N_12594);
nor U12985 (N_12985,N_12542,N_12565);
nor U12986 (N_12986,N_12619,N_12696);
or U12987 (N_12987,N_12699,N_12592);
nor U12988 (N_12988,N_12693,N_12651);
xor U12989 (N_12989,N_12535,N_12631);
and U12990 (N_12990,N_12638,N_12522);
or U12991 (N_12991,N_12620,N_12553);
xor U12992 (N_12992,N_12731,N_12691);
and U12993 (N_12993,N_12539,N_12726);
xor U12994 (N_12994,N_12734,N_12747);
and U12995 (N_12995,N_12539,N_12560);
nor U12996 (N_12996,N_12606,N_12660);
and U12997 (N_12997,N_12608,N_12592);
xnor U12998 (N_12998,N_12515,N_12605);
or U12999 (N_12999,N_12565,N_12595);
or U13000 (N_13000,N_12754,N_12793);
and U13001 (N_13001,N_12896,N_12809);
nor U13002 (N_13002,N_12925,N_12802);
and U13003 (N_13003,N_12782,N_12808);
and U13004 (N_13004,N_12842,N_12970);
nand U13005 (N_13005,N_12982,N_12757);
xor U13006 (N_13006,N_12860,N_12894);
or U13007 (N_13007,N_12822,N_12934);
xor U13008 (N_13008,N_12848,N_12932);
and U13009 (N_13009,N_12920,N_12882);
and U13010 (N_13010,N_12996,N_12886);
nand U13011 (N_13011,N_12951,N_12918);
and U13012 (N_13012,N_12977,N_12993);
nor U13013 (N_13013,N_12928,N_12846);
nor U13014 (N_13014,N_12841,N_12930);
or U13015 (N_13015,N_12967,N_12946);
nand U13016 (N_13016,N_12844,N_12861);
nand U13017 (N_13017,N_12989,N_12881);
or U13018 (N_13018,N_12781,N_12839);
or U13019 (N_13019,N_12883,N_12891);
and U13020 (N_13020,N_12862,N_12807);
xor U13021 (N_13021,N_12922,N_12806);
or U13022 (N_13022,N_12837,N_12800);
nor U13023 (N_13023,N_12903,N_12905);
nand U13024 (N_13024,N_12972,N_12772);
nor U13025 (N_13025,N_12863,N_12816);
nand U13026 (N_13026,N_12798,N_12760);
xor U13027 (N_13027,N_12978,N_12872);
or U13028 (N_13028,N_12824,N_12829);
xor U13029 (N_13029,N_12874,N_12811);
nand U13030 (N_13030,N_12887,N_12799);
xor U13031 (N_13031,N_12937,N_12838);
and U13032 (N_13032,N_12942,N_12777);
or U13033 (N_13033,N_12756,N_12966);
nand U13034 (N_13034,N_12889,N_12865);
nand U13035 (N_13035,N_12955,N_12969);
nand U13036 (N_13036,N_12952,N_12975);
and U13037 (N_13037,N_12884,N_12795);
nor U13038 (N_13038,N_12769,N_12995);
xnor U13039 (N_13039,N_12893,N_12992);
or U13040 (N_13040,N_12752,N_12971);
or U13041 (N_13041,N_12871,N_12927);
and U13042 (N_13042,N_12912,N_12897);
and U13043 (N_13043,N_12876,N_12751);
nand U13044 (N_13044,N_12990,N_12774);
nand U13045 (N_13045,N_12900,N_12999);
nor U13046 (N_13046,N_12771,N_12895);
or U13047 (N_13047,N_12880,N_12787);
nand U13048 (N_13048,N_12941,N_12985);
and U13049 (N_13049,N_12812,N_12849);
or U13050 (N_13050,N_12899,N_12965);
or U13051 (N_13051,N_12898,N_12959);
xor U13052 (N_13052,N_12938,N_12974);
nand U13053 (N_13053,N_12851,N_12916);
xnor U13054 (N_13054,N_12820,N_12796);
xnor U13055 (N_13055,N_12950,N_12909);
nand U13056 (N_13056,N_12758,N_12924);
nor U13057 (N_13057,N_12931,N_12980);
nand U13058 (N_13058,N_12888,N_12998);
or U13059 (N_13059,N_12983,N_12981);
and U13060 (N_13060,N_12908,N_12776);
nand U13061 (N_13061,N_12847,N_12828);
or U13062 (N_13062,N_12929,N_12761);
and U13063 (N_13063,N_12832,N_12853);
and U13064 (N_13064,N_12765,N_12762);
and U13065 (N_13065,N_12814,N_12852);
nor U13066 (N_13066,N_12956,N_12875);
xor U13067 (N_13067,N_12858,N_12767);
xnor U13068 (N_13068,N_12819,N_12773);
nor U13069 (N_13069,N_12783,N_12830);
nand U13070 (N_13070,N_12994,N_12910);
or U13071 (N_13071,N_12854,N_12794);
nor U13072 (N_13072,N_12940,N_12792);
nand U13073 (N_13073,N_12813,N_12919);
nor U13074 (N_13074,N_12788,N_12803);
xor U13075 (N_13075,N_12833,N_12869);
nand U13076 (N_13076,N_12785,N_12789);
nand U13077 (N_13077,N_12836,N_12821);
nor U13078 (N_13078,N_12984,N_12964);
nand U13079 (N_13079,N_12986,N_12921);
xor U13080 (N_13080,N_12759,N_12943);
xor U13081 (N_13081,N_12963,N_12805);
nand U13082 (N_13082,N_12947,N_12823);
or U13083 (N_13083,N_12968,N_12835);
nand U13084 (N_13084,N_12850,N_12763);
and U13085 (N_13085,N_12868,N_12979);
or U13086 (N_13086,N_12917,N_12915);
nand U13087 (N_13087,N_12949,N_12933);
or U13088 (N_13088,N_12945,N_12864);
and U13089 (N_13089,N_12960,N_12834);
nand U13090 (N_13090,N_12775,N_12818);
and U13091 (N_13091,N_12815,N_12810);
xnor U13092 (N_13092,N_12907,N_12840);
xnor U13093 (N_13093,N_12753,N_12825);
or U13094 (N_13094,N_12911,N_12779);
and U13095 (N_13095,N_12866,N_12755);
nand U13096 (N_13096,N_12904,N_12826);
xor U13097 (N_13097,N_12843,N_12879);
xor U13098 (N_13098,N_12991,N_12948);
or U13099 (N_13099,N_12976,N_12855);
and U13100 (N_13100,N_12926,N_12867);
and U13101 (N_13101,N_12801,N_12804);
nand U13102 (N_13102,N_12906,N_12780);
nor U13103 (N_13103,N_12890,N_12797);
nor U13104 (N_13104,N_12957,N_12997);
xor U13105 (N_13105,N_12936,N_12902);
and U13106 (N_13106,N_12750,N_12885);
nand U13107 (N_13107,N_12831,N_12892);
nor U13108 (N_13108,N_12914,N_12944);
nand U13109 (N_13109,N_12786,N_12923);
nor U13110 (N_13110,N_12784,N_12766);
xnor U13111 (N_13111,N_12954,N_12857);
nand U13112 (N_13112,N_12827,N_12973);
or U13113 (N_13113,N_12764,N_12768);
nor U13114 (N_13114,N_12870,N_12961);
xnor U13115 (N_13115,N_12935,N_12913);
nand U13116 (N_13116,N_12878,N_12845);
nand U13117 (N_13117,N_12939,N_12953);
nor U13118 (N_13118,N_12988,N_12901);
nand U13119 (N_13119,N_12873,N_12791);
and U13120 (N_13120,N_12987,N_12856);
and U13121 (N_13121,N_12877,N_12778);
nor U13122 (N_13122,N_12790,N_12958);
nor U13123 (N_13123,N_12817,N_12770);
nor U13124 (N_13124,N_12859,N_12962);
xor U13125 (N_13125,N_12961,N_12755);
or U13126 (N_13126,N_12758,N_12869);
or U13127 (N_13127,N_12934,N_12963);
and U13128 (N_13128,N_12859,N_12986);
or U13129 (N_13129,N_12948,N_12960);
nor U13130 (N_13130,N_12996,N_12875);
nor U13131 (N_13131,N_12809,N_12916);
xnor U13132 (N_13132,N_12795,N_12807);
and U13133 (N_13133,N_12823,N_12864);
or U13134 (N_13134,N_12874,N_12788);
xor U13135 (N_13135,N_12870,N_12896);
and U13136 (N_13136,N_12867,N_12779);
xnor U13137 (N_13137,N_12952,N_12753);
xnor U13138 (N_13138,N_12785,N_12825);
or U13139 (N_13139,N_12832,N_12981);
or U13140 (N_13140,N_12796,N_12827);
or U13141 (N_13141,N_12885,N_12757);
nor U13142 (N_13142,N_12823,N_12911);
nor U13143 (N_13143,N_12962,N_12881);
or U13144 (N_13144,N_12876,N_12862);
nand U13145 (N_13145,N_12815,N_12934);
and U13146 (N_13146,N_12908,N_12758);
nand U13147 (N_13147,N_12959,N_12942);
xor U13148 (N_13148,N_12921,N_12922);
or U13149 (N_13149,N_12813,N_12903);
and U13150 (N_13150,N_12767,N_12825);
nand U13151 (N_13151,N_12897,N_12913);
nand U13152 (N_13152,N_12948,N_12990);
nor U13153 (N_13153,N_12756,N_12853);
nor U13154 (N_13154,N_12933,N_12895);
xor U13155 (N_13155,N_12776,N_12875);
nor U13156 (N_13156,N_12796,N_12777);
and U13157 (N_13157,N_12866,N_12853);
and U13158 (N_13158,N_12780,N_12956);
nand U13159 (N_13159,N_12781,N_12952);
nand U13160 (N_13160,N_12802,N_12883);
nor U13161 (N_13161,N_12793,N_12855);
nand U13162 (N_13162,N_12873,N_12943);
and U13163 (N_13163,N_12893,N_12825);
and U13164 (N_13164,N_12871,N_12945);
xor U13165 (N_13165,N_12973,N_12980);
nand U13166 (N_13166,N_12904,N_12939);
and U13167 (N_13167,N_12969,N_12780);
and U13168 (N_13168,N_12819,N_12850);
xnor U13169 (N_13169,N_12956,N_12837);
and U13170 (N_13170,N_12775,N_12993);
and U13171 (N_13171,N_12856,N_12942);
xnor U13172 (N_13172,N_12848,N_12750);
or U13173 (N_13173,N_12918,N_12828);
nor U13174 (N_13174,N_12888,N_12886);
and U13175 (N_13175,N_12791,N_12838);
xor U13176 (N_13176,N_12872,N_12902);
nor U13177 (N_13177,N_12812,N_12842);
xor U13178 (N_13178,N_12828,N_12786);
nand U13179 (N_13179,N_12783,N_12756);
nand U13180 (N_13180,N_12956,N_12928);
nor U13181 (N_13181,N_12793,N_12924);
nand U13182 (N_13182,N_12864,N_12805);
nand U13183 (N_13183,N_12885,N_12754);
nor U13184 (N_13184,N_12965,N_12896);
nand U13185 (N_13185,N_12827,N_12955);
nand U13186 (N_13186,N_12783,N_12820);
or U13187 (N_13187,N_12935,N_12751);
nor U13188 (N_13188,N_12879,N_12816);
nand U13189 (N_13189,N_12858,N_12805);
nand U13190 (N_13190,N_12800,N_12856);
xnor U13191 (N_13191,N_12780,N_12842);
and U13192 (N_13192,N_12906,N_12850);
or U13193 (N_13193,N_12834,N_12935);
nand U13194 (N_13194,N_12991,N_12931);
or U13195 (N_13195,N_12883,N_12990);
nand U13196 (N_13196,N_12790,N_12887);
xnor U13197 (N_13197,N_12762,N_12918);
nor U13198 (N_13198,N_12818,N_12950);
and U13199 (N_13199,N_12889,N_12754);
or U13200 (N_13200,N_12799,N_12814);
nand U13201 (N_13201,N_12820,N_12798);
xnor U13202 (N_13202,N_12882,N_12788);
nand U13203 (N_13203,N_12831,N_12844);
xor U13204 (N_13204,N_12930,N_12910);
nand U13205 (N_13205,N_12806,N_12973);
or U13206 (N_13206,N_12900,N_12928);
nor U13207 (N_13207,N_12885,N_12835);
nor U13208 (N_13208,N_12927,N_12949);
and U13209 (N_13209,N_12853,N_12962);
and U13210 (N_13210,N_12895,N_12755);
xnor U13211 (N_13211,N_12949,N_12841);
or U13212 (N_13212,N_12823,N_12857);
nand U13213 (N_13213,N_12810,N_12850);
and U13214 (N_13214,N_12902,N_12844);
nor U13215 (N_13215,N_12889,N_12848);
and U13216 (N_13216,N_12971,N_12938);
nand U13217 (N_13217,N_12838,N_12991);
xor U13218 (N_13218,N_12908,N_12972);
xnor U13219 (N_13219,N_12806,N_12809);
nand U13220 (N_13220,N_12813,N_12991);
or U13221 (N_13221,N_12836,N_12911);
or U13222 (N_13222,N_12856,N_12972);
xnor U13223 (N_13223,N_12792,N_12868);
nor U13224 (N_13224,N_12844,N_12890);
nand U13225 (N_13225,N_12793,N_12796);
nand U13226 (N_13226,N_12784,N_12753);
nor U13227 (N_13227,N_12899,N_12903);
and U13228 (N_13228,N_12797,N_12818);
or U13229 (N_13229,N_12857,N_12905);
and U13230 (N_13230,N_12937,N_12944);
or U13231 (N_13231,N_12896,N_12955);
or U13232 (N_13232,N_12931,N_12824);
and U13233 (N_13233,N_12799,N_12902);
nor U13234 (N_13234,N_12816,N_12903);
xnor U13235 (N_13235,N_12785,N_12973);
and U13236 (N_13236,N_12918,N_12812);
and U13237 (N_13237,N_12786,N_12989);
nand U13238 (N_13238,N_12978,N_12797);
xnor U13239 (N_13239,N_12929,N_12939);
nand U13240 (N_13240,N_12861,N_12860);
xor U13241 (N_13241,N_12884,N_12814);
nor U13242 (N_13242,N_12887,N_12961);
nor U13243 (N_13243,N_12806,N_12872);
or U13244 (N_13244,N_12808,N_12936);
and U13245 (N_13245,N_12826,N_12984);
and U13246 (N_13246,N_12813,N_12943);
xnor U13247 (N_13247,N_12888,N_12845);
or U13248 (N_13248,N_12841,N_12819);
nand U13249 (N_13249,N_12976,N_12767);
and U13250 (N_13250,N_13159,N_13035);
xnor U13251 (N_13251,N_13066,N_13201);
or U13252 (N_13252,N_13217,N_13017);
xor U13253 (N_13253,N_13056,N_13040);
nand U13254 (N_13254,N_13146,N_13224);
and U13255 (N_13255,N_13031,N_13178);
xnor U13256 (N_13256,N_13225,N_13108);
and U13257 (N_13257,N_13139,N_13241);
and U13258 (N_13258,N_13230,N_13240);
xor U13259 (N_13259,N_13203,N_13202);
and U13260 (N_13260,N_13106,N_13021);
or U13261 (N_13261,N_13245,N_13174);
xnor U13262 (N_13262,N_13218,N_13175);
xnor U13263 (N_13263,N_13212,N_13052);
and U13264 (N_13264,N_13238,N_13020);
xnor U13265 (N_13265,N_13115,N_13128);
xnor U13266 (N_13266,N_13247,N_13188);
xor U13267 (N_13267,N_13095,N_13064);
or U13268 (N_13268,N_13151,N_13177);
and U13269 (N_13269,N_13135,N_13235);
or U13270 (N_13270,N_13038,N_13029);
nand U13271 (N_13271,N_13185,N_13016);
or U13272 (N_13272,N_13243,N_13169);
xor U13273 (N_13273,N_13087,N_13167);
nor U13274 (N_13274,N_13157,N_13114);
nor U13275 (N_13275,N_13089,N_13024);
and U13276 (N_13276,N_13121,N_13078);
nor U13277 (N_13277,N_13227,N_13098);
and U13278 (N_13278,N_13189,N_13077);
nand U13279 (N_13279,N_13161,N_13007);
nand U13280 (N_13280,N_13136,N_13044);
or U13281 (N_13281,N_13155,N_13194);
nor U13282 (N_13282,N_13062,N_13083);
nor U13283 (N_13283,N_13039,N_13236);
or U13284 (N_13284,N_13242,N_13246);
nand U13285 (N_13285,N_13129,N_13050);
nand U13286 (N_13286,N_13120,N_13216);
and U13287 (N_13287,N_13150,N_13181);
nand U13288 (N_13288,N_13047,N_13075);
nand U13289 (N_13289,N_13099,N_13096);
nand U13290 (N_13290,N_13213,N_13208);
nor U13291 (N_13291,N_13080,N_13112);
or U13292 (N_13292,N_13148,N_13143);
or U13293 (N_13293,N_13109,N_13170);
nor U13294 (N_13294,N_13000,N_13011);
nand U13295 (N_13295,N_13018,N_13063);
xor U13296 (N_13296,N_13204,N_13045);
xnor U13297 (N_13297,N_13195,N_13125);
xor U13298 (N_13298,N_13074,N_13033);
nor U13299 (N_13299,N_13032,N_13207);
nor U13300 (N_13300,N_13184,N_13193);
or U13301 (N_13301,N_13015,N_13059);
nand U13302 (N_13302,N_13061,N_13126);
nor U13303 (N_13303,N_13152,N_13037);
nor U13304 (N_13304,N_13182,N_13168);
nor U13305 (N_13305,N_13090,N_13081);
nand U13306 (N_13306,N_13197,N_13205);
xnor U13307 (N_13307,N_13110,N_13053);
xor U13308 (N_13308,N_13104,N_13231);
xnor U13309 (N_13309,N_13009,N_13117);
or U13310 (N_13310,N_13060,N_13196);
nor U13311 (N_13311,N_13065,N_13093);
nand U13312 (N_13312,N_13226,N_13036);
and U13313 (N_13313,N_13149,N_13012);
nand U13314 (N_13314,N_13048,N_13119);
nand U13315 (N_13315,N_13076,N_13014);
xor U13316 (N_13316,N_13091,N_13237);
or U13317 (N_13317,N_13034,N_13043);
nor U13318 (N_13318,N_13111,N_13123);
nor U13319 (N_13319,N_13141,N_13041);
nand U13320 (N_13320,N_13137,N_13210);
nor U13321 (N_13321,N_13215,N_13232);
nor U13322 (N_13322,N_13191,N_13220);
or U13323 (N_13323,N_13030,N_13122);
nor U13324 (N_13324,N_13082,N_13097);
xnor U13325 (N_13325,N_13166,N_13154);
and U13326 (N_13326,N_13179,N_13228);
or U13327 (N_13327,N_13192,N_13173);
and U13328 (N_13328,N_13249,N_13234);
nand U13329 (N_13329,N_13214,N_13102);
nor U13330 (N_13330,N_13172,N_13134);
and U13331 (N_13331,N_13068,N_13219);
or U13332 (N_13332,N_13142,N_13019);
nor U13333 (N_13333,N_13092,N_13013);
xnor U13334 (N_13334,N_13248,N_13086);
and U13335 (N_13335,N_13131,N_13084);
and U13336 (N_13336,N_13105,N_13107);
nor U13337 (N_13337,N_13164,N_13088);
and U13338 (N_13338,N_13156,N_13163);
and U13339 (N_13339,N_13116,N_13211);
xnor U13340 (N_13340,N_13003,N_13186);
and U13341 (N_13341,N_13070,N_13160);
xnor U13342 (N_13342,N_13100,N_13094);
nor U13343 (N_13343,N_13153,N_13118);
and U13344 (N_13344,N_13171,N_13001);
or U13345 (N_13345,N_13206,N_13002);
and U13346 (N_13346,N_13209,N_13162);
nor U13347 (N_13347,N_13199,N_13057);
and U13348 (N_13348,N_13028,N_13058);
xnor U13349 (N_13349,N_13132,N_13187);
nand U13350 (N_13350,N_13101,N_13190);
xor U13351 (N_13351,N_13055,N_13180);
and U13352 (N_13352,N_13067,N_13026);
nand U13353 (N_13353,N_13023,N_13165);
or U13354 (N_13354,N_13073,N_13005);
nor U13355 (N_13355,N_13071,N_13072);
nor U13356 (N_13356,N_13027,N_13085);
nor U13357 (N_13357,N_13138,N_13221);
nand U13358 (N_13358,N_13176,N_13006);
nor U13359 (N_13359,N_13054,N_13127);
nor U13360 (N_13360,N_13198,N_13049);
and U13361 (N_13361,N_13140,N_13244);
and U13362 (N_13362,N_13103,N_13239);
xnor U13363 (N_13363,N_13069,N_13025);
xnor U13364 (N_13364,N_13223,N_13229);
or U13365 (N_13365,N_13144,N_13113);
or U13366 (N_13366,N_13133,N_13147);
xnor U13367 (N_13367,N_13008,N_13158);
nand U13368 (N_13368,N_13004,N_13042);
or U13369 (N_13369,N_13183,N_13233);
nand U13370 (N_13370,N_13010,N_13022);
nor U13371 (N_13371,N_13145,N_13124);
nand U13372 (N_13372,N_13079,N_13051);
nor U13373 (N_13373,N_13130,N_13200);
nand U13374 (N_13374,N_13046,N_13222);
or U13375 (N_13375,N_13180,N_13113);
nor U13376 (N_13376,N_13009,N_13064);
and U13377 (N_13377,N_13012,N_13225);
and U13378 (N_13378,N_13154,N_13131);
and U13379 (N_13379,N_13226,N_13152);
and U13380 (N_13380,N_13227,N_13084);
xor U13381 (N_13381,N_13019,N_13037);
nor U13382 (N_13382,N_13193,N_13244);
xnor U13383 (N_13383,N_13109,N_13079);
and U13384 (N_13384,N_13005,N_13207);
and U13385 (N_13385,N_13192,N_13225);
and U13386 (N_13386,N_13123,N_13224);
and U13387 (N_13387,N_13157,N_13004);
xor U13388 (N_13388,N_13187,N_13118);
and U13389 (N_13389,N_13021,N_13122);
nor U13390 (N_13390,N_13010,N_13222);
and U13391 (N_13391,N_13127,N_13076);
xor U13392 (N_13392,N_13209,N_13024);
and U13393 (N_13393,N_13213,N_13027);
and U13394 (N_13394,N_13002,N_13216);
nand U13395 (N_13395,N_13049,N_13215);
nor U13396 (N_13396,N_13121,N_13232);
or U13397 (N_13397,N_13136,N_13208);
nor U13398 (N_13398,N_13229,N_13049);
nor U13399 (N_13399,N_13088,N_13001);
xnor U13400 (N_13400,N_13241,N_13124);
xnor U13401 (N_13401,N_13025,N_13154);
and U13402 (N_13402,N_13095,N_13149);
and U13403 (N_13403,N_13056,N_13230);
nor U13404 (N_13404,N_13065,N_13202);
xor U13405 (N_13405,N_13240,N_13161);
nand U13406 (N_13406,N_13177,N_13212);
and U13407 (N_13407,N_13063,N_13132);
xnor U13408 (N_13408,N_13195,N_13076);
nand U13409 (N_13409,N_13043,N_13025);
nor U13410 (N_13410,N_13074,N_13200);
or U13411 (N_13411,N_13079,N_13236);
nand U13412 (N_13412,N_13161,N_13194);
and U13413 (N_13413,N_13061,N_13045);
nand U13414 (N_13414,N_13192,N_13038);
and U13415 (N_13415,N_13002,N_13152);
nor U13416 (N_13416,N_13179,N_13133);
xor U13417 (N_13417,N_13082,N_13049);
and U13418 (N_13418,N_13044,N_13089);
nand U13419 (N_13419,N_13210,N_13116);
xor U13420 (N_13420,N_13102,N_13183);
xnor U13421 (N_13421,N_13196,N_13079);
nand U13422 (N_13422,N_13154,N_13030);
nor U13423 (N_13423,N_13210,N_13002);
nand U13424 (N_13424,N_13202,N_13213);
and U13425 (N_13425,N_13153,N_13240);
or U13426 (N_13426,N_13224,N_13246);
and U13427 (N_13427,N_13209,N_13182);
or U13428 (N_13428,N_13216,N_13145);
nand U13429 (N_13429,N_13139,N_13009);
and U13430 (N_13430,N_13024,N_13003);
xor U13431 (N_13431,N_13139,N_13147);
nor U13432 (N_13432,N_13004,N_13187);
or U13433 (N_13433,N_13218,N_13095);
xnor U13434 (N_13434,N_13013,N_13088);
and U13435 (N_13435,N_13078,N_13084);
xnor U13436 (N_13436,N_13051,N_13073);
xor U13437 (N_13437,N_13033,N_13169);
nand U13438 (N_13438,N_13247,N_13047);
nor U13439 (N_13439,N_13216,N_13060);
and U13440 (N_13440,N_13149,N_13189);
nor U13441 (N_13441,N_13103,N_13044);
nor U13442 (N_13442,N_13215,N_13016);
nand U13443 (N_13443,N_13048,N_13043);
nand U13444 (N_13444,N_13232,N_13095);
and U13445 (N_13445,N_13228,N_13236);
nand U13446 (N_13446,N_13096,N_13119);
nand U13447 (N_13447,N_13052,N_13110);
xnor U13448 (N_13448,N_13241,N_13206);
or U13449 (N_13449,N_13088,N_13089);
nor U13450 (N_13450,N_13108,N_13033);
nand U13451 (N_13451,N_13236,N_13212);
and U13452 (N_13452,N_13048,N_13091);
xor U13453 (N_13453,N_13126,N_13152);
or U13454 (N_13454,N_13039,N_13006);
or U13455 (N_13455,N_13207,N_13172);
nor U13456 (N_13456,N_13213,N_13111);
nor U13457 (N_13457,N_13105,N_13017);
nand U13458 (N_13458,N_13192,N_13020);
or U13459 (N_13459,N_13195,N_13023);
nor U13460 (N_13460,N_13216,N_13097);
and U13461 (N_13461,N_13025,N_13177);
and U13462 (N_13462,N_13164,N_13227);
or U13463 (N_13463,N_13007,N_13115);
nor U13464 (N_13464,N_13100,N_13123);
nand U13465 (N_13465,N_13041,N_13019);
nor U13466 (N_13466,N_13071,N_13125);
xor U13467 (N_13467,N_13221,N_13099);
and U13468 (N_13468,N_13099,N_13114);
xnor U13469 (N_13469,N_13144,N_13244);
or U13470 (N_13470,N_13005,N_13022);
and U13471 (N_13471,N_13129,N_13089);
xnor U13472 (N_13472,N_13191,N_13061);
xnor U13473 (N_13473,N_13135,N_13241);
xor U13474 (N_13474,N_13031,N_13105);
xnor U13475 (N_13475,N_13020,N_13061);
xnor U13476 (N_13476,N_13087,N_13071);
or U13477 (N_13477,N_13208,N_13234);
or U13478 (N_13478,N_13019,N_13029);
and U13479 (N_13479,N_13231,N_13043);
xnor U13480 (N_13480,N_13090,N_13077);
and U13481 (N_13481,N_13237,N_13170);
xor U13482 (N_13482,N_13192,N_13139);
nand U13483 (N_13483,N_13174,N_13029);
xor U13484 (N_13484,N_13168,N_13053);
nand U13485 (N_13485,N_13202,N_13197);
nor U13486 (N_13486,N_13036,N_13185);
xnor U13487 (N_13487,N_13045,N_13019);
xnor U13488 (N_13488,N_13055,N_13240);
xor U13489 (N_13489,N_13183,N_13141);
nand U13490 (N_13490,N_13104,N_13152);
and U13491 (N_13491,N_13233,N_13194);
or U13492 (N_13492,N_13119,N_13092);
nor U13493 (N_13493,N_13249,N_13169);
or U13494 (N_13494,N_13179,N_13200);
nor U13495 (N_13495,N_13173,N_13013);
nand U13496 (N_13496,N_13128,N_13164);
nand U13497 (N_13497,N_13086,N_13206);
nand U13498 (N_13498,N_13180,N_13095);
xnor U13499 (N_13499,N_13222,N_13023);
or U13500 (N_13500,N_13252,N_13346);
and U13501 (N_13501,N_13289,N_13444);
and U13502 (N_13502,N_13463,N_13253);
and U13503 (N_13503,N_13337,N_13474);
nand U13504 (N_13504,N_13469,N_13334);
and U13505 (N_13505,N_13449,N_13448);
and U13506 (N_13506,N_13491,N_13312);
xnor U13507 (N_13507,N_13440,N_13261);
and U13508 (N_13508,N_13255,N_13488);
xnor U13509 (N_13509,N_13303,N_13340);
xor U13510 (N_13510,N_13296,N_13436);
nand U13511 (N_13511,N_13392,N_13386);
or U13512 (N_13512,N_13409,N_13470);
and U13513 (N_13513,N_13356,N_13313);
and U13514 (N_13514,N_13351,N_13357);
nor U13515 (N_13515,N_13472,N_13464);
nand U13516 (N_13516,N_13323,N_13344);
nor U13517 (N_13517,N_13427,N_13426);
or U13518 (N_13518,N_13434,N_13382);
xor U13519 (N_13519,N_13370,N_13264);
and U13520 (N_13520,N_13421,N_13330);
nand U13521 (N_13521,N_13379,N_13499);
nor U13522 (N_13522,N_13481,N_13398);
nand U13523 (N_13523,N_13367,N_13332);
and U13524 (N_13524,N_13494,N_13271);
nor U13525 (N_13525,N_13416,N_13401);
nor U13526 (N_13526,N_13288,N_13305);
nand U13527 (N_13527,N_13453,N_13454);
nor U13528 (N_13528,N_13487,N_13428);
and U13529 (N_13529,N_13433,N_13358);
nand U13530 (N_13530,N_13497,N_13347);
or U13531 (N_13531,N_13399,N_13310);
or U13532 (N_13532,N_13282,N_13402);
nor U13533 (N_13533,N_13269,N_13498);
and U13534 (N_13534,N_13277,N_13394);
or U13535 (N_13535,N_13300,N_13315);
nor U13536 (N_13536,N_13257,N_13293);
xnor U13537 (N_13537,N_13359,N_13423);
and U13538 (N_13538,N_13299,N_13435);
or U13539 (N_13539,N_13405,N_13361);
nor U13540 (N_13540,N_13384,N_13287);
and U13541 (N_13541,N_13281,N_13495);
or U13542 (N_13542,N_13492,N_13383);
or U13543 (N_13543,N_13280,N_13466);
or U13544 (N_13544,N_13286,N_13335);
nand U13545 (N_13545,N_13341,N_13294);
nor U13546 (N_13546,N_13336,N_13459);
nor U13547 (N_13547,N_13302,N_13324);
xnor U13548 (N_13548,N_13429,N_13484);
or U13549 (N_13549,N_13363,N_13420);
xor U13550 (N_13550,N_13489,N_13317);
and U13551 (N_13551,N_13268,N_13397);
xnor U13552 (N_13552,N_13328,N_13365);
and U13553 (N_13553,N_13339,N_13400);
or U13554 (N_13554,N_13283,N_13352);
and U13555 (N_13555,N_13258,N_13276);
xor U13556 (N_13556,N_13417,N_13375);
nor U13557 (N_13557,N_13267,N_13476);
xor U13558 (N_13558,N_13414,N_13331);
and U13559 (N_13559,N_13362,N_13446);
nor U13560 (N_13560,N_13273,N_13290);
or U13561 (N_13561,N_13343,N_13263);
and U13562 (N_13562,N_13298,N_13322);
xor U13563 (N_13563,N_13376,N_13460);
and U13564 (N_13564,N_13393,N_13278);
or U13565 (N_13565,N_13260,N_13285);
xor U13566 (N_13566,N_13430,N_13396);
xnor U13567 (N_13567,N_13471,N_13439);
or U13568 (N_13568,N_13389,N_13274);
and U13569 (N_13569,N_13371,N_13301);
xnor U13570 (N_13570,N_13364,N_13473);
nor U13571 (N_13571,N_13493,N_13490);
or U13572 (N_13572,N_13462,N_13265);
or U13573 (N_13573,N_13441,N_13461);
or U13574 (N_13574,N_13412,N_13411);
xnor U13575 (N_13575,N_13284,N_13374);
xnor U13576 (N_13576,N_13390,N_13377);
nor U13577 (N_13577,N_13348,N_13403);
and U13578 (N_13578,N_13477,N_13445);
and U13579 (N_13579,N_13295,N_13432);
and U13580 (N_13580,N_13329,N_13319);
or U13581 (N_13581,N_13482,N_13372);
xor U13582 (N_13582,N_13483,N_13369);
or U13583 (N_13583,N_13388,N_13431);
nand U13584 (N_13584,N_13304,N_13314);
or U13585 (N_13585,N_13316,N_13422);
and U13586 (N_13586,N_13468,N_13404);
or U13587 (N_13587,N_13478,N_13456);
xor U13588 (N_13588,N_13327,N_13254);
nand U13589 (N_13589,N_13381,N_13408);
xor U13590 (N_13590,N_13425,N_13373);
and U13591 (N_13591,N_13309,N_13378);
and U13592 (N_13592,N_13380,N_13297);
and U13593 (N_13593,N_13424,N_13279);
nand U13594 (N_13594,N_13366,N_13407);
xnor U13595 (N_13595,N_13318,N_13387);
and U13596 (N_13596,N_13272,N_13354);
or U13597 (N_13597,N_13413,N_13262);
or U13598 (N_13598,N_13251,N_13292);
and U13599 (N_13599,N_13368,N_13479);
nand U13600 (N_13600,N_13350,N_13306);
or U13601 (N_13601,N_13486,N_13270);
or U13602 (N_13602,N_13438,N_13475);
or U13603 (N_13603,N_13345,N_13418);
and U13604 (N_13604,N_13485,N_13442);
and U13605 (N_13605,N_13250,N_13452);
and U13606 (N_13606,N_13333,N_13326);
xnor U13607 (N_13607,N_13415,N_13391);
xor U13608 (N_13608,N_13311,N_13320);
or U13609 (N_13609,N_13355,N_13353);
xor U13610 (N_13610,N_13467,N_13451);
nand U13611 (N_13611,N_13266,N_13325);
or U13612 (N_13612,N_13496,N_13256);
xnor U13613 (N_13613,N_13395,N_13308);
xor U13614 (N_13614,N_13457,N_13455);
xnor U13615 (N_13615,N_13480,N_13458);
nand U13616 (N_13616,N_13385,N_13275);
xnor U13617 (N_13617,N_13321,N_13349);
xnor U13618 (N_13618,N_13437,N_13342);
or U13619 (N_13619,N_13443,N_13419);
nand U13620 (N_13620,N_13259,N_13450);
nand U13621 (N_13621,N_13465,N_13447);
nand U13622 (N_13622,N_13410,N_13406);
nor U13623 (N_13623,N_13360,N_13338);
and U13624 (N_13624,N_13307,N_13291);
xor U13625 (N_13625,N_13448,N_13446);
nand U13626 (N_13626,N_13338,N_13419);
nand U13627 (N_13627,N_13342,N_13463);
or U13628 (N_13628,N_13471,N_13415);
xor U13629 (N_13629,N_13361,N_13403);
or U13630 (N_13630,N_13459,N_13472);
or U13631 (N_13631,N_13485,N_13400);
or U13632 (N_13632,N_13479,N_13282);
nor U13633 (N_13633,N_13332,N_13399);
nand U13634 (N_13634,N_13274,N_13497);
xnor U13635 (N_13635,N_13490,N_13424);
or U13636 (N_13636,N_13419,N_13278);
and U13637 (N_13637,N_13396,N_13415);
nor U13638 (N_13638,N_13372,N_13484);
nand U13639 (N_13639,N_13281,N_13292);
xor U13640 (N_13640,N_13432,N_13352);
or U13641 (N_13641,N_13423,N_13269);
xnor U13642 (N_13642,N_13428,N_13455);
nor U13643 (N_13643,N_13444,N_13364);
nand U13644 (N_13644,N_13257,N_13453);
nand U13645 (N_13645,N_13300,N_13253);
or U13646 (N_13646,N_13406,N_13281);
or U13647 (N_13647,N_13410,N_13420);
and U13648 (N_13648,N_13439,N_13472);
nor U13649 (N_13649,N_13251,N_13491);
and U13650 (N_13650,N_13370,N_13467);
nand U13651 (N_13651,N_13407,N_13338);
and U13652 (N_13652,N_13444,N_13282);
or U13653 (N_13653,N_13466,N_13499);
xor U13654 (N_13654,N_13387,N_13488);
nor U13655 (N_13655,N_13403,N_13252);
and U13656 (N_13656,N_13356,N_13372);
and U13657 (N_13657,N_13349,N_13410);
xnor U13658 (N_13658,N_13407,N_13447);
and U13659 (N_13659,N_13347,N_13403);
xor U13660 (N_13660,N_13256,N_13251);
or U13661 (N_13661,N_13497,N_13423);
nand U13662 (N_13662,N_13422,N_13303);
or U13663 (N_13663,N_13366,N_13382);
and U13664 (N_13664,N_13268,N_13408);
xor U13665 (N_13665,N_13359,N_13479);
nand U13666 (N_13666,N_13433,N_13305);
and U13667 (N_13667,N_13465,N_13318);
nor U13668 (N_13668,N_13385,N_13323);
and U13669 (N_13669,N_13469,N_13311);
nor U13670 (N_13670,N_13299,N_13258);
nand U13671 (N_13671,N_13459,N_13404);
nand U13672 (N_13672,N_13259,N_13335);
nand U13673 (N_13673,N_13416,N_13363);
nor U13674 (N_13674,N_13262,N_13265);
and U13675 (N_13675,N_13389,N_13275);
nand U13676 (N_13676,N_13374,N_13470);
xor U13677 (N_13677,N_13252,N_13304);
or U13678 (N_13678,N_13493,N_13440);
and U13679 (N_13679,N_13398,N_13485);
and U13680 (N_13680,N_13337,N_13415);
xor U13681 (N_13681,N_13353,N_13431);
or U13682 (N_13682,N_13456,N_13314);
xnor U13683 (N_13683,N_13401,N_13252);
nor U13684 (N_13684,N_13312,N_13274);
nand U13685 (N_13685,N_13461,N_13353);
xor U13686 (N_13686,N_13291,N_13290);
and U13687 (N_13687,N_13357,N_13486);
nand U13688 (N_13688,N_13351,N_13403);
nand U13689 (N_13689,N_13329,N_13429);
or U13690 (N_13690,N_13398,N_13375);
xor U13691 (N_13691,N_13420,N_13254);
xnor U13692 (N_13692,N_13382,N_13367);
and U13693 (N_13693,N_13421,N_13402);
nand U13694 (N_13694,N_13313,N_13446);
nor U13695 (N_13695,N_13303,N_13286);
or U13696 (N_13696,N_13323,N_13301);
xnor U13697 (N_13697,N_13485,N_13387);
and U13698 (N_13698,N_13358,N_13311);
or U13699 (N_13699,N_13453,N_13350);
or U13700 (N_13700,N_13325,N_13491);
nand U13701 (N_13701,N_13479,N_13428);
and U13702 (N_13702,N_13424,N_13261);
xnor U13703 (N_13703,N_13280,N_13334);
xnor U13704 (N_13704,N_13263,N_13385);
xnor U13705 (N_13705,N_13392,N_13497);
and U13706 (N_13706,N_13491,N_13459);
xor U13707 (N_13707,N_13425,N_13261);
nand U13708 (N_13708,N_13314,N_13400);
and U13709 (N_13709,N_13273,N_13499);
and U13710 (N_13710,N_13256,N_13252);
or U13711 (N_13711,N_13312,N_13461);
nand U13712 (N_13712,N_13477,N_13275);
nand U13713 (N_13713,N_13379,N_13388);
nor U13714 (N_13714,N_13304,N_13499);
nor U13715 (N_13715,N_13487,N_13495);
xor U13716 (N_13716,N_13427,N_13474);
and U13717 (N_13717,N_13289,N_13497);
xnor U13718 (N_13718,N_13371,N_13468);
nand U13719 (N_13719,N_13291,N_13331);
and U13720 (N_13720,N_13288,N_13331);
or U13721 (N_13721,N_13376,N_13255);
xor U13722 (N_13722,N_13477,N_13450);
and U13723 (N_13723,N_13387,N_13402);
nor U13724 (N_13724,N_13326,N_13452);
xor U13725 (N_13725,N_13345,N_13267);
and U13726 (N_13726,N_13372,N_13380);
nor U13727 (N_13727,N_13301,N_13362);
xor U13728 (N_13728,N_13336,N_13479);
nand U13729 (N_13729,N_13258,N_13264);
xnor U13730 (N_13730,N_13361,N_13270);
nand U13731 (N_13731,N_13393,N_13459);
xor U13732 (N_13732,N_13303,N_13477);
xnor U13733 (N_13733,N_13316,N_13443);
xnor U13734 (N_13734,N_13252,N_13347);
and U13735 (N_13735,N_13349,N_13424);
and U13736 (N_13736,N_13321,N_13422);
and U13737 (N_13737,N_13472,N_13421);
nor U13738 (N_13738,N_13310,N_13306);
nor U13739 (N_13739,N_13496,N_13498);
or U13740 (N_13740,N_13313,N_13337);
nand U13741 (N_13741,N_13363,N_13395);
xor U13742 (N_13742,N_13471,N_13297);
or U13743 (N_13743,N_13455,N_13445);
xor U13744 (N_13744,N_13342,N_13360);
nand U13745 (N_13745,N_13360,N_13422);
nand U13746 (N_13746,N_13456,N_13447);
nand U13747 (N_13747,N_13431,N_13390);
nand U13748 (N_13748,N_13292,N_13495);
and U13749 (N_13749,N_13330,N_13496);
xor U13750 (N_13750,N_13658,N_13522);
nand U13751 (N_13751,N_13632,N_13540);
or U13752 (N_13752,N_13686,N_13556);
nand U13753 (N_13753,N_13608,N_13643);
nand U13754 (N_13754,N_13672,N_13718);
nand U13755 (N_13755,N_13655,N_13679);
nand U13756 (N_13756,N_13710,N_13576);
and U13757 (N_13757,N_13558,N_13708);
xor U13758 (N_13758,N_13518,N_13562);
or U13759 (N_13759,N_13692,N_13744);
and U13760 (N_13760,N_13590,N_13728);
or U13761 (N_13761,N_13695,N_13624);
and U13762 (N_13762,N_13694,N_13525);
nand U13763 (N_13763,N_13527,N_13661);
or U13764 (N_13764,N_13603,N_13524);
and U13765 (N_13765,N_13700,N_13572);
and U13766 (N_13766,N_13662,N_13649);
nand U13767 (N_13767,N_13618,N_13668);
or U13768 (N_13768,N_13704,N_13516);
and U13769 (N_13769,N_13610,N_13712);
nor U13770 (N_13770,N_13585,N_13602);
or U13771 (N_13771,N_13507,N_13538);
xnor U13772 (N_13772,N_13663,N_13721);
or U13773 (N_13773,N_13553,N_13521);
or U13774 (N_13774,N_13535,N_13620);
or U13775 (N_13775,N_13641,N_13616);
nand U13776 (N_13776,N_13706,N_13681);
nand U13777 (N_13777,N_13723,N_13564);
nor U13778 (N_13778,N_13554,N_13523);
nand U13779 (N_13779,N_13514,N_13738);
nand U13780 (N_13780,N_13515,N_13628);
or U13781 (N_13781,N_13670,N_13653);
and U13782 (N_13782,N_13683,N_13642);
and U13783 (N_13783,N_13664,N_13536);
and U13784 (N_13784,N_13665,N_13740);
nand U13785 (N_13785,N_13648,N_13598);
or U13786 (N_13786,N_13577,N_13551);
or U13787 (N_13787,N_13715,N_13578);
or U13788 (N_13788,N_13651,N_13594);
and U13789 (N_13789,N_13689,N_13619);
and U13790 (N_13790,N_13592,N_13702);
nor U13791 (N_13791,N_13501,N_13621);
nand U13792 (N_13792,N_13749,N_13505);
or U13793 (N_13793,N_13506,N_13720);
nand U13794 (N_13794,N_13543,N_13609);
and U13795 (N_13795,N_13529,N_13705);
nor U13796 (N_13796,N_13605,N_13550);
or U13797 (N_13797,N_13588,N_13682);
and U13798 (N_13798,N_13617,N_13526);
xnor U13799 (N_13799,N_13688,N_13659);
or U13800 (N_13800,N_13500,N_13511);
nor U13801 (N_13801,N_13560,N_13656);
and U13802 (N_13802,N_13690,N_13549);
nand U13803 (N_13803,N_13719,N_13697);
and U13804 (N_13804,N_13508,N_13680);
nor U13805 (N_13805,N_13532,N_13513);
nand U13806 (N_13806,N_13504,N_13623);
or U13807 (N_13807,N_13583,N_13735);
nor U13808 (N_13808,N_13555,N_13650);
and U13809 (N_13809,N_13584,N_13547);
xnor U13810 (N_13810,N_13646,N_13737);
xor U13811 (N_13811,N_13636,N_13579);
nand U13812 (N_13812,N_13630,N_13745);
or U13813 (N_13813,N_13716,N_13746);
or U13814 (N_13814,N_13559,N_13582);
or U13815 (N_13815,N_13509,N_13729);
or U13816 (N_13816,N_13569,N_13546);
nor U13817 (N_13817,N_13652,N_13742);
xor U13818 (N_13818,N_13666,N_13595);
or U13819 (N_13819,N_13713,N_13600);
xnor U13820 (N_13820,N_13685,N_13732);
nand U13821 (N_13821,N_13667,N_13520);
nor U13822 (N_13822,N_13635,N_13698);
and U13823 (N_13823,N_13565,N_13727);
or U13824 (N_13824,N_13596,N_13519);
and U13825 (N_13825,N_13613,N_13517);
xor U13826 (N_13826,N_13601,N_13539);
xor U13827 (N_13827,N_13530,N_13731);
and U13828 (N_13828,N_13726,N_13677);
and U13829 (N_13829,N_13587,N_13589);
nor U13830 (N_13830,N_13612,N_13730);
nand U13831 (N_13831,N_13674,N_13510);
xor U13832 (N_13832,N_13736,N_13627);
nand U13833 (N_13833,N_13638,N_13599);
nand U13834 (N_13834,N_13678,N_13671);
xnor U13835 (N_13835,N_13574,N_13639);
and U13836 (N_13836,N_13633,N_13631);
and U13837 (N_13837,N_13542,N_13673);
and U13838 (N_13838,N_13657,N_13724);
and U13839 (N_13839,N_13586,N_13591);
xnor U13840 (N_13840,N_13687,N_13733);
nand U13841 (N_13841,N_13552,N_13645);
nor U13842 (N_13842,N_13725,N_13676);
nand U13843 (N_13843,N_13566,N_13570);
nand U13844 (N_13844,N_13614,N_13544);
xor U13845 (N_13845,N_13699,N_13714);
nor U13846 (N_13846,N_13640,N_13644);
nand U13847 (N_13847,N_13561,N_13573);
nor U13848 (N_13848,N_13563,N_13545);
xnor U13849 (N_13849,N_13597,N_13548);
nand U13850 (N_13850,N_13611,N_13626);
nor U13851 (N_13851,N_13647,N_13534);
nor U13852 (N_13852,N_13581,N_13537);
and U13853 (N_13853,N_13625,N_13528);
xor U13854 (N_13854,N_13568,N_13660);
and U13855 (N_13855,N_13615,N_13739);
and U13856 (N_13856,N_13593,N_13575);
nor U13857 (N_13857,N_13709,N_13684);
and U13858 (N_13858,N_13654,N_13701);
and U13859 (N_13859,N_13696,N_13669);
nor U13860 (N_13860,N_13691,N_13747);
xnor U13861 (N_13861,N_13541,N_13567);
nor U13862 (N_13862,N_13748,N_13717);
xnor U13863 (N_13863,N_13604,N_13622);
and U13864 (N_13864,N_13734,N_13571);
xor U13865 (N_13865,N_13741,N_13503);
and U13866 (N_13866,N_13743,N_13711);
nand U13867 (N_13867,N_13557,N_13512);
or U13868 (N_13868,N_13607,N_13606);
and U13869 (N_13869,N_13580,N_13634);
nand U13870 (N_13870,N_13502,N_13703);
or U13871 (N_13871,N_13693,N_13533);
nand U13872 (N_13872,N_13707,N_13637);
xor U13873 (N_13873,N_13722,N_13675);
xnor U13874 (N_13874,N_13531,N_13629);
nand U13875 (N_13875,N_13713,N_13652);
nor U13876 (N_13876,N_13641,N_13729);
xor U13877 (N_13877,N_13641,N_13518);
nand U13878 (N_13878,N_13721,N_13556);
nand U13879 (N_13879,N_13622,N_13567);
xnor U13880 (N_13880,N_13553,N_13526);
xor U13881 (N_13881,N_13736,N_13598);
xor U13882 (N_13882,N_13539,N_13663);
nor U13883 (N_13883,N_13501,N_13664);
and U13884 (N_13884,N_13689,N_13600);
nor U13885 (N_13885,N_13555,N_13602);
and U13886 (N_13886,N_13611,N_13565);
nor U13887 (N_13887,N_13514,N_13596);
nand U13888 (N_13888,N_13607,N_13583);
or U13889 (N_13889,N_13646,N_13626);
nor U13890 (N_13890,N_13729,N_13606);
xnor U13891 (N_13891,N_13704,N_13576);
nand U13892 (N_13892,N_13602,N_13535);
or U13893 (N_13893,N_13608,N_13576);
xor U13894 (N_13894,N_13582,N_13669);
xnor U13895 (N_13895,N_13712,N_13619);
xor U13896 (N_13896,N_13528,N_13554);
or U13897 (N_13897,N_13560,N_13630);
and U13898 (N_13898,N_13508,N_13643);
nand U13899 (N_13899,N_13650,N_13702);
or U13900 (N_13900,N_13698,N_13661);
or U13901 (N_13901,N_13543,N_13544);
and U13902 (N_13902,N_13550,N_13537);
xnor U13903 (N_13903,N_13580,N_13538);
and U13904 (N_13904,N_13719,N_13560);
xnor U13905 (N_13905,N_13699,N_13728);
or U13906 (N_13906,N_13740,N_13717);
nand U13907 (N_13907,N_13518,N_13581);
xnor U13908 (N_13908,N_13656,N_13519);
nor U13909 (N_13909,N_13685,N_13515);
nor U13910 (N_13910,N_13538,N_13564);
or U13911 (N_13911,N_13697,N_13510);
and U13912 (N_13912,N_13590,N_13518);
or U13913 (N_13913,N_13591,N_13691);
nor U13914 (N_13914,N_13605,N_13505);
xnor U13915 (N_13915,N_13650,N_13528);
or U13916 (N_13916,N_13671,N_13636);
nand U13917 (N_13917,N_13716,N_13563);
nand U13918 (N_13918,N_13539,N_13638);
nor U13919 (N_13919,N_13740,N_13558);
or U13920 (N_13920,N_13749,N_13534);
nand U13921 (N_13921,N_13675,N_13506);
and U13922 (N_13922,N_13746,N_13612);
xor U13923 (N_13923,N_13609,N_13516);
or U13924 (N_13924,N_13710,N_13644);
nand U13925 (N_13925,N_13596,N_13537);
nand U13926 (N_13926,N_13712,N_13731);
and U13927 (N_13927,N_13542,N_13633);
nand U13928 (N_13928,N_13665,N_13660);
nor U13929 (N_13929,N_13515,N_13524);
and U13930 (N_13930,N_13648,N_13673);
nand U13931 (N_13931,N_13551,N_13570);
and U13932 (N_13932,N_13594,N_13590);
xnor U13933 (N_13933,N_13716,N_13598);
xor U13934 (N_13934,N_13669,N_13713);
or U13935 (N_13935,N_13613,N_13700);
xor U13936 (N_13936,N_13655,N_13512);
nand U13937 (N_13937,N_13654,N_13502);
xor U13938 (N_13938,N_13695,N_13616);
or U13939 (N_13939,N_13669,N_13717);
or U13940 (N_13940,N_13631,N_13712);
or U13941 (N_13941,N_13592,N_13683);
and U13942 (N_13942,N_13559,N_13503);
and U13943 (N_13943,N_13601,N_13695);
nor U13944 (N_13944,N_13582,N_13521);
or U13945 (N_13945,N_13541,N_13616);
nor U13946 (N_13946,N_13572,N_13696);
nor U13947 (N_13947,N_13688,N_13661);
nand U13948 (N_13948,N_13502,N_13535);
or U13949 (N_13949,N_13524,N_13658);
nor U13950 (N_13950,N_13613,N_13524);
and U13951 (N_13951,N_13557,N_13735);
nor U13952 (N_13952,N_13528,N_13713);
xnor U13953 (N_13953,N_13619,N_13531);
or U13954 (N_13954,N_13520,N_13610);
nor U13955 (N_13955,N_13535,N_13578);
nand U13956 (N_13956,N_13552,N_13598);
nand U13957 (N_13957,N_13508,N_13682);
or U13958 (N_13958,N_13742,N_13709);
nor U13959 (N_13959,N_13537,N_13643);
nand U13960 (N_13960,N_13516,N_13656);
and U13961 (N_13961,N_13548,N_13635);
nand U13962 (N_13962,N_13506,N_13688);
nand U13963 (N_13963,N_13550,N_13711);
or U13964 (N_13964,N_13524,N_13620);
xor U13965 (N_13965,N_13689,N_13660);
and U13966 (N_13966,N_13690,N_13686);
nand U13967 (N_13967,N_13593,N_13662);
nor U13968 (N_13968,N_13626,N_13669);
and U13969 (N_13969,N_13578,N_13635);
xor U13970 (N_13970,N_13738,N_13716);
nor U13971 (N_13971,N_13614,N_13588);
nand U13972 (N_13972,N_13610,N_13552);
xnor U13973 (N_13973,N_13664,N_13713);
nand U13974 (N_13974,N_13581,N_13668);
and U13975 (N_13975,N_13522,N_13734);
nand U13976 (N_13976,N_13597,N_13620);
nand U13977 (N_13977,N_13714,N_13522);
or U13978 (N_13978,N_13643,N_13676);
xor U13979 (N_13979,N_13529,N_13731);
and U13980 (N_13980,N_13716,N_13542);
nand U13981 (N_13981,N_13626,N_13676);
and U13982 (N_13982,N_13560,N_13638);
nor U13983 (N_13983,N_13623,N_13581);
nor U13984 (N_13984,N_13538,N_13634);
or U13985 (N_13985,N_13588,N_13656);
nand U13986 (N_13986,N_13524,N_13746);
xnor U13987 (N_13987,N_13541,N_13634);
xnor U13988 (N_13988,N_13739,N_13747);
and U13989 (N_13989,N_13695,N_13725);
nor U13990 (N_13990,N_13713,N_13674);
xnor U13991 (N_13991,N_13585,N_13674);
and U13992 (N_13992,N_13618,N_13685);
or U13993 (N_13993,N_13644,N_13568);
nand U13994 (N_13994,N_13620,N_13623);
nor U13995 (N_13995,N_13698,N_13532);
and U13996 (N_13996,N_13747,N_13574);
or U13997 (N_13997,N_13575,N_13678);
nand U13998 (N_13998,N_13513,N_13577);
and U13999 (N_13999,N_13648,N_13722);
and U14000 (N_14000,N_13856,N_13981);
nor U14001 (N_14001,N_13886,N_13927);
xor U14002 (N_14002,N_13782,N_13804);
nor U14003 (N_14003,N_13789,N_13817);
or U14004 (N_14004,N_13982,N_13956);
and U14005 (N_14005,N_13987,N_13903);
nor U14006 (N_14006,N_13858,N_13781);
nor U14007 (N_14007,N_13904,N_13831);
or U14008 (N_14008,N_13890,N_13780);
and U14009 (N_14009,N_13756,N_13821);
nand U14010 (N_14010,N_13928,N_13941);
nand U14011 (N_14011,N_13899,N_13964);
nand U14012 (N_14012,N_13971,N_13773);
nand U14013 (N_14013,N_13994,N_13888);
or U14014 (N_14014,N_13812,N_13960);
xnor U14015 (N_14015,N_13834,N_13753);
nor U14016 (N_14016,N_13957,N_13949);
xnor U14017 (N_14017,N_13998,N_13900);
and U14018 (N_14018,N_13792,N_13860);
or U14019 (N_14019,N_13879,N_13986);
or U14020 (N_14020,N_13922,N_13800);
nor U14021 (N_14021,N_13881,N_13865);
nor U14022 (N_14022,N_13952,N_13861);
nand U14023 (N_14023,N_13754,N_13823);
or U14024 (N_14024,N_13958,N_13912);
and U14025 (N_14025,N_13828,N_13791);
nand U14026 (N_14026,N_13947,N_13961);
nand U14027 (N_14027,N_13822,N_13778);
and U14028 (N_14028,N_13959,N_13850);
and U14029 (N_14029,N_13925,N_13917);
nor U14030 (N_14030,N_13783,N_13931);
xor U14031 (N_14031,N_13825,N_13776);
or U14032 (N_14032,N_13936,N_13852);
and U14033 (N_14033,N_13965,N_13762);
or U14034 (N_14034,N_13975,N_13833);
or U14035 (N_14035,N_13909,N_13761);
nor U14036 (N_14036,N_13871,N_13832);
or U14037 (N_14037,N_13955,N_13836);
nor U14038 (N_14038,N_13970,N_13851);
xnor U14039 (N_14039,N_13914,N_13877);
xnor U14040 (N_14040,N_13862,N_13884);
nor U14041 (N_14041,N_13784,N_13854);
nor U14042 (N_14042,N_13967,N_13802);
xor U14043 (N_14043,N_13777,N_13973);
or U14044 (N_14044,N_13905,N_13793);
xor U14045 (N_14045,N_13842,N_13990);
nand U14046 (N_14046,N_13966,N_13902);
and U14047 (N_14047,N_13924,N_13787);
or U14048 (N_14048,N_13840,N_13993);
nand U14049 (N_14049,N_13995,N_13807);
xor U14050 (N_14050,N_13979,N_13846);
xnor U14051 (N_14051,N_13989,N_13760);
xnor U14052 (N_14052,N_13953,N_13808);
nor U14053 (N_14053,N_13794,N_13894);
or U14054 (N_14054,N_13750,N_13863);
and U14055 (N_14055,N_13797,N_13878);
or U14056 (N_14056,N_13887,N_13870);
xnor U14057 (N_14057,N_13991,N_13882);
nor U14058 (N_14058,N_13873,N_13770);
xnor U14059 (N_14059,N_13942,N_13830);
and U14060 (N_14060,N_13765,N_13849);
nor U14061 (N_14061,N_13757,N_13795);
nor U14062 (N_14062,N_13885,N_13923);
xor U14063 (N_14063,N_13977,N_13997);
nand U14064 (N_14064,N_13940,N_13968);
nor U14065 (N_14065,N_13908,N_13768);
xor U14066 (N_14066,N_13813,N_13837);
or U14067 (N_14067,N_13875,N_13946);
or U14068 (N_14068,N_13751,N_13829);
nand U14069 (N_14069,N_13847,N_13932);
nand U14070 (N_14070,N_13896,N_13859);
and U14071 (N_14071,N_13866,N_13788);
and U14072 (N_14072,N_13857,N_13996);
nor U14073 (N_14073,N_13944,N_13818);
or U14074 (N_14074,N_13880,N_13868);
and U14075 (N_14075,N_13992,N_13867);
nand U14076 (N_14076,N_13926,N_13892);
nor U14077 (N_14077,N_13848,N_13939);
nand U14078 (N_14078,N_13816,N_13893);
and U14079 (N_14079,N_13938,N_13843);
nand U14080 (N_14080,N_13930,N_13937);
nor U14081 (N_14081,N_13916,N_13838);
xor U14082 (N_14082,N_13824,N_13948);
or U14083 (N_14083,N_13972,N_13820);
nand U14084 (N_14084,N_13911,N_13898);
or U14085 (N_14085,N_13872,N_13811);
or U14086 (N_14086,N_13920,N_13901);
nand U14087 (N_14087,N_13855,N_13771);
nor U14088 (N_14088,N_13988,N_13767);
nor U14089 (N_14089,N_13976,N_13889);
nand U14090 (N_14090,N_13853,N_13766);
nand U14091 (N_14091,N_13999,N_13951);
and U14092 (N_14092,N_13985,N_13984);
or U14093 (N_14093,N_13803,N_13906);
or U14094 (N_14094,N_13775,N_13798);
xnor U14095 (N_14095,N_13950,N_13796);
or U14096 (N_14096,N_13913,N_13839);
nor U14097 (N_14097,N_13769,N_13963);
xor U14098 (N_14098,N_13815,N_13758);
and U14099 (N_14099,N_13919,N_13819);
xnor U14100 (N_14100,N_13895,N_13845);
nor U14101 (N_14101,N_13772,N_13763);
or U14102 (N_14102,N_13826,N_13945);
nand U14103 (N_14103,N_13921,N_13910);
xnor U14104 (N_14104,N_13980,N_13810);
nor U14105 (N_14105,N_13790,N_13786);
and U14106 (N_14106,N_13799,N_13809);
nor U14107 (N_14107,N_13814,N_13915);
or U14108 (N_14108,N_13983,N_13907);
xnor U14109 (N_14109,N_13978,N_13954);
nor U14110 (N_14110,N_13943,N_13869);
xor U14111 (N_14111,N_13806,N_13805);
and U14112 (N_14112,N_13779,N_13874);
nand U14113 (N_14113,N_13935,N_13801);
xor U14114 (N_14114,N_13929,N_13755);
and U14115 (N_14115,N_13876,N_13962);
nand U14116 (N_14116,N_13764,N_13827);
nor U14117 (N_14117,N_13752,N_13774);
nand U14118 (N_14118,N_13841,N_13864);
and U14119 (N_14119,N_13891,N_13918);
xor U14120 (N_14120,N_13969,N_13974);
nor U14121 (N_14121,N_13759,N_13897);
xor U14122 (N_14122,N_13934,N_13835);
or U14123 (N_14123,N_13933,N_13883);
or U14124 (N_14124,N_13844,N_13785);
and U14125 (N_14125,N_13777,N_13912);
xor U14126 (N_14126,N_13915,N_13902);
and U14127 (N_14127,N_13764,N_13979);
nand U14128 (N_14128,N_13891,N_13781);
xnor U14129 (N_14129,N_13813,N_13909);
nand U14130 (N_14130,N_13892,N_13893);
xor U14131 (N_14131,N_13809,N_13858);
or U14132 (N_14132,N_13856,N_13912);
and U14133 (N_14133,N_13776,N_13878);
or U14134 (N_14134,N_13906,N_13959);
and U14135 (N_14135,N_13994,N_13995);
nor U14136 (N_14136,N_13806,N_13961);
nand U14137 (N_14137,N_13872,N_13806);
xnor U14138 (N_14138,N_13952,N_13776);
nand U14139 (N_14139,N_13853,N_13918);
nor U14140 (N_14140,N_13899,N_13854);
nor U14141 (N_14141,N_13800,N_13826);
and U14142 (N_14142,N_13941,N_13764);
nor U14143 (N_14143,N_13817,N_13947);
nand U14144 (N_14144,N_13988,N_13832);
nor U14145 (N_14145,N_13869,N_13933);
nand U14146 (N_14146,N_13792,N_13865);
or U14147 (N_14147,N_13953,N_13979);
nand U14148 (N_14148,N_13885,N_13848);
nor U14149 (N_14149,N_13803,N_13994);
or U14150 (N_14150,N_13965,N_13992);
and U14151 (N_14151,N_13990,N_13963);
and U14152 (N_14152,N_13925,N_13774);
xnor U14153 (N_14153,N_13898,N_13815);
nand U14154 (N_14154,N_13937,N_13835);
or U14155 (N_14155,N_13935,N_13866);
and U14156 (N_14156,N_13754,N_13957);
nor U14157 (N_14157,N_13852,N_13903);
nor U14158 (N_14158,N_13775,N_13887);
and U14159 (N_14159,N_13964,N_13786);
xnor U14160 (N_14160,N_13861,N_13976);
or U14161 (N_14161,N_13952,N_13830);
xor U14162 (N_14162,N_13968,N_13894);
nand U14163 (N_14163,N_13848,N_13824);
or U14164 (N_14164,N_13990,N_13852);
nand U14165 (N_14165,N_13756,N_13797);
xnor U14166 (N_14166,N_13800,N_13854);
nor U14167 (N_14167,N_13894,N_13829);
nand U14168 (N_14168,N_13940,N_13800);
nand U14169 (N_14169,N_13817,N_13860);
xnor U14170 (N_14170,N_13986,N_13790);
or U14171 (N_14171,N_13974,N_13906);
nor U14172 (N_14172,N_13920,N_13762);
xnor U14173 (N_14173,N_13824,N_13840);
or U14174 (N_14174,N_13910,N_13887);
or U14175 (N_14175,N_13768,N_13867);
nand U14176 (N_14176,N_13994,N_13999);
nand U14177 (N_14177,N_13922,N_13896);
and U14178 (N_14178,N_13995,N_13915);
or U14179 (N_14179,N_13929,N_13766);
nor U14180 (N_14180,N_13762,N_13808);
or U14181 (N_14181,N_13824,N_13826);
xnor U14182 (N_14182,N_13864,N_13839);
and U14183 (N_14183,N_13909,N_13964);
nand U14184 (N_14184,N_13912,N_13875);
and U14185 (N_14185,N_13906,N_13915);
and U14186 (N_14186,N_13778,N_13951);
xor U14187 (N_14187,N_13866,N_13923);
nor U14188 (N_14188,N_13998,N_13828);
nand U14189 (N_14189,N_13924,N_13969);
and U14190 (N_14190,N_13977,N_13940);
or U14191 (N_14191,N_13965,N_13932);
or U14192 (N_14192,N_13881,N_13783);
and U14193 (N_14193,N_13879,N_13975);
or U14194 (N_14194,N_13812,N_13931);
nor U14195 (N_14195,N_13906,N_13935);
or U14196 (N_14196,N_13897,N_13980);
and U14197 (N_14197,N_13912,N_13955);
nand U14198 (N_14198,N_13825,N_13920);
or U14199 (N_14199,N_13971,N_13758);
xor U14200 (N_14200,N_13819,N_13824);
and U14201 (N_14201,N_13911,N_13917);
xor U14202 (N_14202,N_13931,N_13909);
xnor U14203 (N_14203,N_13919,N_13871);
xnor U14204 (N_14204,N_13782,N_13790);
and U14205 (N_14205,N_13796,N_13822);
or U14206 (N_14206,N_13880,N_13923);
and U14207 (N_14207,N_13959,N_13813);
nand U14208 (N_14208,N_13812,N_13822);
nor U14209 (N_14209,N_13811,N_13788);
nand U14210 (N_14210,N_13805,N_13907);
nand U14211 (N_14211,N_13796,N_13976);
xnor U14212 (N_14212,N_13759,N_13877);
nand U14213 (N_14213,N_13773,N_13801);
or U14214 (N_14214,N_13961,N_13841);
xor U14215 (N_14215,N_13780,N_13790);
nand U14216 (N_14216,N_13941,N_13874);
nand U14217 (N_14217,N_13904,N_13766);
and U14218 (N_14218,N_13766,N_13991);
nor U14219 (N_14219,N_13868,N_13823);
xor U14220 (N_14220,N_13898,N_13984);
and U14221 (N_14221,N_13931,N_13920);
nand U14222 (N_14222,N_13772,N_13784);
nor U14223 (N_14223,N_13988,N_13940);
and U14224 (N_14224,N_13792,N_13958);
or U14225 (N_14225,N_13990,N_13824);
and U14226 (N_14226,N_13874,N_13824);
or U14227 (N_14227,N_13920,N_13783);
nor U14228 (N_14228,N_13859,N_13903);
or U14229 (N_14229,N_13911,N_13899);
or U14230 (N_14230,N_13989,N_13759);
xnor U14231 (N_14231,N_13882,N_13778);
nor U14232 (N_14232,N_13989,N_13833);
nor U14233 (N_14233,N_13887,N_13919);
nand U14234 (N_14234,N_13764,N_13777);
and U14235 (N_14235,N_13993,N_13838);
and U14236 (N_14236,N_13782,N_13846);
and U14237 (N_14237,N_13830,N_13757);
xor U14238 (N_14238,N_13902,N_13835);
nor U14239 (N_14239,N_13969,N_13868);
nor U14240 (N_14240,N_13939,N_13794);
xor U14241 (N_14241,N_13998,N_13947);
nand U14242 (N_14242,N_13773,N_13777);
xnor U14243 (N_14243,N_13973,N_13946);
xor U14244 (N_14244,N_13925,N_13967);
or U14245 (N_14245,N_13874,N_13983);
xor U14246 (N_14246,N_13952,N_13918);
nor U14247 (N_14247,N_13883,N_13911);
nor U14248 (N_14248,N_13922,N_13936);
or U14249 (N_14249,N_13941,N_13905);
nor U14250 (N_14250,N_14089,N_14215);
or U14251 (N_14251,N_14153,N_14232);
xnor U14252 (N_14252,N_14130,N_14131);
xor U14253 (N_14253,N_14043,N_14228);
and U14254 (N_14254,N_14021,N_14243);
xor U14255 (N_14255,N_14079,N_14219);
and U14256 (N_14256,N_14247,N_14206);
or U14257 (N_14257,N_14036,N_14155);
nor U14258 (N_14258,N_14193,N_14007);
nand U14259 (N_14259,N_14248,N_14004);
or U14260 (N_14260,N_14188,N_14109);
or U14261 (N_14261,N_14046,N_14172);
nor U14262 (N_14262,N_14108,N_14121);
nand U14263 (N_14263,N_14018,N_14017);
nand U14264 (N_14264,N_14047,N_14045);
nor U14265 (N_14265,N_14071,N_14103);
xnor U14266 (N_14266,N_14239,N_14015);
or U14267 (N_14267,N_14023,N_14191);
nor U14268 (N_14268,N_14222,N_14008);
xnor U14269 (N_14269,N_14226,N_14100);
or U14270 (N_14270,N_14236,N_14106);
and U14271 (N_14271,N_14126,N_14068);
or U14272 (N_14272,N_14218,N_14069);
xor U14273 (N_14273,N_14177,N_14167);
or U14274 (N_14274,N_14154,N_14245);
xnor U14275 (N_14275,N_14065,N_14234);
nor U14276 (N_14276,N_14088,N_14115);
nor U14277 (N_14277,N_14037,N_14164);
nand U14278 (N_14278,N_14011,N_14180);
or U14279 (N_14279,N_14000,N_14129);
or U14280 (N_14280,N_14022,N_14246);
and U14281 (N_14281,N_14210,N_14159);
xor U14282 (N_14282,N_14146,N_14102);
nor U14283 (N_14283,N_14173,N_14050);
nand U14284 (N_14284,N_14145,N_14211);
or U14285 (N_14285,N_14196,N_14113);
nand U14286 (N_14286,N_14151,N_14161);
xor U14287 (N_14287,N_14052,N_14162);
xnor U14288 (N_14288,N_14158,N_14064);
nor U14289 (N_14289,N_14181,N_14095);
nand U14290 (N_14290,N_14117,N_14214);
or U14291 (N_14291,N_14074,N_14090);
or U14292 (N_14292,N_14168,N_14148);
or U14293 (N_14293,N_14066,N_14092);
xor U14294 (N_14294,N_14012,N_14224);
xor U14295 (N_14295,N_14030,N_14152);
nor U14296 (N_14296,N_14216,N_14205);
xnor U14297 (N_14297,N_14078,N_14237);
xnor U14298 (N_14298,N_14060,N_14054);
or U14299 (N_14299,N_14203,N_14067);
or U14300 (N_14300,N_14122,N_14133);
and U14301 (N_14301,N_14024,N_14002);
or U14302 (N_14302,N_14099,N_14005);
nor U14303 (N_14303,N_14166,N_14040);
or U14304 (N_14304,N_14141,N_14231);
xor U14305 (N_14305,N_14233,N_14116);
xnor U14306 (N_14306,N_14031,N_14199);
nor U14307 (N_14307,N_14170,N_14213);
xor U14308 (N_14308,N_14077,N_14132);
xnor U14309 (N_14309,N_14020,N_14128);
nor U14310 (N_14310,N_14042,N_14197);
and U14311 (N_14311,N_14134,N_14016);
xnor U14312 (N_14312,N_14013,N_14186);
nand U14313 (N_14313,N_14104,N_14096);
nor U14314 (N_14314,N_14073,N_14220);
nand U14315 (N_14315,N_14144,N_14194);
or U14316 (N_14316,N_14135,N_14192);
nor U14317 (N_14317,N_14072,N_14178);
or U14318 (N_14318,N_14217,N_14125);
xor U14319 (N_14319,N_14059,N_14080);
nand U14320 (N_14320,N_14185,N_14183);
xnor U14321 (N_14321,N_14142,N_14204);
or U14322 (N_14322,N_14070,N_14003);
xor U14323 (N_14323,N_14179,N_14034);
and U14324 (N_14324,N_14147,N_14190);
nor U14325 (N_14325,N_14163,N_14001);
nand U14326 (N_14326,N_14086,N_14051);
nand U14327 (N_14327,N_14063,N_14111);
nor U14328 (N_14328,N_14143,N_14087);
and U14329 (N_14329,N_14014,N_14165);
nor U14330 (N_14330,N_14249,N_14238);
nand U14331 (N_14331,N_14140,N_14057);
nand U14332 (N_14332,N_14082,N_14019);
xnor U14333 (N_14333,N_14184,N_14058);
and U14334 (N_14334,N_14105,N_14160);
xnor U14335 (N_14335,N_14195,N_14028);
nand U14336 (N_14336,N_14171,N_14235);
and U14337 (N_14337,N_14107,N_14094);
or U14338 (N_14338,N_14061,N_14201);
xnor U14339 (N_14339,N_14027,N_14029);
and U14340 (N_14340,N_14055,N_14174);
nand U14341 (N_14341,N_14053,N_14229);
nand U14342 (N_14342,N_14032,N_14048);
xnor U14343 (N_14343,N_14150,N_14056);
xnor U14344 (N_14344,N_14025,N_14227);
nand U14345 (N_14345,N_14200,N_14049);
nand U14346 (N_14346,N_14026,N_14081);
nor U14347 (N_14347,N_14176,N_14223);
or U14348 (N_14348,N_14212,N_14118);
nor U14349 (N_14349,N_14189,N_14207);
or U14350 (N_14350,N_14169,N_14038);
and U14351 (N_14351,N_14009,N_14242);
xnor U14352 (N_14352,N_14230,N_14138);
nand U14353 (N_14353,N_14208,N_14084);
or U14354 (N_14354,N_14137,N_14225);
nor U14355 (N_14355,N_14175,N_14098);
xor U14356 (N_14356,N_14119,N_14075);
and U14357 (N_14357,N_14209,N_14123);
and U14358 (N_14358,N_14033,N_14241);
and U14359 (N_14359,N_14006,N_14091);
xnor U14360 (N_14360,N_14101,N_14062);
or U14361 (N_14361,N_14083,N_14187);
or U14362 (N_14362,N_14112,N_14085);
nor U14363 (N_14363,N_14127,N_14110);
and U14364 (N_14364,N_14157,N_14139);
nand U14365 (N_14365,N_14035,N_14149);
or U14366 (N_14366,N_14041,N_14156);
xnor U14367 (N_14367,N_14244,N_14010);
nor U14368 (N_14368,N_14182,N_14240);
and U14369 (N_14369,N_14039,N_14221);
or U14370 (N_14370,N_14097,N_14124);
nand U14371 (N_14371,N_14076,N_14136);
or U14372 (N_14372,N_14120,N_14044);
and U14373 (N_14373,N_14198,N_14114);
or U14374 (N_14374,N_14202,N_14093);
nand U14375 (N_14375,N_14069,N_14015);
nor U14376 (N_14376,N_14249,N_14109);
and U14377 (N_14377,N_14020,N_14040);
or U14378 (N_14378,N_14233,N_14007);
nor U14379 (N_14379,N_14132,N_14230);
xnor U14380 (N_14380,N_14098,N_14168);
xnor U14381 (N_14381,N_14205,N_14238);
or U14382 (N_14382,N_14147,N_14065);
nor U14383 (N_14383,N_14089,N_14180);
or U14384 (N_14384,N_14129,N_14221);
nor U14385 (N_14385,N_14054,N_14206);
nor U14386 (N_14386,N_14222,N_14111);
nor U14387 (N_14387,N_14006,N_14145);
nand U14388 (N_14388,N_14048,N_14121);
nor U14389 (N_14389,N_14123,N_14079);
or U14390 (N_14390,N_14174,N_14212);
nand U14391 (N_14391,N_14235,N_14054);
nand U14392 (N_14392,N_14061,N_14234);
and U14393 (N_14393,N_14043,N_14160);
xor U14394 (N_14394,N_14082,N_14079);
xor U14395 (N_14395,N_14044,N_14236);
xnor U14396 (N_14396,N_14122,N_14227);
xor U14397 (N_14397,N_14080,N_14087);
xor U14398 (N_14398,N_14217,N_14157);
nand U14399 (N_14399,N_14227,N_14207);
and U14400 (N_14400,N_14158,N_14187);
and U14401 (N_14401,N_14054,N_14027);
or U14402 (N_14402,N_14131,N_14139);
nand U14403 (N_14403,N_14065,N_14103);
xnor U14404 (N_14404,N_14201,N_14127);
and U14405 (N_14405,N_14059,N_14187);
nand U14406 (N_14406,N_14132,N_14043);
nor U14407 (N_14407,N_14175,N_14066);
nor U14408 (N_14408,N_14105,N_14141);
or U14409 (N_14409,N_14224,N_14055);
xnor U14410 (N_14410,N_14174,N_14023);
xor U14411 (N_14411,N_14213,N_14220);
nand U14412 (N_14412,N_14078,N_14094);
or U14413 (N_14413,N_14179,N_14215);
or U14414 (N_14414,N_14077,N_14178);
nand U14415 (N_14415,N_14114,N_14236);
nand U14416 (N_14416,N_14127,N_14208);
xor U14417 (N_14417,N_14134,N_14169);
nand U14418 (N_14418,N_14196,N_14044);
and U14419 (N_14419,N_14165,N_14069);
nor U14420 (N_14420,N_14213,N_14112);
nor U14421 (N_14421,N_14169,N_14063);
or U14422 (N_14422,N_14070,N_14118);
or U14423 (N_14423,N_14076,N_14131);
nand U14424 (N_14424,N_14147,N_14066);
nor U14425 (N_14425,N_14246,N_14146);
xnor U14426 (N_14426,N_14244,N_14236);
or U14427 (N_14427,N_14134,N_14115);
xor U14428 (N_14428,N_14183,N_14237);
nand U14429 (N_14429,N_14088,N_14075);
and U14430 (N_14430,N_14005,N_14167);
nand U14431 (N_14431,N_14249,N_14154);
and U14432 (N_14432,N_14172,N_14237);
nand U14433 (N_14433,N_14039,N_14203);
xnor U14434 (N_14434,N_14157,N_14123);
or U14435 (N_14435,N_14070,N_14221);
nand U14436 (N_14436,N_14021,N_14029);
nand U14437 (N_14437,N_14009,N_14116);
and U14438 (N_14438,N_14122,N_14027);
and U14439 (N_14439,N_14013,N_14178);
nor U14440 (N_14440,N_14124,N_14047);
nor U14441 (N_14441,N_14127,N_14042);
nor U14442 (N_14442,N_14246,N_14072);
xor U14443 (N_14443,N_14093,N_14105);
or U14444 (N_14444,N_14092,N_14117);
and U14445 (N_14445,N_14090,N_14247);
nand U14446 (N_14446,N_14188,N_14036);
and U14447 (N_14447,N_14200,N_14036);
nor U14448 (N_14448,N_14120,N_14215);
nor U14449 (N_14449,N_14231,N_14015);
or U14450 (N_14450,N_14011,N_14179);
and U14451 (N_14451,N_14003,N_14010);
and U14452 (N_14452,N_14137,N_14106);
xnor U14453 (N_14453,N_14096,N_14064);
nor U14454 (N_14454,N_14189,N_14072);
nor U14455 (N_14455,N_14216,N_14032);
and U14456 (N_14456,N_14139,N_14146);
or U14457 (N_14457,N_14223,N_14047);
or U14458 (N_14458,N_14132,N_14183);
xor U14459 (N_14459,N_14199,N_14125);
and U14460 (N_14460,N_14072,N_14127);
and U14461 (N_14461,N_14244,N_14019);
and U14462 (N_14462,N_14158,N_14045);
xor U14463 (N_14463,N_14096,N_14050);
nand U14464 (N_14464,N_14176,N_14045);
xnor U14465 (N_14465,N_14227,N_14156);
nand U14466 (N_14466,N_14001,N_14008);
or U14467 (N_14467,N_14247,N_14201);
or U14468 (N_14468,N_14037,N_14097);
nand U14469 (N_14469,N_14147,N_14021);
or U14470 (N_14470,N_14248,N_14113);
or U14471 (N_14471,N_14199,N_14059);
nor U14472 (N_14472,N_14187,N_14065);
or U14473 (N_14473,N_14081,N_14225);
nor U14474 (N_14474,N_14020,N_14071);
and U14475 (N_14475,N_14216,N_14035);
nor U14476 (N_14476,N_14195,N_14220);
nor U14477 (N_14477,N_14238,N_14184);
or U14478 (N_14478,N_14003,N_14124);
xor U14479 (N_14479,N_14210,N_14071);
xor U14480 (N_14480,N_14142,N_14169);
nor U14481 (N_14481,N_14240,N_14090);
nor U14482 (N_14482,N_14057,N_14218);
or U14483 (N_14483,N_14214,N_14249);
xor U14484 (N_14484,N_14076,N_14086);
and U14485 (N_14485,N_14038,N_14235);
or U14486 (N_14486,N_14240,N_14077);
and U14487 (N_14487,N_14161,N_14157);
nor U14488 (N_14488,N_14071,N_14234);
or U14489 (N_14489,N_14154,N_14091);
nor U14490 (N_14490,N_14023,N_14086);
nor U14491 (N_14491,N_14210,N_14244);
nand U14492 (N_14492,N_14228,N_14021);
nand U14493 (N_14493,N_14006,N_14018);
and U14494 (N_14494,N_14192,N_14137);
nor U14495 (N_14495,N_14198,N_14192);
nor U14496 (N_14496,N_14140,N_14183);
and U14497 (N_14497,N_14203,N_14180);
nor U14498 (N_14498,N_14195,N_14119);
nand U14499 (N_14499,N_14007,N_14211);
xnor U14500 (N_14500,N_14487,N_14473);
and U14501 (N_14501,N_14355,N_14392);
nand U14502 (N_14502,N_14422,N_14388);
xnor U14503 (N_14503,N_14403,N_14409);
xnor U14504 (N_14504,N_14449,N_14333);
and U14505 (N_14505,N_14306,N_14380);
and U14506 (N_14506,N_14457,N_14419);
or U14507 (N_14507,N_14300,N_14498);
nand U14508 (N_14508,N_14485,N_14253);
or U14509 (N_14509,N_14413,N_14338);
nand U14510 (N_14510,N_14254,N_14384);
nor U14511 (N_14511,N_14421,N_14370);
or U14512 (N_14512,N_14321,N_14359);
or U14513 (N_14513,N_14378,N_14488);
xnor U14514 (N_14514,N_14381,N_14279);
nand U14515 (N_14515,N_14336,N_14373);
or U14516 (N_14516,N_14299,N_14434);
xnor U14517 (N_14517,N_14453,N_14448);
or U14518 (N_14518,N_14353,N_14414);
and U14519 (N_14519,N_14286,N_14343);
xnor U14520 (N_14520,N_14447,N_14404);
nand U14521 (N_14521,N_14314,N_14364);
xor U14522 (N_14522,N_14301,N_14346);
nand U14523 (N_14523,N_14436,N_14400);
and U14524 (N_14524,N_14397,N_14308);
and U14525 (N_14525,N_14461,N_14455);
nand U14526 (N_14526,N_14291,N_14426);
nand U14527 (N_14527,N_14357,N_14389);
nand U14528 (N_14528,N_14264,N_14270);
nor U14529 (N_14529,N_14294,N_14372);
nand U14530 (N_14530,N_14425,N_14385);
nor U14531 (N_14531,N_14307,N_14444);
xnor U14532 (N_14532,N_14273,N_14474);
or U14533 (N_14533,N_14258,N_14324);
xnor U14534 (N_14534,N_14458,N_14491);
and U14535 (N_14535,N_14399,N_14496);
and U14536 (N_14536,N_14340,N_14477);
nand U14537 (N_14537,N_14309,N_14433);
or U14538 (N_14538,N_14467,N_14313);
nor U14539 (N_14539,N_14437,N_14280);
and U14540 (N_14540,N_14420,N_14416);
nor U14541 (N_14541,N_14328,N_14311);
or U14542 (N_14542,N_14302,N_14315);
or U14543 (N_14543,N_14483,N_14395);
xnor U14544 (N_14544,N_14350,N_14326);
or U14545 (N_14545,N_14450,N_14263);
and U14546 (N_14546,N_14495,N_14452);
or U14547 (N_14547,N_14480,N_14482);
nor U14548 (N_14548,N_14466,N_14494);
xor U14549 (N_14549,N_14289,N_14362);
nor U14550 (N_14550,N_14470,N_14354);
or U14551 (N_14551,N_14337,N_14440);
and U14552 (N_14552,N_14410,N_14391);
xnor U14553 (N_14553,N_14316,N_14411);
and U14554 (N_14554,N_14429,N_14464);
and U14555 (N_14555,N_14435,N_14298);
and U14556 (N_14556,N_14481,N_14278);
nor U14557 (N_14557,N_14405,N_14342);
and U14558 (N_14558,N_14454,N_14261);
and U14559 (N_14559,N_14369,N_14292);
nor U14560 (N_14560,N_14438,N_14368);
and U14561 (N_14561,N_14347,N_14323);
or U14562 (N_14562,N_14250,N_14281);
nor U14563 (N_14563,N_14296,N_14351);
nor U14564 (N_14564,N_14257,N_14352);
nor U14565 (N_14565,N_14265,N_14382);
and U14566 (N_14566,N_14327,N_14312);
nor U14567 (N_14567,N_14423,N_14325);
nor U14568 (N_14568,N_14430,N_14432);
and U14569 (N_14569,N_14360,N_14462);
and U14570 (N_14570,N_14304,N_14418);
nor U14571 (N_14571,N_14365,N_14428);
xor U14572 (N_14572,N_14318,N_14492);
or U14573 (N_14573,N_14406,N_14468);
or U14574 (N_14574,N_14376,N_14417);
and U14575 (N_14575,N_14377,N_14431);
and U14576 (N_14576,N_14288,N_14387);
and U14577 (N_14577,N_14490,N_14374);
and U14578 (N_14578,N_14489,N_14478);
xnor U14579 (N_14579,N_14259,N_14402);
or U14580 (N_14580,N_14275,N_14442);
nand U14581 (N_14581,N_14460,N_14266);
nor U14582 (N_14582,N_14272,N_14331);
nor U14583 (N_14583,N_14441,N_14349);
nor U14584 (N_14584,N_14356,N_14484);
xor U14585 (N_14585,N_14335,N_14366);
nand U14586 (N_14586,N_14295,N_14398);
nand U14587 (N_14587,N_14251,N_14396);
or U14588 (N_14588,N_14443,N_14363);
or U14589 (N_14589,N_14297,N_14394);
and U14590 (N_14590,N_14282,N_14329);
xor U14591 (N_14591,N_14317,N_14290);
xor U14592 (N_14592,N_14320,N_14322);
or U14593 (N_14593,N_14277,N_14268);
nor U14594 (N_14594,N_14285,N_14367);
xnor U14595 (N_14595,N_14439,N_14472);
or U14596 (N_14596,N_14479,N_14358);
xor U14597 (N_14597,N_14471,N_14283);
nand U14598 (N_14598,N_14424,N_14255);
and U14599 (N_14599,N_14345,N_14319);
xnor U14600 (N_14600,N_14341,N_14256);
nand U14601 (N_14601,N_14260,N_14390);
or U14602 (N_14602,N_14348,N_14475);
xnor U14603 (N_14603,N_14493,N_14284);
nor U14604 (N_14604,N_14271,N_14386);
xnor U14605 (N_14605,N_14427,N_14371);
and U14606 (N_14606,N_14446,N_14303);
xor U14607 (N_14607,N_14252,N_14407);
nand U14608 (N_14608,N_14456,N_14274);
and U14609 (N_14609,N_14465,N_14332);
or U14610 (N_14610,N_14344,N_14401);
or U14611 (N_14611,N_14334,N_14361);
or U14612 (N_14612,N_14379,N_14486);
nor U14613 (N_14613,N_14305,N_14408);
and U14614 (N_14614,N_14287,N_14476);
nor U14615 (N_14615,N_14393,N_14262);
nand U14616 (N_14616,N_14497,N_14499);
and U14617 (N_14617,N_14269,N_14463);
or U14618 (N_14618,N_14276,N_14330);
and U14619 (N_14619,N_14445,N_14412);
xnor U14620 (N_14620,N_14469,N_14375);
and U14621 (N_14621,N_14451,N_14459);
or U14622 (N_14622,N_14293,N_14339);
and U14623 (N_14623,N_14267,N_14383);
xor U14624 (N_14624,N_14310,N_14415);
nand U14625 (N_14625,N_14307,N_14470);
and U14626 (N_14626,N_14280,N_14274);
xor U14627 (N_14627,N_14315,N_14329);
nand U14628 (N_14628,N_14372,N_14492);
nand U14629 (N_14629,N_14268,N_14318);
xor U14630 (N_14630,N_14355,N_14283);
nor U14631 (N_14631,N_14296,N_14377);
and U14632 (N_14632,N_14455,N_14446);
nand U14633 (N_14633,N_14250,N_14450);
xor U14634 (N_14634,N_14468,N_14422);
or U14635 (N_14635,N_14316,N_14385);
nand U14636 (N_14636,N_14372,N_14400);
and U14637 (N_14637,N_14334,N_14258);
nand U14638 (N_14638,N_14476,N_14405);
nor U14639 (N_14639,N_14321,N_14361);
or U14640 (N_14640,N_14256,N_14336);
nand U14641 (N_14641,N_14477,N_14490);
nor U14642 (N_14642,N_14253,N_14333);
xnor U14643 (N_14643,N_14371,N_14265);
or U14644 (N_14644,N_14414,N_14423);
nor U14645 (N_14645,N_14278,N_14469);
nor U14646 (N_14646,N_14295,N_14336);
xnor U14647 (N_14647,N_14402,N_14420);
nand U14648 (N_14648,N_14336,N_14429);
nand U14649 (N_14649,N_14286,N_14419);
xor U14650 (N_14650,N_14330,N_14490);
and U14651 (N_14651,N_14251,N_14279);
nand U14652 (N_14652,N_14279,N_14412);
nor U14653 (N_14653,N_14341,N_14321);
and U14654 (N_14654,N_14334,N_14358);
xnor U14655 (N_14655,N_14288,N_14276);
nor U14656 (N_14656,N_14479,N_14447);
or U14657 (N_14657,N_14471,N_14277);
nor U14658 (N_14658,N_14302,N_14415);
nand U14659 (N_14659,N_14490,N_14434);
and U14660 (N_14660,N_14385,N_14312);
xnor U14661 (N_14661,N_14381,N_14457);
or U14662 (N_14662,N_14282,N_14430);
or U14663 (N_14663,N_14355,N_14386);
xnor U14664 (N_14664,N_14305,N_14389);
xor U14665 (N_14665,N_14265,N_14256);
and U14666 (N_14666,N_14254,N_14478);
nor U14667 (N_14667,N_14418,N_14400);
and U14668 (N_14668,N_14383,N_14295);
nand U14669 (N_14669,N_14406,N_14301);
and U14670 (N_14670,N_14355,N_14347);
xnor U14671 (N_14671,N_14320,N_14318);
and U14672 (N_14672,N_14420,N_14320);
nand U14673 (N_14673,N_14344,N_14394);
and U14674 (N_14674,N_14353,N_14371);
and U14675 (N_14675,N_14380,N_14360);
and U14676 (N_14676,N_14303,N_14388);
nor U14677 (N_14677,N_14379,N_14496);
or U14678 (N_14678,N_14357,N_14358);
xor U14679 (N_14679,N_14480,N_14352);
or U14680 (N_14680,N_14461,N_14347);
and U14681 (N_14681,N_14417,N_14390);
xnor U14682 (N_14682,N_14262,N_14412);
nor U14683 (N_14683,N_14363,N_14412);
xor U14684 (N_14684,N_14456,N_14284);
nand U14685 (N_14685,N_14444,N_14284);
nand U14686 (N_14686,N_14445,N_14443);
xnor U14687 (N_14687,N_14352,N_14371);
or U14688 (N_14688,N_14354,N_14293);
nor U14689 (N_14689,N_14349,N_14315);
and U14690 (N_14690,N_14451,N_14303);
and U14691 (N_14691,N_14271,N_14480);
xnor U14692 (N_14692,N_14393,N_14480);
and U14693 (N_14693,N_14347,N_14338);
and U14694 (N_14694,N_14342,N_14307);
xnor U14695 (N_14695,N_14271,N_14461);
xnor U14696 (N_14696,N_14350,N_14261);
and U14697 (N_14697,N_14389,N_14283);
or U14698 (N_14698,N_14365,N_14357);
and U14699 (N_14699,N_14284,N_14315);
or U14700 (N_14700,N_14314,N_14403);
nor U14701 (N_14701,N_14267,N_14435);
and U14702 (N_14702,N_14489,N_14441);
nor U14703 (N_14703,N_14419,N_14384);
xor U14704 (N_14704,N_14267,N_14449);
and U14705 (N_14705,N_14472,N_14481);
nand U14706 (N_14706,N_14252,N_14415);
nor U14707 (N_14707,N_14342,N_14326);
or U14708 (N_14708,N_14368,N_14381);
nand U14709 (N_14709,N_14268,N_14322);
xor U14710 (N_14710,N_14406,N_14275);
or U14711 (N_14711,N_14385,N_14309);
nor U14712 (N_14712,N_14284,N_14265);
or U14713 (N_14713,N_14453,N_14470);
nand U14714 (N_14714,N_14316,N_14430);
and U14715 (N_14715,N_14469,N_14258);
nand U14716 (N_14716,N_14260,N_14476);
xor U14717 (N_14717,N_14406,N_14325);
and U14718 (N_14718,N_14493,N_14426);
nor U14719 (N_14719,N_14327,N_14406);
nor U14720 (N_14720,N_14458,N_14420);
nand U14721 (N_14721,N_14315,N_14303);
nand U14722 (N_14722,N_14453,N_14258);
and U14723 (N_14723,N_14370,N_14486);
nor U14724 (N_14724,N_14258,N_14302);
and U14725 (N_14725,N_14255,N_14459);
nand U14726 (N_14726,N_14430,N_14322);
nand U14727 (N_14727,N_14322,N_14284);
xor U14728 (N_14728,N_14308,N_14467);
xor U14729 (N_14729,N_14297,N_14469);
and U14730 (N_14730,N_14275,N_14293);
and U14731 (N_14731,N_14418,N_14362);
nor U14732 (N_14732,N_14466,N_14450);
or U14733 (N_14733,N_14392,N_14484);
nor U14734 (N_14734,N_14480,N_14301);
or U14735 (N_14735,N_14278,N_14316);
xnor U14736 (N_14736,N_14427,N_14375);
or U14737 (N_14737,N_14496,N_14483);
nand U14738 (N_14738,N_14399,N_14278);
and U14739 (N_14739,N_14274,N_14296);
xnor U14740 (N_14740,N_14377,N_14438);
or U14741 (N_14741,N_14484,N_14480);
and U14742 (N_14742,N_14360,N_14252);
nand U14743 (N_14743,N_14364,N_14312);
and U14744 (N_14744,N_14483,N_14374);
xor U14745 (N_14745,N_14375,N_14277);
nor U14746 (N_14746,N_14341,N_14311);
and U14747 (N_14747,N_14433,N_14419);
nor U14748 (N_14748,N_14343,N_14482);
and U14749 (N_14749,N_14298,N_14470);
nand U14750 (N_14750,N_14571,N_14662);
and U14751 (N_14751,N_14732,N_14536);
and U14752 (N_14752,N_14739,N_14721);
nor U14753 (N_14753,N_14741,N_14592);
and U14754 (N_14754,N_14646,N_14747);
or U14755 (N_14755,N_14688,N_14595);
and U14756 (N_14756,N_14645,N_14722);
or U14757 (N_14757,N_14594,N_14587);
xnor U14758 (N_14758,N_14748,N_14535);
nor U14759 (N_14759,N_14672,N_14541);
or U14760 (N_14760,N_14519,N_14548);
xor U14761 (N_14761,N_14614,N_14681);
or U14762 (N_14762,N_14575,N_14708);
nor U14763 (N_14763,N_14635,N_14532);
and U14764 (N_14764,N_14524,N_14656);
or U14765 (N_14765,N_14690,N_14619);
xor U14766 (N_14766,N_14648,N_14731);
nand U14767 (N_14767,N_14627,N_14668);
nand U14768 (N_14768,N_14559,N_14572);
nor U14769 (N_14769,N_14704,N_14523);
or U14770 (N_14770,N_14637,N_14634);
and U14771 (N_14771,N_14584,N_14706);
and U14772 (N_14772,N_14736,N_14604);
nor U14773 (N_14773,N_14629,N_14724);
or U14774 (N_14774,N_14566,N_14598);
nand U14775 (N_14775,N_14676,N_14577);
nand U14776 (N_14776,N_14581,N_14638);
or U14777 (N_14777,N_14539,N_14544);
nor U14778 (N_14778,N_14625,N_14679);
or U14779 (N_14779,N_14596,N_14683);
nand U14780 (N_14780,N_14710,N_14616);
xnor U14781 (N_14781,N_14583,N_14685);
xnor U14782 (N_14782,N_14602,N_14609);
nor U14783 (N_14783,N_14529,N_14699);
xor U14784 (N_14784,N_14586,N_14737);
xor U14785 (N_14785,N_14564,N_14511);
or U14786 (N_14786,N_14590,N_14563);
or U14787 (N_14787,N_14723,N_14597);
nor U14788 (N_14788,N_14654,N_14743);
nand U14789 (N_14789,N_14703,N_14749);
nor U14790 (N_14790,N_14503,N_14745);
nor U14791 (N_14791,N_14684,N_14658);
nor U14792 (N_14792,N_14502,N_14660);
xor U14793 (N_14793,N_14555,N_14601);
xnor U14794 (N_14794,N_14647,N_14702);
nor U14795 (N_14795,N_14517,N_14593);
nand U14796 (N_14796,N_14508,N_14666);
nor U14797 (N_14797,N_14667,N_14578);
or U14798 (N_14798,N_14669,N_14697);
nand U14799 (N_14799,N_14533,N_14514);
nor U14800 (N_14800,N_14714,N_14695);
nor U14801 (N_14801,N_14500,N_14530);
nor U14802 (N_14802,N_14692,N_14650);
nand U14803 (N_14803,N_14557,N_14554);
xor U14804 (N_14804,N_14506,N_14611);
and U14805 (N_14805,N_14623,N_14726);
nor U14806 (N_14806,N_14691,N_14639);
or U14807 (N_14807,N_14591,N_14513);
nand U14808 (N_14808,N_14678,N_14733);
nand U14809 (N_14809,N_14633,N_14653);
nor U14810 (N_14810,N_14610,N_14527);
xor U14811 (N_14811,N_14700,N_14607);
and U14812 (N_14812,N_14716,N_14644);
xor U14813 (N_14813,N_14715,N_14580);
and U14814 (N_14814,N_14713,N_14738);
nor U14815 (N_14815,N_14556,N_14568);
xor U14816 (N_14816,N_14657,N_14664);
xnor U14817 (N_14817,N_14576,N_14661);
or U14818 (N_14818,N_14665,N_14522);
xnor U14819 (N_14819,N_14670,N_14735);
or U14820 (N_14820,N_14728,N_14573);
or U14821 (N_14821,N_14674,N_14632);
xnor U14822 (N_14822,N_14649,N_14680);
nand U14823 (N_14823,N_14641,N_14547);
nor U14824 (N_14824,N_14542,N_14707);
and U14825 (N_14825,N_14520,N_14620);
or U14826 (N_14826,N_14725,N_14574);
or U14827 (N_14827,N_14677,N_14570);
or U14828 (N_14828,N_14552,N_14505);
nand U14829 (N_14829,N_14562,N_14603);
nor U14830 (N_14830,N_14501,N_14746);
xnor U14831 (N_14831,N_14663,N_14551);
nand U14832 (N_14832,N_14567,N_14531);
and U14833 (N_14833,N_14673,N_14553);
or U14834 (N_14834,N_14613,N_14585);
xor U14835 (N_14835,N_14642,N_14682);
nor U14836 (N_14836,N_14510,N_14512);
and U14837 (N_14837,N_14705,N_14526);
and U14838 (N_14838,N_14693,N_14742);
nand U14839 (N_14839,N_14655,N_14694);
and U14840 (N_14840,N_14640,N_14558);
or U14841 (N_14841,N_14525,N_14617);
xnor U14842 (N_14842,N_14729,N_14621);
or U14843 (N_14843,N_14675,N_14636);
and U14844 (N_14844,N_14744,N_14588);
or U14845 (N_14845,N_14615,N_14631);
nand U14846 (N_14846,N_14712,N_14569);
xnor U14847 (N_14847,N_14540,N_14516);
xor U14848 (N_14848,N_14720,N_14734);
or U14849 (N_14849,N_14671,N_14698);
nand U14850 (N_14850,N_14696,N_14606);
and U14851 (N_14851,N_14652,N_14622);
nor U14852 (N_14852,N_14579,N_14509);
and U14853 (N_14853,N_14727,N_14719);
or U14854 (N_14854,N_14624,N_14521);
xor U14855 (N_14855,N_14630,N_14560);
and U14856 (N_14856,N_14565,N_14628);
or U14857 (N_14857,N_14686,N_14717);
and U14858 (N_14858,N_14550,N_14730);
xor U14859 (N_14859,N_14651,N_14599);
nor U14860 (N_14860,N_14605,N_14537);
and U14861 (N_14861,N_14709,N_14549);
nand U14862 (N_14862,N_14518,N_14543);
and U14863 (N_14863,N_14507,N_14687);
nand U14864 (N_14864,N_14589,N_14689);
xnor U14865 (N_14865,N_14643,N_14608);
and U14866 (N_14866,N_14612,N_14659);
nand U14867 (N_14867,N_14740,N_14701);
nand U14868 (N_14868,N_14538,N_14718);
and U14869 (N_14869,N_14546,N_14515);
and U14870 (N_14870,N_14504,N_14626);
xnor U14871 (N_14871,N_14561,N_14582);
and U14872 (N_14872,N_14600,N_14534);
nand U14873 (N_14873,N_14545,N_14528);
or U14874 (N_14874,N_14711,N_14618);
nor U14875 (N_14875,N_14662,N_14608);
nand U14876 (N_14876,N_14675,N_14683);
nor U14877 (N_14877,N_14514,N_14704);
xor U14878 (N_14878,N_14549,N_14644);
xor U14879 (N_14879,N_14644,N_14690);
nand U14880 (N_14880,N_14576,N_14645);
or U14881 (N_14881,N_14743,N_14587);
and U14882 (N_14882,N_14738,N_14638);
and U14883 (N_14883,N_14743,N_14516);
xor U14884 (N_14884,N_14570,N_14552);
xnor U14885 (N_14885,N_14739,N_14723);
or U14886 (N_14886,N_14681,N_14604);
nor U14887 (N_14887,N_14608,N_14592);
or U14888 (N_14888,N_14567,N_14550);
and U14889 (N_14889,N_14685,N_14689);
xnor U14890 (N_14890,N_14689,N_14746);
nand U14891 (N_14891,N_14515,N_14721);
xnor U14892 (N_14892,N_14549,N_14605);
xnor U14893 (N_14893,N_14551,N_14692);
nand U14894 (N_14894,N_14747,N_14724);
nor U14895 (N_14895,N_14736,N_14702);
or U14896 (N_14896,N_14589,N_14732);
xnor U14897 (N_14897,N_14681,N_14541);
or U14898 (N_14898,N_14618,N_14719);
nand U14899 (N_14899,N_14705,N_14667);
and U14900 (N_14900,N_14741,N_14605);
nand U14901 (N_14901,N_14574,N_14642);
and U14902 (N_14902,N_14559,N_14566);
or U14903 (N_14903,N_14612,N_14580);
and U14904 (N_14904,N_14701,N_14663);
or U14905 (N_14905,N_14580,N_14641);
nor U14906 (N_14906,N_14714,N_14541);
nor U14907 (N_14907,N_14513,N_14567);
xor U14908 (N_14908,N_14725,N_14697);
nand U14909 (N_14909,N_14708,N_14658);
nor U14910 (N_14910,N_14691,N_14707);
xor U14911 (N_14911,N_14571,N_14678);
xnor U14912 (N_14912,N_14715,N_14700);
nor U14913 (N_14913,N_14517,N_14658);
and U14914 (N_14914,N_14563,N_14728);
and U14915 (N_14915,N_14523,N_14593);
nand U14916 (N_14916,N_14673,N_14639);
nor U14917 (N_14917,N_14517,N_14642);
and U14918 (N_14918,N_14541,N_14668);
nand U14919 (N_14919,N_14514,N_14631);
or U14920 (N_14920,N_14749,N_14645);
and U14921 (N_14921,N_14722,N_14546);
xor U14922 (N_14922,N_14554,N_14686);
and U14923 (N_14923,N_14573,N_14592);
and U14924 (N_14924,N_14713,N_14555);
xnor U14925 (N_14925,N_14707,N_14692);
and U14926 (N_14926,N_14710,N_14727);
nor U14927 (N_14927,N_14552,N_14577);
nor U14928 (N_14928,N_14745,N_14559);
and U14929 (N_14929,N_14747,N_14592);
and U14930 (N_14930,N_14693,N_14668);
xor U14931 (N_14931,N_14573,N_14714);
and U14932 (N_14932,N_14714,N_14662);
or U14933 (N_14933,N_14581,N_14544);
and U14934 (N_14934,N_14679,N_14704);
nor U14935 (N_14935,N_14649,N_14664);
or U14936 (N_14936,N_14554,N_14590);
xnor U14937 (N_14937,N_14510,N_14658);
and U14938 (N_14938,N_14586,N_14718);
nor U14939 (N_14939,N_14550,N_14691);
nand U14940 (N_14940,N_14684,N_14555);
nor U14941 (N_14941,N_14725,N_14584);
nor U14942 (N_14942,N_14718,N_14500);
nand U14943 (N_14943,N_14656,N_14588);
xor U14944 (N_14944,N_14642,N_14673);
xor U14945 (N_14945,N_14724,N_14597);
nor U14946 (N_14946,N_14636,N_14505);
nand U14947 (N_14947,N_14608,N_14701);
xnor U14948 (N_14948,N_14708,N_14649);
or U14949 (N_14949,N_14618,N_14543);
xnor U14950 (N_14950,N_14733,N_14651);
or U14951 (N_14951,N_14618,N_14622);
nor U14952 (N_14952,N_14562,N_14574);
or U14953 (N_14953,N_14503,N_14657);
or U14954 (N_14954,N_14687,N_14558);
or U14955 (N_14955,N_14539,N_14564);
and U14956 (N_14956,N_14626,N_14543);
nor U14957 (N_14957,N_14583,N_14514);
nand U14958 (N_14958,N_14608,N_14699);
nand U14959 (N_14959,N_14739,N_14719);
nor U14960 (N_14960,N_14523,N_14587);
and U14961 (N_14961,N_14520,N_14642);
nand U14962 (N_14962,N_14669,N_14512);
nor U14963 (N_14963,N_14637,N_14613);
xor U14964 (N_14964,N_14731,N_14536);
and U14965 (N_14965,N_14733,N_14564);
nand U14966 (N_14966,N_14562,N_14697);
or U14967 (N_14967,N_14625,N_14676);
nor U14968 (N_14968,N_14680,N_14659);
or U14969 (N_14969,N_14714,N_14703);
or U14970 (N_14970,N_14562,N_14571);
and U14971 (N_14971,N_14599,N_14645);
xor U14972 (N_14972,N_14710,N_14672);
nor U14973 (N_14973,N_14626,N_14570);
nor U14974 (N_14974,N_14678,N_14511);
and U14975 (N_14975,N_14667,N_14580);
nor U14976 (N_14976,N_14681,N_14517);
nand U14977 (N_14977,N_14657,N_14587);
or U14978 (N_14978,N_14653,N_14706);
and U14979 (N_14979,N_14714,N_14745);
nand U14980 (N_14980,N_14618,N_14697);
nor U14981 (N_14981,N_14599,N_14720);
and U14982 (N_14982,N_14744,N_14648);
or U14983 (N_14983,N_14641,N_14636);
or U14984 (N_14984,N_14601,N_14523);
or U14985 (N_14985,N_14539,N_14526);
nor U14986 (N_14986,N_14611,N_14698);
xnor U14987 (N_14987,N_14697,N_14591);
xor U14988 (N_14988,N_14601,N_14645);
nand U14989 (N_14989,N_14651,N_14681);
nand U14990 (N_14990,N_14598,N_14514);
or U14991 (N_14991,N_14737,N_14500);
xor U14992 (N_14992,N_14535,N_14609);
nor U14993 (N_14993,N_14626,N_14531);
xnor U14994 (N_14994,N_14688,N_14661);
xor U14995 (N_14995,N_14529,N_14571);
or U14996 (N_14996,N_14646,N_14633);
nand U14997 (N_14997,N_14565,N_14579);
or U14998 (N_14998,N_14689,N_14732);
xnor U14999 (N_14999,N_14732,N_14686);
xnor UO_0 (O_0,N_14837,N_14929);
and UO_1 (O_1,N_14806,N_14923);
xnor UO_2 (O_2,N_14792,N_14771);
nor UO_3 (O_3,N_14832,N_14803);
or UO_4 (O_4,N_14753,N_14796);
nor UO_5 (O_5,N_14779,N_14920);
and UO_6 (O_6,N_14919,N_14988);
and UO_7 (O_7,N_14958,N_14894);
and UO_8 (O_8,N_14788,N_14862);
nand UO_9 (O_9,N_14835,N_14883);
xnor UO_10 (O_10,N_14888,N_14915);
xor UO_11 (O_11,N_14933,N_14943);
nand UO_12 (O_12,N_14909,N_14847);
nand UO_13 (O_13,N_14899,N_14926);
xor UO_14 (O_14,N_14893,N_14900);
nor UO_15 (O_15,N_14995,N_14793);
or UO_16 (O_16,N_14831,N_14782);
nand UO_17 (O_17,N_14986,N_14874);
xor UO_18 (O_18,N_14754,N_14829);
or UO_19 (O_19,N_14800,N_14759);
nor UO_20 (O_20,N_14872,N_14844);
nand UO_21 (O_21,N_14853,N_14934);
xor UO_22 (O_22,N_14777,N_14983);
or UO_23 (O_23,N_14839,N_14811);
or UO_24 (O_24,N_14869,N_14886);
and UO_25 (O_25,N_14968,N_14815);
xnor UO_26 (O_26,N_14816,N_14980);
xnor UO_27 (O_27,N_14921,N_14845);
nor UO_28 (O_28,N_14973,N_14780);
xnor UO_29 (O_29,N_14996,N_14967);
nor UO_30 (O_30,N_14972,N_14812);
and UO_31 (O_31,N_14767,N_14808);
xor UO_32 (O_32,N_14965,N_14964);
nand UO_33 (O_33,N_14783,N_14963);
nand UO_34 (O_34,N_14945,N_14804);
nand UO_35 (O_35,N_14957,N_14838);
or UO_36 (O_36,N_14914,N_14764);
or UO_37 (O_37,N_14758,N_14757);
nand UO_38 (O_38,N_14798,N_14992);
nand UO_39 (O_39,N_14998,N_14877);
xnor UO_40 (O_40,N_14828,N_14931);
nor UO_41 (O_41,N_14850,N_14867);
nand UO_42 (O_42,N_14940,N_14953);
nand UO_43 (O_43,N_14858,N_14876);
nor UO_44 (O_44,N_14810,N_14820);
and UO_45 (O_45,N_14917,N_14834);
xor UO_46 (O_46,N_14941,N_14781);
and UO_47 (O_47,N_14807,N_14994);
nand UO_48 (O_48,N_14773,N_14855);
or UO_49 (O_49,N_14954,N_14903);
nand UO_50 (O_50,N_14885,N_14814);
nand UO_51 (O_51,N_14763,N_14993);
and UO_52 (O_52,N_14916,N_14956);
and UO_53 (O_53,N_14962,N_14982);
nor UO_54 (O_54,N_14969,N_14866);
or UO_55 (O_55,N_14813,N_14880);
xnor UO_56 (O_56,N_14774,N_14786);
or UO_57 (O_57,N_14787,N_14827);
nand UO_58 (O_58,N_14930,N_14790);
and UO_59 (O_59,N_14922,N_14906);
nor UO_60 (O_60,N_14889,N_14991);
xor UO_61 (O_61,N_14939,N_14784);
nand UO_62 (O_62,N_14960,N_14971);
and UO_63 (O_63,N_14805,N_14868);
and UO_64 (O_64,N_14821,N_14842);
or UO_65 (O_65,N_14825,N_14822);
xnor UO_66 (O_66,N_14852,N_14951);
and UO_67 (O_67,N_14979,N_14762);
xor UO_68 (O_68,N_14794,N_14830);
xor UO_69 (O_69,N_14947,N_14890);
and UO_70 (O_70,N_14823,N_14959);
and UO_71 (O_71,N_14775,N_14978);
nor UO_72 (O_72,N_14949,N_14878);
or UO_73 (O_73,N_14857,N_14975);
or UO_74 (O_74,N_14881,N_14824);
xor UO_75 (O_75,N_14818,N_14836);
and UO_76 (O_76,N_14799,N_14769);
nand UO_77 (O_77,N_14879,N_14750);
xnor UO_78 (O_78,N_14860,N_14896);
nand UO_79 (O_79,N_14887,N_14752);
nand UO_80 (O_80,N_14948,N_14895);
xnor UO_81 (O_81,N_14849,N_14801);
and UO_82 (O_82,N_14802,N_14841);
xnor UO_83 (O_83,N_14952,N_14976);
nand UO_84 (O_84,N_14864,N_14809);
and UO_85 (O_85,N_14851,N_14999);
nand UO_86 (O_86,N_14913,N_14974);
nand UO_87 (O_87,N_14755,N_14950);
xnor UO_88 (O_88,N_14846,N_14756);
nand UO_89 (O_89,N_14901,N_14891);
or UO_90 (O_90,N_14840,N_14843);
nor UO_91 (O_91,N_14932,N_14912);
and UO_92 (O_92,N_14861,N_14768);
nand UO_93 (O_93,N_14776,N_14785);
xnor UO_94 (O_94,N_14770,N_14977);
or UO_95 (O_95,N_14910,N_14875);
nand UO_96 (O_96,N_14791,N_14772);
and UO_97 (O_97,N_14936,N_14865);
nand UO_98 (O_98,N_14984,N_14863);
xor UO_99 (O_99,N_14942,N_14927);
nor UO_100 (O_100,N_14856,N_14826);
or UO_101 (O_101,N_14897,N_14989);
nand UO_102 (O_102,N_14817,N_14870);
nor UO_103 (O_103,N_14766,N_14797);
and UO_104 (O_104,N_14981,N_14938);
or UO_105 (O_105,N_14937,N_14902);
xor UO_106 (O_106,N_14898,N_14907);
or UO_107 (O_107,N_14751,N_14997);
or UO_108 (O_108,N_14990,N_14848);
nor UO_109 (O_109,N_14873,N_14987);
nand UO_110 (O_110,N_14778,N_14911);
or UO_111 (O_111,N_14918,N_14884);
xor UO_112 (O_112,N_14985,N_14905);
nand UO_113 (O_113,N_14760,N_14795);
and UO_114 (O_114,N_14955,N_14854);
and UO_115 (O_115,N_14904,N_14946);
nand UO_116 (O_116,N_14761,N_14882);
and UO_117 (O_117,N_14833,N_14859);
or UO_118 (O_118,N_14928,N_14925);
xnor UO_119 (O_119,N_14924,N_14789);
and UO_120 (O_120,N_14892,N_14908);
or UO_121 (O_121,N_14961,N_14765);
xnor UO_122 (O_122,N_14871,N_14935);
xnor UO_123 (O_123,N_14819,N_14944);
or UO_124 (O_124,N_14970,N_14966);
nand UO_125 (O_125,N_14902,N_14965);
or UO_126 (O_126,N_14977,N_14773);
and UO_127 (O_127,N_14942,N_14874);
xnor UO_128 (O_128,N_14814,N_14937);
nor UO_129 (O_129,N_14962,N_14923);
and UO_130 (O_130,N_14892,N_14995);
or UO_131 (O_131,N_14860,N_14952);
nand UO_132 (O_132,N_14832,N_14835);
nand UO_133 (O_133,N_14892,N_14842);
or UO_134 (O_134,N_14843,N_14818);
xor UO_135 (O_135,N_14994,N_14898);
or UO_136 (O_136,N_14822,N_14873);
nand UO_137 (O_137,N_14955,N_14784);
and UO_138 (O_138,N_14923,N_14876);
and UO_139 (O_139,N_14972,N_14907);
nor UO_140 (O_140,N_14989,N_14895);
nor UO_141 (O_141,N_14763,N_14860);
and UO_142 (O_142,N_14853,N_14915);
and UO_143 (O_143,N_14869,N_14770);
nor UO_144 (O_144,N_14959,N_14936);
or UO_145 (O_145,N_14838,N_14883);
or UO_146 (O_146,N_14900,N_14956);
nand UO_147 (O_147,N_14887,N_14902);
nor UO_148 (O_148,N_14808,N_14765);
nand UO_149 (O_149,N_14812,N_14833);
and UO_150 (O_150,N_14817,N_14981);
xor UO_151 (O_151,N_14862,N_14890);
nor UO_152 (O_152,N_14970,N_14792);
xnor UO_153 (O_153,N_14775,N_14867);
nor UO_154 (O_154,N_14904,N_14753);
xnor UO_155 (O_155,N_14910,N_14983);
nand UO_156 (O_156,N_14891,N_14859);
or UO_157 (O_157,N_14842,N_14838);
nor UO_158 (O_158,N_14799,N_14958);
nor UO_159 (O_159,N_14851,N_14932);
or UO_160 (O_160,N_14971,N_14779);
nor UO_161 (O_161,N_14893,N_14951);
nand UO_162 (O_162,N_14839,N_14790);
nor UO_163 (O_163,N_14760,N_14752);
nand UO_164 (O_164,N_14826,N_14922);
and UO_165 (O_165,N_14859,N_14863);
or UO_166 (O_166,N_14983,N_14960);
nand UO_167 (O_167,N_14979,N_14760);
nor UO_168 (O_168,N_14869,N_14991);
and UO_169 (O_169,N_14929,N_14918);
xor UO_170 (O_170,N_14950,N_14930);
xnor UO_171 (O_171,N_14867,N_14812);
or UO_172 (O_172,N_14865,N_14972);
xor UO_173 (O_173,N_14776,N_14829);
xor UO_174 (O_174,N_14750,N_14912);
xor UO_175 (O_175,N_14950,N_14896);
nor UO_176 (O_176,N_14941,N_14955);
and UO_177 (O_177,N_14899,N_14821);
and UO_178 (O_178,N_14981,N_14812);
and UO_179 (O_179,N_14954,N_14988);
nand UO_180 (O_180,N_14865,N_14822);
and UO_181 (O_181,N_14786,N_14955);
xnor UO_182 (O_182,N_14869,N_14913);
and UO_183 (O_183,N_14783,N_14981);
nand UO_184 (O_184,N_14877,N_14983);
or UO_185 (O_185,N_14791,N_14930);
or UO_186 (O_186,N_14965,N_14878);
nand UO_187 (O_187,N_14960,N_14772);
nand UO_188 (O_188,N_14890,N_14785);
nand UO_189 (O_189,N_14776,N_14937);
or UO_190 (O_190,N_14929,N_14887);
or UO_191 (O_191,N_14946,N_14751);
or UO_192 (O_192,N_14870,N_14960);
xor UO_193 (O_193,N_14814,N_14794);
xnor UO_194 (O_194,N_14958,N_14971);
and UO_195 (O_195,N_14915,N_14809);
or UO_196 (O_196,N_14807,N_14993);
xnor UO_197 (O_197,N_14886,N_14940);
nor UO_198 (O_198,N_14877,N_14857);
and UO_199 (O_199,N_14912,N_14858);
nor UO_200 (O_200,N_14879,N_14892);
nor UO_201 (O_201,N_14900,N_14807);
nor UO_202 (O_202,N_14874,N_14880);
or UO_203 (O_203,N_14797,N_14760);
nor UO_204 (O_204,N_14912,N_14998);
nor UO_205 (O_205,N_14874,N_14790);
and UO_206 (O_206,N_14807,N_14984);
or UO_207 (O_207,N_14923,N_14930);
xor UO_208 (O_208,N_14879,N_14969);
xnor UO_209 (O_209,N_14800,N_14986);
xor UO_210 (O_210,N_14938,N_14773);
or UO_211 (O_211,N_14885,N_14983);
xnor UO_212 (O_212,N_14954,N_14884);
nor UO_213 (O_213,N_14873,N_14833);
nand UO_214 (O_214,N_14899,N_14962);
nand UO_215 (O_215,N_14914,N_14896);
nor UO_216 (O_216,N_14787,N_14854);
xnor UO_217 (O_217,N_14862,N_14986);
and UO_218 (O_218,N_14826,N_14752);
and UO_219 (O_219,N_14769,N_14960);
nor UO_220 (O_220,N_14769,N_14827);
or UO_221 (O_221,N_14996,N_14930);
nor UO_222 (O_222,N_14807,N_14828);
xnor UO_223 (O_223,N_14965,N_14831);
nand UO_224 (O_224,N_14975,N_14866);
xor UO_225 (O_225,N_14786,N_14868);
nor UO_226 (O_226,N_14931,N_14909);
or UO_227 (O_227,N_14952,N_14834);
nand UO_228 (O_228,N_14972,N_14941);
and UO_229 (O_229,N_14948,N_14992);
or UO_230 (O_230,N_14953,N_14760);
or UO_231 (O_231,N_14850,N_14954);
and UO_232 (O_232,N_14865,N_14832);
nor UO_233 (O_233,N_14911,N_14809);
and UO_234 (O_234,N_14762,N_14856);
xor UO_235 (O_235,N_14916,N_14866);
xor UO_236 (O_236,N_14869,N_14841);
nor UO_237 (O_237,N_14768,N_14818);
and UO_238 (O_238,N_14937,N_14886);
nor UO_239 (O_239,N_14751,N_14811);
nor UO_240 (O_240,N_14757,N_14890);
and UO_241 (O_241,N_14889,N_14883);
xnor UO_242 (O_242,N_14834,N_14845);
and UO_243 (O_243,N_14763,N_14882);
or UO_244 (O_244,N_14970,N_14861);
nand UO_245 (O_245,N_14828,N_14843);
or UO_246 (O_246,N_14856,N_14995);
or UO_247 (O_247,N_14922,N_14889);
or UO_248 (O_248,N_14909,N_14930);
and UO_249 (O_249,N_14881,N_14804);
and UO_250 (O_250,N_14937,N_14793);
xor UO_251 (O_251,N_14842,N_14924);
nor UO_252 (O_252,N_14881,N_14765);
nor UO_253 (O_253,N_14768,N_14878);
nor UO_254 (O_254,N_14980,N_14884);
xnor UO_255 (O_255,N_14783,N_14830);
nand UO_256 (O_256,N_14961,N_14777);
and UO_257 (O_257,N_14839,N_14827);
xor UO_258 (O_258,N_14763,N_14892);
nand UO_259 (O_259,N_14903,N_14826);
nor UO_260 (O_260,N_14936,N_14766);
and UO_261 (O_261,N_14964,N_14979);
and UO_262 (O_262,N_14796,N_14868);
or UO_263 (O_263,N_14789,N_14939);
or UO_264 (O_264,N_14859,N_14766);
nor UO_265 (O_265,N_14759,N_14939);
and UO_266 (O_266,N_14792,N_14805);
nand UO_267 (O_267,N_14766,N_14853);
or UO_268 (O_268,N_14883,N_14912);
xnor UO_269 (O_269,N_14838,N_14836);
and UO_270 (O_270,N_14757,N_14913);
or UO_271 (O_271,N_14766,N_14999);
nand UO_272 (O_272,N_14991,N_14768);
xnor UO_273 (O_273,N_14754,N_14915);
or UO_274 (O_274,N_14754,N_14846);
or UO_275 (O_275,N_14774,N_14966);
or UO_276 (O_276,N_14934,N_14815);
and UO_277 (O_277,N_14862,N_14951);
nand UO_278 (O_278,N_14866,N_14955);
nor UO_279 (O_279,N_14823,N_14822);
xor UO_280 (O_280,N_14874,N_14814);
or UO_281 (O_281,N_14995,N_14834);
and UO_282 (O_282,N_14990,N_14832);
and UO_283 (O_283,N_14812,N_14946);
nor UO_284 (O_284,N_14848,N_14997);
or UO_285 (O_285,N_14840,N_14932);
or UO_286 (O_286,N_14845,N_14843);
nand UO_287 (O_287,N_14918,N_14764);
xnor UO_288 (O_288,N_14890,N_14989);
xnor UO_289 (O_289,N_14892,N_14992);
and UO_290 (O_290,N_14829,N_14945);
xor UO_291 (O_291,N_14887,N_14890);
and UO_292 (O_292,N_14794,N_14917);
nor UO_293 (O_293,N_14803,N_14897);
nand UO_294 (O_294,N_14812,N_14937);
nor UO_295 (O_295,N_14765,N_14759);
or UO_296 (O_296,N_14756,N_14913);
or UO_297 (O_297,N_14938,N_14912);
nor UO_298 (O_298,N_14869,N_14937);
and UO_299 (O_299,N_14788,N_14917);
nand UO_300 (O_300,N_14941,N_14786);
nor UO_301 (O_301,N_14969,N_14834);
or UO_302 (O_302,N_14988,N_14930);
nor UO_303 (O_303,N_14948,N_14809);
nor UO_304 (O_304,N_14777,N_14752);
nand UO_305 (O_305,N_14957,N_14969);
or UO_306 (O_306,N_14910,N_14828);
or UO_307 (O_307,N_14766,N_14963);
xnor UO_308 (O_308,N_14985,N_14829);
or UO_309 (O_309,N_14912,N_14761);
and UO_310 (O_310,N_14847,N_14871);
xor UO_311 (O_311,N_14846,N_14917);
and UO_312 (O_312,N_14783,N_14841);
or UO_313 (O_313,N_14809,N_14975);
xor UO_314 (O_314,N_14841,N_14954);
or UO_315 (O_315,N_14848,N_14864);
nand UO_316 (O_316,N_14984,N_14985);
and UO_317 (O_317,N_14866,N_14953);
and UO_318 (O_318,N_14991,N_14756);
nand UO_319 (O_319,N_14975,N_14786);
nor UO_320 (O_320,N_14913,N_14987);
nor UO_321 (O_321,N_14906,N_14896);
nand UO_322 (O_322,N_14951,N_14928);
nor UO_323 (O_323,N_14809,N_14844);
or UO_324 (O_324,N_14841,N_14776);
xnor UO_325 (O_325,N_14968,N_14997);
and UO_326 (O_326,N_14751,N_14799);
xnor UO_327 (O_327,N_14953,N_14893);
xor UO_328 (O_328,N_14959,N_14902);
or UO_329 (O_329,N_14816,N_14941);
and UO_330 (O_330,N_14961,N_14885);
and UO_331 (O_331,N_14923,N_14961);
or UO_332 (O_332,N_14774,N_14798);
nor UO_333 (O_333,N_14751,N_14837);
or UO_334 (O_334,N_14904,N_14775);
xnor UO_335 (O_335,N_14878,N_14844);
or UO_336 (O_336,N_14996,N_14801);
or UO_337 (O_337,N_14919,N_14755);
nand UO_338 (O_338,N_14963,N_14801);
or UO_339 (O_339,N_14863,N_14755);
nor UO_340 (O_340,N_14997,N_14867);
and UO_341 (O_341,N_14767,N_14758);
and UO_342 (O_342,N_14964,N_14995);
xor UO_343 (O_343,N_14901,N_14766);
or UO_344 (O_344,N_14761,N_14991);
and UO_345 (O_345,N_14868,N_14854);
or UO_346 (O_346,N_14871,N_14823);
xor UO_347 (O_347,N_14943,N_14828);
and UO_348 (O_348,N_14854,N_14786);
nand UO_349 (O_349,N_14975,N_14973);
and UO_350 (O_350,N_14806,N_14869);
and UO_351 (O_351,N_14893,N_14884);
nor UO_352 (O_352,N_14865,N_14930);
and UO_353 (O_353,N_14953,N_14977);
nand UO_354 (O_354,N_14978,N_14847);
nand UO_355 (O_355,N_14940,N_14844);
xor UO_356 (O_356,N_14788,N_14987);
or UO_357 (O_357,N_14910,N_14795);
nor UO_358 (O_358,N_14766,N_14897);
nor UO_359 (O_359,N_14973,N_14960);
and UO_360 (O_360,N_14856,N_14816);
or UO_361 (O_361,N_14921,N_14968);
nand UO_362 (O_362,N_14762,N_14940);
xnor UO_363 (O_363,N_14904,N_14891);
and UO_364 (O_364,N_14939,N_14762);
nand UO_365 (O_365,N_14894,N_14800);
nor UO_366 (O_366,N_14920,N_14975);
xor UO_367 (O_367,N_14874,N_14806);
or UO_368 (O_368,N_14819,N_14991);
or UO_369 (O_369,N_14923,N_14826);
nand UO_370 (O_370,N_14992,N_14876);
and UO_371 (O_371,N_14761,N_14903);
and UO_372 (O_372,N_14994,N_14856);
nor UO_373 (O_373,N_14761,N_14939);
or UO_374 (O_374,N_14992,N_14973);
nand UO_375 (O_375,N_14927,N_14800);
nand UO_376 (O_376,N_14936,N_14796);
and UO_377 (O_377,N_14798,N_14867);
or UO_378 (O_378,N_14950,N_14953);
and UO_379 (O_379,N_14780,N_14768);
and UO_380 (O_380,N_14882,N_14758);
xor UO_381 (O_381,N_14845,N_14939);
nor UO_382 (O_382,N_14799,N_14831);
and UO_383 (O_383,N_14975,N_14869);
and UO_384 (O_384,N_14847,N_14797);
nor UO_385 (O_385,N_14799,N_14821);
nor UO_386 (O_386,N_14848,N_14752);
xnor UO_387 (O_387,N_14822,N_14987);
nor UO_388 (O_388,N_14764,N_14770);
and UO_389 (O_389,N_14977,N_14989);
xnor UO_390 (O_390,N_14972,N_14893);
nand UO_391 (O_391,N_14961,N_14919);
and UO_392 (O_392,N_14979,N_14962);
nand UO_393 (O_393,N_14763,N_14761);
and UO_394 (O_394,N_14841,N_14834);
and UO_395 (O_395,N_14884,N_14841);
xor UO_396 (O_396,N_14970,N_14765);
nor UO_397 (O_397,N_14970,N_14881);
or UO_398 (O_398,N_14955,N_14893);
or UO_399 (O_399,N_14822,N_14938);
nor UO_400 (O_400,N_14992,N_14950);
xnor UO_401 (O_401,N_14751,N_14764);
or UO_402 (O_402,N_14907,N_14754);
and UO_403 (O_403,N_14853,N_14840);
nand UO_404 (O_404,N_14752,N_14831);
or UO_405 (O_405,N_14816,N_14908);
and UO_406 (O_406,N_14893,N_14965);
xnor UO_407 (O_407,N_14803,N_14954);
xnor UO_408 (O_408,N_14961,N_14957);
nor UO_409 (O_409,N_14851,N_14964);
or UO_410 (O_410,N_14842,N_14754);
nor UO_411 (O_411,N_14776,N_14883);
and UO_412 (O_412,N_14908,N_14930);
or UO_413 (O_413,N_14926,N_14769);
and UO_414 (O_414,N_14858,N_14910);
xor UO_415 (O_415,N_14990,N_14954);
nor UO_416 (O_416,N_14852,N_14796);
nand UO_417 (O_417,N_14885,N_14990);
nor UO_418 (O_418,N_14857,N_14978);
nor UO_419 (O_419,N_14926,N_14808);
and UO_420 (O_420,N_14815,N_14888);
nand UO_421 (O_421,N_14755,N_14925);
xor UO_422 (O_422,N_14776,N_14885);
nand UO_423 (O_423,N_14991,N_14770);
and UO_424 (O_424,N_14960,N_14953);
nor UO_425 (O_425,N_14755,N_14935);
nor UO_426 (O_426,N_14918,N_14974);
xnor UO_427 (O_427,N_14845,N_14987);
or UO_428 (O_428,N_14962,N_14844);
nor UO_429 (O_429,N_14896,N_14999);
or UO_430 (O_430,N_14757,N_14835);
or UO_431 (O_431,N_14780,N_14827);
nand UO_432 (O_432,N_14829,N_14804);
or UO_433 (O_433,N_14932,N_14817);
and UO_434 (O_434,N_14867,N_14962);
nand UO_435 (O_435,N_14756,N_14781);
or UO_436 (O_436,N_14980,N_14793);
nand UO_437 (O_437,N_14969,N_14907);
or UO_438 (O_438,N_14914,N_14859);
or UO_439 (O_439,N_14879,N_14883);
and UO_440 (O_440,N_14766,N_14837);
nor UO_441 (O_441,N_14905,N_14761);
nand UO_442 (O_442,N_14879,N_14895);
and UO_443 (O_443,N_14777,N_14795);
or UO_444 (O_444,N_14883,N_14866);
nor UO_445 (O_445,N_14868,N_14979);
xor UO_446 (O_446,N_14754,N_14833);
or UO_447 (O_447,N_14797,N_14918);
xor UO_448 (O_448,N_14948,N_14923);
nor UO_449 (O_449,N_14818,N_14922);
nand UO_450 (O_450,N_14895,N_14913);
nor UO_451 (O_451,N_14978,N_14958);
nand UO_452 (O_452,N_14877,N_14791);
nand UO_453 (O_453,N_14974,N_14757);
and UO_454 (O_454,N_14813,N_14938);
or UO_455 (O_455,N_14954,N_14882);
nand UO_456 (O_456,N_14813,N_14774);
xor UO_457 (O_457,N_14872,N_14956);
or UO_458 (O_458,N_14933,N_14884);
xor UO_459 (O_459,N_14978,N_14844);
xnor UO_460 (O_460,N_14866,N_14798);
nor UO_461 (O_461,N_14920,N_14987);
nand UO_462 (O_462,N_14780,N_14898);
nand UO_463 (O_463,N_14895,N_14975);
nand UO_464 (O_464,N_14840,N_14760);
and UO_465 (O_465,N_14768,N_14947);
nor UO_466 (O_466,N_14760,N_14900);
nand UO_467 (O_467,N_14948,N_14896);
or UO_468 (O_468,N_14761,N_14819);
nand UO_469 (O_469,N_14789,N_14869);
xor UO_470 (O_470,N_14836,N_14865);
or UO_471 (O_471,N_14904,N_14943);
nor UO_472 (O_472,N_14897,N_14928);
or UO_473 (O_473,N_14837,N_14893);
xnor UO_474 (O_474,N_14946,N_14834);
nand UO_475 (O_475,N_14890,N_14941);
nor UO_476 (O_476,N_14935,N_14836);
and UO_477 (O_477,N_14837,N_14950);
nor UO_478 (O_478,N_14900,N_14797);
and UO_479 (O_479,N_14835,N_14870);
nand UO_480 (O_480,N_14922,N_14834);
and UO_481 (O_481,N_14756,N_14877);
xnor UO_482 (O_482,N_14966,N_14823);
and UO_483 (O_483,N_14867,N_14899);
nor UO_484 (O_484,N_14965,N_14807);
and UO_485 (O_485,N_14917,N_14807);
nand UO_486 (O_486,N_14941,N_14892);
nand UO_487 (O_487,N_14970,N_14867);
xnor UO_488 (O_488,N_14970,N_14781);
nor UO_489 (O_489,N_14850,N_14933);
nand UO_490 (O_490,N_14754,N_14792);
nor UO_491 (O_491,N_14764,N_14981);
or UO_492 (O_492,N_14953,N_14782);
nand UO_493 (O_493,N_14818,N_14772);
or UO_494 (O_494,N_14994,N_14947);
nor UO_495 (O_495,N_14886,N_14916);
nand UO_496 (O_496,N_14875,N_14760);
nor UO_497 (O_497,N_14926,N_14871);
nor UO_498 (O_498,N_14752,N_14936);
xor UO_499 (O_499,N_14996,N_14960);
nor UO_500 (O_500,N_14935,N_14892);
or UO_501 (O_501,N_14810,N_14759);
xor UO_502 (O_502,N_14830,N_14828);
nor UO_503 (O_503,N_14793,N_14927);
xor UO_504 (O_504,N_14956,N_14844);
xor UO_505 (O_505,N_14932,N_14994);
nand UO_506 (O_506,N_14939,N_14892);
nand UO_507 (O_507,N_14844,N_14790);
nor UO_508 (O_508,N_14819,N_14838);
and UO_509 (O_509,N_14946,N_14769);
xnor UO_510 (O_510,N_14777,N_14979);
xnor UO_511 (O_511,N_14857,N_14862);
nor UO_512 (O_512,N_14857,N_14753);
nand UO_513 (O_513,N_14833,N_14843);
nand UO_514 (O_514,N_14751,N_14777);
nor UO_515 (O_515,N_14975,N_14877);
xnor UO_516 (O_516,N_14916,N_14998);
or UO_517 (O_517,N_14871,N_14939);
or UO_518 (O_518,N_14869,N_14963);
or UO_519 (O_519,N_14860,N_14854);
nor UO_520 (O_520,N_14853,N_14961);
nand UO_521 (O_521,N_14892,N_14962);
xnor UO_522 (O_522,N_14887,N_14781);
nand UO_523 (O_523,N_14824,N_14977);
or UO_524 (O_524,N_14761,N_14776);
or UO_525 (O_525,N_14862,N_14883);
and UO_526 (O_526,N_14930,N_14882);
nor UO_527 (O_527,N_14946,N_14925);
or UO_528 (O_528,N_14957,N_14809);
nor UO_529 (O_529,N_14837,N_14944);
and UO_530 (O_530,N_14967,N_14909);
nand UO_531 (O_531,N_14915,N_14865);
nand UO_532 (O_532,N_14949,N_14776);
or UO_533 (O_533,N_14911,N_14804);
nand UO_534 (O_534,N_14935,N_14875);
and UO_535 (O_535,N_14913,N_14855);
nor UO_536 (O_536,N_14805,N_14798);
nand UO_537 (O_537,N_14800,N_14849);
or UO_538 (O_538,N_14845,N_14943);
xor UO_539 (O_539,N_14827,N_14794);
and UO_540 (O_540,N_14843,N_14821);
or UO_541 (O_541,N_14881,N_14823);
nand UO_542 (O_542,N_14821,N_14871);
nand UO_543 (O_543,N_14868,N_14985);
nand UO_544 (O_544,N_14873,N_14997);
and UO_545 (O_545,N_14835,N_14955);
nor UO_546 (O_546,N_14851,N_14842);
and UO_547 (O_547,N_14898,N_14784);
or UO_548 (O_548,N_14850,N_14862);
xnor UO_549 (O_549,N_14942,N_14989);
xnor UO_550 (O_550,N_14951,N_14963);
or UO_551 (O_551,N_14904,N_14959);
or UO_552 (O_552,N_14752,N_14935);
or UO_553 (O_553,N_14943,N_14928);
or UO_554 (O_554,N_14806,N_14750);
and UO_555 (O_555,N_14801,N_14967);
or UO_556 (O_556,N_14876,N_14852);
or UO_557 (O_557,N_14808,N_14875);
nor UO_558 (O_558,N_14886,N_14979);
or UO_559 (O_559,N_14824,N_14808);
nor UO_560 (O_560,N_14830,N_14965);
or UO_561 (O_561,N_14769,N_14813);
nand UO_562 (O_562,N_14798,N_14829);
nand UO_563 (O_563,N_14839,N_14794);
or UO_564 (O_564,N_14851,N_14803);
nand UO_565 (O_565,N_14756,N_14786);
and UO_566 (O_566,N_14789,N_14919);
nand UO_567 (O_567,N_14842,N_14879);
nor UO_568 (O_568,N_14860,N_14994);
and UO_569 (O_569,N_14988,N_14831);
xor UO_570 (O_570,N_14821,N_14908);
xor UO_571 (O_571,N_14776,N_14789);
or UO_572 (O_572,N_14954,N_14839);
nor UO_573 (O_573,N_14845,N_14813);
nand UO_574 (O_574,N_14895,N_14884);
nand UO_575 (O_575,N_14822,N_14985);
xnor UO_576 (O_576,N_14874,N_14807);
nor UO_577 (O_577,N_14863,N_14881);
or UO_578 (O_578,N_14879,N_14971);
nand UO_579 (O_579,N_14817,N_14997);
nand UO_580 (O_580,N_14758,N_14917);
xor UO_581 (O_581,N_14774,N_14999);
or UO_582 (O_582,N_14876,N_14966);
nor UO_583 (O_583,N_14918,N_14767);
xnor UO_584 (O_584,N_14881,N_14858);
or UO_585 (O_585,N_14888,N_14775);
nand UO_586 (O_586,N_14817,N_14783);
nor UO_587 (O_587,N_14991,N_14902);
nor UO_588 (O_588,N_14827,N_14896);
and UO_589 (O_589,N_14869,N_14962);
or UO_590 (O_590,N_14800,N_14970);
xor UO_591 (O_591,N_14768,N_14924);
nor UO_592 (O_592,N_14949,N_14866);
and UO_593 (O_593,N_14936,N_14799);
nor UO_594 (O_594,N_14914,N_14986);
or UO_595 (O_595,N_14942,N_14820);
xor UO_596 (O_596,N_14786,N_14856);
nor UO_597 (O_597,N_14804,N_14823);
and UO_598 (O_598,N_14914,N_14816);
nand UO_599 (O_599,N_14849,N_14851);
nor UO_600 (O_600,N_14844,N_14958);
nand UO_601 (O_601,N_14801,N_14794);
nand UO_602 (O_602,N_14832,N_14868);
and UO_603 (O_603,N_14875,N_14967);
nor UO_604 (O_604,N_14872,N_14870);
xnor UO_605 (O_605,N_14862,N_14908);
nor UO_606 (O_606,N_14872,N_14851);
xnor UO_607 (O_607,N_14782,N_14932);
and UO_608 (O_608,N_14981,N_14961);
nor UO_609 (O_609,N_14796,N_14853);
or UO_610 (O_610,N_14808,N_14987);
nand UO_611 (O_611,N_14957,N_14966);
nand UO_612 (O_612,N_14878,N_14882);
or UO_613 (O_613,N_14815,N_14932);
nand UO_614 (O_614,N_14857,N_14956);
xor UO_615 (O_615,N_14840,N_14841);
and UO_616 (O_616,N_14866,N_14896);
nand UO_617 (O_617,N_14768,N_14916);
and UO_618 (O_618,N_14857,N_14764);
and UO_619 (O_619,N_14837,N_14770);
nor UO_620 (O_620,N_14922,N_14959);
or UO_621 (O_621,N_14945,N_14981);
and UO_622 (O_622,N_14943,N_14753);
nand UO_623 (O_623,N_14991,N_14924);
nor UO_624 (O_624,N_14941,N_14854);
and UO_625 (O_625,N_14993,N_14926);
xnor UO_626 (O_626,N_14996,N_14752);
xor UO_627 (O_627,N_14792,N_14939);
nor UO_628 (O_628,N_14812,N_14888);
nor UO_629 (O_629,N_14996,N_14813);
nor UO_630 (O_630,N_14904,N_14927);
nor UO_631 (O_631,N_14923,N_14973);
nor UO_632 (O_632,N_14831,N_14998);
nand UO_633 (O_633,N_14817,N_14926);
and UO_634 (O_634,N_14806,N_14767);
and UO_635 (O_635,N_14872,N_14906);
nand UO_636 (O_636,N_14931,N_14918);
nor UO_637 (O_637,N_14962,N_14778);
xnor UO_638 (O_638,N_14914,N_14932);
nand UO_639 (O_639,N_14842,N_14891);
nor UO_640 (O_640,N_14973,N_14752);
nand UO_641 (O_641,N_14811,N_14855);
nand UO_642 (O_642,N_14972,N_14822);
nand UO_643 (O_643,N_14802,N_14867);
xor UO_644 (O_644,N_14848,N_14889);
nor UO_645 (O_645,N_14895,N_14880);
xnor UO_646 (O_646,N_14818,N_14763);
xor UO_647 (O_647,N_14762,N_14924);
xnor UO_648 (O_648,N_14808,N_14846);
nand UO_649 (O_649,N_14921,N_14971);
and UO_650 (O_650,N_14890,N_14790);
nand UO_651 (O_651,N_14977,N_14928);
nand UO_652 (O_652,N_14792,N_14929);
xor UO_653 (O_653,N_14758,N_14853);
and UO_654 (O_654,N_14973,N_14884);
xor UO_655 (O_655,N_14894,N_14987);
and UO_656 (O_656,N_14828,N_14936);
and UO_657 (O_657,N_14892,N_14898);
and UO_658 (O_658,N_14841,N_14823);
nand UO_659 (O_659,N_14967,N_14750);
xnor UO_660 (O_660,N_14881,N_14788);
or UO_661 (O_661,N_14812,N_14996);
or UO_662 (O_662,N_14769,N_14816);
xor UO_663 (O_663,N_14787,N_14959);
nand UO_664 (O_664,N_14879,N_14998);
or UO_665 (O_665,N_14753,N_14998);
xnor UO_666 (O_666,N_14950,N_14946);
and UO_667 (O_667,N_14908,N_14858);
or UO_668 (O_668,N_14907,N_14949);
nor UO_669 (O_669,N_14872,N_14882);
xnor UO_670 (O_670,N_14954,N_14910);
nand UO_671 (O_671,N_14950,N_14979);
and UO_672 (O_672,N_14863,N_14941);
and UO_673 (O_673,N_14895,N_14858);
nand UO_674 (O_674,N_14970,N_14838);
and UO_675 (O_675,N_14904,N_14978);
nor UO_676 (O_676,N_14804,N_14998);
nand UO_677 (O_677,N_14828,N_14946);
nand UO_678 (O_678,N_14953,N_14832);
xnor UO_679 (O_679,N_14819,N_14884);
xor UO_680 (O_680,N_14868,N_14896);
nor UO_681 (O_681,N_14977,N_14838);
and UO_682 (O_682,N_14877,N_14884);
nor UO_683 (O_683,N_14908,N_14830);
and UO_684 (O_684,N_14910,N_14861);
nand UO_685 (O_685,N_14846,N_14922);
nand UO_686 (O_686,N_14953,N_14872);
xnor UO_687 (O_687,N_14839,N_14775);
or UO_688 (O_688,N_14946,N_14786);
xnor UO_689 (O_689,N_14791,N_14973);
or UO_690 (O_690,N_14887,N_14917);
nand UO_691 (O_691,N_14843,N_14856);
xnor UO_692 (O_692,N_14792,N_14896);
nor UO_693 (O_693,N_14875,N_14920);
nor UO_694 (O_694,N_14803,N_14772);
and UO_695 (O_695,N_14945,N_14780);
xnor UO_696 (O_696,N_14999,N_14863);
nor UO_697 (O_697,N_14947,N_14971);
nor UO_698 (O_698,N_14939,N_14760);
nand UO_699 (O_699,N_14910,N_14881);
and UO_700 (O_700,N_14770,N_14994);
xnor UO_701 (O_701,N_14897,N_14753);
and UO_702 (O_702,N_14876,N_14995);
and UO_703 (O_703,N_14908,N_14814);
nand UO_704 (O_704,N_14905,N_14841);
or UO_705 (O_705,N_14950,N_14842);
nand UO_706 (O_706,N_14908,N_14985);
xnor UO_707 (O_707,N_14815,N_14949);
nand UO_708 (O_708,N_14789,N_14945);
and UO_709 (O_709,N_14771,N_14871);
and UO_710 (O_710,N_14882,N_14753);
nand UO_711 (O_711,N_14849,N_14811);
or UO_712 (O_712,N_14788,N_14805);
nand UO_713 (O_713,N_14870,N_14907);
xor UO_714 (O_714,N_14846,N_14942);
xor UO_715 (O_715,N_14797,N_14866);
or UO_716 (O_716,N_14968,N_14961);
nor UO_717 (O_717,N_14975,N_14847);
nor UO_718 (O_718,N_14828,N_14959);
or UO_719 (O_719,N_14940,N_14957);
nor UO_720 (O_720,N_14774,N_14875);
nor UO_721 (O_721,N_14836,N_14800);
or UO_722 (O_722,N_14811,N_14892);
and UO_723 (O_723,N_14903,N_14965);
and UO_724 (O_724,N_14878,N_14813);
or UO_725 (O_725,N_14851,N_14782);
nor UO_726 (O_726,N_14855,N_14849);
nand UO_727 (O_727,N_14963,N_14996);
nor UO_728 (O_728,N_14848,N_14886);
xnor UO_729 (O_729,N_14912,N_14751);
nand UO_730 (O_730,N_14900,N_14945);
xor UO_731 (O_731,N_14903,N_14774);
and UO_732 (O_732,N_14879,N_14853);
or UO_733 (O_733,N_14773,N_14784);
nor UO_734 (O_734,N_14953,N_14870);
and UO_735 (O_735,N_14822,N_14894);
nand UO_736 (O_736,N_14809,N_14837);
nand UO_737 (O_737,N_14843,N_14880);
and UO_738 (O_738,N_14866,N_14950);
nor UO_739 (O_739,N_14830,N_14773);
nor UO_740 (O_740,N_14849,N_14985);
nand UO_741 (O_741,N_14971,N_14846);
nand UO_742 (O_742,N_14953,N_14954);
xnor UO_743 (O_743,N_14839,N_14764);
nor UO_744 (O_744,N_14772,N_14884);
xor UO_745 (O_745,N_14838,N_14790);
nand UO_746 (O_746,N_14976,N_14956);
or UO_747 (O_747,N_14991,N_14873);
and UO_748 (O_748,N_14820,N_14842);
xor UO_749 (O_749,N_14788,N_14905);
nor UO_750 (O_750,N_14819,N_14902);
nor UO_751 (O_751,N_14962,N_14802);
or UO_752 (O_752,N_14766,N_14895);
nor UO_753 (O_753,N_14839,N_14799);
and UO_754 (O_754,N_14910,N_14859);
and UO_755 (O_755,N_14764,N_14983);
nand UO_756 (O_756,N_14860,N_14964);
and UO_757 (O_757,N_14893,N_14802);
or UO_758 (O_758,N_14780,N_14871);
or UO_759 (O_759,N_14949,N_14807);
xnor UO_760 (O_760,N_14928,N_14780);
and UO_761 (O_761,N_14890,N_14763);
nor UO_762 (O_762,N_14848,N_14896);
nand UO_763 (O_763,N_14935,N_14924);
or UO_764 (O_764,N_14994,N_14865);
and UO_765 (O_765,N_14841,N_14877);
and UO_766 (O_766,N_14851,N_14897);
or UO_767 (O_767,N_14753,N_14843);
nand UO_768 (O_768,N_14972,N_14984);
and UO_769 (O_769,N_14941,N_14855);
nor UO_770 (O_770,N_14822,N_14820);
and UO_771 (O_771,N_14775,N_14963);
nand UO_772 (O_772,N_14869,N_14839);
or UO_773 (O_773,N_14767,N_14803);
nor UO_774 (O_774,N_14967,N_14991);
nor UO_775 (O_775,N_14775,N_14977);
or UO_776 (O_776,N_14849,N_14936);
nor UO_777 (O_777,N_14931,N_14886);
and UO_778 (O_778,N_14987,N_14979);
nor UO_779 (O_779,N_14894,N_14809);
nor UO_780 (O_780,N_14763,N_14811);
or UO_781 (O_781,N_14867,N_14991);
nor UO_782 (O_782,N_14872,N_14914);
xnor UO_783 (O_783,N_14947,N_14820);
xnor UO_784 (O_784,N_14893,N_14949);
nor UO_785 (O_785,N_14766,N_14986);
xor UO_786 (O_786,N_14777,N_14910);
xnor UO_787 (O_787,N_14754,N_14961);
and UO_788 (O_788,N_14950,N_14835);
or UO_789 (O_789,N_14861,N_14829);
nor UO_790 (O_790,N_14959,N_14850);
nor UO_791 (O_791,N_14890,N_14874);
nor UO_792 (O_792,N_14829,N_14931);
xnor UO_793 (O_793,N_14867,N_14763);
and UO_794 (O_794,N_14805,N_14770);
nand UO_795 (O_795,N_14831,N_14999);
and UO_796 (O_796,N_14913,N_14911);
xor UO_797 (O_797,N_14914,N_14978);
or UO_798 (O_798,N_14759,N_14932);
and UO_799 (O_799,N_14786,N_14853);
and UO_800 (O_800,N_14886,N_14814);
or UO_801 (O_801,N_14766,N_14794);
nand UO_802 (O_802,N_14887,N_14963);
xor UO_803 (O_803,N_14976,N_14773);
or UO_804 (O_804,N_14908,N_14849);
and UO_805 (O_805,N_14986,N_14987);
and UO_806 (O_806,N_14909,N_14996);
nor UO_807 (O_807,N_14925,N_14824);
nor UO_808 (O_808,N_14942,N_14893);
and UO_809 (O_809,N_14819,N_14790);
xnor UO_810 (O_810,N_14893,N_14988);
nand UO_811 (O_811,N_14874,N_14751);
nand UO_812 (O_812,N_14935,N_14973);
and UO_813 (O_813,N_14889,N_14872);
or UO_814 (O_814,N_14917,N_14929);
nand UO_815 (O_815,N_14811,N_14843);
and UO_816 (O_816,N_14851,N_14911);
nor UO_817 (O_817,N_14759,N_14850);
nand UO_818 (O_818,N_14812,N_14794);
or UO_819 (O_819,N_14889,N_14851);
nor UO_820 (O_820,N_14840,N_14988);
nand UO_821 (O_821,N_14843,N_14773);
xor UO_822 (O_822,N_14787,N_14934);
and UO_823 (O_823,N_14817,N_14831);
xor UO_824 (O_824,N_14932,N_14946);
nand UO_825 (O_825,N_14930,N_14983);
nor UO_826 (O_826,N_14841,N_14993);
nand UO_827 (O_827,N_14981,N_14969);
or UO_828 (O_828,N_14775,N_14966);
nor UO_829 (O_829,N_14765,N_14835);
nor UO_830 (O_830,N_14865,N_14923);
xor UO_831 (O_831,N_14878,N_14922);
xor UO_832 (O_832,N_14771,N_14885);
xor UO_833 (O_833,N_14755,N_14883);
and UO_834 (O_834,N_14969,N_14922);
or UO_835 (O_835,N_14868,N_14916);
and UO_836 (O_836,N_14825,N_14846);
xnor UO_837 (O_837,N_14892,N_14882);
nor UO_838 (O_838,N_14767,N_14939);
nand UO_839 (O_839,N_14878,N_14792);
xnor UO_840 (O_840,N_14774,N_14881);
and UO_841 (O_841,N_14853,N_14837);
or UO_842 (O_842,N_14751,N_14769);
nand UO_843 (O_843,N_14822,N_14783);
nand UO_844 (O_844,N_14934,N_14990);
xor UO_845 (O_845,N_14928,N_14889);
nor UO_846 (O_846,N_14819,N_14925);
nand UO_847 (O_847,N_14806,N_14982);
or UO_848 (O_848,N_14983,N_14875);
nor UO_849 (O_849,N_14801,N_14837);
nand UO_850 (O_850,N_14956,N_14920);
nor UO_851 (O_851,N_14944,N_14917);
or UO_852 (O_852,N_14956,N_14751);
nand UO_853 (O_853,N_14760,N_14941);
nand UO_854 (O_854,N_14957,N_14897);
xnor UO_855 (O_855,N_14789,N_14997);
and UO_856 (O_856,N_14778,N_14997);
and UO_857 (O_857,N_14875,N_14834);
and UO_858 (O_858,N_14844,N_14854);
or UO_859 (O_859,N_14916,N_14853);
nor UO_860 (O_860,N_14831,N_14824);
xnor UO_861 (O_861,N_14802,N_14973);
nor UO_862 (O_862,N_14825,N_14784);
xnor UO_863 (O_863,N_14823,N_14985);
or UO_864 (O_864,N_14903,N_14947);
nand UO_865 (O_865,N_14781,N_14808);
xor UO_866 (O_866,N_14771,N_14809);
and UO_867 (O_867,N_14807,N_14855);
or UO_868 (O_868,N_14754,N_14757);
or UO_869 (O_869,N_14925,N_14949);
xnor UO_870 (O_870,N_14968,N_14880);
or UO_871 (O_871,N_14845,N_14782);
and UO_872 (O_872,N_14865,N_14850);
nand UO_873 (O_873,N_14990,N_14776);
and UO_874 (O_874,N_14920,N_14810);
nand UO_875 (O_875,N_14931,N_14754);
or UO_876 (O_876,N_14860,N_14796);
nand UO_877 (O_877,N_14951,N_14968);
nor UO_878 (O_878,N_14890,N_14891);
or UO_879 (O_879,N_14750,N_14867);
nor UO_880 (O_880,N_14888,N_14940);
nand UO_881 (O_881,N_14882,N_14879);
or UO_882 (O_882,N_14805,N_14931);
xnor UO_883 (O_883,N_14975,N_14912);
and UO_884 (O_884,N_14909,N_14852);
nor UO_885 (O_885,N_14791,N_14858);
and UO_886 (O_886,N_14994,N_14883);
nor UO_887 (O_887,N_14777,N_14764);
or UO_888 (O_888,N_14843,N_14927);
nand UO_889 (O_889,N_14792,N_14874);
nor UO_890 (O_890,N_14960,N_14886);
xor UO_891 (O_891,N_14842,N_14922);
xor UO_892 (O_892,N_14779,N_14942);
or UO_893 (O_893,N_14935,N_14918);
and UO_894 (O_894,N_14859,N_14836);
nor UO_895 (O_895,N_14998,N_14888);
or UO_896 (O_896,N_14894,N_14975);
nand UO_897 (O_897,N_14927,N_14802);
and UO_898 (O_898,N_14943,N_14789);
or UO_899 (O_899,N_14933,N_14848);
and UO_900 (O_900,N_14829,N_14807);
nor UO_901 (O_901,N_14795,N_14939);
and UO_902 (O_902,N_14820,N_14916);
nand UO_903 (O_903,N_14877,N_14858);
or UO_904 (O_904,N_14754,N_14956);
or UO_905 (O_905,N_14888,N_14961);
nor UO_906 (O_906,N_14971,N_14982);
nand UO_907 (O_907,N_14934,N_14929);
or UO_908 (O_908,N_14966,N_14943);
and UO_909 (O_909,N_14975,N_14879);
or UO_910 (O_910,N_14794,N_14927);
or UO_911 (O_911,N_14954,N_14782);
nor UO_912 (O_912,N_14932,N_14858);
or UO_913 (O_913,N_14937,N_14788);
nand UO_914 (O_914,N_14970,N_14962);
xor UO_915 (O_915,N_14758,N_14983);
or UO_916 (O_916,N_14998,N_14841);
nor UO_917 (O_917,N_14882,N_14844);
and UO_918 (O_918,N_14795,N_14889);
nor UO_919 (O_919,N_14985,N_14926);
and UO_920 (O_920,N_14825,N_14971);
xnor UO_921 (O_921,N_14869,N_14828);
nand UO_922 (O_922,N_14970,N_14997);
or UO_923 (O_923,N_14786,N_14777);
or UO_924 (O_924,N_14874,N_14826);
or UO_925 (O_925,N_14864,N_14774);
xor UO_926 (O_926,N_14783,N_14756);
and UO_927 (O_927,N_14882,N_14895);
xor UO_928 (O_928,N_14934,N_14948);
nand UO_929 (O_929,N_14905,N_14878);
xor UO_930 (O_930,N_14788,N_14901);
and UO_931 (O_931,N_14811,N_14900);
nand UO_932 (O_932,N_14984,N_14870);
xnor UO_933 (O_933,N_14943,N_14838);
and UO_934 (O_934,N_14828,N_14994);
and UO_935 (O_935,N_14950,N_14942);
nand UO_936 (O_936,N_14882,N_14828);
or UO_937 (O_937,N_14902,N_14877);
and UO_938 (O_938,N_14868,N_14902);
and UO_939 (O_939,N_14902,N_14757);
nor UO_940 (O_940,N_14762,N_14899);
and UO_941 (O_941,N_14796,N_14801);
or UO_942 (O_942,N_14868,N_14913);
nand UO_943 (O_943,N_14919,N_14780);
nor UO_944 (O_944,N_14960,N_14854);
xor UO_945 (O_945,N_14893,N_14898);
nor UO_946 (O_946,N_14782,N_14854);
or UO_947 (O_947,N_14876,N_14766);
and UO_948 (O_948,N_14978,N_14846);
nor UO_949 (O_949,N_14950,N_14989);
nor UO_950 (O_950,N_14792,N_14872);
nand UO_951 (O_951,N_14889,N_14925);
nor UO_952 (O_952,N_14926,N_14976);
nor UO_953 (O_953,N_14865,N_14770);
and UO_954 (O_954,N_14815,N_14981);
and UO_955 (O_955,N_14808,N_14871);
or UO_956 (O_956,N_14947,N_14963);
xor UO_957 (O_957,N_14905,N_14754);
nor UO_958 (O_958,N_14974,N_14975);
nand UO_959 (O_959,N_14956,N_14832);
xnor UO_960 (O_960,N_14802,N_14798);
and UO_961 (O_961,N_14949,N_14964);
or UO_962 (O_962,N_14895,N_14855);
and UO_963 (O_963,N_14826,N_14954);
or UO_964 (O_964,N_14772,N_14885);
nor UO_965 (O_965,N_14775,N_14897);
nand UO_966 (O_966,N_14923,N_14787);
nand UO_967 (O_967,N_14944,N_14886);
nor UO_968 (O_968,N_14869,N_14992);
nand UO_969 (O_969,N_14900,N_14910);
xnor UO_970 (O_970,N_14805,N_14872);
or UO_971 (O_971,N_14772,N_14851);
or UO_972 (O_972,N_14884,N_14771);
xor UO_973 (O_973,N_14879,N_14984);
or UO_974 (O_974,N_14815,N_14891);
nand UO_975 (O_975,N_14869,N_14781);
nor UO_976 (O_976,N_14910,N_14836);
nand UO_977 (O_977,N_14778,N_14764);
and UO_978 (O_978,N_14816,N_14890);
or UO_979 (O_979,N_14961,N_14905);
or UO_980 (O_980,N_14888,N_14855);
nand UO_981 (O_981,N_14945,N_14826);
nand UO_982 (O_982,N_14987,N_14892);
or UO_983 (O_983,N_14786,N_14776);
or UO_984 (O_984,N_14753,N_14823);
nor UO_985 (O_985,N_14944,N_14953);
nor UO_986 (O_986,N_14862,N_14990);
xor UO_987 (O_987,N_14983,N_14751);
and UO_988 (O_988,N_14930,N_14822);
and UO_989 (O_989,N_14795,N_14995);
nand UO_990 (O_990,N_14834,N_14815);
nor UO_991 (O_991,N_14835,N_14838);
or UO_992 (O_992,N_14888,N_14925);
nand UO_993 (O_993,N_14897,N_14837);
and UO_994 (O_994,N_14832,N_14918);
xor UO_995 (O_995,N_14962,N_14990);
xor UO_996 (O_996,N_14864,N_14996);
nand UO_997 (O_997,N_14952,N_14790);
nand UO_998 (O_998,N_14969,N_14947);
and UO_999 (O_999,N_14841,N_14769);
nand UO_1000 (O_1000,N_14856,N_14986);
and UO_1001 (O_1001,N_14754,N_14832);
xor UO_1002 (O_1002,N_14807,N_14826);
nor UO_1003 (O_1003,N_14939,N_14797);
or UO_1004 (O_1004,N_14892,N_14815);
nor UO_1005 (O_1005,N_14857,N_14848);
xnor UO_1006 (O_1006,N_14795,N_14902);
xor UO_1007 (O_1007,N_14814,N_14800);
xor UO_1008 (O_1008,N_14930,N_14893);
and UO_1009 (O_1009,N_14991,N_14960);
or UO_1010 (O_1010,N_14943,N_14896);
and UO_1011 (O_1011,N_14986,N_14866);
nand UO_1012 (O_1012,N_14773,N_14865);
nor UO_1013 (O_1013,N_14891,N_14922);
and UO_1014 (O_1014,N_14970,N_14833);
or UO_1015 (O_1015,N_14919,N_14761);
or UO_1016 (O_1016,N_14925,N_14857);
nand UO_1017 (O_1017,N_14776,N_14846);
and UO_1018 (O_1018,N_14776,N_14945);
nor UO_1019 (O_1019,N_14910,N_14773);
nand UO_1020 (O_1020,N_14920,N_14825);
or UO_1021 (O_1021,N_14789,N_14842);
nor UO_1022 (O_1022,N_14764,N_14758);
or UO_1023 (O_1023,N_14932,N_14786);
nand UO_1024 (O_1024,N_14811,N_14961);
xnor UO_1025 (O_1025,N_14949,N_14939);
xor UO_1026 (O_1026,N_14990,N_14935);
and UO_1027 (O_1027,N_14822,N_14826);
xor UO_1028 (O_1028,N_14798,N_14904);
nand UO_1029 (O_1029,N_14942,N_14775);
nor UO_1030 (O_1030,N_14939,N_14837);
nand UO_1031 (O_1031,N_14946,N_14776);
nand UO_1032 (O_1032,N_14891,N_14801);
xor UO_1033 (O_1033,N_14794,N_14779);
nor UO_1034 (O_1034,N_14990,N_14906);
or UO_1035 (O_1035,N_14887,N_14879);
nor UO_1036 (O_1036,N_14792,N_14766);
or UO_1037 (O_1037,N_14850,N_14992);
nor UO_1038 (O_1038,N_14779,N_14944);
xnor UO_1039 (O_1039,N_14870,N_14783);
or UO_1040 (O_1040,N_14816,N_14855);
or UO_1041 (O_1041,N_14928,N_14903);
and UO_1042 (O_1042,N_14818,N_14801);
nand UO_1043 (O_1043,N_14978,N_14788);
and UO_1044 (O_1044,N_14774,N_14819);
and UO_1045 (O_1045,N_14766,N_14955);
and UO_1046 (O_1046,N_14987,N_14862);
and UO_1047 (O_1047,N_14756,N_14807);
nor UO_1048 (O_1048,N_14802,N_14999);
nand UO_1049 (O_1049,N_14991,N_14995);
or UO_1050 (O_1050,N_14973,N_14759);
nor UO_1051 (O_1051,N_14902,N_14901);
xor UO_1052 (O_1052,N_14861,N_14965);
nor UO_1053 (O_1053,N_14778,N_14931);
and UO_1054 (O_1054,N_14755,N_14804);
and UO_1055 (O_1055,N_14985,N_14846);
nand UO_1056 (O_1056,N_14888,N_14919);
nor UO_1057 (O_1057,N_14817,N_14972);
nand UO_1058 (O_1058,N_14793,N_14812);
nand UO_1059 (O_1059,N_14844,N_14786);
xnor UO_1060 (O_1060,N_14959,N_14907);
nor UO_1061 (O_1061,N_14952,N_14996);
nor UO_1062 (O_1062,N_14764,N_14826);
nor UO_1063 (O_1063,N_14787,N_14783);
nor UO_1064 (O_1064,N_14818,N_14908);
nand UO_1065 (O_1065,N_14928,N_14789);
and UO_1066 (O_1066,N_14855,N_14841);
nand UO_1067 (O_1067,N_14923,N_14812);
and UO_1068 (O_1068,N_14908,N_14771);
and UO_1069 (O_1069,N_14800,N_14857);
nand UO_1070 (O_1070,N_14968,N_14999);
xnor UO_1071 (O_1071,N_14850,N_14912);
xor UO_1072 (O_1072,N_14845,N_14811);
nor UO_1073 (O_1073,N_14750,N_14864);
or UO_1074 (O_1074,N_14989,N_14976);
nor UO_1075 (O_1075,N_14971,N_14830);
and UO_1076 (O_1076,N_14815,N_14873);
and UO_1077 (O_1077,N_14861,N_14815);
or UO_1078 (O_1078,N_14915,N_14841);
and UO_1079 (O_1079,N_14775,N_14831);
xor UO_1080 (O_1080,N_14920,N_14895);
xor UO_1081 (O_1081,N_14806,N_14786);
and UO_1082 (O_1082,N_14918,N_14960);
nand UO_1083 (O_1083,N_14998,N_14825);
nor UO_1084 (O_1084,N_14753,N_14776);
or UO_1085 (O_1085,N_14983,N_14933);
nand UO_1086 (O_1086,N_14981,N_14787);
nand UO_1087 (O_1087,N_14771,N_14939);
nor UO_1088 (O_1088,N_14789,N_14761);
nand UO_1089 (O_1089,N_14865,N_14880);
and UO_1090 (O_1090,N_14962,N_14773);
xor UO_1091 (O_1091,N_14936,N_14794);
nor UO_1092 (O_1092,N_14971,N_14750);
and UO_1093 (O_1093,N_14779,N_14830);
nand UO_1094 (O_1094,N_14943,N_14905);
xor UO_1095 (O_1095,N_14874,N_14996);
xnor UO_1096 (O_1096,N_14938,N_14952);
nor UO_1097 (O_1097,N_14977,N_14930);
or UO_1098 (O_1098,N_14833,N_14918);
nand UO_1099 (O_1099,N_14773,N_14897);
or UO_1100 (O_1100,N_14791,N_14845);
nand UO_1101 (O_1101,N_14916,N_14787);
or UO_1102 (O_1102,N_14892,N_14900);
and UO_1103 (O_1103,N_14886,N_14779);
xor UO_1104 (O_1104,N_14879,N_14829);
and UO_1105 (O_1105,N_14858,N_14756);
or UO_1106 (O_1106,N_14945,N_14956);
nor UO_1107 (O_1107,N_14818,N_14925);
nand UO_1108 (O_1108,N_14996,N_14781);
and UO_1109 (O_1109,N_14897,N_14939);
or UO_1110 (O_1110,N_14876,N_14751);
nor UO_1111 (O_1111,N_14897,N_14835);
or UO_1112 (O_1112,N_14980,N_14806);
nor UO_1113 (O_1113,N_14935,N_14778);
xor UO_1114 (O_1114,N_14920,N_14852);
nor UO_1115 (O_1115,N_14763,N_14978);
nor UO_1116 (O_1116,N_14942,N_14761);
or UO_1117 (O_1117,N_14868,N_14901);
and UO_1118 (O_1118,N_14802,N_14966);
nor UO_1119 (O_1119,N_14781,N_14780);
and UO_1120 (O_1120,N_14802,N_14809);
nand UO_1121 (O_1121,N_14960,N_14893);
nor UO_1122 (O_1122,N_14915,N_14805);
and UO_1123 (O_1123,N_14943,N_14862);
nor UO_1124 (O_1124,N_14762,N_14878);
nand UO_1125 (O_1125,N_14805,N_14966);
or UO_1126 (O_1126,N_14853,N_14986);
nand UO_1127 (O_1127,N_14885,N_14952);
and UO_1128 (O_1128,N_14907,N_14977);
nand UO_1129 (O_1129,N_14753,N_14869);
and UO_1130 (O_1130,N_14867,N_14858);
xnor UO_1131 (O_1131,N_14929,N_14933);
or UO_1132 (O_1132,N_14813,N_14952);
nor UO_1133 (O_1133,N_14751,N_14893);
nor UO_1134 (O_1134,N_14950,N_14961);
and UO_1135 (O_1135,N_14822,N_14871);
nand UO_1136 (O_1136,N_14963,N_14926);
and UO_1137 (O_1137,N_14987,N_14904);
xnor UO_1138 (O_1138,N_14814,N_14931);
nand UO_1139 (O_1139,N_14787,N_14910);
and UO_1140 (O_1140,N_14952,N_14828);
or UO_1141 (O_1141,N_14768,N_14845);
xnor UO_1142 (O_1142,N_14954,N_14899);
xnor UO_1143 (O_1143,N_14981,N_14858);
or UO_1144 (O_1144,N_14886,N_14841);
nor UO_1145 (O_1145,N_14845,N_14780);
nand UO_1146 (O_1146,N_14775,N_14774);
xnor UO_1147 (O_1147,N_14950,N_14943);
nand UO_1148 (O_1148,N_14926,N_14851);
and UO_1149 (O_1149,N_14981,N_14806);
nand UO_1150 (O_1150,N_14854,N_14999);
nand UO_1151 (O_1151,N_14940,N_14890);
xnor UO_1152 (O_1152,N_14808,N_14841);
or UO_1153 (O_1153,N_14923,N_14960);
xor UO_1154 (O_1154,N_14954,N_14894);
nand UO_1155 (O_1155,N_14847,N_14873);
or UO_1156 (O_1156,N_14850,N_14962);
nor UO_1157 (O_1157,N_14942,N_14804);
nand UO_1158 (O_1158,N_14804,N_14752);
xor UO_1159 (O_1159,N_14968,N_14800);
or UO_1160 (O_1160,N_14930,N_14793);
and UO_1161 (O_1161,N_14973,N_14950);
nor UO_1162 (O_1162,N_14838,N_14907);
nor UO_1163 (O_1163,N_14870,N_14757);
and UO_1164 (O_1164,N_14900,N_14995);
nand UO_1165 (O_1165,N_14818,N_14777);
and UO_1166 (O_1166,N_14943,N_14918);
or UO_1167 (O_1167,N_14891,N_14778);
or UO_1168 (O_1168,N_14820,N_14965);
nand UO_1169 (O_1169,N_14798,N_14756);
or UO_1170 (O_1170,N_14795,N_14963);
or UO_1171 (O_1171,N_14771,N_14965);
nand UO_1172 (O_1172,N_14947,N_14793);
nand UO_1173 (O_1173,N_14828,N_14768);
nor UO_1174 (O_1174,N_14918,N_14874);
nor UO_1175 (O_1175,N_14790,N_14880);
xnor UO_1176 (O_1176,N_14914,N_14801);
and UO_1177 (O_1177,N_14780,N_14954);
xnor UO_1178 (O_1178,N_14964,N_14915);
or UO_1179 (O_1179,N_14827,N_14786);
nor UO_1180 (O_1180,N_14875,N_14784);
nand UO_1181 (O_1181,N_14880,N_14860);
nand UO_1182 (O_1182,N_14830,N_14818);
xnor UO_1183 (O_1183,N_14826,N_14819);
nand UO_1184 (O_1184,N_14863,N_14777);
and UO_1185 (O_1185,N_14952,N_14797);
nor UO_1186 (O_1186,N_14901,N_14780);
and UO_1187 (O_1187,N_14872,N_14962);
or UO_1188 (O_1188,N_14878,N_14924);
nand UO_1189 (O_1189,N_14838,N_14753);
and UO_1190 (O_1190,N_14952,N_14857);
nor UO_1191 (O_1191,N_14778,N_14863);
xnor UO_1192 (O_1192,N_14951,N_14894);
nor UO_1193 (O_1193,N_14823,N_14814);
nor UO_1194 (O_1194,N_14946,N_14975);
nor UO_1195 (O_1195,N_14818,N_14996);
xnor UO_1196 (O_1196,N_14778,N_14865);
nor UO_1197 (O_1197,N_14850,N_14960);
and UO_1198 (O_1198,N_14831,N_14943);
nor UO_1199 (O_1199,N_14901,N_14873);
and UO_1200 (O_1200,N_14825,N_14885);
nand UO_1201 (O_1201,N_14808,N_14805);
nand UO_1202 (O_1202,N_14838,N_14786);
xnor UO_1203 (O_1203,N_14929,N_14919);
nand UO_1204 (O_1204,N_14920,N_14804);
nand UO_1205 (O_1205,N_14766,N_14858);
nor UO_1206 (O_1206,N_14823,N_14802);
nand UO_1207 (O_1207,N_14759,N_14760);
nand UO_1208 (O_1208,N_14868,N_14811);
or UO_1209 (O_1209,N_14990,N_14964);
nand UO_1210 (O_1210,N_14801,N_14942);
nand UO_1211 (O_1211,N_14763,N_14962);
or UO_1212 (O_1212,N_14954,N_14976);
or UO_1213 (O_1213,N_14837,N_14943);
nor UO_1214 (O_1214,N_14833,N_14865);
nor UO_1215 (O_1215,N_14775,N_14819);
nand UO_1216 (O_1216,N_14953,N_14851);
or UO_1217 (O_1217,N_14833,N_14976);
or UO_1218 (O_1218,N_14930,N_14944);
and UO_1219 (O_1219,N_14922,N_14832);
nand UO_1220 (O_1220,N_14757,N_14930);
nor UO_1221 (O_1221,N_14970,N_14936);
nand UO_1222 (O_1222,N_14918,N_14992);
xor UO_1223 (O_1223,N_14819,N_14802);
nand UO_1224 (O_1224,N_14898,N_14855);
nand UO_1225 (O_1225,N_14864,N_14976);
nand UO_1226 (O_1226,N_14892,N_14925);
xor UO_1227 (O_1227,N_14948,N_14898);
nor UO_1228 (O_1228,N_14930,N_14839);
nor UO_1229 (O_1229,N_14891,N_14989);
and UO_1230 (O_1230,N_14921,N_14866);
nor UO_1231 (O_1231,N_14784,N_14978);
nand UO_1232 (O_1232,N_14962,N_14769);
or UO_1233 (O_1233,N_14827,N_14879);
and UO_1234 (O_1234,N_14874,N_14795);
and UO_1235 (O_1235,N_14971,N_14915);
and UO_1236 (O_1236,N_14875,N_14962);
nor UO_1237 (O_1237,N_14947,N_14761);
nor UO_1238 (O_1238,N_14798,N_14772);
or UO_1239 (O_1239,N_14812,N_14795);
or UO_1240 (O_1240,N_14954,N_14798);
or UO_1241 (O_1241,N_14813,N_14892);
and UO_1242 (O_1242,N_14896,N_14979);
and UO_1243 (O_1243,N_14928,N_14817);
xnor UO_1244 (O_1244,N_14764,N_14848);
and UO_1245 (O_1245,N_14839,N_14911);
or UO_1246 (O_1246,N_14907,N_14908);
nor UO_1247 (O_1247,N_14936,N_14858);
nor UO_1248 (O_1248,N_14968,N_14803);
nand UO_1249 (O_1249,N_14927,N_14782);
nor UO_1250 (O_1250,N_14753,N_14913);
nor UO_1251 (O_1251,N_14828,N_14863);
nand UO_1252 (O_1252,N_14838,N_14956);
nand UO_1253 (O_1253,N_14893,N_14848);
and UO_1254 (O_1254,N_14787,N_14782);
and UO_1255 (O_1255,N_14895,N_14870);
nor UO_1256 (O_1256,N_14789,N_14768);
or UO_1257 (O_1257,N_14890,N_14829);
nand UO_1258 (O_1258,N_14913,N_14850);
nor UO_1259 (O_1259,N_14851,N_14840);
and UO_1260 (O_1260,N_14801,N_14846);
xnor UO_1261 (O_1261,N_14846,N_14911);
or UO_1262 (O_1262,N_14994,N_14964);
xor UO_1263 (O_1263,N_14954,N_14771);
nand UO_1264 (O_1264,N_14873,N_14860);
nand UO_1265 (O_1265,N_14893,N_14932);
and UO_1266 (O_1266,N_14923,N_14789);
or UO_1267 (O_1267,N_14820,N_14783);
or UO_1268 (O_1268,N_14925,N_14880);
or UO_1269 (O_1269,N_14883,N_14957);
or UO_1270 (O_1270,N_14996,N_14926);
nor UO_1271 (O_1271,N_14780,N_14765);
nor UO_1272 (O_1272,N_14943,N_14785);
or UO_1273 (O_1273,N_14964,N_14989);
and UO_1274 (O_1274,N_14994,N_14879);
or UO_1275 (O_1275,N_14901,N_14770);
nor UO_1276 (O_1276,N_14751,N_14827);
nor UO_1277 (O_1277,N_14968,N_14994);
xnor UO_1278 (O_1278,N_14948,N_14813);
and UO_1279 (O_1279,N_14756,N_14909);
nand UO_1280 (O_1280,N_14832,N_14875);
xor UO_1281 (O_1281,N_14843,N_14892);
or UO_1282 (O_1282,N_14761,N_14804);
and UO_1283 (O_1283,N_14814,N_14981);
or UO_1284 (O_1284,N_14855,N_14944);
nor UO_1285 (O_1285,N_14868,N_14754);
nand UO_1286 (O_1286,N_14752,N_14970);
and UO_1287 (O_1287,N_14963,N_14826);
and UO_1288 (O_1288,N_14911,N_14756);
nand UO_1289 (O_1289,N_14840,N_14768);
nand UO_1290 (O_1290,N_14898,N_14966);
nand UO_1291 (O_1291,N_14961,N_14817);
nand UO_1292 (O_1292,N_14949,N_14843);
nand UO_1293 (O_1293,N_14939,N_14872);
xnor UO_1294 (O_1294,N_14881,N_14962);
xor UO_1295 (O_1295,N_14938,N_14815);
xor UO_1296 (O_1296,N_14980,N_14799);
nor UO_1297 (O_1297,N_14892,N_14833);
nor UO_1298 (O_1298,N_14999,N_14958);
or UO_1299 (O_1299,N_14831,N_14820);
xor UO_1300 (O_1300,N_14866,N_14910);
xnor UO_1301 (O_1301,N_14930,N_14847);
nor UO_1302 (O_1302,N_14964,N_14854);
nor UO_1303 (O_1303,N_14896,N_14883);
and UO_1304 (O_1304,N_14773,N_14984);
nand UO_1305 (O_1305,N_14955,N_14857);
xor UO_1306 (O_1306,N_14892,N_14787);
and UO_1307 (O_1307,N_14968,N_14925);
nand UO_1308 (O_1308,N_14843,N_14995);
nand UO_1309 (O_1309,N_14855,N_14774);
and UO_1310 (O_1310,N_14948,N_14956);
nand UO_1311 (O_1311,N_14947,N_14924);
or UO_1312 (O_1312,N_14978,N_14811);
or UO_1313 (O_1313,N_14994,N_14773);
or UO_1314 (O_1314,N_14875,N_14801);
xnor UO_1315 (O_1315,N_14917,N_14892);
nor UO_1316 (O_1316,N_14837,N_14942);
nand UO_1317 (O_1317,N_14954,N_14912);
nor UO_1318 (O_1318,N_14813,N_14916);
xnor UO_1319 (O_1319,N_14797,N_14950);
and UO_1320 (O_1320,N_14893,N_14804);
or UO_1321 (O_1321,N_14944,N_14996);
nand UO_1322 (O_1322,N_14828,N_14866);
nor UO_1323 (O_1323,N_14999,N_14830);
xor UO_1324 (O_1324,N_14935,N_14940);
and UO_1325 (O_1325,N_14981,N_14867);
or UO_1326 (O_1326,N_14877,N_14761);
xor UO_1327 (O_1327,N_14894,N_14927);
xor UO_1328 (O_1328,N_14915,N_14814);
nand UO_1329 (O_1329,N_14923,N_14978);
nor UO_1330 (O_1330,N_14916,N_14992);
nand UO_1331 (O_1331,N_14996,N_14889);
and UO_1332 (O_1332,N_14930,N_14981);
nor UO_1333 (O_1333,N_14784,N_14918);
nand UO_1334 (O_1334,N_14753,N_14918);
nand UO_1335 (O_1335,N_14889,N_14960);
and UO_1336 (O_1336,N_14983,N_14925);
xor UO_1337 (O_1337,N_14758,N_14975);
nor UO_1338 (O_1338,N_14896,N_14853);
nor UO_1339 (O_1339,N_14864,N_14960);
nand UO_1340 (O_1340,N_14955,N_14794);
or UO_1341 (O_1341,N_14882,N_14764);
nand UO_1342 (O_1342,N_14778,N_14881);
nor UO_1343 (O_1343,N_14900,N_14894);
nor UO_1344 (O_1344,N_14846,N_14887);
nand UO_1345 (O_1345,N_14811,N_14821);
nor UO_1346 (O_1346,N_14933,N_14949);
xor UO_1347 (O_1347,N_14944,N_14985);
and UO_1348 (O_1348,N_14795,N_14918);
nand UO_1349 (O_1349,N_14850,N_14888);
xor UO_1350 (O_1350,N_14877,N_14893);
nor UO_1351 (O_1351,N_14874,N_14952);
nand UO_1352 (O_1352,N_14832,N_14925);
nand UO_1353 (O_1353,N_14947,N_14950);
and UO_1354 (O_1354,N_14847,N_14750);
and UO_1355 (O_1355,N_14787,N_14811);
and UO_1356 (O_1356,N_14798,N_14857);
and UO_1357 (O_1357,N_14988,N_14869);
nand UO_1358 (O_1358,N_14818,N_14994);
or UO_1359 (O_1359,N_14895,N_14842);
xor UO_1360 (O_1360,N_14998,N_14788);
xnor UO_1361 (O_1361,N_14832,N_14936);
xor UO_1362 (O_1362,N_14789,N_14958);
or UO_1363 (O_1363,N_14794,N_14802);
nand UO_1364 (O_1364,N_14886,N_14755);
xnor UO_1365 (O_1365,N_14993,N_14793);
nand UO_1366 (O_1366,N_14928,N_14937);
and UO_1367 (O_1367,N_14838,N_14759);
and UO_1368 (O_1368,N_14904,N_14771);
and UO_1369 (O_1369,N_14842,N_14904);
or UO_1370 (O_1370,N_14928,N_14948);
or UO_1371 (O_1371,N_14773,N_14975);
nand UO_1372 (O_1372,N_14842,N_14896);
nor UO_1373 (O_1373,N_14832,N_14785);
or UO_1374 (O_1374,N_14996,N_14900);
and UO_1375 (O_1375,N_14875,N_14786);
nand UO_1376 (O_1376,N_14860,N_14941);
and UO_1377 (O_1377,N_14952,N_14907);
nor UO_1378 (O_1378,N_14793,N_14813);
nand UO_1379 (O_1379,N_14939,N_14916);
nor UO_1380 (O_1380,N_14919,N_14771);
or UO_1381 (O_1381,N_14764,N_14841);
nor UO_1382 (O_1382,N_14807,N_14870);
xor UO_1383 (O_1383,N_14958,N_14802);
or UO_1384 (O_1384,N_14919,N_14979);
or UO_1385 (O_1385,N_14880,N_14949);
and UO_1386 (O_1386,N_14812,N_14977);
nand UO_1387 (O_1387,N_14878,N_14862);
xnor UO_1388 (O_1388,N_14954,N_14754);
and UO_1389 (O_1389,N_14791,N_14984);
nand UO_1390 (O_1390,N_14753,N_14835);
nor UO_1391 (O_1391,N_14965,N_14910);
and UO_1392 (O_1392,N_14790,N_14810);
nand UO_1393 (O_1393,N_14980,N_14852);
nand UO_1394 (O_1394,N_14904,N_14870);
or UO_1395 (O_1395,N_14856,N_14782);
or UO_1396 (O_1396,N_14796,N_14779);
and UO_1397 (O_1397,N_14871,N_14954);
xor UO_1398 (O_1398,N_14771,N_14758);
nor UO_1399 (O_1399,N_14907,N_14786);
xnor UO_1400 (O_1400,N_14881,N_14932);
nand UO_1401 (O_1401,N_14868,N_14799);
nand UO_1402 (O_1402,N_14958,N_14752);
or UO_1403 (O_1403,N_14789,N_14826);
and UO_1404 (O_1404,N_14862,N_14898);
or UO_1405 (O_1405,N_14770,N_14868);
or UO_1406 (O_1406,N_14834,N_14884);
and UO_1407 (O_1407,N_14870,N_14943);
nor UO_1408 (O_1408,N_14975,N_14885);
and UO_1409 (O_1409,N_14768,N_14812);
nor UO_1410 (O_1410,N_14987,N_14923);
nand UO_1411 (O_1411,N_14991,N_14820);
nand UO_1412 (O_1412,N_14803,N_14814);
or UO_1413 (O_1413,N_14846,N_14894);
nand UO_1414 (O_1414,N_14977,N_14782);
or UO_1415 (O_1415,N_14943,N_14798);
nand UO_1416 (O_1416,N_14842,N_14899);
nor UO_1417 (O_1417,N_14917,N_14987);
nand UO_1418 (O_1418,N_14763,N_14952);
nor UO_1419 (O_1419,N_14801,N_14989);
or UO_1420 (O_1420,N_14955,N_14831);
nor UO_1421 (O_1421,N_14854,N_14893);
or UO_1422 (O_1422,N_14812,N_14926);
nor UO_1423 (O_1423,N_14750,N_14972);
nor UO_1424 (O_1424,N_14859,N_14795);
xnor UO_1425 (O_1425,N_14999,N_14804);
nor UO_1426 (O_1426,N_14927,N_14862);
xnor UO_1427 (O_1427,N_14958,N_14882);
xnor UO_1428 (O_1428,N_14797,N_14898);
and UO_1429 (O_1429,N_14787,N_14948);
nor UO_1430 (O_1430,N_14894,N_14956);
nor UO_1431 (O_1431,N_14865,N_14767);
and UO_1432 (O_1432,N_14904,N_14810);
and UO_1433 (O_1433,N_14990,N_14871);
xnor UO_1434 (O_1434,N_14896,N_14903);
or UO_1435 (O_1435,N_14977,N_14994);
and UO_1436 (O_1436,N_14752,N_14839);
xor UO_1437 (O_1437,N_14863,N_14808);
or UO_1438 (O_1438,N_14768,N_14863);
xor UO_1439 (O_1439,N_14893,N_14760);
nor UO_1440 (O_1440,N_14981,N_14988);
nor UO_1441 (O_1441,N_14998,N_14819);
and UO_1442 (O_1442,N_14979,N_14839);
or UO_1443 (O_1443,N_14885,N_14928);
and UO_1444 (O_1444,N_14753,N_14756);
nor UO_1445 (O_1445,N_14759,N_14870);
nand UO_1446 (O_1446,N_14920,N_14925);
nor UO_1447 (O_1447,N_14938,N_14881);
nand UO_1448 (O_1448,N_14755,N_14850);
nand UO_1449 (O_1449,N_14889,N_14881);
nor UO_1450 (O_1450,N_14902,N_14838);
nand UO_1451 (O_1451,N_14941,N_14919);
and UO_1452 (O_1452,N_14912,N_14760);
nor UO_1453 (O_1453,N_14828,N_14908);
nand UO_1454 (O_1454,N_14866,N_14809);
nor UO_1455 (O_1455,N_14952,N_14850);
xnor UO_1456 (O_1456,N_14988,N_14794);
and UO_1457 (O_1457,N_14849,N_14976);
nor UO_1458 (O_1458,N_14782,N_14779);
nor UO_1459 (O_1459,N_14910,N_14831);
xnor UO_1460 (O_1460,N_14953,N_14958);
xnor UO_1461 (O_1461,N_14778,N_14803);
xnor UO_1462 (O_1462,N_14906,N_14838);
or UO_1463 (O_1463,N_14967,N_14834);
nand UO_1464 (O_1464,N_14783,N_14931);
or UO_1465 (O_1465,N_14867,N_14859);
and UO_1466 (O_1466,N_14828,N_14892);
and UO_1467 (O_1467,N_14907,N_14976);
xnor UO_1468 (O_1468,N_14937,N_14995);
or UO_1469 (O_1469,N_14961,N_14867);
nand UO_1470 (O_1470,N_14950,N_14924);
nor UO_1471 (O_1471,N_14822,N_14879);
nand UO_1472 (O_1472,N_14849,N_14886);
and UO_1473 (O_1473,N_14919,N_14902);
nor UO_1474 (O_1474,N_14938,N_14950);
nor UO_1475 (O_1475,N_14828,N_14835);
or UO_1476 (O_1476,N_14971,N_14883);
xor UO_1477 (O_1477,N_14883,N_14785);
and UO_1478 (O_1478,N_14958,N_14759);
xnor UO_1479 (O_1479,N_14935,N_14929);
xor UO_1480 (O_1480,N_14862,N_14928);
and UO_1481 (O_1481,N_14876,N_14851);
nor UO_1482 (O_1482,N_14920,N_14864);
xnor UO_1483 (O_1483,N_14992,N_14879);
xnor UO_1484 (O_1484,N_14771,N_14853);
or UO_1485 (O_1485,N_14887,N_14806);
and UO_1486 (O_1486,N_14750,N_14780);
xnor UO_1487 (O_1487,N_14993,N_14957);
nand UO_1488 (O_1488,N_14993,N_14880);
nand UO_1489 (O_1489,N_14839,N_14934);
xor UO_1490 (O_1490,N_14892,N_14758);
nand UO_1491 (O_1491,N_14809,N_14976);
nand UO_1492 (O_1492,N_14969,N_14852);
or UO_1493 (O_1493,N_14856,N_14917);
nor UO_1494 (O_1494,N_14859,N_14898);
nand UO_1495 (O_1495,N_14991,N_14940);
nand UO_1496 (O_1496,N_14853,N_14808);
nand UO_1497 (O_1497,N_14955,N_14882);
nor UO_1498 (O_1498,N_14957,N_14815);
xor UO_1499 (O_1499,N_14808,N_14918);
nor UO_1500 (O_1500,N_14896,N_14858);
nand UO_1501 (O_1501,N_14958,N_14952);
nand UO_1502 (O_1502,N_14764,N_14809);
xnor UO_1503 (O_1503,N_14853,N_14817);
xor UO_1504 (O_1504,N_14831,N_14768);
and UO_1505 (O_1505,N_14883,N_14750);
nand UO_1506 (O_1506,N_14972,N_14870);
and UO_1507 (O_1507,N_14926,N_14905);
xnor UO_1508 (O_1508,N_14975,N_14812);
nor UO_1509 (O_1509,N_14802,N_14763);
and UO_1510 (O_1510,N_14798,N_14770);
or UO_1511 (O_1511,N_14894,N_14938);
or UO_1512 (O_1512,N_14792,N_14942);
nand UO_1513 (O_1513,N_14817,N_14849);
nor UO_1514 (O_1514,N_14979,N_14965);
nor UO_1515 (O_1515,N_14824,N_14924);
xnor UO_1516 (O_1516,N_14971,N_14914);
or UO_1517 (O_1517,N_14863,N_14899);
and UO_1518 (O_1518,N_14931,N_14893);
nand UO_1519 (O_1519,N_14978,N_14821);
or UO_1520 (O_1520,N_14828,N_14912);
nor UO_1521 (O_1521,N_14951,N_14789);
xnor UO_1522 (O_1522,N_14933,N_14926);
nor UO_1523 (O_1523,N_14783,N_14925);
nor UO_1524 (O_1524,N_14978,N_14773);
nand UO_1525 (O_1525,N_14967,N_14896);
or UO_1526 (O_1526,N_14761,N_14863);
and UO_1527 (O_1527,N_14873,N_14794);
and UO_1528 (O_1528,N_14998,N_14893);
or UO_1529 (O_1529,N_14770,N_14871);
xor UO_1530 (O_1530,N_14921,N_14855);
nand UO_1531 (O_1531,N_14805,N_14857);
nor UO_1532 (O_1532,N_14769,N_14950);
xnor UO_1533 (O_1533,N_14949,N_14830);
nand UO_1534 (O_1534,N_14754,N_14906);
nor UO_1535 (O_1535,N_14862,N_14977);
or UO_1536 (O_1536,N_14824,N_14772);
nor UO_1537 (O_1537,N_14912,N_14764);
or UO_1538 (O_1538,N_14854,N_14961);
xor UO_1539 (O_1539,N_14899,N_14778);
nor UO_1540 (O_1540,N_14895,N_14863);
nor UO_1541 (O_1541,N_14915,N_14803);
xor UO_1542 (O_1542,N_14858,N_14815);
nand UO_1543 (O_1543,N_14988,N_14942);
xor UO_1544 (O_1544,N_14803,N_14950);
and UO_1545 (O_1545,N_14879,N_14846);
and UO_1546 (O_1546,N_14770,N_14998);
or UO_1547 (O_1547,N_14972,N_14894);
xnor UO_1548 (O_1548,N_14760,N_14962);
nor UO_1549 (O_1549,N_14978,N_14761);
xor UO_1550 (O_1550,N_14872,N_14838);
nor UO_1551 (O_1551,N_14958,N_14803);
or UO_1552 (O_1552,N_14752,N_14986);
xor UO_1553 (O_1553,N_14973,N_14889);
xor UO_1554 (O_1554,N_14763,N_14901);
or UO_1555 (O_1555,N_14840,N_14890);
or UO_1556 (O_1556,N_14964,N_14868);
or UO_1557 (O_1557,N_14798,N_14969);
xnor UO_1558 (O_1558,N_14982,N_14860);
xnor UO_1559 (O_1559,N_14903,N_14921);
or UO_1560 (O_1560,N_14822,N_14913);
or UO_1561 (O_1561,N_14885,N_14967);
and UO_1562 (O_1562,N_14862,N_14777);
or UO_1563 (O_1563,N_14837,N_14857);
xnor UO_1564 (O_1564,N_14861,N_14972);
xor UO_1565 (O_1565,N_14823,N_14911);
nor UO_1566 (O_1566,N_14831,N_14948);
nand UO_1567 (O_1567,N_14942,N_14889);
nor UO_1568 (O_1568,N_14880,N_14899);
nor UO_1569 (O_1569,N_14992,N_14858);
nor UO_1570 (O_1570,N_14817,N_14830);
and UO_1571 (O_1571,N_14876,N_14909);
and UO_1572 (O_1572,N_14973,N_14927);
nor UO_1573 (O_1573,N_14988,N_14848);
nor UO_1574 (O_1574,N_14916,N_14794);
nand UO_1575 (O_1575,N_14913,N_14962);
xnor UO_1576 (O_1576,N_14911,N_14773);
nand UO_1577 (O_1577,N_14858,N_14879);
nand UO_1578 (O_1578,N_14804,N_14763);
and UO_1579 (O_1579,N_14877,N_14919);
nor UO_1580 (O_1580,N_14770,N_14765);
xnor UO_1581 (O_1581,N_14932,N_14820);
or UO_1582 (O_1582,N_14751,N_14886);
xnor UO_1583 (O_1583,N_14828,N_14856);
and UO_1584 (O_1584,N_14779,N_14792);
and UO_1585 (O_1585,N_14895,N_14891);
nand UO_1586 (O_1586,N_14857,N_14936);
nor UO_1587 (O_1587,N_14833,N_14947);
nand UO_1588 (O_1588,N_14945,N_14757);
and UO_1589 (O_1589,N_14945,N_14917);
xnor UO_1590 (O_1590,N_14825,N_14844);
or UO_1591 (O_1591,N_14842,N_14769);
nor UO_1592 (O_1592,N_14814,N_14822);
xnor UO_1593 (O_1593,N_14815,N_14878);
or UO_1594 (O_1594,N_14855,N_14922);
xnor UO_1595 (O_1595,N_14830,N_14845);
and UO_1596 (O_1596,N_14848,N_14755);
and UO_1597 (O_1597,N_14968,N_14947);
nor UO_1598 (O_1598,N_14796,N_14913);
and UO_1599 (O_1599,N_14945,N_14994);
nand UO_1600 (O_1600,N_14949,N_14790);
or UO_1601 (O_1601,N_14849,N_14807);
or UO_1602 (O_1602,N_14856,N_14929);
nand UO_1603 (O_1603,N_14823,N_14936);
and UO_1604 (O_1604,N_14940,N_14767);
and UO_1605 (O_1605,N_14977,N_14917);
xor UO_1606 (O_1606,N_14881,N_14950);
nor UO_1607 (O_1607,N_14934,N_14972);
and UO_1608 (O_1608,N_14832,N_14812);
nor UO_1609 (O_1609,N_14815,N_14978);
and UO_1610 (O_1610,N_14924,N_14942);
nor UO_1611 (O_1611,N_14954,N_14938);
nand UO_1612 (O_1612,N_14797,N_14985);
nand UO_1613 (O_1613,N_14801,N_14912);
nand UO_1614 (O_1614,N_14791,N_14780);
xnor UO_1615 (O_1615,N_14761,N_14941);
and UO_1616 (O_1616,N_14989,N_14752);
xnor UO_1617 (O_1617,N_14804,N_14924);
nor UO_1618 (O_1618,N_14814,N_14796);
xnor UO_1619 (O_1619,N_14910,N_14785);
nor UO_1620 (O_1620,N_14764,N_14955);
xnor UO_1621 (O_1621,N_14863,N_14878);
xnor UO_1622 (O_1622,N_14844,N_14921);
nand UO_1623 (O_1623,N_14814,N_14807);
nand UO_1624 (O_1624,N_14755,N_14763);
nor UO_1625 (O_1625,N_14774,N_14764);
or UO_1626 (O_1626,N_14982,N_14787);
and UO_1627 (O_1627,N_14769,N_14902);
nand UO_1628 (O_1628,N_14997,N_14963);
nand UO_1629 (O_1629,N_14986,N_14831);
xor UO_1630 (O_1630,N_14811,N_14785);
or UO_1631 (O_1631,N_14766,N_14967);
and UO_1632 (O_1632,N_14909,N_14965);
nand UO_1633 (O_1633,N_14753,N_14979);
and UO_1634 (O_1634,N_14959,N_14933);
nor UO_1635 (O_1635,N_14988,N_14776);
and UO_1636 (O_1636,N_14861,N_14846);
and UO_1637 (O_1637,N_14792,N_14845);
nor UO_1638 (O_1638,N_14930,N_14848);
or UO_1639 (O_1639,N_14906,N_14842);
and UO_1640 (O_1640,N_14872,N_14871);
or UO_1641 (O_1641,N_14765,N_14800);
nor UO_1642 (O_1642,N_14886,N_14808);
nor UO_1643 (O_1643,N_14848,N_14948);
and UO_1644 (O_1644,N_14832,N_14777);
and UO_1645 (O_1645,N_14895,N_14865);
or UO_1646 (O_1646,N_14877,N_14941);
or UO_1647 (O_1647,N_14928,N_14751);
xnor UO_1648 (O_1648,N_14878,N_14824);
xnor UO_1649 (O_1649,N_14939,N_14995);
or UO_1650 (O_1650,N_14937,N_14780);
and UO_1651 (O_1651,N_14883,N_14878);
nor UO_1652 (O_1652,N_14822,N_14872);
or UO_1653 (O_1653,N_14779,N_14993);
and UO_1654 (O_1654,N_14932,N_14978);
or UO_1655 (O_1655,N_14841,N_14937);
nand UO_1656 (O_1656,N_14807,N_14920);
nand UO_1657 (O_1657,N_14786,N_14956);
nor UO_1658 (O_1658,N_14989,N_14906);
nand UO_1659 (O_1659,N_14874,N_14886);
nor UO_1660 (O_1660,N_14943,N_14977);
nand UO_1661 (O_1661,N_14780,N_14867);
and UO_1662 (O_1662,N_14929,N_14985);
xnor UO_1663 (O_1663,N_14977,N_14950);
nor UO_1664 (O_1664,N_14880,N_14835);
xor UO_1665 (O_1665,N_14954,N_14874);
nor UO_1666 (O_1666,N_14991,N_14888);
and UO_1667 (O_1667,N_14950,N_14955);
nor UO_1668 (O_1668,N_14845,N_14770);
nand UO_1669 (O_1669,N_14952,N_14947);
or UO_1670 (O_1670,N_14950,N_14802);
and UO_1671 (O_1671,N_14930,N_14760);
xnor UO_1672 (O_1672,N_14858,N_14768);
nand UO_1673 (O_1673,N_14924,N_14944);
xor UO_1674 (O_1674,N_14956,N_14756);
nand UO_1675 (O_1675,N_14877,N_14927);
or UO_1676 (O_1676,N_14877,N_14838);
or UO_1677 (O_1677,N_14762,N_14919);
nand UO_1678 (O_1678,N_14899,N_14907);
or UO_1679 (O_1679,N_14926,N_14827);
or UO_1680 (O_1680,N_14756,N_14995);
nand UO_1681 (O_1681,N_14938,N_14918);
xor UO_1682 (O_1682,N_14785,N_14864);
nor UO_1683 (O_1683,N_14936,N_14885);
xor UO_1684 (O_1684,N_14877,N_14795);
or UO_1685 (O_1685,N_14833,N_14841);
or UO_1686 (O_1686,N_14942,N_14974);
or UO_1687 (O_1687,N_14873,N_14963);
or UO_1688 (O_1688,N_14968,N_14765);
nor UO_1689 (O_1689,N_14767,N_14887);
or UO_1690 (O_1690,N_14814,N_14768);
or UO_1691 (O_1691,N_14919,N_14807);
nor UO_1692 (O_1692,N_14844,N_14960);
or UO_1693 (O_1693,N_14889,N_14936);
nand UO_1694 (O_1694,N_14946,N_14805);
nand UO_1695 (O_1695,N_14994,N_14881);
nor UO_1696 (O_1696,N_14960,N_14992);
nor UO_1697 (O_1697,N_14894,N_14928);
nand UO_1698 (O_1698,N_14861,N_14898);
and UO_1699 (O_1699,N_14949,N_14827);
or UO_1700 (O_1700,N_14774,N_14773);
nand UO_1701 (O_1701,N_14952,N_14757);
or UO_1702 (O_1702,N_14898,N_14926);
xor UO_1703 (O_1703,N_14915,N_14901);
and UO_1704 (O_1704,N_14966,N_14998);
nand UO_1705 (O_1705,N_14854,N_14862);
nor UO_1706 (O_1706,N_14895,N_14862);
nor UO_1707 (O_1707,N_14816,N_14903);
nor UO_1708 (O_1708,N_14954,N_14958);
and UO_1709 (O_1709,N_14985,N_14901);
nor UO_1710 (O_1710,N_14809,N_14808);
nand UO_1711 (O_1711,N_14913,N_14887);
nor UO_1712 (O_1712,N_14916,N_14755);
xor UO_1713 (O_1713,N_14883,N_14975);
xnor UO_1714 (O_1714,N_14757,N_14866);
xnor UO_1715 (O_1715,N_14772,N_14799);
xnor UO_1716 (O_1716,N_14765,N_14958);
or UO_1717 (O_1717,N_14912,N_14904);
xor UO_1718 (O_1718,N_14920,N_14848);
nor UO_1719 (O_1719,N_14992,N_14947);
or UO_1720 (O_1720,N_14791,N_14963);
nand UO_1721 (O_1721,N_14855,N_14852);
nand UO_1722 (O_1722,N_14949,N_14940);
and UO_1723 (O_1723,N_14785,N_14808);
xnor UO_1724 (O_1724,N_14766,N_14863);
and UO_1725 (O_1725,N_14847,N_14820);
nor UO_1726 (O_1726,N_14775,N_14887);
nor UO_1727 (O_1727,N_14998,N_14872);
nor UO_1728 (O_1728,N_14949,N_14868);
xnor UO_1729 (O_1729,N_14851,N_14996);
xnor UO_1730 (O_1730,N_14929,N_14772);
nor UO_1731 (O_1731,N_14783,N_14916);
nand UO_1732 (O_1732,N_14842,N_14952);
and UO_1733 (O_1733,N_14796,N_14971);
nor UO_1734 (O_1734,N_14975,N_14796);
xor UO_1735 (O_1735,N_14835,N_14895);
nand UO_1736 (O_1736,N_14884,N_14805);
nor UO_1737 (O_1737,N_14970,N_14926);
xnor UO_1738 (O_1738,N_14841,N_14929);
xnor UO_1739 (O_1739,N_14818,N_14770);
nand UO_1740 (O_1740,N_14888,N_14783);
xor UO_1741 (O_1741,N_14851,N_14991);
nand UO_1742 (O_1742,N_14844,N_14883);
nand UO_1743 (O_1743,N_14814,N_14928);
and UO_1744 (O_1744,N_14979,N_14997);
nor UO_1745 (O_1745,N_14921,N_14982);
and UO_1746 (O_1746,N_14787,N_14776);
nand UO_1747 (O_1747,N_14801,N_14906);
nor UO_1748 (O_1748,N_14801,N_14868);
xor UO_1749 (O_1749,N_14906,N_14996);
nand UO_1750 (O_1750,N_14875,N_14765);
nand UO_1751 (O_1751,N_14852,N_14836);
or UO_1752 (O_1752,N_14972,N_14789);
and UO_1753 (O_1753,N_14779,N_14907);
xnor UO_1754 (O_1754,N_14913,N_14773);
nand UO_1755 (O_1755,N_14972,N_14982);
nand UO_1756 (O_1756,N_14770,N_14763);
nor UO_1757 (O_1757,N_14777,N_14833);
or UO_1758 (O_1758,N_14979,N_14841);
nand UO_1759 (O_1759,N_14803,N_14824);
or UO_1760 (O_1760,N_14942,N_14944);
and UO_1761 (O_1761,N_14885,N_14848);
xnor UO_1762 (O_1762,N_14793,N_14891);
nand UO_1763 (O_1763,N_14775,N_14936);
and UO_1764 (O_1764,N_14857,N_14963);
xnor UO_1765 (O_1765,N_14811,N_14796);
nand UO_1766 (O_1766,N_14768,N_14802);
nor UO_1767 (O_1767,N_14813,N_14814);
xor UO_1768 (O_1768,N_14949,N_14983);
and UO_1769 (O_1769,N_14898,N_14953);
and UO_1770 (O_1770,N_14947,N_14789);
nand UO_1771 (O_1771,N_14801,N_14790);
and UO_1772 (O_1772,N_14763,N_14946);
nor UO_1773 (O_1773,N_14969,N_14848);
xnor UO_1774 (O_1774,N_14988,N_14992);
xor UO_1775 (O_1775,N_14761,N_14859);
and UO_1776 (O_1776,N_14834,N_14930);
or UO_1777 (O_1777,N_14818,N_14946);
and UO_1778 (O_1778,N_14782,N_14840);
xor UO_1779 (O_1779,N_14985,N_14826);
and UO_1780 (O_1780,N_14984,N_14922);
or UO_1781 (O_1781,N_14766,N_14983);
xnor UO_1782 (O_1782,N_14814,N_14932);
xor UO_1783 (O_1783,N_14762,N_14764);
or UO_1784 (O_1784,N_14960,N_14756);
xor UO_1785 (O_1785,N_14883,N_14991);
and UO_1786 (O_1786,N_14996,N_14880);
xor UO_1787 (O_1787,N_14891,N_14832);
xnor UO_1788 (O_1788,N_14863,N_14898);
nand UO_1789 (O_1789,N_14922,N_14841);
nand UO_1790 (O_1790,N_14831,N_14854);
or UO_1791 (O_1791,N_14948,N_14916);
nand UO_1792 (O_1792,N_14851,N_14829);
nor UO_1793 (O_1793,N_14781,N_14857);
nor UO_1794 (O_1794,N_14950,N_14952);
nand UO_1795 (O_1795,N_14963,N_14911);
or UO_1796 (O_1796,N_14853,N_14784);
nor UO_1797 (O_1797,N_14901,N_14890);
nand UO_1798 (O_1798,N_14895,N_14814);
nand UO_1799 (O_1799,N_14896,N_14971);
or UO_1800 (O_1800,N_14986,N_14758);
or UO_1801 (O_1801,N_14831,N_14973);
xnor UO_1802 (O_1802,N_14840,N_14892);
and UO_1803 (O_1803,N_14946,N_14801);
nor UO_1804 (O_1804,N_14818,N_14846);
or UO_1805 (O_1805,N_14909,N_14884);
nor UO_1806 (O_1806,N_14990,N_14946);
and UO_1807 (O_1807,N_14946,N_14850);
nor UO_1808 (O_1808,N_14786,N_14998);
xnor UO_1809 (O_1809,N_14967,N_14914);
and UO_1810 (O_1810,N_14896,N_14763);
and UO_1811 (O_1811,N_14897,N_14949);
and UO_1812 (O_1812,N_14776,N_14800);
xnor UO_1813 (O_1813,N_14856,N_14998);
and UO_1814 (O_1814,N_14759,N_14794);
nor UO_1815 (O_1815,N_14833,N_14890);
nand UO_1816 (O_1816,N_14797,N_14933);
xnor UO_1817 (O_1817,N_14796,N_14923);
and UO_1818 (O_1818,N_14950,N_14813);
nand UO_1819 (O_1819,N_14899,N_14808);
xnor UO_1820 (O_1820,N_14944,N_14891);
xor UO_1821 (O_1821,N_14952,N_14931);
and UO_1822 (O_1822,N_14885,N_14892);
nand UO_1823 (O_1823,N_14881,N_14786);
and UO_1824 (O_1824,N_14918,N_14912);
and UO_1825 (O_1825,N_14911,N_14777);
or UO_1826 (O_1826,N_14841,N_14768);
and UO_1827 (O_1827,N_14911,N_14866);
or UO_1828 (O_1828,N_14911,N_14858);
xor UO_1829 (O_1829,N_14876,N_14804);
nor UO_1830 (O_1830,N_14855,N_14795);
and UO_1831 (O_1831,N_14800,N_14780);
and UO_1832 (O_1832,N_14967,N_14957);
xnor UO_1833 (O_1833,N_14778,N_14877);
or UO_1834 (O_1834,N_14791,N_14921);
nand UO_1835 (O_1835,N_14930,N_14855);
nand UO_1836 (O_1836,N_14900,N_14796);
nor UO_1837 (O_1837,N_14916,N_14751);
xnor UO_1838 (O_1838,N_14907,N_14755);
and UO_1839 (O_1839,N_14790,N_14976);
xnor UO_1840 (O_1840,N_14809,N_14904);
nor UO_1841 (O_1841,N_14887,N_14811);
and UO_1842 (O_1842,N_14791,N_14757);
and UO_1843 (O_1843,N_14780,N_14925);
and UO_1844 (O_1844,N_14769,N_14923);
nor UO_1845 (O_1845,N_14856,N_14898);
xor UO_1846 (O_1846,N_14940,N_14814);
and UO_1847 (O_1847,N_14792,N_14890);
nand UO_1848 (O_1848,N_14976,N_14851);
and UO_1849 (O_1849,N_14832,N_14850);
or UO_1850 (O_1850,N_14753,N_14830);
nor UO_1851 (O_1851,N_14750,N_14845);
xnor UO_1852 (O_1852,N_14800,N_14845);
xnor UO_1853 (O_1853,N_14768,N_14801);
or UO_1854 (O_1854,N_14772,N_14802);
nand UO_1855 (O_1855,N_14977,N_14985);
nand UO_1856 (O_1856,N_14805,N_14781);
and UO_1857 (O_1857,N_14779,N_14832);
xnor UO_1858 (O_1858,N_14790,N_14850);
xnor UO_1859 (O_1859,N_14871,N_14992);
nand UO_1860 (O_1860,N_14795,N_14803);
and UO_1861 (O_1861,N_14799,N_14859);
nand UO_1862 (O_1862,N_14807,N_14856);
or UO_1863 (O_1863,N_14858,N_14849);
xnor UO_1864 (O_1864,N_14963,N_14932);
and UO_1865 (O_1865,N_14926,N_14839);
or UO_1866 (O_1866,N_14881,N_14766);
or UO_1867 (O_1867,N_14978,N_14856);
and UO_1868 (O_1868,N_14869,N_14812);
and UO_1869 (O_1869,N_14929,N_14966);
and UO_1870 (O_1870,N_14829,N_14811);
nand UO_1871 (O_1871,N_14995,N_14867);
and UO_1872 (O_1872,N_14886,N_14999);
nand UO_1873 (O_1873,N_14782,N_14770);
xnor UO_1874 (O_1874,N_14819,N_14896);
xor UO_1875 (O_1875,N_14899,N_14965);
nand UO_1876 (O_1876,N_14847,N_14902);
and UO_1877 (O_1877,N_14846,N_14949);
nand UO_1878 (O_1878,N_14816,N_14841);
nor UO_1879 (O_1879,N_14936,N_14904);
nand UO_1880 (O_1880,N_14989,N_14849);
nand UO_1881 (O_1881,N_14765,N_14858);
and UO_1882 (O_1882,N_14915,N_14948);
and UO_1883 (O_1883,N_14812,N_14893);
xnor UO_1884 (O_1884,N_14987,N_14869);
nand UO_1885 (O_1885,N_14901,N_14967);
nor UO_1886 (O_1886,N_14866,N_14890);
nor UO_1887 (O_1887,N_14909,N_14825);
xor UO_1888 (O_1888,N_14791,N_14762);
nor UO_1889 (O_1889,N_14982,N_14936);
and UO_1890 (O_1890,N_14976,N_14867);
or UO_1891 (O_1891,N_14963,N_14845);
nor UO_1892 (O_1892,N_14977,N_14992);
nand UO_1893 (O_1893,N_14808,N_14941);
nand UO_1894 (O_1894,N_14768,N_14957);
nand UO_1895 (O_1895,N_14790,N_14908);
or UO_1896 (O_1896,N_14894,N_14854);
or UO_1897 (O_1897,N_14973,N_14797);
and UO_1898 (O_1898,N_14809,N_14789);
or UO_1899 (O_1899,N_14935,N_14950);
nor UO_1900 (O_1900,N_14793,N_14841);
or UO_1901 (O_1901,N_14942,N_14885);
and UO_1902 (O_1902,N_14901,N_14935);
xor UO_1903 (O_1903,N_14761,N_14807);
nor UO_1904 (O_1904,N_14752,N_14786);
nor UO_1905 (O_1905,N_14897,N_14894);
and UO_1906 (O_1906,N_14863,N_14854);
nor UO_1907 (O_1907,N_14865,N_14818);
or UO_1908 (O_1908,N_14943,N_14824);
nor UO_1909 (O_1909,N_14799,N_14917);
or UO_1910 (O_1910,N_14958,N_14968);
xnor UO_1911 (O_1911,N_14823,N_14902);
and UO_1912 (O_1912,N_14918,N_14867);
nor UO_1913 (O_1913,N_14922,N_14779);
nor UO_1914 (O_1914,N_14860,N_14769);
nor UO_1915 (O_1915,N_14985,N_14927);
xnor UO_1916 (O_1916,N_14799,N_14794);
or UO_1917 (O_1917,N_14933,N_14757);
and UO_1918 (O_1918,N_14819,N_14864);
or UO_1919 (O_1919,N_14968,N_14809);
nand UO_1920 (O_1920,N_14839,N_14958);
xor UO_1921 (O_1921,N_14754,N_14891);
nor UO_1922 (O_1922,N_14874,N_14985);
or UO_1923 (O_1923,N_14837,N_14957);
nand UO_1924 (O_1924,N_14962,N_14796);
nand UO_1925 (O_1925,N_14941,N_14948);
and UO_1926 (O_1926,N_14844,N_14764);
and UO_1927 (O_1927,N_14993,N_14765);
xor UO_1928 (O_1928,N_14862,N_14900);
xnor UO_1929 (O_1929,N_14838,N_14910);
nor UO_1930 (O_1930,N_14799,N_14810);
nand UO_1931 (O_1931,N_14767,N_14863);
xor UO_1932 (O_1932,N_14891,N_14959);
xnor UO_1933 (O_1933,N_14866,N_14939);
and UO_1934 (O_1934,N_14941,N_14753);
or UO_1935 (O_1935,N_14966,N_14968);
or UO_1936 (O_1936,N_14897,N_14941);
and UO_1937 (O_1937,N_14873,N_14810);
nor UO_1938 (O_1938,N_14961,N_14776);
nand UO_1939 (O_1939,N_14839,N_14989);
and UO_1940 (O_1940,N_14942,N_14936);
xor UO_1941 (O_1941,N_14795,N_14876);
and UO_1942 (O_1942,N_14839,N_14936);
and UO_1943 (O_1943,N_14779,N_14962);
and UO_1944 (O_1944,N_14815,N_14860);
xor UO_1945 (O_1945,N_14973,N_14882);
and UO_1946 (O_1946,N_14943,N_14915);
nor UO_1947 (O_1947,N_14968,N_14767);
nand UO_1948 (O_1948,N_14758,N_14812);
or UO_1949 (O_1949,N_14947,N_14839);
nand UO_1950 (O_1950,N_14968,N_14946);
xnor UO_1951 (O_1951,N_14993,N_14894);
nand UO_1952 (O_1952,N_14968,N_14760);
nor UO_1953 (O_1953,N_14954,N_14764);
or UO_1954 (O_1954,N_14966,N_14840);
and UO_1955 (O_1955,N_14759,N_14786);
xor UO_1956 (O_1956,N_14760,N_14929);
nand UO_1957 (O_1957,N_14999,N_14764);
or UO_1958 (O_1958,N_14975,N_14999);
xor UO_1959 (O_1959,N_14921,N_14851);
and UO_1960 (O_1960,N_14923,N_14907);
xnor UO_1961 (O_1961,N_14855,N_14851);
nor UO_1962 (O_1962,N_14960,N_14888);
xor UO_1963 (O_1963,N_14993,N_14929);
nor UO_1964 (O_1964,N_14851,N_14861);
nand UO_1965 (O_1965,N_14884,N_14755);
nand UO_1966 (O_1966,N_14944,N_14906);
or UO_1967 (O_1967,N_14921,N_14965);
or UO_1968 (O_1968,N_14790,N_14812);
xor UO_1969 (O_1969,N_14921,N_14901);
or UO_1970 (O_1970,N_14908,N_14946);
nor UO_1971 (O_1971,N_14807,N_14911);
nand UO_1972 (O_1972,N_14996,N_14955);
or UO_1973 (O_1973,N_14896,N_14753);
nand UO_1974 (O_1974,N_14903,N_14813);
nor UO_1975 (O_1975,N_14997,N_14915);
or UO_1976 (O_1976,N_14988,N_14839);
xor UO_1977 (O_1977,N_14935,N_14776);
and UO_1978 (O_1978,N_14940,N_14904);
xnor UO_1979 (O_1979,N_14770,N_14756);
and UO_1980 (O_1980,N_14856,N_14984);
nand UO_1981 (O_1981,N_14891,N_14933);
or UO_1982 (O_1982,N_14882,N_14807);
nor UO_1983 (O_1983,N_14936,N_14837);
or UO_1984 (O_1984,N_14983,N_14870);
or UO_1985 (O_1985,N_14860,N_14932);
and UO_1986 (O_1986,N_14925,N_14998);
nor UO_1987 (O_1987,N_14765,N_14810);
xor UO_1988 (O_1988,N_14756,N_14834);
and UO_1989 (O_1989,N_14825,N_14853);
nor UO_1990 (O_1990,N_14982,N_14958);
xnor UO_1991 (O_1991,N_14958,N_14981);
and UO_1992 (O_1992,N_14877,N_14944);
nand UO_1993 (O_1993,N_14938,N_14762);
or UO_1994 (O_1994,N_14934,N_14826);
xnor UO_1995 (O_1995,N_14929,N_14814);
xor UO_1996 (O_1996,N_14811,N_14846);
nand UO_1997 (O_1997,N_14777,N_14955);
nand UO_1998 (O_1998,N_14879,N_14796);
nand UO_1999 (O_1999,N_14900,N_14791);
endmodule