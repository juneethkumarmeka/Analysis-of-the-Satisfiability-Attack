module basic_1500_15000_2000_100_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_108,In_18);
and U1 (N_1,In_393,In_1391);
or U2 (N_2,In_1149,In_1006);
and U3 (N_3,In_193,In_4);
nand U4 (N_4,In_36,In_1104);
or U5 (N_5,In_863,In_1403);
xnor U6 (N_6,In_630,In_284);
xor U7 (N_7,In_1323,In_770);
or U8 (N_8,In_1260,In_41);
nand U9 (N_9,In_678,In_49);
xor U10 (N_10,In_268,In_800);
nand U11 (N_11,In_973,In_166);
or U12 (N_12,In_703,In_240);
nand U13 (N_13,In_173,In_62);
or U14 (N_14,In_199,In_402);
or U15 (N_15,In_12,In_263);
and U16 (N_16,In_1175,In_100);
nand U17 (N_17,In_386,In_436);
nor U18 (N_18,In_232,In_326);
xnor U19 (N_19,In_1032,In_1350);
and U20 (N_20,In_242,In_1045);
and U21 (N_21,In_1455,In_471);
or U22 (N_22,In_1127,In_1272);
nor U23 (N_23,In_744,In_843);
xor U24 (N_24,In_374,In_321);
and U25 (N_25,In_717,In_702);
xor U26 (N_26,In_1282,In_559);
and U27 (N_27,In_1141,In_459);
nor U28 (N_28,In_90,In_535);
nor U29 (N_29,In_767,In_1340);
xor U30 (N_30,In_1178,In_1367);
xnor U31 (N_31,In_1203,In_575);
nand U32 (N_32,In_328,In_146);
and U33 (N_33,In_668,In_747);
xnor U34 (N_34,In_430,In_635);
nor U35 (N_35,In_434,In_327);
or U36 (N_36,In_1366,In_296);
xnor U37 (N_37,In_130,In_388);
xor U38 (N_38,In_316,In_71);
or U39 (N_39,In_1486,In_214);
nand U40 (N_40,In_615,In_1316);
nor U41 (N_41,In_174,In_1448);
xnor U42 (N_42,In_1472,In_239);
xor U43 (N_43,In_1173,In_1189);
and U44 (N_44,In_475,In_845);
or U45 (N_45,In_506,In_19);
nor U46 (N_46,In_503,In_1137);
and U47 (N_47,In_330,In_289);
xor U48 (N_48,In_291,In_1090);
and U49 (N_49,In_213,In_589);
or U50 (N_50,In_1204,In_1462);
xnor U51 (N_51,In_496,In_743);
or U52 (N_52,In_68,In_377);
and U53 (N_53,In_354,In_1491);
and U54 (N_54,In_1479,In_387);
and U55 (N_55,In_206,In_1264);
or U56 (N_56,In_711,In_482);
nand U57 (N_57,In_456,In_1093);
nand U58 (N_58,In_105,In_912);
nor U59 (N_59,In_1481,In_990);
nor U60 (N_60,In_1330,In_860);
nand U61 (N_61,In_1099,In_523);
and U62 (N_62,In_865,In_1430);
xor U63 (N_63,In_833,In_1466);
nand U64 (N_64,In_93,In_489);
and U65 (N_65,In_350,In_1125);
nor U66 (N_66,In_1091,In_264);
nor U67 (N_67,In_835,In_1123);
xor U68 (N_68,In_247,In_141);
xor U69 (N_69,In_2,In_1290);
or U70 (N_70,In_1201,In_437);
nor U71 (N_71,In_188,In_723);
nand U72 (N_72,In_182,In_1014);
nor U73 (N_73,In_161,In_1103);
and U74 (N_74,In_1413,In_1028);
nor U75 (N_75,In_510,In_1400);
nand U76 (N_76,In_1305,In_1256);
and U77 (N_77,In_604,In_372);
nor U78 (N_78,In_352,In_447);
and U79 (N_79,In_902,In_844);
or U80 (N_80,In_94,In_1136);
nor U81 (N_81,In_574,In_1012);
nor U82 (N_82,In_917,In_39);
or U83 (N_83,In_1301,In_1478);
nand U84 (N_84,In_820,In_585);
nor U85 (N_85,In_907,In_850);
nor U86 (N_86,In_1306,In_935);
and U87 (N_87,In_204,In_925);
nand U88 (N_88,In_1075,In_207);
nand U89 (N_89,In_1388,In_362);
xnor U90 (N_90,In_281,In_1037);
nand U91 (N_91,In_157,In_1026);
xor U92 (N_92,In_519,In_889);
or U93 (N_93,In_1176,In_1051);
and U94 (N_94,In_1434,In_722);
nor U95 (N_95,In_265,In_558);
xnor U96 (N_96,In_632,In_353);
or U97 (N_97,In_254,In_1474);
or U98 (N_98,In_1346,In_772);
nor U99 (N_99,In_339,In_177);
nand U100 (N_100,In_60,In_1420);
or U101 (N_101,In_701,In_989);
or U102 (N_102,In_883,In_1296);
or U103 (N_103,In_672,In_652);
xnor U104 (N_104,In_915,In_922);
or U105 (N_105,In_298,In_1345);
xnor U106 (N_106,In_1022,In_1036);
and U107 (N_107,In_861,In_1067);
xor U108 (N_108,In_826,In_1143);
or U109 (N_109,In_1440,In_1182);
nand U110 (N_110,In_1092,In_1321);
xnor U111 (N_111,In_187,In_1038);
or U112 (N_112,In_412,In_588);
and U113 (N_113,In_1184,In_584);
or U114 (N_114,In_195,In_155);
or U115 (N_115,In_964,In_137);
and U116 (N_116,In_745,In_86);
and U117 (N_117,In_1179,In_244);
nor U118 (N_118,In_966,In_501);
and U119 (N_119,In_34,In_746);
nand U120 (N_120,In_101,In_1213);
nor U121 (N_121,In_949,In_1432);
nor U122 (N_122,In_295,In_1168);
and U123 (N_123,In_662,In_719);
and U124 (N_124,In_1490,In_453);
nand U125 (N_125,In_78,In_158);
nand U126 (N_126,In_822,In_555);
nand U127 (N_127,In_901,In_572);
nor U128 (N_128,In_655,In_764);
nor U129 (N_129,In_971,In_293);
and U130 (N_130,In_1236,In_646);
and U131 (N_131,In_56,In_151);
and U132 (N_132,In_1473,In_356);
or U133 (N_133,In_1154,In_1102);
xor U134 (N_134,In_563,In_1110);
and U135 (N_135,In_470,In_910);
nand U136 (N_136,In_836,In_58);
nand U137 (N_137,In_346,In_761);
or U138 (N_138,In_677,In_618);
or U139 (N_139,In_325,In_680);
nand U140 (N_140,In_391,In_1202);
nor U141 (N_141,In_540,In_1132);
nor U142 (N_142,In_1342,In_817);
nor U143 (N_143,In_537,In_382);
and U144 (N_144,In_1331,In_120);
and U145 (N_145,In_939,In_418);
nor U146 (N_146,In_53,In_385);
and U147 (N_147,In_444,In_806);
xnor U148 (N_148,In_895,In_867);
nand U149 (N_149,In_492,In_787);
xnor U150 (N_150,In_1198,In_938);
xor U151 (N_151,In_1445,N_101);
or U152 (N_152,In_116,In_241);
nand U153 (N_153,In_408,In_682);
nand U154 (N_154,In_288,In_621);
or U155 (N_155,In_319,In_696);
and U156 (N_156,In_786,In_890);
nand U157 (N_157,In_469,In_999);
xnor U158 (N_158,In_439,In_721);
nand U159 (N_159,In_927,In_600);
nand U160 (N_160,N_123,In_1057);
nor U161 (N_161,In_1109,N_84);
nor U162 (N_162,In_169,In_376);
xnor U163 (N_163,In_892,In_28);
xnor U164 (N_164,In_790,In_1197);
xnor U165 (N_165,In_1389,In_1218);
or U166 (N_166,In_428,In_760);
or U167 (N_167,In_64,In_1114);
xnor U168 (N_168,In_340,In_733);
xnor U169 (N_169,In_258,N_113);
nor U170 (N_170,N_70,In_70);
xor U171 (N_171,In_950,In_1356);
nand U172 (N_172,In_753,In_961);
xor U173 (N_173,In_716,In_1021);
nand U174 (N_174,In_499,In_1436);
nor U175 (N_175,In_1053,In_566);
xor U176 (N_176,N_61,In_1464);
nor U177 (N_177,In_958,In_335);
or U178 (N_178,N_37,In_410);
nand U179 (N_179,N_114,In_1191);
and U180 (N_180,In_171,In_421);
nor U181 (N_181,In_490,In_583);
and U182 (N_182,In_923,In_875);
or U183 (N_183,In_72,In_567);
nand U184 (N_184,N_99,In_879);
or U185 (N_185,In_888,In_323);
nor U186 (N_186,In_838,In_612);
nand U187 (N_187,In_1263,In_368);
or U188 (N_188,N_33,In_1159);
or U189 (N_189,N_82,In_1039);
nor U190 (N_190,In_67,In_1031);
nand U191 (N_191,In_311,In_1374);
nand U192 (N_192,In_507,In_33);
nand U193 (N_193,In_1292,In_688);
and U194 (N_194,In_96,In_107);
or U195 (N_195,In_314,In_128);
and U196 (N_196,In_683,In_1378);
or U197 (N_197,In_1415,In_1054);
and U198 (N_198,In_1461,N_135);
and U199 (N_199,In_1344,In_1207);
or U200 (N_200,N_18,In_653);
nor U201 (N_201,In_739,In_262);
nand U202 (N_202,In_715,In_1327);
xor U203 (N_203,In_1369,N_65);
xnor U204 (N_204,In_952,In_934);
nor U205 (N_205,In_134,In_1365);
xor U206 (N_206,In_1371,In_570);
xnor U207 (N_207,N_133,In_1497);
or U208 (N_208,In_32,In_1223);
nand U209 (N_209,In_564,N_108);
nand U210 (N_210,In_1253,In_243);
or U211 (N_211,In_1337,In_216);
xnor U212 (N_212,In_361,In_527);
nor U213 (N_213,In_1181,In_9);
and U214 (N_214,N_14,In_568);
nand U215 (N_215,In_266,In_705);
nand U216 (N_216,In_579,In_183);
nor U217 (N_217,In_980,In_616);
nor U218 (N_218,In_1397,In_797);
or U219 (N_219,In_360,In_426);
or U220 (N_220,In_409,In_1465);
nand U221 (N_221,In_1111,In_752);
and U222 (N_222,In_468,In_776);
xnor U223 (N_223,In_606,N_80);
xor U224 (N_224,In_549,In_82);
nor U225 (N_225,In_1112,N_69);
xnor U226 (N_226,In_846,In_1442);
nor U227 (N_227,In_365,In_275);
or U228 (N_228,In_1452,In_348);
nor U229 (N_229,In_903,N_68);
and U230 (N_230,In_1108,In_127);
xor U231 (N_231,In_455,In_1435);
nand U232 (N_232,In_164,N_98);
nand U233 (N_233,In_248,In_525);
or U234 (N_234,N_125,In_272);
nand U235 (N_235,In_399,In_1082);
nor U236 (N_236,In_1254,In_1412);
or U237 (N_237,In_176,In_200);
and U238 (N_238,In_231,In_40);
nor U239 (N_239,In_286,In_740);
nand U240 (N_240,In_1240,In_109);
nand U241 (N_241,In_1360,In_598);
xnor U242 (N_242,In_1250,In_1244);
nand U243 (N_243,In_123,In_947);
xnor U244 (N_244,In_31,In_756);
nand U245 (N_245,In_650,In_643);
nand U246 (N_246,In_942,In_909);
nand U247 (N_247,In_819,In_550);
xnor U248 (N_248,In_156,N_110);
nand U249 (N_249,In_1252,In_417);
or U250 (N_250,In_1237,In_1120);
and U251 (N_251,In_1382,In_792);
xnor U252 (N_252,In_1208,In_748);
or U253 (N_253,In_1152,N_74);
or U254 (N_254,In_255,In_789);
nand U255 (N_255,In_1105,In_429);
and U256 (N_256,In_74,N_109);
nor U257 (N_257,In_1401,In_1251);
or U258 (N_258,In_1482,In_61);
nor U259 (N_259,In_698,In_225);
or U260 (N_260,In_1018,In_1193);
or U261 (N_261,N_36,In_957);
xnor U262 (N_262,N_0,N_11);
xor U263 (N_263,In_1089,In_103);
nor U264 (N_264,In_461,In_675);
nand U265 (N_265,In_1439,N_50);
and U266 (N_266,In_1106,In_636);
or U267 (N_267,N_54,In_1171);
and U268 (N_268,In_331,N_87);
or U269 (N_269,In_687,In_29);
or U270 (N_270,In_147,In_1122);
nor U271 (N_271,In_900,In_593);
nor U272 (N_272,In_1096,In_638);
and U273 (N_273,In_344,In_818);
xor U274 (N_274,N_20,In_42);
nor U275 (N_275,N_105,In_341);
nand U276 (N_276,In_1144,In_642);
or U277 (N_277,In_1329,In_738);
or U278 (N_278,In_106,In_1271);
or U279 (N_279,In_245,In_977);
nor U280 (N_280,In_114,In_1424);
or U281 (N_281,N_141,In_706);
and U282 (N_282,In_1278,In_420);
nor U283 (N_283,In_1395,N_126);
nor U284 (N_284,In_956,In_1081);
or U285 (N_285,In_1229,In_1315);
nand U286 (N_286,In_1079,In_926);
nand U287 (N_287,In_918,In_1158);
and U288 (N_288,In_1310,In_1161);
or U289 (N_289,In_1381,In_153);
and U290 (N_290,In_1243,In_500);
or U291 (N_291,In_1196,In_608);
xnor U292 (N_292,In_394,In_477);
nand U293 (N_293,In_369,In_186);
or U294 (N_294,In_1476,In_948);
nand U295 (N_295,N_95,In_138);
nand U296 (N_296,In_508,In_1140);
xor U297 (N_297,In_75,In_857);
and U298 (N_298,In_1273,In_1027);
nor U299 (N_299,In_92,N_134);
xor U300 (N_300,In_951,In_343);
nor U301 (N_301,N_144,In_357);
nor U302 (N_302,In_491,N_232);
xnor U303 (N_303,In_85,N_272);
or U304 (N_304,N_287,In_887);
xnor U305 (N_305,In_389,In_778);
or U306 (N_306,In_367,In_985);
nor U307 (N_307,In_140,In_1024);
xnor U308 (N_308,N_143,In_5);
xor U309 (N_309,In_839,In_665);
and U310 (N_310,In_1133,In_1078);
nand U311 (N_311,In_801,In_342);
or U312 (N_312,In_390,In_661);
and U313 (N_313,In_1239,In_1084);
xnor U314 (N_314,In_152,In_1370);
nor U315 (N_315,In_472,In_407);
or U316 (N_316,N_154,N_67);
nand U317 (N_317,In_269,In_1107);
nand U318 (N_318,In_828,In_253);
nor U319 (N_319,In_1097,In_1390);
and U320 (N_320,In_984,In_1469);
and U321 (N_321,In_230,In_1499);
nand U322 (N_322,N_234,N_103);
or U323 (N_323,In_1048,N_56);
and U324 (N_324,In_222,N_63);
xnor U325 (N_325,In_279,N_10);
nor U326 (N_326,In_1146,N_111);
nand U327 (N_327,N_5,N_224);
and U328 (N_328,In_1285,In_1309);
xnor U329 (N_329,In_679,In_415);
xor U330 (N_330,N_2,In_118);
xor U331 (N_331,In_513,N_83);
nand U332 (N_332,In_592,In_1319);
or U333 (N_333,In_227,N_137);
or U334 (N_334,In_1281,In_609);
and U335 (N_335,In_1157,In_1080);
or U336 (N_336,N_210,In_1328);
nand U337 (N_337,In_929,In_751);
nand U338 (N_338,In_37,N_241);
xnor U339 (N_339,In_924,N_278);
xnor U340 (N_340,In_87,In_1494);
nor U341 (N_341,In_1368,N_157);
nand U342 (N_342,In_611,In_941);
nor U343 (N_343,In_553,In_280);
nand U344 (N_344,In_788,N_259);
xor U345 (N_345,In_6,In_1066);
and U346 (N_346,In_1165,In_656);
nand U347 (N_347,In_1072,In_26);
and U348 (N_348,In_277,In_476);
and U349 (N_349,In_710,N_77);
nand U350 (N_350,In_795,N_79);
xnor U351 (N_351,In_414,In_1206);
nand U352 (N_352,In_1386,In_59);
or U353 (N_353,N_299,N_91);
and U354 (N_354,In_866,In_781);
nand U355 (N_355,In_400,In_1020);
xnor U356 (N_356,In_965,In_1227);
nand U357 (N_357,In_1405,In_763);
nor U358 (N_358,In_310,N_88);
nand U359 (N_359,N_21,In_66);
xnor U360 (N_360,In_853,In_1270);
xnor U361 (N_361,In_460,In_271);
nand U362 (N_362,In_16,In_1302);
nor U363 (N_363,In_992,In_465);
and U364 (N_364,N_274,In_1393);
and U365 (N_365,In_596,In_700);
and U366 (N_366,In_932,In_1005);
xnor U367 (N_367,In_986,N_51);
nand U368 (N_368,In_1069,In_1186);
nand U369 (N_369,In_397,In_228);
nand U370 (N_370,N_41,In_1164);
xnor U371 (N_371,In_505,N_60);
and U372 (N_372,N_185,In_560);
xor U373 (N_373,In_921,In_35);
nand U374 (N_374,In_97,In_270);
nand U375 (N_375,N_212,In_79);
nor U376 (N_376,In_842,In_991);
or U377 (N_377,In_395,N_8);
xnor U378 (N_378,In_11,In_1467);
nand U379 (N_379,In_1194,In_483);
nand U380 (N_380,In_725,In_1334);
nor U381 (N_381,In_457,N_151);
and U382 (N_382,In_1129,N_44);
nand U383 (N_383,In_1100,In_919);
and U384 (N_384,In_520,In_1190);
and U385 (N_385,In_1284,In_1447);
nor U386 (N_386,N_213,In_1353);
nand U387 (N_387,In_774,In_1289);
or U388 (N_388,In_749,N_120);
nor U389 (N_389,In_994,In_1364);
nand U390 (N_390,In_690,In_132);
or U391 (N_391,In_282,In_1457);
and U392 (N_392,In_1279,In_1362);
nand U393 (N_393,In_1118,In_1459);
xnor U394 (N_394,In_773,N_257);
and U395 (N_395,In_547,In_813);
xnor U396 (N_396,N_22,In_22);
xor U397 (N_397,In_815,In_46);
xnor U398 (N_398,In_165,In_1333);
and U399 (N_399,In_734,In_684);
xor U400 (N_400,N_225,In_113);
or U401 (N_401,In_1493,In_518);
nand U402 (N_402,In_1219,In_1180);
xnor U403 (N_403,In_1347,In_855);
xnor U404 (N_404,In_851,In_234);
nand U405 (N_405,N_184,In_996);
or U406 (N_406,In_336,N_81);
nor U407 (N_407,In_237,N_169);
nand U408 (N_408,In_1052,In_1433);
xnor U409 (N_409,In_260,In_304);
nand U410 (N_410,N_24,In_1291);
nand U411 (N_411,In_180,In_849);
nor U412 (N_412,In_1117,In_904);
and U413 (N_413,In_333,In_48);
or U414 (N_414,In_283,In_112);
and U415 (N_415,In_17,N_260);
xnor U416 (N_416,N_261,In_1349);
or U417 (N_417,In_381,In_590);
and U418 (N_418,In_7,In_673);
or U419 (N_419,In_65,In_181);
xor U420 (N_420,In_494,In_27);
nand U421 (N_421,In_308,In_15);
nor U422 (N_422,In_1308,In_1148);
nor U423 (N_423,In_561,In_1343);
nand U424 (N_424,In_1384,In_1062);
or U425 (N_425,In_1394,In_91);
or U426 (N_426,In_1453,In_1267);
and U427 (N_427,In_897,N_34);
nand U428 (N_428,In_1485,In_287);
or U429 (N_429,N_127,N_40);
and U430 (N_430,In_478,In_1409);
and U431 (N_431,In_775,N_186);
xnor U432 (N_432,In_1417,In_63);
nand U433 (N_433,In_824,In_98);
or U434 (N_434,In_1408,N_228);
xor U435 (N_435,In_1242,In_198);
nand U436 (N_436,In_51,In_102);
nor U437 (N_437,In_1139,In_435);
or U438 (N_438,N_17,N_211);
xnor U439 (N_439,In_969,In_623);
xnor U440 (N_440,In_614,In_913);
nand U441 (N_441,N_238,In_1088);
nand U442 (N_442,N_90,In_783);
xor U443 (N_443,In_963,In_1317);
nor U444 (N_444,In_210,In_1399);
nor U445 (N_445,In_1142,In_730);
nand U446 (N_446,In_306,In_663);
or U447 (N_447,In_1225,In_396);
or U448 (N_448,In_576,In_1003);
nand U449 (N_449,In_619,In_1443);
xnor U450 (N_450,N_258,N_214);
and U451 (N_451,In_955,In_968);
and U452 (N_452,In_697,In_552);
nand U453 (N_453,In_975,In_1046);
xnor U454 (N_454,In_516,In_562);
or U455 (N_455,N_436,N_30);
nor U456 (N_456,In_398,In_647);
and U457 (N_457,In_1313,N_128);
nand U458 (N_458,In_868,In_1115);
and U459 (N_459,N_226,N_97);
xor U460 (N_460,In_1380,N_422);
nand U461 (N_461,In_256,In_724);
nand U462 (N_462,In_755,N_136);
nor U463 (N_463,N_75,N_118);
nand U464 (N_464,In_631,In_908);
or U465 (N_465,N_330,N_271);
nand U466 (N_466,N_310,N_156);
and U467 (N_467,N_198,N_178);
or U468 (N_468,In_45,In_754);
xor U469 (N_469,In_1422,In_823);
nand U470 (N_470,In_168,N_161);
and U471 (N_471,N_367,In_1150);
xnor U472 (N_472,In_273,In_834);
nand U473 (N_473,In_274,In_1247);
nor U474 (N_474,In_595,In_840);
and U475 (N_475,In_1454,N_243);
or U476 (N_476,N_404,N_316);
nand U477 (N_477,In_610,In_1217);
xnor U478 (N_478,In_1221,In_766);
nand U479 (N_479,N_216,In_832);
xor U480 (N_480,In_150,N_48);
nand U481 (N_481,In_143,In_873);
xnor U482 (N_482,In_148,In_758);
nand U483 (N_483,In_315,In_580);
and U484 (N_484,In_983,In_704);
nor U485 (N_485,In_937,N_155);
or U486 (N_486,In_674,In_1354);
and U487 (N_487,In_856,In_886);
nor U488 (N_488,In_714,In_285);
and U489 (N_489,In_312,In_1451);
nand U490 (N_490,In_1456,In_1475);
nand U491 (N_491,In_424,In_829);
and U492 (N_492,In_626,In_1121);
or U493 (N_493,In_959,In_962);
xor U494 (N_494,In_205,N_195);
nand U495 (N_495,N_78,N_240);
nand U496 (N_496,N_396,N_313);
and U497 (N_497,In_451,In_1318);
nor U498 (N_498,N_376,In_104);
nand U499 (N_499,In_486,In_617);
xor U500 (N_500,N_388,In_495);
and U501 (N_501,In_1410,N_117);
nor U502 (N_502,N_239,In_1268);
nor U503 (N_503,In_149,In_586);
nor U504 (N_504,N_369,In_1352);
nor U505 (N_505,N_409,N_339);
xor U506 (N_506,In_765,In_1293);
xnor U507 (N_507,In_1177,N_405);
and U508 (N_508,In_737,In_1322);
nand U509 (N_509,In_422,In_463);
or U510 (N_510,In_1257,In_1460);
or U511 (N_511,In_1232,N_307);
and U512 (N_512,In_742,N_431);
xnor U513 (N_513,In_14,In_115);
xor U514 (N_514,N_275,In_1372);
nor U515 (N_515,In_124,In_1283);
and U516 (N_516,N_315,In_1163);
and U517 (N_517,In_648,In_1147);
nand U518 (N_518,In_1063,N_85);
xnor U519 (N_519,In_154,In_1245);
xnor U520 (N_520,In_144,In_811);
or U521 (N_521,In_762,In_178);
nor U522 (N_522,N_252,N_28);
nor U523 (N_523,In_1009,In_1423);
and U524 (N_524,In_139,In_179);
or U525 (N_525,In_1138,N_235);
or U526 (N_526,N_132,N_361);
nand U527 (N_527,N_229,In_882);
xnor U528 (N_528,In_1419,In_629);
xor U529 (N_529,N_406,In_324);
xnor U530 (N_530,In_305,In_194);
and U531 (N_531,N_177,N_222);
or U532 (N_532,In_1280,In_443);
xnor U533 (N_533,In_874,In_1);
and U534 (N_534,In_809,In_261);
nor U535 (N_535,N_251,In_557);
or U536 (N_536,In_645,N_153);
nor U537 (N_537,N_130,In_1269);
or U538 (N_538,In_364,In_329);
nand U539 (N_539,N_182,In_89);
xor U540 (N_540,In_1017,In_976);
and U541 (N_541,N_276,In_603);
xnor U542 (N_542,N_39,In_911);
nand U543 (N_543,N_264,In_1043);
and U544 (N_544,In_332,In_175);
and U545 (N_545,In_514,In_110);
and U546 (N_546,In_884,In_1070);
nand U547 (N_547,In_594,In_1297);
and U548 (N_548,N_236,In_1261);
or U549 (N_549,In_1004,N_398);
nand U550 (N_550,In_1226,In_235);
nand U551 (N_551,In_1162,In_664);
xnor U552 (N_552,In_821,In_693);
xor U553 (N_553,N_352,In_779);
or U554 (N_554,In_474,In_57);
nand U555 (N_555,N_140,In_551);
xnor U556 (N_556,In_1116,In_202);
nand U557 (N_557,In_1307,N_223);
xor U558 (N_558,In_55,In_1392);
or U559 (N_559,In_1348,In_1426);
and U560 (N_560,In_1056,In_1418);
nand U561 (N_561,N_331,In_449);
and U562 (N_562,N_104,In_933);
xor U563 (N_563,N_385,In_1230);
and U564 (N_564,N_73,In_1463);
nand U565 (N_565,In_1200,In_218);
nor U566 (N_566,N_233,In_1113);
and U567 (N_567,In_681,In_542);
xnor U568 (N_568,In_10,N_372);
xnor U569 (N_569,N_415,In_1013);
and U570 (N_570,N_300,In_1166);
nor U571 (N_571,N_148,N_200);
xor U572 (N_572,In_1276,N_303);
nand U573 (N_573,In_208,In_521);
xor U574 (N_574,In_658,N_138);
and U575 (N_575,N_344,In_1458);
nor U576 (N_576,In_1029,In_223);
nor U577 (N_577,In_1019,In_1216);
nor U578 (N_578,In_442,N_298);
and U579 (N_579,In_299,In_257);
xnor U580 (N_580,N_269,In_1047);
xnor U581 (N_581,In_1205,In_0);
nand U582 (N_582,In_1259,N_384);
xnor U583 (N_583,N_89,In_498);
or U584 (N_584,In_432,In_1135);
and U585 (N_585,N_250,In_1130);
and U586 (N_586,In_1059,In_509);
or U587 (N_587,In_111,In_318);
nor U588 (N_588,In_914,In_359);
nor U589 (N_589,In_526,N_242);
xnor U590 (N_590,N_449,In_802);
nor U591 (N_591,In_1085,In_458);
nor U592 (N_592,N_428,In_201);
nor U593 (N_593,In_1498,In_219);
nor U594 (N_594,N_382,N_267);
nand U595 (N_595,In_872,In_718);
nor U596 (N_596,N_435,In_38);
or U597 (N_597,N_438,In_267);
nand U598 (N_598,In_1355,N_266);
or U599 (N_599,N_4,N_311);
nor U600 (N_600,N_489,N_463);
nand U601 (N_601,N_338,In_1396);
nand U602 (N_602,In_995,In_862);
xor U603 (N_603,N_552,N_230);
or U604 (N_604,N_529,N_35);
and U605 (N_605,In_1304,In_20);
or U606 (N_606,N_343,In_898);
nor U607 (N_607,In_726,In_294);
nor U608 (N_608,In_1324,In_338);
or U609 (N_609,N_183,N_254);
nor U610 (N_610,In_881,N_395);
xor U611 (N_611,N_49,In_1437);
xnor U612 (N_612,N_393,N_12);
xor U613 (N_613,N_255,In_1294);
nand U614 (N_614,N_473,In_1170);
and U615 (N_615,N_6,N_197);
nor U616 (N_616,N_55,N_172);
nand U617 (N_617,In_1049,In_309);
nand U618 (N_618,N_444,N_558);
xor U619 (N_619,N_187,In_1220);
or U620 (N_620,In_569,In_480);
and U621 (N_621,In_1375,N_470);
and U622 (N_622,In_1224,N_53);
nand U623 (N_623,N_64,N_568);
nand U624 (N_624,In_259,In_358);
nand U625 (N_625,N_554,In_1083);
and U626 (N_626,In_854,N_306);
nand U627 (N_627,In_847,N_547);
and U628 (N_628,In_73,In_1449);
nand U629 (N_629,N_349,N_327);
nor U630 (N_630,N_440,In_142);
xor U631 (N_631,In_226,N_9);
nor U632 (N_632,In_1298,N_326);
and U633 (N_633,In_1341,N_534);
nand U634 (N_634,In_211,In_167);
or U635 (N_635,In_1030,N_500);
or U636 (N_636,N_32,In_906);
nor U637 (N_637,N_478,In_713);
nand U638 (N_638,In_639,In_184);
nor U639 (N_639,In_1266,In_896);
xor U640 (N_640,In_1233,N_439);
or U641 (N_641,N_504,In_159);
or U642 (N_642,In_649,In_366);
xnor U643 (N_643,In_1055,N_196);
xor U644 (N_644,N_121,In_1094);
nor U645 (N_645,N_468,In_633);
and U646 (N_646,N_180,In_1438);
nor U647 (N_647,In_21,In_709);
and U648 (N_648,N_383,In_1071);
nand U649 (N_649,In_121,In_1040);
and U650 (N_650,N_479,In_1489);
xor U651 (N_651,In_782,N_163);
xnor U652 (N_652,In_539,In_864);
and U653 (N_653,In_481,N_485);
xor U654 (N_654,In_858,In_548);
nor U655 (N_655,N_588,N_417);
xnor U656 (N_656,N_496,In_423);
or U657 (N_657,In_708,N_205);
or U658 (N_658,N_540,In_597);
nor U659 (N_659,In_1383,N_513);
and U660 (N_660,N_451,In_667);
and U661 (N_661,N_375,In_431);
or U662 (N_662,N_555,In_1320);
or U663 (N_663,N_447,N_204);
nor U664 (N_664,In_689,N_284);
xor U665 (N_665,In_290,In_848);
or U666 (N_666,N_47,In_784);
or U667 (N_667,N_107,In_1361);
and U668 (N_668,N_493,N_392);
xnor U669 (N_669,N_556,N_515);
xnor U670 (N_670,In_1425,In_1287);
and U671 (N_671,N_481,N_290);
xor U672 (N_672,In_307,In_810);
and U673 (N_673,In_692,In_1077);
or U674 (N_674,N_166,N_486);
xor U675 (N_675,In_533,N_57);
xor U676 (N_676,N_593,In_351);
nor U677 (N_677,In_1358,In_467);
nor U678 (N_678,N_551,In_654);
and U679 (N_679,N_206,In_1185);
and U680 (N_680,N_594,In_1235);
or U681 (N_681,N_592,In_172);
nand U682 (N_682,N_159,N_215);
xor U683 (N_683,In_757,N_333);
xor U684 (N_684,In_808,In_448);
and U685 (N_685,In_416,N_270);
or U686 (N_686,N_371,N_368);
nor U687 (N_687,N_58,In_735);
nor U688 (N_688,N_301,In_345);
and U689 (N_689,In_8,N_319);
or U690 (N_690,In_163,N_576);
xor U691 (N_691,In_1058,In_972);
nand U692 (N_692,N_469,In_1275);
xnor U693 (N_693,In_946,In_54);
or U694 (N_694,In_349,In_591);
nor U695 (N_695,In_403,N_459);
xnor U696 (N_696,In_885,In_920);
and U697 (N_697,N_221,In_1007);
xor U698 (N_698,In_727,N_190);
nor U699 (N_699,In_798,N_541);
or U700 (N_700,In_1025,N_418);
nand U701 (N_701,N_505,N_199);
and U702 (N_702,In_185,N_354);
nand U703 (N_703,In_1199,In_799);
or U704 (N_704,N_346,In_1487);
nor U705 (N_705,N_129,In_515);
nand U706 (N_706,N_509,In_1215);
nand U707 (N_707,In_1188,In_1145);
xnor U708 (N_708,In_869,In_841);
nor U709 (N_709,In_76,N_571);
or U710 (N_710,N_93,In_466);
or U711 (N_711,In_493,N_389);
nor U712 (N_712,In_300,In_373);
xor U713 (N_713,In_404,N_227);
xor U714 (N_714,In_1325,N_573);
and U715 (N_715,N_297,N_66);
or U716 (N_716,N_176,N_191);
xnor U717 (N_717,N_546,N_420);
and U718 (N_718,In_129,In_728);
nor U719 (N_719,In_1044,N_173);
and U720 (N_720,In_276,N_345);
and U721 (N_721,In_512,N_45);
xor U722 (N_722,N_579,In_1000);
nor U723 (N_723,N_525,In_571);
nor U724 (N_724,In_967,N_441);
and U725 (N_725,N_362,N_302);
nor U726 (N_726,In_3,N_209);
and U727 (N_727,N_374,In_250);
and U728 (N_728,N_160,N_181);
or U729 (N_729,In_1061,In_313);
nand U730 (N_730,In_1450,N_483);
xor U731 (N_731,In_522,In_974);
nand U732 (N_732,N_570,N_502);
and U733 (N_733,In_624,In_1131);
nand U734 (N_734,In_462,N_150);
xor U735 (N_735,N_399,In_625);
nand U736 (N_736,N_429,In_587);
nand U737 (N_737,In_543,In_1153);
xor U738 (N_738,N_201,In_536);
nand U739 (N_739,N_208,In_190);
xnor U740 (N_740,In_383,In_406);
and U741 (N_741,N_194,In_859);
and U742 (N_742,N_562,In_1295);
xor U743 (N_743,In_1488,N_419);
xnor U744 (N_744,N_432,In_928);
nor U745 (N_745,N_475,In_601);
xnor U746 (N_746,N_179,In_1480);
or U747 (N_747,In_1495,In_43);
nor U748 (N_748,N_380,N_407);
nor U749 (N_749,In_233,In_1484);
and U750 (N_750,N_461,N_640);
or U751 (N_751,N_739,In_905);
nor U752 (N_752,N_585,In_1387);
xnor U753 (N_753,N_437,N_320);
nor U754 (N_754,N_580,In_796);
nor U755 (N_755,In_803,N_743);
and U756 (N_756,In_712,In_464);
nor U757 (N_757,In_292,N_714);
and U758 (N_758,In_1335,N_46);
xor U759 (N_759,In_1444,In_1496);
nand U760 (N_760,N_709,N_59);
or U761 (N_761,N_564,In_825);
or U762 (N_762,In_651,N_336);
nor U763 (N_763,In_1041,In_916);
nand U764 (N_764,N_604,In_669);
and U765 (N_765,N_321,N_426);
and U766 (N_766,In_880,N_644);
nor U767 (N_767,N_411,N_445);
xor U768 (N_768,In_1470,N_676);
xor U769 (N_769,In_998,In_1068);
and U770 (N_770,In_930,N_619);
and U771 (N_771,In_1314,N_503);
nand U772 (N_772,In_807,In_487);
xor U773 (N_773,N_693,N_387);
xnor U774 (N_774,N_657,In_221);
nand U775 (N_775,N_625,N_582);
nand U776 (N_776,N_390,In_1477);
nand U777 (N_777,In_657,In_189);
xnor U778 (N_778,N_702,N_561);
and U779 (N_779,N_377,N_304);
and U780 (N_780,N_328,In_1169);
nor U781 (N_781,N_660,N_427);
nor U782 (N_782,N_581,In_1008);
or U783 (N_783,N_749,In_162);
nor U784 (N_784,N_188,In_220);
nor U785 (N_785,N_711,In_769);
xnor U786 (N_786,In_1156,In_249);
or U787 (N_787,In_433,N_62);
xnor U788 (N_788,N_102,N_730);
nand U789 (N_789,In_538,N_724);
nor U790 (N_790,In_1172,N_495);
nand U791 (N_791,In_77,N_710);
or U792 (N_792,N_231,N_379);
nand U793 (N_793,N_434,In_982);
or U794 (N_794,N_543,N_597);
and U795 (N_795,In_852,In_1023);
nand U796 (N_796,In_1286,In_686);
nor U797 (N_797,N_174,N_612);
or U798 (N_798,In_1002,In_830);
nand U799 (N_799,In_347,N_747);
nor U800 (N_800,In_135,N_146);
and U801 (N_801,In_1402,N_507);
nor U802 (N_802,N_165,N_624);
and U803 (N_803,N_457,N_536);
xor U804 (N_804,N_560,In_528);
nand U805 (N_805,In_122,N_262);
nor U806 (N_806,In_891,In_1134);
and U807 (N_807,N_296,N_247);
or U808 (N_808,In_1228,N_618);
nand U809 (N_809,In_1187,N_590);
or U810 (N_810,N_279,In_827);
and U811 (N_811,In_750,In_970);
or U812 (N_812,In_1241,In_452);
xnor U813 (N_813,N_591,N_678);
and U814 (N_814,N_292,In_640);
or U815 (N_815,In_1332,In_80);
nand U816 (N_816,N_355,N_425);
xnor U817 (N_817,N_707,In_454);
nand U818 (N_818,In_979,In_805);
nand U819 (N_819,N_701,N_689);
or U820 (N_820,N_413,N_498);
or U821 (N_821,N_263,In_804);
nor U822 (N_822,In_731,N_549);
xor U823 (N_823,N_589,In_497);
nor U824 (N_824,In_613,N_453);
or U825 (N_825,In_602,N_96);
nor U826 (N_826,In_160,N_677);
nor U827 (N_827,In_1064,N_23);
nor U828 (N_828,N_484,N_480);
and U829 (N_829,N_715,In_1411);
or U830 (N_830,N_577,N_706);
nor U831 (N_831,In_337,In_940);
and U832 (N_832,In_953,In_741);
or U833 (N_833,N_340,In_1124);
nand U834 (N_834,N_13,N_654);
nor U835 (N_835,In_1404,N_43);
nor U836 (N_836,In_1336,N_687);
or U837 (N_837,In_1431,In_694);
nor U838 (N_838,In_488,N_537);
or U839 (N_839,N_351,N_520);
nand U840 (N_840,N_682,In_1311);
nand U841 (N_841,In_945,N_595);
nor U842 (N_842,N_673,In_899);
and U843 (N_843,N_639,In_729);
and U844 (N_844,N_220,N_293);
or U845 (N_845,N_716,In_581);
xor U846 (N_846,In_1167,In_126);
or U847 (N_847,In_99,N_635);
xnor U848 (N_848,N_309,In_1446);
nand U849 (N_849,N_416,N_521);
xnor U850 (N_850,In_1128,N_465);
xor U851 (N_851,In_720,In_427);
xnor U852 (N_852,In_1160,In_1211);
and U853 (N_853,In_215,N_658);
or U854 (N_854,In_573,N_544);
and U855 (N_855,N_466,N_288);
xnor U856 (N_856,N_16,In_425);
xnor U857 (N_857,In_303,N_601);
xor U858 (N_858,N_289,In_392);
nor U859 (N_859,N_516,N_674);
nor U860 (N_860,In_1016,In_517);
nand U861 (N_861,N_717,In_47);
xor U862 (N_862,In_1231,In_1119);
xnor U863 (N_863,N_578,In_380);
nand U864 (N_864,In_212,N_421);
xnor U865 (N_865,In_837,N_189);
nand U866 (N_866,N_285,N_586);
xor U867 (N_867,N_566,N_718);
or U868 (N_868,In_831,In_1209);
nand U869 (N_869,N_528,N_628);
and U870 (N_870,In_1312,N_219);
or U871 (N_871,N_685,N_72);
nand U872 (N_872,N_647,N_688);
or U873 (N_873,N_116,N_740);
nand U874 (N_874,N_695,In_246);
nor U875 (N_875,N_203,N_280);
or U876 (N_876,In_622,N_248);
and U877 (N_877,In_95,In_768);
or U878 (N_878,N_508,In_1299);
and U879 (N_879,N_735,In_785);
xor U880 (N_880,In_217,In_666);
or U881 (N_881,In_1428,In_943);
xor U882 (N_882,N_450,N_665);
xnor U883 (N_883,In_544,N_670);
and U884 (N_884,N_337,N_605);
or U885 (N_885,In_556,N_611);
nor U886 (N_886,N_268,N_666);
nand U887 (N_887,N_145,N_410);
xnor U888 (N_888,N_175,N_630);
and U889 (N_889,In_1076,N_472);
or U890 (N_890,In_987,N_423);
and U891 (N_891,N_664,N_697);
or U892 (N_892,In_69,In_484);
nor U893 (N_893,In_438,In_577);
nor U894 (N_894,N_699,N_686);
nor U895 (N_895,N_27,N_402);
or U896 (N_896,N_655,N_572);
nand U897 (N_897,In_405,N_638);
nand U898 (N_898,N_139,N_490);
nor U899 (N_899,In_530,In_1065);
nor U900 (N_900,N_893,N_94);
and U901 (N_901,In_1074,N_412);
or U902 (N_902,N_518,N_829);
nand U903 (N_903,In_411,In_413);
xnor U904 (N_904,In_524,N_342);
and U905 (N_905,N_733,In_83);
nand U906 (N_906,In_627,N_728);
or U907 (N_907,N_820,In_320);
and U908 (N_908,N_768,N_510);
and U909 (N_909,N_646,N_734);
and U910 (N_910,In_145,In_229);
nor U911 (N_911,N_499,N_804);
and U912 (N_912,N_642,N_827);
or U913 (N_913,N_874,N_522);
nand U914 (N_914,N_249,N_632);
xnor U915 (N_915,In_791,N_603);
nor U916 (N_916,N_899,In_52);
and U917 (N_917,N_786,N_863);
nor U918 (N_918,In_81,N_631);
or U919 (N_919,N_629,N_364);
and U920 (N_920,In_379,N_855);
xnor U921 (N_921,N_858,N_782);
and U922 (N_922,In_1087,N_667);
xor U923 (N_923,N_896,N_870);
xor U924 (N_924,N_645,In_814);
and U925 (N_925,N_851,In_620);
xnor U926 (N_926,In_1015,N_790);
nand U927 (N_927,N_753,N_759);
nand U928 (N_928,In_1262,N_723);
nor U929 (N_929,In_1471,In_1379);
nand U930 (N_930,N_776,N_325);
xor U931 (N_931,N_680,In_670);
nor U932 (N_932,N_626,N_849);
and U933 (N_933,N_365,N_669);
xnor U934 (N_934,N_621,In_954);
or U935 (N_935,In_378,In_13);
and U936 (N_936,N_700,In_978);
xor U937 (N_937,In_473,N_841);
and U938 (N_938,N_443,N_796);
or U939 (N_939,N_791,N_442);
xor U940 (N_940,N_291,N_550);
nor U941 (N_941,N_771,N_567);
or U942 (N_942,N_1,In_960);
or U943 (N_943,N_652,In_1429);
or U944 (N_944,N_890,In_125);
xor U945 (N_945,In_981,In_671);
xor U946 (N_946,In_532,N_816);
nor U947 (N_947,In_1101,In_794);
and U948 (N_948,N_857,N_524);
xor U949 (N_949,N_462,N_487);
xor U950 (N_950,In_203,N_888);
nor U951 (N_951,N_778,In_1246);
xor U952 (N_952,N_773,In_793);
and U953 (N_953,N_868,N_775);
nor U954 (N_954,In_301,In_988);
xnor U955 (N_955,In_334,N_312);
nand U956 (N_956,N_828,N_844);
and U957 (N_957,N_643,In_1414);
and U958 (N_958,N_634,N_602);
and U959 (N_959,In_565,N_381);
or U960 (N_960,N_757,In_660);
xnor U961 (N_961,N_704,N_732);
nand U962 (N_962,N_553,N_633);
xnor U963 (N_963,N_722,N_785);
nand U964 (N_964,N_770,N_830);
and U965 (N_965,In_1385,N_454);
nor U966 (N_966,N_476,N_683);
or U967 (N_967,In_1338,In_685);
xor U968 (N_968,N_836,N_391);
and U969 (N_969,In_197,N_864);
and U970 (N_970,In_355,N_891);
and U971 (N_971,N_853,N_265);
or U972 (N_972,N_506,N_519);
xor U973 (N_973,N_671,N_763);
and U974 (N_974,N_171,N_878);
or U975 (N_975,N_147,In_1035);
xnor U976 (N_976,In_1373,N_897);
xnor U977 (N_977,N_350,N_523);
and U978 (N_978,In_531,N_52);
or U979 (N_979,N_358,N_780);
nor U980 (N_980,N_672,N_663);
nand U981 (N_981,N_124,N_318);
and U982 (N_982,N_653,N_356);
xor U983 (N_983,In_871,N_661);
nand U984 (N_984,In_117,N_862);
or U985 (N_985,N_871,N_861);
or U986 (N_986,N_885,N_684);
nand U987 (N_987,In_780,N_826);
or U988 (N_988,N_668,N_115);
and U989 (N_989,N_737,N_401);
xnor U990 (N_990,N_323,N_295);
xnor U991 (N_991,N_378,N_744);
and U992 (N_992,N_876,N_867);
and U993 (N_993,In_997,In_1249);
xor U994 (N_994,In_1010,In_545);
nand U995 (N_995,In_1155,N_531);
and U996 (N_996,N_758,N_712);
nor U997 (N_997,In_1126,N_777);
and U998 (N_998,N_881,In_1060);
or U999 (N_999,In_192,N_207);
or U1000 (N_1000,In_371,In_1326);
or U1001 (N_1001,N_810,N_840);
xnor U1002 (N_1002,N_641,In_1073);
xor U1003 (N_1003,N_256,In_1300);
xnor U1004 (N_1004,In_1359,N_458);
or U1005 (N_1005,N_802,In_502);
nor U1006 (N_1006,In_1407,N_852);
xor U1007 (N_1007,N_341,In_322);
and U1008 (N_1008,N_741,N_363);
and U1009 (N_1009,N_281,N_681);
nor U1010 (N_1010,N_822,N_394);
nor U1011 (N_1011,In_1192,In_1303);
nand U1012 (N_1012,In_1398,N_886);
nand U1013 (N_1013,N_889,In_251);
and U1014 (N_1014,N_535,N_755);
xor U1015 (N_1015,In_24,N_623);
or U1016 (N_1016,N_149,N_526);
nand U1017 (N_1017,N_477,N_895);
and U1018 (N_1018,N_756,In_419);
and U1019 (N_1019,N_565,N_636);
nor U1020 (N_1020,N_497,In_1086);
xor U1021 (N_1021,N_808,N_26);
xor U1022 (N_1022,N_823,N_659);
or U1023 (N_1023,N_620,In_1427);
and U1024 (N_1024,In_363,N_282);
or U1025 (N_1025,N_729,In_637);
or U1026 (N_1026,N_656,N_71);
or U1027 (N_1027,In_878,N_847);
nand U1028 (N_1028,N_488,N_584);
xnor U1029 (N_1029,N_456,N_42);
nand U1030 (N_1030,N_801,N_703);
and U1031 (N_1031,N_170,N_15);
and U1032 (N_1032,N_86,N_814);
xor U1033 (N_1033,In_252,N_277);
nor U1034 (N_1034,N_217,In_1238);
and U1035 (N_1035,N_152,N_839);
nor U1036 (N_1036,N_599,N_548);
xor U1037 (N_1037,N_679,N_569);
xor U1038 (N_1038,N_736,In_224);
nor U1039 (N_1039,In_1339,N_332);
and U1040 (N_1040,N_348,N_882);
nor U1041 (N_1041,N_542,N_784);
or U1042 (N_1042,N_731,In_691);
nor U1043 (N_1043,N_781,N_769);
and U1044 (N_1044,In_1098,N_799);
and U1045 (N_1045,N_334,N_244);
nand U1046 (N_1046,N_798,N_446);
and U1047 (N_1047,N_807,N_408);
xnor U1048 (N_1048,In_1222,N_583);
nand U1049 (N_1049,N_617,In_1441);
xor U1050 (N_1050,N_575,N_875);
or U1051 (N_1051,In_88,N_1024);
or U1052 (N_1052,N_850,In_816);
xor U1053 (N_1053,N_846,N_794);
nand U1054 (N_1054,N_953,N_373);
and U1055 (N_1055,N_910,N_1011);
nor U1056 (N_1056,N_648,N_539);
or U1057 (N_1057,In_1095,In_931);
nor U1058 (N_1058,N_866,In_732);
xor U1059 (N_1059,N_961,N_954);
and U1060 (N_1060,N_944,N_779);
xor U1061 (N_1061,N_237,N_905);
nand U1062 (N_1062,N_609,N_1020);
or U1063 (N_1063,N_860,N_727);
xor U1064 (N_1064,N_939,In_1033);
or U1065 (N_1065,N_514,N_246);
or U1066 (N_1066,N_112,N_811);
xnor U1067 (N_1067,N_517,N_698);
or U1068 (N_1068,N_158,N_983);
nor U1069 (N_1069,N_662,In_936);
and U1070 (N_1070,N_1025,In_534);
and U1071 (N_1071,In_1034,In_759);
nor U1072 (N_1072,In_445,N_936);
nor U1073 (N_1073,N_696,In_1151);
and U1074 (N_1074,N_922,In_1011);
xnor U1075 (N_1075,N_692,N_433);
nand U1076 (N_1076,N_911,In_30);
and U1077 (N_1077,N_452,N_883);
or U1078 (N_1078,N_965,N_958);
nor U1079 (N_1079,In_707,N_976);
xor U1080 (N_1080,N_1049,N_990);
nor U1081 (N_1081,N_787,N_809);
nor U1082 (N_1082,N_748,In_1265);
and U1083 (N_1083,N_360,N_253);
nor U1084 (N_1084,N_106,N_973);
or U1085 (N_1085,In_641,N_29);
nand U1086 (N_1086,N_813,N_848);
nand U1087 (N_1087,N_766,N_596);
nand U1088 (N_1088,N_218,In_1214);
or U1089 (N_1089,In_1001,N_869);
or U1090 (N_1090,N_752,N_598);
nor U1091 (N_1091,N_783,In_695);
xnor U1092 (N_1092,N_474,N_430);
nand U1093 (N_1093,In_25,In_23);
nor U1094 (N_1094,N_397,N_819);
nand U1095 (N_1095,N_941,In_699);
and U1096 (N_1096,N_386,N_987);
or U1097 (N_1097,N_795,In_1357);
nor U1098 (N_1098,N_806,N_538);
nor U1099 (N_1099,N_651,N_545);
xnor U1100 (N_1100,In_944,N_1041);
nor U1101 (N_1101,N_824,N_963);
or U1102 (N_1102,N_19,In_384);
or U1103 (N_1103,N_995,In_771);
nor U1104 (N_1104,In_1274,In_554);
or U1105 (N_1105,In_136,N_400);
and U1106 (N_1106,N_832,N_1014);
and U1107 (N_1107,In_870,N_800);
nand U1108 (N_1108,N_600,N_721);
or U1109 (N_1109,N_788,N_713);
xnor U1110 (N_1110,N_511,N_119);
and U1111 (N_1111,In_209,N_843);
or U1112 (N_1112,N_563,In_736);
nor U1113 (N_1113,In_511,N_984);
nor U1114 (N_1114,In_777,N_455);
nor U1115 (N_1115,N_940,N_957);
nand U1116 (N_1116,N_329,N_835);
or U1117 (N_1117,N_719,N_131);
nor U1118 (N_1118,N_532,N_879);
and U1119 (N_1119,N_616,N_968);
xnor U1120 (N_1120,In_236,N_812);
xnor U1121 (N_1121,N_322,N_915);
xor U1122 (N_1122,N_909,In_1050);
nand U1123 (N_1123,N_1012,N_986);
xor U1124 (N_1124,N_245,N_193);
or U1125 (N_1125,In_676,N_1045);
nor U1126 (N_1126,N_738,N_366);
xor U1127 (N_1127,N_1046,N_357);
or U1128 (N_1128,In_893,In_1421);
xnor U1129 (N_1129,N_950,N_948);
or U1130 (N_1130,N_971,N_1003);
xnor U1131 (N_1131,N_1048,In_644);
nor U1132 (N_1132,N_873,N_792);
xnor U1133 (N_1133,N_694,N_1007);
nand U1134 (N_1134,In_634,N_720);
or U1135 (N_1135,N_613,N_762);
and U1136 (N_1136,N_913,In_44);
nand U1137 (N_1137,In_119,N_1035);
nor U1138 (N_1138,In_1183,N_1047);
xor U1139 (N_1139,N_979,N_833);
nand U1140 (N_1140,N_76,N_559);
xor U1141 (N_1141,N_904,N_649);
or U1142 (N_1142,N_1008,N_482);
nand U1143 (N_1143,In_450,N_1009);
xor U1144 (N_1144,N_494,N_750);
nand U1145 (N_1145,N_906,N_614);
nand U1146 (N_1146,N_1013,N_1031);
nor U1147 (N_1147,N_167,In_1212);
nand U1148 (N_1148,N_467,In_546);
nor U1149 (N_1149,N_774,N_607);
or U1150 (N_1150,N_938,N_1000);
nor U1151 (N_1151,N_821,N_308);
and U1152 (N_1152,N_912,N_1021);
nand U1153 (N_1153,N_142,N_1027);
or U1154 (N_1154,In_278,N_900);
nand U1155 (N_1155,In_993,N_865);
and U1156 (N_1156,N_854,N_347);
nor U1157 (N_1157,N_608,N_1043);
xnor U1158 (N_1158,N_980,N_92);
xnor U1159 (N_1159,N_916,N_932);
and U1160 (N_1160,N_925,N_974);
nand U1161 (N_1161,N_805,N_448);
nor U1162 (N_1162,In_894,In_302);
nand U1163 (N_1163,N_1036,In_1483);
or U1164 (N_1164,In_812,N_959);
and U1165 (N_1165,In_599,N_923);
nor U1166 (N_1166,N_746,N_998);
xnor U1167 (N_1167,N_877,N_924);
nor U1168 (N_1168,In_1248,N_880);
or U1169 (N_1169,N_742,N_370);
nor U1170 (N_1170,N_492,N_918);
nor U1171 (N_1171,N_1018,N_937);
or U1172 (N_1172,In_170,N_902);
and U1173 (N_1173,In_1174,N_981);
nor U1174 (N_1174,N_464,N_754);
or U1175 (N_1175,N_803,N_745);
nand U1176 (N_1176,N_294,In_504);
or U1177 (N_1177,N_533,N_859);
xnor U1178 (N_1178,N_930,N_901);
and U1179 (N_1179,N_690,N_970);
nand U1180 (N_1180,In_1406,N_7);
xnor U1181 (N_1181,N_929,N_927);
or U1182 (N_1182,In_1468,N_772);
and U1183 (N_1183,N_837,N_985);
nor U1184 (N_1184,N_817,N_917);
or U1185 (N_1185,N_992,N_892);
and U1186 (N_1186,N_991,N_993);
or U1187 (N_1187,N_825,In_375);
or U1188 (N_1188,N_491,In_479);
nor U1189 (N_1189,N_946,N_1002);
and U1190 (N_1190,N_1006,In_607);
or U1191 (N_1191,In_1195,N_872);
or U1192 (N_1192,N_38,In_1255);
and U1193 (N_1193,N_831,N_920);
xor U1194 (N_1194,N_994,N_164);
and U1195 (N_1195,N_972,In_133);
nor U1196 (N_1196,N_815,In_1277);
and U1197 (N_1197,N_1030,N_1023);
and U1198 (N_1198,N_928,N_914);
nand U1199 (N_1199,N_314,N_943);
and U1200 (N_1200,N_1129,N_1004);
or U1201 (N_1201,N_1123,N_1016);
xnor U1202 (N_1202,N_955,N_997);
and U1203 (N_1203,N_1101,N_1090);
xnor U1204 (N_1204,N_1142,N_1166);
nand U1205 (N_1205,N_1195,N_1116);
or U1206 (N_1206,N_760,N_926);
nor U1207 (N_1207,In_191,N_1130);
nor U1208 (N_1208,N_622,N_1125);
xor U1209 (N_1209,N_1079,N_708);
nand U1210 (N_1210,N_1120,N_1115);
and U1211 (N_1211,N_949,N_1033);
or U1212 (N_1212,N_1022,N_962);
or U1213 (N_1213,N_162,N_856);
nor U1214 (N_1214,N_1183,N_471);
nand U1215 (N_1215,N_691,N_919);
or U1216 (N_1216,N_1122,N_1155);
xnor U1217 (N_1217,N_627,N_1039);
and U1218 (N_1218,N_705,N_1105);
and U1219 (N_1219,N_122,N_1073);
nand U1220 (N_1220,N_610,N_1065);
nor U1221 (N_1221,N_1095,N_1177);
or U1222 (N_1222,N_637,N_1051);
nor U1223 (N_1223,N_1067,N_1188);
and U1224 (N_1224,In_446,N_887);
nor U1225 (N_1225,N_1159,N_764);
nor U1226 (N_1226,N_25,N_1179);
xnor U1227 (N_1227,N_1121,N_1174);
nor U1228 (N_1228,N_1133,N_767);
xor U1229 (N_1229,N_999,N_1141);
nor U1230 (N_1230,In_317,N_1182);
nor U1231 (N_1231,N_1102,N_907);
or U1232 (N_1232,N_1199,N_1088);
nor U1233 (N_1233,N_1042,N_615);
xor U1234 (N_1234,N_359,In_541);
nor U1235 (N_1235,N_3,N_1153);
nor U1236 (N_1236,N_1143,N_1157);
or U1237 (N_1237,N_1059,N_530);
nor U1238 (N_1238,In_605,In_50);
nor U1239 (N_1239,N_975,N_1185);
xnor U1240 (N_1240,N_414,N_818);
nor U1241 (N_1241,N_964,N_1098);
and U1242 (N_1242,N_168,In_440);
nand U1243 (N_1243,N_1107,N_1072);
nand U1244 (N_1244,N_1032,N_903);
xnor U1245 (N_1245,In_370,In_1258);
and U1246 (N_1246,N_951,N_1171);
xnor U1247 (N_1247,In_84,N_1147);
nor U1248 (N_1248,N_1158,N_1063);
xnor U1249 (N_1249,N_1162,N_1053);
and U1250 (N_1250,N_1001,N_898);
or U1251 (N_1251,N_1092,N_1167);
nor U1252 (N_1252,N_1112,N_1074);
nor U1253 (N_1253,N_202,N_1138);
nor U1254 (N_1254,N_935,N_789);
or U1255 (N_1255,In_877,N_1198);
nor U1256 (N_1256,N_1113,N_403);
xor U1257 (N_1257,N_1170,N_1019);
or U1258 (N_1258,In_196,N_1194);
xor U1259 (N_1259,In_659,N_982);
or U1260 (N_1260,N_1103,N_1058);
nor U1261 (N_1261,N_353,In_1234);
xor U1262 (N_1262,In_578,In_1377);
nor U1263 (N_1263,N_1144,N_1061);
or U1264 (N_1264,N_650,N_1178);
xnor U1265 (N_1265,N_1081,N_1069);
and U1266 (N_1266,N_1137,N_1068);
and U1267 (N_1267,N_1131,N_996);
or U1268 (N_1268,N_675,N_977);
nor U1269 (N_1269,N_934,In_441);
and U1270 (N_1270,N_960,N_1111);
nor U1271 (N_1271,In_1288,N_1034);
nor U1272 (N_1272,N_1064,N_305);
xnor U1273 (N_1273,In_529,N_1165);
nor U1274 (N_1274,N_1151,N_1082);
or U1275 (N_1275,N_1091,N_1117);
or U1276 (N_1276,N_1028,In_401);
nor U1277 (N_1277,N_969,N_989);
xor U1278 (N_1278,N_1128,N_1100);
or U1279 (N_1279,N_942,N_1163);
or U1280 (N_1280,N_947,N_31);
nor U1281 (N_1281,N_1037,N_894);
or U1282 (N_1282,N_1168,N_1134);
and U1283 (N_1283,N_1057,N_1191);
nor U1284 (N_1284,N_751,N_838);
or U1285 (N_1285,N_1118,N_1089);
and U1286 (N_1286,N_1005,N_1093);
xnor U1287 (N_1287,N_1124,N_1148);
nor U1288 (N_1288,N_1062,N_1094);
xnor U1289 (N_1289,N_1017,N_1075);
xnor U1290 (N_1290,In_1351,N_1193);
xnor U1291 (N_1291,N_1040,N_1126);
and U1292 (N_1292,N_1096,N_1139);
nor U1293 (N_1293,N_512,N_527);
nand U1294 (N_1294,In_876,N_1060);
nor U1295 (N_1295,N_1026,N_1110);
xnor U1296 (N_1296,N_1106,In_1210);
nor U1297 (N_1297,N_574,In_582);
or U1298 (N_1298,In_1376,N_1169);
nor U1299 (N_1299,N_931,In_297);
xnor U1300 (N_1300,N_283,N_1071);
and U1301 (N_1301,N_1173,N_1149);
xor U1302 (N_1302,N_726,N_1085);
nand U1303 (N_1303,N_286,N_884);
and U1304 (N_1304,N_1083,N_1135);
nor U1305 (N_1305,N_1189,N_1187);
or U1306 (N_1306,N_1186,N_1087);
xor U1307 (N_1307,N_1010,N_1119);
and U1308 (N_1308,N_1197,N_956);
or U1309 (N_1309,N_1181,N_1161);
or U1310 (N_1310,N_1196,N_725);
xnor U1311 (N_1311,In_131,N_945);
or U1312 (N_1312,N_1052,N_1164);
xor U1313 (N_1313,N_834,N_1156);
or U1314 (N_1314,N_1086,N_1175);
nor U1315 (N_1315,N_1160,N_933);
nand U1316 (N_1316,In_485,N_1066);
nor U1317 (N_1317,N_273,N_1104);
or U1318 (N_1318,N_1146,N_1180);
nand U1319 (N_1319,N_1127,N_1145);
xnor U1320 (N_1320,N_921,N_1150);
and U1321 (N_1321,N_1114,N_793);
or U1322 (N_1322,N_845,N_1056);
nor U1323 (N_1323,N_335,N_1097);
nand U1324 (N_1324,N_324,N_1190);
xor U1325 (N_1325,N_1078,N_1184);
and U1326 (N_1326,N_1084,N_952);
nor U1327 (N_1327,N_424,N_988);
and U1328 (N_1328,N_1154,N_1029);
nand U1329 (N_1329,N_1152,N_765);
or U1330 (N_1330,N_501,N_1132);
nor U1331 (N_1331,N_460,N_966);
or U1332 (N_1332,N_317,N_1099);
or U1333 (N_1333,N_1109,N_1055);
or U1334 (N_1334,N_842,N_1070);
xnor U1335 (N_1335,N_1108,N_1176);
nor U1336 (N_1336,N_761,N_1192);
nand U1337 (N_1337,N_908,N_1077);
nor U1338 (N_1338,N_192,N_1076);
and U1339 (N_1339,N_797,In_1042);
and U1340 (N_1340,In_1416,N_1044);
and U1341 (N_1341,N_1050,N_587);
and U1342 (N_1342,N_1136,N_1038);
and U1343 (N_1343,N_1015,N_100);
and U1344 (N_1344,N_1140,N_1172);
or U1345 (N_1345,N_557,In_628);
nor U1346 (N_1346,N_978,N_967);
and U1347 (N_1347,In_1492,In_1363);
and U1348 (N_1348,N_606,In_238);
or U1349 (N_1349,N_1054,N_1080);
nand U1350 (N_1350,N_1212,N_1333);
nor U1351 (N_1351,N_1302,N_1255);
nand U1352 (N_1352,N_1233,N_1214);
or U1353 (N_1353,N_1304,N_1329);
nor U1354 (N_1354,N_1340,N_1344);
nand U1355 (N_1355,N_1232,N_1262);
xnor U1356 (N_1356,N_1237,N_1349);
and U1357 (N_1357,N_1245,N_1338);
or U1358 (N_1358,N_1253,N_1322);
xnor U1359 (N_1359,N_1246,N_1226);
nor U1360 (N_1360,N_1293,N_1336);
or U1361 (N_1361,N_1308,N_1321);
nand U1362 (N_1362,N_1201,N_1292);
nand U1363 (N_1363,N_1238,N_1263);
nand U1364 (N_1364,N_1217,N_1317);
nand U1365 (N_1365,N_1240,N_1231);
and U1366 (N_1366,N_1346,N_1319);
and U1367 (N_1367,N_1347,N_1331);
xor U1368 (N_1368,N_1256,N_1229);
xnor U1369 (N_1369,N_1290,N_1258);
or U1370 (N_1370,N_1328,N_1264);
nor U1371 (N_1371,N_1320,N_1247);
or U1372 (N_1372,N_1330,N_1297);
nor U1373 (N_1373,N_1335,N_1224);
nor U1374 (N_1374,N_1342,N_1220);
or U1375 (N_1375,N_1339,N_1326);
or U1376 (N_1376,N_1236,N_1307);
or U1377 (N_1377,N_1209,N_1306);
or U1378 (N_1378,N_1267,N_1222);
nand U1379 (N_1379,N_1341,N_1218);
nand U1380 (N_1380,N_1219,N_1273);
xnor U1381 (N_1381,N_1289,N_1227);
nand U1382 (N_1382,N_1301,N_1310);
or U1383 (N_1383,N_1343,N_1332);
xor U1384 (N_1384,N_1295,N_1239);
xnor U1385 (N_1385,N_1287,N_1313);
and U1386 (N_1386,N_1327,N_1210);
xor U1387 (N_1387,N_1337,N_1325);
and U1388 (N_1388,N_1270,N_1316);
nand U1389 (N_1389,N_1276,N_1211);
nand U1390 (N_1390,N_1282,N_1235);
and U1391 (N_1391,N_1266,N_1241);
nor U1392 (N_1392,N_1348,N_1285);
and U1393 (N_1393,N_1294,N_1206);
or U1394 (N_1394,N_1334,N_1268);
nor U1395 (N_1395,N_1234,N_1265);
nand U1396 (N_1396,N_1252,N_1323);
or U1397 (N_1397,N_1281,N_1284);
and U1398 (N_1398,N_1205,N_1223);
and U1399 (N_1399,N_1261,N_1260);
and U1400 (N_1400,N_1251,N_1280);
or U1401 (N_1401,N_1202,N_1208);
or U1402 (N_1402,N_1269,N_1291);
nand U1403 (N_1403,N_1216,N_1272);
nor U1404 (N_1404,N_1300,N_1324);
nor U1405 (N_1405,N_1345,N_1225);
xnor U1406 (N_1406,N_1315,N_1303);
nor U1407 (N_1407,N_1215,N_1228);
or U1408 (N_1408,N_1296,N_1299);
and U1409 (N_1409,N_1203,N_1277);
xnor U1410 (N_1410,N_1257,N_1283);
nor U1411 (N_1411,N_1249,N_1242);
nand U1412 (N_1412,N_1311,N_1275);
nand U1413 (N_1413,N_1221,N_1271);
and U1414 (N_1414,N_1250,N_1230);
nand U1415 (N_1415,N_1254,N_1279);
xor U1416 (N_1416,N_1286,N_1278);
or U1417 (N_1417,N_1288,N_1244);
and U1418 (N_1418,N_1248,N_1314);
nand U1419 (N_1419,N_1243,N_1312);
xor U1420 (N_1420,N_1200,N_1213);
nor U1421 (N_1421,N_1207,N_1318);
and U1422 (N_1422,N_1274,N_1259);
and U1423 (N_1423,N_1298,N_1305);
or U1424 (N_1424,N_1204,N_1309);
or U1425 (N_1425,N_1324,N_1297);
xor U1426 (N_1426,N_1255,N_1279);
xor U1427 (N_1427,N_1300,N_1253);
or U1428 (N_1428,N_1271,N_1262);
or U1429 (N_1429,N_1243,N_1208);
nand U1430 (N_1430,N_1253,N_1254);
xnor U1431 (N_1431,N_1283,N_1267);
or U1432 (N_1432,N_1213,N_1344);
xnor U1433 (N_1433,N_1298,N_1292);
nand U1434 (N_1434,N_1307,N_1232);
nor U1435 (N_1435,N_1244,N_1251);
nor U1436 (N_1436,N_1253,N_1245);
or U1437 (N_1437,N_1339,N_1243);
or U1438 (N_1438,N_1298,N_1277);
nor U1439 (N_1439,N_1294,N_1347);
xor U1440 (N_1440,N_1225,N_1335);
and U1441 (N_1441,N_1324,N_1341);
xnor U1442 (N_1442,N_1288,N_1320);
and U1443 (N_1443,N_1326,N_1205);
and U1444 (N_1444,N_1219,N_1314);
xor U1445 (N_1445,N_1303,N_1207);
nand U1446 (N_1446,N_1281,N_1210);
and U1447 (N_1447,N_1286,N_1291);
nor U1448 (N_1448,N_1200,N_1348);
or U1449 (N_1449,N_1223,N_1277);
xor U1450 (N_1450,N_1328,N_1274);
nor U1451 (N_1451,N_1214,N_1338);
nand U1452 (N_1452,N_1340,N_1208);
or U1453 (N_1453,N_1259,N_1278);
nand U1454 (N_1454,N_1271,N_1316);
nor U1455 (N_1455,N_1228,N_1325);
or U1456 (N_1456,N_1329,N_1225);
and U1457 (N_1457,N_1238,N_1264);
xnor U1458 (N_1458,N_1273,N_1318);
xnor U1459 (N_1459,N_1308,N_1326);
nor U1460 (N_1460,N_1345,N_1337);
nor U1461 (N_1461,N_1228,N_1229);
xor U1462 (N_1462,N_1280,N_1209);
and U1463 (N_1463,N_1224,N_1257);
or U1464 (N_1464,N_1329,N_1246);
nand U1465 (N_1465,N_1340,N_1206);
and U1466 (N_1466,N_1299,N_1346);
nor U1467 (N_1467,N_1334,N_1224);
and U1468 (N_1468,N_1307,N_1267);
nor U1469 (N_1469,N_1266,N_1276);
nor U1470 (N_1470,N_1212,N_1290);
or U1471 (N_1471,N_1260,N_1270);
and U1472 (N_1472,N_1244,N_1322);
nor U1473 (N_1473,N_1253,N_1220);
nor U1474 (N_1474,N_1290,N_1205);
nand U1475 (N_1475,N_1269,N_1258);
and U1476 (N_1476,N_1297,N_1259);
and U1477 (N_1477,N_1284,N_1261);
nand U1478 (N_1478,N_1207,N_1257);
nor U1479 (N_1479,N_1254,N_1269);
nand U1480 (N_1480,N_1257,N_1273);
or U1481 (N_1481,N_1303,N_1214);
and U1482 (N_1482,N_1322,N_1225);
and U1483 (N_1483,N_1320,N_1294);
nand U1484 (N_1484,N_1207,N_1256);
and U1485 (N_1485,N_1251,N_1320);
and U1486 (N_1486,N_1291,N_1328);
or U1487 (N_1487,N_1282,N_1341);
or U1488 (N_1488,N_1293,N_1222);
xnor U1489 (N_1489,N_1225,N_1271);
and U1490 (N_1490,N_1228,N_1201);
or U1491 (N_1491,N_1313,N_1251);
and U1492 (N_1492,N_1338,N_1263);
xor U1493 (N_1493,N_1280,N_1284);
xor U1494 (N_1494,N_1298,N_1249);
nand U1495 (N_1495,N_1211,N_1210);
nor U1496 (N_1496,N_1290,N_1281);
nor U1497 (N_1497,N_1201,N_1299);
nor U1498 (N_1498,N_1304,N_1331);
or U1499 (N_1499,N_1283,N_1304);
or U1500 (N_1500,N_1479,N_1418);
xnor U1501 (N_1501,N_1357,N_1455);
and U1502 (N_1502,N_1411,N_1497);
and U1503 (N_1503,N_1358,N_1382);
nand U1504 (N_1504,N_1463,N_1424);
nor U1505 (N_1505,N_1498,N_1428);
or U1506 (N_1506,N_1448,N_1452);
and U1507 (N_1507,N_1400,N_1480);
xor U1508 (N_1508,N_1457,N_1364);
xnor U1509 (N_1509,N_1441,N_1461);
or U1510 (N_1510,N_1392,N_1354);
and U1511 (N_1511,N_1467,N_1446);
nor U1512 (N_1512,N_1360,N_1359);
nor U1513 (N_1513,N_1485,N_1389);
or U1514 (N_1514,N_1414,N_1372);
nor U1515 (N_1515,N_1491,N_1397);
or U1516 (N_1516,N_1390,N_1366);
or U1517 (N_1517,N_1406,N_1384);
and U1518 (N_1518,N_1427,N_1496);
xor U1519 (N_1519,N_1477,N_1368);
nor U1520 (N_1520,N_1399,N_1379);
and U1521 (N_1521,N_1432,N_1425);
or U1522 (N_1522,N_1429,N_1373);
xor U1523 (N_1523,N_1458,N_1493);
or U1524 (N_1524,N_1492,N_1470);
and U1525 (N_1525,N_1464,N_1468);
or U1526 (N_1526,N_1421,N_1356);
nand U1527 (N_1527,N_1473,N_1495);
xor U1528 (N_1528,N_1405,N_1436);
nand U1529 (N_1529,N_1404,N_1462);
nor U1530 (N_1530,N_1499,N_1365);
nand U1531 (N_1531,N_1444,N_1361);
nor U1532 (N_1532,N_1430,N_1385);
xnor U1533 (N_1533,N_1393,N_1383);
nor U1534 (N_1534,N_1387,N_1442);
xnor U1535 (N_1535,N_1370,N_1434);
xor U1536 (N_1536,N_1386,N_1410);
nor U1537 (N_1537,N_1409,N_1435);
or U1538 (N_1538,N_1433,N_1471);
nor U1539 (N_1539,N_1417,N_1466);
and U1540 (N_1540,N_1391,N_1402);
and U1541 (N_1541,N_1419,N_1460);
and U1542 (N_1542,N_1403,N_1423);
nand U1543 (N_1543,N_1380,N_1367);
nand U1544 (N_1544,N_1353,N_1355);
nand U1545 (N_1545,N_1447,N_1396);
nand U1546 (N_1546,N_1431,N_1453);
nand U1547 (N_1547,N_1352,N_1478);
and U1548 (N_1548,N_1440,N_1490);
or U1549 (N_1549,N_1487,N_1413);
or U1550 (N_1550,N_1476,N_1420);
xnor U1551 (N_1551,N_1443,N_1451);
nand U1552 (N_1552,N_1472,N_1351);
nor U1553 (N_1553,N_1456,N_1489);
nand U1554 (N_1554,N_1450,N_1474);
or U1555 (N_1555,N_1376,N_1375);
xor U1556 (N_1556,N_1454,N_1494);
and U1557 (N_1557,N_1416,N_1395);
nor U1558 (N_1558,N_1377,N_1449);
nor U1559 (N_1559,N_1437,N_1407);
xor U1560 (N_1560,N_1381,N_1481);
nand U1561 (N_1561,N_1484,N_1415);
nand U1562 (N_1562,N_1388,N_1369);
nand U1563 (N_1563,N_1362,N_1398);
nand U1564 (N_1564,N_1488,N_1482);
and U1565 (N_1565,N_1378,N_1475);
or U1566 (N_1566,N_1408,N_1422);
xor U1567 (N_1567,N_1426,N_1486);
and U1568 (N_1568,N_1394,N_1469);
xor U1569 (N_1569,N_1483,N_1459);
xor U1570 (N_1570,N_1445,N_1438);
xor U1571 (N_1571,N_1401,N_1439);
xor U1572 (N_1572,N_1350,N_1412);
and U1573 (N_1573,N_1465,N_1374);
or U1574 (N_1574,N_1363,N_1371);
nor U1575 (N_1575,N_1463,N_1490);
and U1576 (N_1576,N_1364,N_1352);
nor U1577 (N_1577,N_1358,N_1495);
nor U1578 (N_1578,N_1498,N_1363);
or U1579 (N_1579,N_1397,N_1480);
and U1580 (N_1580,N_1472,N_1497);
nor U1581 (N_1581,N_1362,N_1477);
nand U1582 (N_1582,N_1424,N_1356);
nand U1583 (N_1583,N_1409,N_1382);
or U1584 (N_1584,N_1408,N_1351);
or U1585 (N_1585,N_1411,N_1453);
nor U1586 (N_1586,N_1382,N_1456);
or U1587 (N_1587,N_1381,N_1359);
xor U1588 (N_1588,N_1420,N_1493);
nor U1589 (N_1589,N_1460,N_1413);
or U1590 (N_1590,N_1393,N_1402);
and U1591 (N_1591,N_1411,N_1387);
xnor U1592 (N_1592,N_1369,N_1475);
nor U1593 (N_1593,N_1483,N_1369);
or U1594 (N_1594,N_1421,N_1405);
nand U1595 (N_1595,N_1387,N_1375);
and U1596 (N_1596,N_1439,N_1358);
or U1597 (N_1597,N_1393,N_1424);
and U1598 (N_1598,N_1444,N_1460);
xnor U1599 (N_1599,N_1477,N_1380);
xnor U1600 (N_1600,N_1472,N_1467);
nor U1601 (N_1601,N_1494,N_1492);
or U1602 (N_1602,N_1400,N_1424);
or U1603 (N_1603,N_1405,N_1439);
or U1604 (N_1604,N_1365,N_1351);
or U1605 (N_1605,N_1370,N_1435);
nor U1606 (N_1606,N_1432,N_1428);
nor U1607 (N_1607,N_1485,N_1351);
and U1608 (N_1608,N_1406,N_1492);
nand U1609 (N_1609,N_1449,N_1381);
and U1610 (N_1610,N_1475,N_1445);
xnor U1611 (N_1611,N_1368,N_1365);
or U1612 (N_1612,N_1469,N_1478);
and U1613 (N_1613,N_1471,N_1421);
xor U1614 (N_1614,N_1354,N_1362);
nand U1615 (N_1615,N_1477,N_1397);
and U1616 (N_1616,N_1381,N_1360);
and U1617 (N_1617,N_1450,N_1444);
nor U1618 (N_1618,N_1373,N_1439);
xor U1619 (N_1619,N_1455,N_1386);
xor U1620 (N_1620,N_1380,N_1474);
nor U1621 (N_1621,N_1453,N_1440);
nor U1622 (N_1622,N_1455,N_1471);
nand U1623 (N_1623,N_1426,N_1461);
nor U1624 (N_1624,N_1353,N_1477);
nor U1625 (N_1625,N_1410,N_1459);
nand U1626 (N_1626,N_1489,N_1447);
nand U1627 (N_1627,N_1353,N_1427);
nor U1628 (N_1628,N_1406,N_1388);
xnor U1629 (N_1629,N_1431,N_1352);
xor U1630 (N_1630,N_1362,N_1481);
xor U1631 (N_1631,N_1378,N_1352);
and U1632 (N_1632,N_1378,N_1460);
and U1633 (N_1633,N_1458,N_1473);
and U1634 (N_1634,N_1388,N_1471);
and U1635 (N_1635,N_1436,N_1499);
nand U1636 (N_1636,N_1481,N_1351);
xor U1637 (N_1637,N_1357,N_1475);
and U1638 (N_1638,N_1487,N_1477);
or U1639 (N_1639,N_1456,N_1472);
and U1640 (N_1640,N_1439,N_1402);
nor U1641 (N_1641,N_1359,N_1409);
or U1642 (N_1642,N_1388,N_1476);
or U1643 (N_1643,N_1462,N_1355);
and U1644 (N_1644,N_1373,N_1492);
xnor U1645 (N_1645,N_1436,N_1475);
or U1646 (N_1646,N_1487,N_1492);
nand U1647 (N_1647,N_1492,N_1410);
and U1648 (N_1648,N_1389,N_1372);
nand U1649 (N_1649,N_1437,N_1423);
nor U1650 (N_1650,N_1524,N_1534);
xor U1651 (N_1651,N_1633,N_1646);
nor U1652 (N_1652,N_1559,N_1502);
nor U1653 (N_1653,N_1576,N_1512);
nor U1654 (N_1654,N_1574,N_1507);
or U1655 (N_1655,N_1552,N_1506);
nand U1656 (N_1656,N_1583,N_1518);
nor U1657 (N_1657,N_1644,N_1551);
or U1658 (N_1658,N_1515,N_1571);
nor U1659 (N_1659,N_1604,N_1620);
nand U1660 (N_1660,N_1636,N_1596);
or U1661 (N_1661,N_1626,N_1527);
nand U1662 (N_1662,N_1594,N_1614);
and U1663 (N_1663,N_1532,N_1643);
nor U1664 (N_1664,N_1549,N_1537);
xor U1665 (N_1665,N_1582,N_1631);
or U1666 (N_1666,N_1589,N_1569);
nor U1667 (N_1667,N_1553,N_1611);
and U1668 (N_1668,N_1557,N_1516);
nor U1669 (N_1669,N_1531,N_1560);
nor U1670 (N_1670,N_1641,N_1529);
and U1671 (N_1671,N_1555,N_1615);
or U1672 (N_1672,N_1592,N_1563);
xor U1673 (N_1673,N_1562,N_1606);
xnor U1674 (N_1674,N_1639,N_1522);
or U1675 (N_1675,N_1547,N_1610);
and U1676 (N_1676,N_1586,N_1587);
or U1677 (N_1677,N_1588,N_1509);
nor U1678 (N_1678,N_1541,N_1600);
xnor U1679 (N_1679,N_1558,N_1623);
nor U1680 (N_1680,N_1621,N_1580);
and U1681 (N_1681,N_1536,N_1649);
nand U1682 (N_1682,N_1591,N_1573);
and U1683 (N_1683,N_1567,N_1540);
nor U1684 (N_1684,N_1629,N_1533);
xor U1685 (N_1685,N_1564,N_1519);
nor U1686 (N_1686,N_1544,N_1648);
and U1687 (N_1687,N_1622,N_1616);
nor U1688 (N_1688,N_1538,N_1548);
and U1689 (N_1689,N_1513,N_1550);
or U1690 (N_1690,N_1647,N_1598);
xnor U1691 (N_1691,N_1561,N_1572);
xnor U1692 (N_1692,N_1546,N_1505);
or U1693 (N_1693,N_1595,N_1632);
nor U1694 (N_1694,N_1638,N_1637);
xor U1695 (N_1695,N_1617,N_1618);
or U1696 (N_1696,N_1503,N_1630);
and U1697 (N_1697,N_1517,N_1526);
nand U1698 (N_1698,N_1508,N_1543);
xnor U1699 (N_1699,N_1528,N_1575);
and U1700 (N_1700,N_1578,N_1599);
xnor U1701 (N_1701,N_1613,N_1584);
xor U1702 (N_1702,N_1510,N_1634);
xnor U1703 (N_1703,N_1642,N_1521);
nor U1704 (N_1704,N_1570,N_1514);
and U1705 (N_1705,N_1627,N_1504);
nor U1706 (N_1706,N_1590,N_1605);
nor U1707 (N_1707,N_1568,N_1593);
xnor U1708 (N_1708,N_1597,N_1556);
xnor U1709 (N_1709,N_1523,N_1554);
nor U1710 (N_1710,N_1609,N_1525);
and U1711 (N_1711,N_1500,N_1585);
xnor U1712 (N_1712,N_1530,N_1539);
or U1713 (N_1713,N_1535,N_1581);
nor U1714 (N_1714,N_1566,N_1628);
xor U1715 (N_1715,N_1619,N_1511);
nand U1716 (N_1716,N_1603,N_1601);
xor U1717 (N_1717,N_1625,N_1520);
xor U1718 (N_1718,N_1579,N_1602);
xor U1719 (N_1719,N_1577,N_1612);
and U1720 (N_1720,N_1635,N_1542);
or U1721 (N_1721,N_1501,N_1607);
xor U1722 (N_1722,N_1645,N_1545);
xor U1723 (N_1723,N_1608,N_1640);
nand U1724 (N_1724,N_1624,N_1565);
xor U1725 (N_1725,N_1572,N_1558);
nand U1726 (N_1726,N_1555,N_1560);
nand U1727 (N_1727,N_1618,N_1552);
xnor U1728 (N_1728,N_1540,N_1607);
xor U1729 (N_1729,N_1564,N_1588);
nor U1730 (N_1730,N_1604,N_1637);
xor U1731 (N_1731,N_1601,N_1599);
or U1732 (N_1732,N_1573,N_1623);
or U1733 (N_1733,N_1512,N_1563);
xnor U1734 (N_1734,N_1620,N_1556);
nor U1735 (N_1735,N_1520,N_1598);
xnor U1736 (N_1736,N_1606,N_1594);
and U1737 (N_1737,N_1520,N_1500);
nor U1738 (N_1738,N_1616,N_1578);
nand U1739 (N_1739,N_1555,N_1539);
or U1740 (N_1740,N_1607,N_1640);
nand U1741 (N_1741,N_1596,N_1645);
or U1742 (N_1742,N_1520,N_1589);
nand U1743 (N_1743,N_1576,N_1619);
xor U1744 (N_1744,N_1632,N_1526);
xnor U1745 (N_1745,N_1541,N_1626);
xnor U1746 (N_1746,N_1532,N_1612);
nor U1747 (N_1747,N_1539,N_1631);
xnor U1748 (N_1748,N_1649,N_1524);
nor U1749 (N_1749,N_1532,N_1588);
and U1750 (N_1750,N_1581,N_1525);
and U1751 (N_1751,N_1635,N_1639);
xnor U1752 (N_1752,N_1646,N_1641);
xnor U1753 (N_1753,N_1606,N_1618);
and U1754 (N_1754,N_1619,N_1512);
and U1755 (N_1755,N_1557,N_1605);
nand U1756 (N_1756,N_1523,N_1516);
xnor U1757 (N_1757,N_1563,N_1608);
xor U1758 (N_1758,N_1583,N_1546);
or U1759 (N_1759,N_1544,N_1565);
xor U1760 (N_1760,N_1521,N_1602);
xnor U1761 (N_1761,N_1551,N_1509);
nand U1762 (N_1762,N_1520,N_1512);
nand U1763 (N_1763,N_1586,N_1570);
or U1764 (N_1764,N_1639,N_1511);
xor U1765 (N_1765,N_1563,N_1529);
nor U1766 (N_1766,N_1531,N_1624);
or U1767 (N_1767,N_1556,N_1583);
nand U1768 (N_1768,N_1575,N_1560);
xnor U1769 (N_1769,N_1550,N_1571);
and U1770 (N_1770,N_1630,N_1547);
or U1771 (N_1771,N_1512,N_1575);
and U1772 (N_1772,N_1566,N_1609);
and U1773 (N_1773,N_1648,N_1596);
nor U1774 (N_1774,N_1554,N_1582);
and U1775 (N_1775,N_1638,N_1531);
nand U1776 (N_1776,N_1571,N_1591);
nor U1777 (N_1777,N_1589,N_1537);
and U1778 (N_1778,N_1647,N_1631);
nand U1779 (N_1779,N_1500,N_1628);
or U1780 (N_1780,N_1619,N_1565);
and U1781 (N_1781,N_1591,N_1579);
nor U1782 (N_1782,N_1546,N_1580);
nand U1783 (N_1783,N_1578,N_1568);
and U1784 (N_1784,N_1611,N_1502);
xor U1785 (N_1785,N_1596,N_1557);
or U1786 (N_1786,N_1570,N_1648);
or U1787 (N_1787,N_1624,N_1526);
or U1788 (N_1788,N_1548,N_1522);
nor U1789 (N_1789,N_1587,N_1636);
and U1790 (N_1790,N_1615,N_1550);
nor U1791 (N_1791,N_1624,N_1516);
nand U1792 (N_1792,N_1549,N_1620);
nor U1793 (N_1793,N_1570,N_1522);
or U1794 (N_1794,N_1542,N_1565);
or U1795 (N_1795,N_1528,N_1594);
nor U1796 (N_1796,N_1587,N_1643);
xnor U1797 (N_1797,N_1594,N_1526);
or U1798 (N_1798,N_1511,N_1503);
and U1799 (N_1799,N_1515,N_1501);
xor U1800 (N_1800,N_1717,N_1751);
nor U1801 (N_1801,N_1707,N_1711);
nor U1802 (N_1802,N_1738,N_1785);
nor U1803 (N_1803,N_1752,N_1715);
and U1804 (N_1804,N_1680,N_1788);
xnor U1805 (N_1805,N_1676,N_1696);
xor U1806 (N_1806,N_1710,N_1749);
and U1807 (N_1807,N_1661,N_1678);
or U1808 (N_1808,N_1779,N_1699);
xnor U1809 (N_1809,N_1768,N_1669);
and U1810 (N_1810,N_1700,N_1798);
or U1811 (N_1811,N_1697,N_1683);
or U1812 (N_1812,N_1784,N_1730);
xnor U1813 (N_1813,N_1652,N_1688);
xnor U1814 (N_1814,N_1681,N_1799);
xor U1815 (N_1815,N_1761,N_1735);
or U1816 (N_1816,N_1775,N_1682);
or U1817 (N_1817,N_1684,N_1698);
or U1818 (N_1818,N_1674,N_1757);
nor U1819 (N_1819,N_1767,N_1745);
or U1820 (N_1820,N_1693,N_1706);
nor U1821 (N_1821,N_1703,N_1662);
nor U1822 (N_1822,N_1748,N_1694);
nand U1823 (N_1823,N_1763,N_1685);
and U1824 (N_1824,N_1650,N_1721);
nor U1825 (N_1825,N_1781,N_1732);
xor U1826 (N_1826,N_1714,N_1769);
and U1827 (N_1827,N_1764,N_1789);
xnor U1828 (N_1828,N_1720,N_1754);
nor U1829 (N_1829,N_1667,N_1737);
or U1830 (N_1830,N_1759,N_1744);
and U1831 (N_1831,N_1670,N_1786);
or U1832 (N_1832,N_1672,N_1651);
nor U1833 (N_1833,N_1731,N_1762);
xnor U1834 (N_1834,N_1687,N_1690);
nor U1835 (N_1835,N_1760,N_1774);
xnor U1836 (N_1836,N_1666,N_1782);
nand U1837 (N_1837,N_1664,N_1770);
nand U1838 (N_1838,N_1713,N_1691);
nand U1839 (N_1839,N_1655,N_1692);
xor U1840 (N_1840,N_1658,N_1704);
and U1841 (N_1841,N_1716,N_1709);
and U1842 (N_1842,N_1665,N_1743);
and U1843 (N_1843,N_1728,N_1657);
xor U1844 (N_1844,N_1755,N_1695);
xnor U1845 (N_1845,N_1772,N_1705);
nor U1846 (N_1846,N_1736,N_1747);
nand U1847 (N_1847,N_1773,N_1719);
nor U1848 (N_1848,N_1724,N_1727);
or U1849 (N_1849,N_1780,N_1712);
or U1850 (N_1850,N_1689,N_1701);
nand U1851 (N_1851,N_1659,N_1702);
nand U1852 (N_1852,N_1742,N_1668);
or U1853 (N_1853,N_1766,N_1734);
and U1854 (N_1854,N_1797,N_1758);
and U1855 (N_1855,N_1741,N_1787);
xnor U1856 (N_1856,N_1790,N_1723);
and U1857 (N_1857,N_1795,N_1756);
nor U1858 (N_1858,N_1776,N_1793);
nand U1859 (N_1859,N_1739,N_1708);
and U1860 (N_1860,N_1722,N_1673);
nand U1861 (N_1861,N_1753,N_1725);
or U1862 (N_1862,N_1718,N_1740);
or U1863 (N_1863,N_1792,N_1677);
xnor U1864 (N_1864,N_1794,N_1796);
nand U1865 (N_1865,N_1729,N_1675);
and U1866 (N_1866,N_1679,N_1660);
nand U1867 (N_1867,N_1654,N_1791);
nand U1868 (N_1868,N_1671,N_1765);
nand U1869 (N_1869,N_1750,N_1778);
or U1870 (N_1870,N_1783,N_1771);
nand U1871 (N_1871,N_1746,N_1777);
and U1872 (N_1872,N_1653,N_1686);
xor U1873 (N_1873,N_1726,N_1733);
xnor U1874 (N_1874,N_1656,N_1663);
and U1875 (N_1875,N_1785,N_1661);
or U1876 (N_1876,N_1670,N_1660);
xor U1877 (N_1877,N_1774,N_1653);
nand U1878 (N_1878,N_1775,N_1736);
and U1879 (N_1879,N_1775,N_1750);
xnor U1880 (N_1880,N_1792,N_1762);
or U1881 (N_1881,N_1758,N_1693);
or U1882 (N_1882,N_1790,N_1756);
nand U1883 (N_1883,N_1669,N_1660);
and U1884 (N_1884,N_1768,N_1744);
xnor U1885 (N_1885,N_1709,N_1772);
nand U1886 (N_1886,N_1716,N_1733);
nand U1887 (N_1887,N_1701,N_1663);
or U1888 (N_1888,N_1765,N_1790);
and U1889 (N_1889,N_1668,N_1733);
xnor U1890 (N_1890,N_1744,N_1709);
and U1891 (N_1891,N_1797,N_1720);
xor U1892 (N_1892,N_1686,N_1764);
nor U1893 (N_1893,N_1739,N_1721);
or U1894 (N_1894,N_1755,N_1761);
nor U1895 (N_1895,N_1706,N_1738);
or U1896 (N_1896,N_1734,N_1768);
or U1897 (N_1897,N_1751,N_1799);
nor U1898 (N_1898,N_1749,N_1685);
xor U1899 (N_1899,N_1760,N_1667);
or U1900 (N_1900,N_1686,N_1750);
or U1901 (N_1901,N_1706,N_1737);
nand U1902 (N_1902,N_1787,N_1727);
and U1903 (N_1903,N_1708,N_1704);
or U1904 (N_1904,N_1689,N_1729);
and U1905 (N_1905,N_1689,N_1776);
xnor U1906 (N_1906,N_1696,N_1792);
or U1907 (N_1907,N_1711,N_1685);
nand U1908 (N_1908,N_1700,N_1695);
and U1909 (N_1909,N_1706,N_1650);
xnor U1910 (N_1910,N_1708,N_1752);
nor U1911 (N_1911,N_1666,N_1694);
or U1912 (N_1912,N_1732,N_1714);
xor U1913 (N_1913,N_1746,N_1775);
xnor U1914 (N_1914,N_1655,N_1679);
nand U1915 (N_1915,N_1686,N_1700);
nand U1916 (N_1916,N_1757,N_1754);
nand U1917 (N_1917,N_1684,N_1681);
or U1918 (N_1918,N_1798,N_1790);
or U1919 (N_1919,N_1678,N_1675);
and U1920 (N_1920,N_1705,N_1752);
nand U1921 (N_1921,N_1712,N_1681);
nand U1922 (N_1922,N_1784,N_1717);
xnor U1923 (N_1923,N_1796,N_1735);
nand U1924 (N_1924,N_1655,N_1772);
nor U1925 (N_1925,N_1795,N_1650);
or U1926 (N_1926,N_1715,N_1739);
or U1927 (N_1927,N_1695,N_1660);
nor U1928 (N_1928,N_1685,N_1732);
xor U1929 (N_1929,N_1666,N_1659);
and U1930 (N_1930,N_1796,N_1729);
and U1931 (N_1931,N_1735,N_1793);
nand U1932 (N_1932,N_1745,N_1792);
nand U1933 (N_1933,N_1663,N_1672);
nand U1934 (N_1934,N_1690,N_1666);
nor U1935 (N_1935,N_1769,N_1731);
xnor U1936 (N_1936,N_1765,N_1697);
nor U1937 (N_1937,N_1671,N_1676);
nand U1938 (N_1938,N_1791,N_1690);
nor U1939 (N_1939,N_1763,N_1656);
and U1940 (N_1940,N_1668,N_1794);
or U1941 (N_1941,N_1656,N_1714);
nor U1942 (N_1942,N_1736,N_1716);
nor U1943 (N_1943,N_1659,N_1671);
nor U1944 (N_1944,N_1776,N_1748);
xnor U1945 (N_1945,N_1773,N_1792);
or U1946 (N_1946,N_1780,N_1665);
nand U1947 (N_1947,N_1725,N_1711);
nor U1948 (N_1948,N_1750,N_1781);
and U1949 (N_1949,N_1772,N_1725);
nand U1950 (N_1950,N_1853,N_1841);
nand U1951 (N_1951,N_1864,N_1870);
and U1952 (N_1952,N_1839,N_1922);
xnor U1953 (N_1953,N_1923,N_1867);
xor U1954 (N_1954,N_1859,N_1918);
nand U1955 (N_1955,N_1822,N_1944);
nor U1956 (N_1956,N_1818,N_1847);
nand U1957 (N_1957,N_1879,N_1926);
xnor U1958 (N_1958,N_1802,N_1803);
and U1959 (N_1959,N_1825,N_1929);
xor U1960 (N_1960,N_1851,N_1908);
and U1961 (N_1961,N_1895,N_1899);
nand U1962 (N_1962,N_1804,N_1927);
xnor U1963 (N_1963,N_1887,N_1925);
nor U1964 (N_1964,N_1811,N_1857);
or U1965 (N_1965,N_1903,N_1850);
and U1966 (N_1966,N_1801,N_1936);
and U1967 (N_1967,N_1932,N_1844);
xnor U1968 (N_1968,N_1917,N_1894);
and U1969 (N_1969,N_1835,N_1838);
nor U1970 (N_1970,N_1933,N_1840);
nand U1971 (N_1971,N_1860,N_1837);
and U1972 (N_1972,N_1947,N_1884);
nand U1973 (N_1973,N_1872,N_1883);
and U1974 (N_1974,N_1814,N_1821);
nor U1975 (N_1975,N_1916,N_1866);
or U1976 (N_1976,N_1800,N_1858);
nor U1977 (N_1977,N_1827,N_1924);
xnor U1978 (N_1978,N_1831,N_1901);
nand U1979 (N_1979,N_1808,N_1896);
xnor U1980 (N_1980,N_1824,N_1942);
nand U1981 (N_1981,N_1873,N_1910);
nor U1982 (N_1982,N_1941,N_1888);
nand U1983 (N_1983,N_1930,N_1928);
and U1984 (N_1984,N_1919,N_1865);
or U1985 (N_1985,N_1931,N_1855);
nand U1986 (N_1986,N_1875,N_1845);
or U1987 (N_1987,N_1815,N_1921);
or U1988 (N_1988,N_1880,N_1876);
xor U1989 (N_1989,N_1836,N_1809);
or U1990 (N_1990,N_1909,N_1939);
or U1991 (N_1991,N_1823,N_1878);
and U1992 (N_1992,N_1907,N_1849);
nor U1993 (N_1993,N_1877,N_1861);
nor U1994 (N_1994,N_1934,N_1937);
and U1995 (N_1995,N_1885,N_1897);
or U1996 (N_1996,N_1830,N_1900);
or U1997 (N_1997,N_1805,N_1829);
nor U1998 (N_1998,N_1882,N_1946);
or U1999 (N_1999,N_1920,N_1826);
nand U2000 (N_2000,N_1890,N_1945);
and U2001 (N_2001,N_1812,N_1869);
nand U2002 (N_2002,N_1856,N_1886);
and U2003 (N_2003,N_1898,N_1820);
nor U2004 (N_2004,N_1846,N_1843);
xor U2005 (N_2005,N_1911,N_1863);
and U2006 (N_2006,N_1913,N_1943);
xor U2007 (N_2007,N_1832,N_1813);
xnor U2008 (N_2008,N_1938,N_1891);
and U2009 (N_2009,N_1852,N_1806);
nor U2010 (N_2010,N_1819,N_1807);
or U2011 (N_2011,N_1834,N_1828);
nand U2012 (N_2012,N_1868,N_1940);
nor U2013 (N_2013,N_1848,N_1881);
nand U2014 (N_2014,N_1862,N_1889);
nor U2015 (N_2015,N_1810,N_1904);
nor U2016 (N_2016,N_1854,N_1833);
nand U2017 (N_2017,N_1915,N_1905);
xnor U2018 (N_2018,N_1892,N_1817);
or U2019 (N_2019,N_1816,N_1902);
nand U2020 (N_2020,N_1949,N_1874);
nor U2021 (N_2021,N_1893,N_1906);
nor U2022 (N_2022,N_1871,N_1948);
nor U2023 (N_2023,N_1842,N_1912);
nand U2024 (N_2024,N_1935,N_1914);
and U2025 (N_2025,N_1831,N_1820);
and U2026 (N_2026,N_1841,N_1861);
and U2027 (N_2027,N_1803,N_1880);
nand U2028 (N_2028,N_1881,N_1851);
nor U2029 (N_2029,N_1907,N_1933);
nor U2030 (N_2030,N_1903,N_1908);
nor U2031 (N_2031,N_1906,N_1866);
nand U2032 (N_2032,N_1880,N_1889);
nand U2033 (N_2033,N_1944,N_1915);
and U2034 (N_2034,N_1890,N_1850);
or U2035 (N_2035,N_1859,N_1938);
xnor U2036 (N_2036,N_1833,N_1903);
nor U2037 (N_2037,N_1869,N_1935);
or U2038 (N_2038,N_1870,N_1817);
or U2039 (N_2039,N_1814,N_1815);
nor U2040 (N_2040,N_1826,N_1900);
nand U2041 (N_2041,N_1946,N_1825);
or U2042 (N_2042,N_1801,N_1905);
xnor U2043 (N_2043,N_1859,N_1929);
nand U2044 (N_2044,N_1862,N_1802);
and U2045 (N_2045,N_1939,N_1881);
xor U2046 (N_2046,N_1868,N_1900);
or U2047 (N_2047,N_1946,N_1875);
or U2048 (N_2048,N_1928,N_1909);
or U2049 (N_2049,N_1919,N_1838);
nor U2050 (N_2050,N_1857,N_1881);
xnor U2051 (N_2051,N_1810,N_1828);
or U2052 (N_2052,N_1931,N_1812);
or U2053 (N_2053,N_1894,N_1893);
nand U2054 (N_2054,N_1928,N_1853);
nand U2055 (N_2055,N_1887,N_1946);
and U2056 (N_2056,N_1826,N_1848);
xor U2057 (N_2057,N_1911,N_1927);
nand U2058 (N_2058,N_1824,N_1895);
or U2059 (N_2059,N_1913,N_1869);
or U2060 (N_2060,N_1817,N_1857);
xor U2061 (N_2061,N_1910,N_1866);
or U2062 (N_2062,N_1811,N_1898);
nand U2063 (N_2063,N_1920,N_1814);
xnor U2064 (N_2064,N_1857,N_1902);
nand U2065 (N_2065,N_1810,N_1917);
or U2066 (N_2066,N_1846,N_1877);
or U2067 (N_2067,N_1861,N_1837);
and U2068 (N_2068,N_1949,N_1854);
or U2069 (N_2069,N_1830,N_1808);
and U2070 (N_2070,N_1853,N_1846);
or U2071 (N_2071,N_1905,N_1856);
nand U2072 (N_2072,N_1878,N_1837);
and U2073 (N_2073,N_1881,N_1947);
or U2074 (N_2074,N_1863,N_1818);
nand U2075 (N_2075,N_1918,N_1945);
or U2076 (N_2076,N_1925,N_1829);
xor U2077 (N_2077,N_1943,N_1815);
and U2078 (N_2078,N_1818,N_1882);
nand U2079 (N_2079,N_1832,N_1819);
and U2080 (N_2080,N_1917,N_1893);
and U2081 (N_2081,N_1929,N_1900);
or U2082 (N_2082,N_1939,N_1928);
xor U2083 (N_2083,N_1890,N_1915);
nor U2084 (N_2084,N_1948,N_1855);
xor U2085 (N_2085,N_1894,N_1911);
and U2086 (N_2086,N_1930,N_1866);
nor U2087 (N_2087,N_1812,N_1866);
nor U2088 (N_2088,N_1850,N_1808);
or U2089 (N_2089,N_1931,N_1821);
or U2090 (N_2090,N_1948,N_1844);
nand U2091 (N_2091,N_1856,N_1910);
nor U2092 (N_2092,N_1856,N_1812);
or U2093 (N_2093,N_1884,N_1848);
xor U2094 (N_2094,N_1849,N_1930);
nand U2095 (N_2095,N_1825,N_1914);
or U2096 (N_2096,N_1870,N_1854);
or U2097 (N_2097,N_1924,N_1923);
nor U2098 (N_2098,N_1802,N_1916);
xnor U2099 (N_2099,N_1880,N_1828);
and U2100 (N_2100,N_1994,N_2000);
nand U2101 (N_2101,N_1972,N_2095);
or U2102 (N_2102,N_2033,N_2021);
nor U2103 (N_2103,N_2020,N_2097);
or U2104 (N_2104,N_1985,N_2010);
or U2105 (N_2105,N_2098,N_2091);
nor U2106 (N_2106,N_2052,N_1998);
xnor U2107 (N_2107,N_2083,N_2040);
nand U2108 (N_2108,N_2069,N_2049);
nand U2109 (N_2109,N_1959,N_2096);
nor U2110 (N_2110,N_1986,N_2047);
or U2111 (N_2111,N_2067,N_2012);
or U2112 (N_2112,N_2022,N_2023);
and U2113 (N_2113,N_2080,N_1979);
xor U2114 (N_2114,N_1957,N_1955);
or U2115 (N_2115,N_2076,N_2066);
or U2116 (N_2116,N_1964,N_1951);
or U2117 (N_2117,N_2015,N_2082);
or U2118 (N_2118,N_1963,N_2054);
nand U2119 (N_2119,N_2058,N_1976);
nor U2120 (N_2120,N_2072,N_2075);
xor U2121 (N_2121,N_2070,N_2034);
nand U2122 (N_2122,N_1973,N_2053);
xnor U2123 (N_2123,N_1974,N_2043);
nor U2124 (N_2124,N_1961,N_2050);
and U2125 (N_2125,N_2019,N_2088);
and U2126 (N_2126,N_2090,N_2099);
nand U2127 (N_2127,N_2041,N_1960);
nor U2128 (N_2128,N_2078,N_2077);
or U2129 (N_2129,N_1980,N_1990);
and U2130 (N_2130,N_2046,N_2042);
nand U2131 (N_2131,N_1958,N_2079);
or U2132 (N_2132,N_2029,N_1954);
nor U2133 (N_2133,N_2026,N_1962);
xor U2134 (N_2134,N_2051,N_2065);
and U2135 (N_2135,N_2045,N_2039);
xor U2136 (N_2136,N_1978,N_2089);
xnor U2137 (N_2137,N_2009,N_1956);
nand U2138 (N_2138,N_2037,N_1996);
or U2139 (N_2139,N_2087,N_2063);
xnor U2140 (N_2140,N_2017,N_2030);
nand U2141 (N_2141,N_2094,N_2036);
and U2142 (N_2142,N_2024,N_2084);
xnor U2143 (N_2143,N_2048,N_2055);
nand U2144 (N_2144,N_1995,N_1966);
or U2145 (N_2145,N_1982,N_2064);
nand U2146 (N_2146,N_2018,N_2086);
xnor U2147 (N_2147,N_2008,N_2092);
and U2148 (N_2148,N_2073,N_2014);
or U2149 (N_2149,N_2093,N_1971);
nand U2150 (N_2150,N_1987,N_1983);
or U2151 (N_2151,N_2011,N_1988);
nand U2152 (N_2152,N_2005,N_1992);
nand U2153 (N_2153,N_2001,N_1968);
nor U2154 (N_2154,N_1952,N_1989);
and U2155 (N_2155,N_2081,N_2071);
and U2156 (N_2156,N_2013,N_2025);
xnor U2157 (N_2157,N_2074,N_1969);
nor U2158 (N_2158,N_2056,N_2027);
or U2159 (N_2159,N_2003,N_2062);
and U2160 (N_2160,N_2007,N_1999);
or U2161 (N_2161,N_1991,N_1984);
nor U2162 (N_2162,N_2004,N_2032);
xnor U2163 (N_2163,N_1981,N_2068);
and U2164 (N_2164,N_2061,N_2059);
nand U2165 (N_2165,N_1993,N_2057);
nand U2166 (N_2166,N_2016,N_1977);
nand U2167 (N_2167,N_1967,N_1953);
and U2168 (N_2168,N_2060,N_2002);
xor U2169 (N_2169,N_2028,N_2085);
and U2170 (N_2170,N_1997,N_2031);
or U2171 (N_2171,N_2038,N_1975);
or U2172 (N_2172,N_1970,N_2035);
and U2173 (N_2173,N_2044,N_2006);
xor U2174 (N_2174,N_1965,N_1950);
nand U2175 (N_2175,N_2057,N_1979);
nor U2176 (N_2176,N_2053,N_2008);
or U2177 (N_2177,N_1950,N_2050);
nor U2178 (N_2178,N_2067,N_1981);
nor U2179 (N_2179,N_2030,N_2027);
and U2180 (N_2180,N_2080,N_2021);
and U2181 (N_2181,N_2084,N_1962);
nor U2182 (N_2182,N_2064,N_2077);
xor U2183 (N_2183,N_1976,N_2053);
and U2184 (N_2184,N_2007,N_2086);
xor U2185 (N_2185,N_1966,N_2094);
nand U2186 (N_2186,N_2039,N_2030);
xor U2187 (N_2187,N_1959,N_2072);
xnor U2188 (N_2188,N_2019,N_2056);
xor U2189 (N_2189,N_1976,N_2012);
and U2190 (N_2190,N_2048,N_1955);
xor U2191 (N_2191,N_2089,N_2042);
and U2192 (N_2192,N_2006,N_2013);
or U2193 (N_2193,N_2062,N_2065);
xor U2194 (N_2194,N_1983,N_2092);
or U2195 (N_2195,N_2027,N_2061);
nand U2196 (N_2196,N_2063,N_2022);
nand U2197 (N_2197,N_1973,N_2028);
or U2198 (N_2198,N_1995,N_2017);
or U2199 (N_2199,N_2068,N_1970);
nor U2200 (N_2200,N_2039,N_1981);
or U2201 (N_2201,N_2002,N_2061);
or U2202 (N_2202,N_2045,N_1973);
nor U2203 (N_2203,N_2034,N_2020);
nor U2204 (N_2204,N_2026,N_2092);
nor U2205 (N_2205,N_2080,N_1975);
nor U2206 (N_2206,N_2000,N_1998);
and U2207 (N_2207,N_2032,N_2016);
nand U2208 (N_2208,N_2022,N_2098);
nand U2209 (N_2209,N_2085,N_2045);
or U2210 (N_2210,N_2046,N_2055);
xor U2211 (N_2211,N_1964,N_2057);
nand U2212 (N_2212,N_1983,N_1967);
xor U2213 (N_2213,N_2049,N_1985);
and U2214 (N_2214,N_1963,N_1998);
or U2215 (N_2215,N_2004,N_2005);
nor U2216 (N_2216,N_2005,N_2055);
nand U2217 (N_2217,N_2072,N_2017);
nor U2218 (N_2218,N_1951,N_2028);
nand U2219 (N_2219,N_2098,N_1961);
nand U2220 (N_2220,N_1977,N_2075);
nand U2221 (N_2221,N_2007,N_2075);
nor U2222 (N_2222,N_2095,N_2074);
nor U2223 (N_2223,N_2039,N_1953);
xnor U2224 (N_2224,N_2096,N_2071);
and U2225 (N_2225,N_2040,N_1989);
or U2226 (N_2226,N_2032,N_1975);
and U2227 (N_2227,N_2044,N_1971);
xor U2228 (N_2228,N_2031,N_1988);
or U2229 (N_2229,N_2039,N_1963);
xnor U2230 (N_2230,N_1966,N_2059);
nor U2231 (N_2231,N_2066,N_1980);
and U2232 (N_2232,N_2046,N_2096);
nor U2233 (N_2233,N_1954,N_1975);
xnor U2234 (N_2234,N_2054,N_2044);
and U2235 (N_2235,N_2032,N_2027);
nand U2236 (N_2236,N_2034,N_2097);
and U2237 (N_2237,N_2047,N_2050);
nand U2238 (N_2238,N_1975,N_2007);
xnor U2239 (N_2239,N_2075,N_2029);
xor U2240 (N_2240,N_2029,N_2069);
nand U2241 (N_2241,N_2001,N_1973);
and U2242 (N_2242,N_2092,N_2016);
and U2243 (N_2243,N_1963,N_2033);
xor U2244 (N_2244,N_1996,N_1969);
or U2245 (N_2245,N_2032,N_1993);
xor U2246 (N_2246,N_1985,N_2075);
xor U2247 (N_2247,N_2019,N_2087);
or U2248 (N_2248,N_2033,N_2068);
or U2249 (N_2249,N_2037,N_2099);
xor U2250 (N_2250,N_2142,N_2209);
or U2251 (N_2251,N_2163,N_2235);
nor U2252 (N_2252,N_2245,N_2109);
xnor U2253 (N_2253,N_2225,N_2205);
xor U2254 (N_2254,N_2110,N_2137);
and U2255 (N_2255,N_2100,N_2114);
nor U2256 (N_2256,N_2227,N_2189);
xor U2257 (N_2257,N_2155,N_2102);
or U2258 (N_2258,N_2204,N_2150);
nor U2259 (N_2259,N_2238,N_2215);
or U2260 (N_2260,N_2219,N_2246);
and U2261 (N_2261,N_2240,N_2221);
xor U2262 (N_2262,N_2218,N_2122);
nand U2263 (N_2263,N_2113,N_2191);
and U2264 (N_2264,N_2217,N_2171);
nor U2265 (N_2265,N_2186,N_2201);
and U2266 (N_2266,N_2115,N_2117);
or U2267 (N_2267,N_2212,N_2139);
nor U2268 (N_2268,N_2210,N_2168);
nand U2269 (N_2269,N_2241,N_2220);
and U2270 (N_2270,N_2222,N_2148);
nor U2271 (N_2271,N_2161,N_2199);
and U2272 (N_2272,N_2140,N_2124);
and U2273 (N_2273,N_2120,N_2133);
or U2274 (N_2274,N_2123,N_2211);
nor U2275 (N_2275,N_2159,N_2182);
and U2276 (N_2276,N_2118,N_2213);
nand U2277 (N_2277,N_2248,N_2107);
nand U2278 (N_2278,N_2188,N_2242);
or U2279 (N_2279,N_2207,N_2237);
xnor U2280 (N_2280,N_2156,N_2170);
or U2281 (N_2281,N_2190,N_2176);
xnor U2282 (N_2282,N_2145,N_2144);
xnor U2283 (N_2283,N_2138,N_2141);
or U2284 (N_2284,N_2152,N_2174);
and U2285 (N_2285,N_2125,N_2206);
or U2286 (N_2286,N_2194,N_2127);
or U2287 (N_2287,N_2180,N_2214);
nor U2288 (N_2288,N_2160,N_2166);
or U2289 (N_2289,N_2177,N_2126);
and U2290 (N_2290,N_2165,N_2105);
nor U2291 (N_2291,N_2224,N_2169);
and U2292 (N_2292,N_2149,N_2184);
and U2293 (N_2293,N_2193,N_2185);
or U2294 (N_2294,N_2147,N_2173);
nor U2295 (N_2295,N_2249,N_2121);
xnor U2296 (N_2296,N_2231,N_2196);
xnor U2297 (N_2297,N_2197,N_2244);
nand U2298 (N_2298,N_2223,N_2129);
and U2299 (N_2299,N_2132,N_2181);
nor U2300 (N_2300,N_2228,N_2106);
nand U2301 (N_2301,N_2130,N_2172);
or U2302 (N_2302,N_2128,N_2146);
nor U2303 (N_2303,N_2154,N_2153);
or U2304 (N_2304,N_2136,N_2157);
or U2305 (N_2305,N_2103,N_2178);
and U2306 (N_2306,N_2195,N_2175);
nand U2307 (N_2307,N_2101,N_2111);
or U2308 (N_2308,N_2229,N_2208);
or U2309 (N_2309,N_2202,N_2192);
xor U2310 (N_2310,N_2183,N_2230);
or U2311 (N_2311,N_2104,N_2134);
and U2312 (N_2312,N_2216,N_2162);
nor U2313 (N_2313,N_2232,N_2131);
nor U2314 (N_2314,N_2234,N_2243);
nand U2315 (N_2315,N_2151,N_2239);
or U2316 (N_2316,N_2143,N_2187);
and U2317 (N_2317,N_2112,N_2179);
nand U2318 (N_2318,N_2247,N_2158);
and U2319 (N_2319,N_2198,N_2203);
nand U2320 (N_2320,N_2236,N_2116);
xor U2321 (N_2321,N_2119,N_2226);
xor U2322 (N_2322,N_2135,N_2233);
nor U2323 (N_2323,N_2200,N_2167);
or U2324 (N_2324,N_2164,N_2108);
xnor U2325 (N_2325,N_2187,N_2216);
and U2326 (N_2326,N_2249,N_2228);
and U2327 (N_2327,N_2188,N_2141);
and U2328 (N_2328,N_2197,N_2126);
and U2329 (N_2329,N_2168,N_2242);
and U2330 (N_2330,N_2104,N_2167);
nor U2331 (N_2331,N_2120,N_2110);
nand U2332 (N_2332,N_2170,N_2178);
or U2333 (N_2333,N_2190,N_2183);
xor U2334 (N_2334,N_2225,N_2101);
nand U2335 (N_2335,N_2208,N_2216);
xnor U2336 (N_2336,N_2150,N_2118);
nor U2337 (N_2337,N_2165,N_2216);
and U2338 (N_2338,N_2165,N_2134);
nand U2339 (N_2339,N_2241,N_2155);
and U2340 (N_2340,N_2240,N_2214);
nand U2341 (N_2341,N_2111,N_2159);
or U2342 (N_2342,N_2239,N_2124);
and U2343 (N_2343,N_2183,N_2238);
or U2344 (N_2344,N_2219,N_2120);
xnor U2345 (N_2345,N_2186,N_2248);
or U2346 (N_2346,N_2132,N_2102);
nand U2347 (N_2347,N_2137,N_2156);
and U2348 (N_2348,N_2125,N_2224);
nand U2349 (N_2349,N_2213,N_2141);
xor U2350 (N_2350,N_2104,N_2242);
nor U2351 (N_2351,N_2153,N_2115);
and U2352 (N_2352,N_2154,N_2208);
or U2353 (N_2353,N_2225,N_2210);
nand U2354 (N_2354,N_2226,N_2158);
xnor U2355 (N_2355,N_2191,N_2162);
nand U2356 (N_2356,N_2242,N_2161);
nand U2357 (N_2357,N_2176,N_2209);
nand U2358 (N_2358,N_2158,N_2232);
and U2359 (N_2359,N_2115,N_2217);
nand U2360 (N_2360,N_2216,N_2203);
nor U2361 (N_2361,N_2236,N_2192);
and U2362 (N_2362,N_2196,N_2176);
or U2363 (N_2363,N_2128,N_2204);
or U2364 (N_2364,N_2152,N_2121);
and U2365 (N_2365,N_2110,N_2127);
nand U2366 (N_2366,N_2103,N_2197);
or U2367 (N_2367,N_2117,N_2102);
nor U2368 (N_2368,N_2224,N_2153);
and U2369 (N_2369,N_2126,N_2118);
xnor U2370 (N_2370,N_2226,N_2203);
or U2371 (N_2371,N_2204,N_2191);
and U2372 (N_2372,N_2137,N_2136);
or U2373 (N_2373,N_2222,N_2130);
and U2374 (N_2374,N_2118,N_2155);
nand U2375 (N_2375,N_2230,N_2147);
nor U2376 (N_2376,N_2178,N_2208);
or U2377 (N_2377,N_2139,N_2156);
or U2378 (N_2378,N_2199,N_2207);
or U2379 (N_2379,N_2213,N_2131);
xor U2380 (N_2380,N_2182,N_2219);
and U2381 (N_2381,N_2129,N_2228);
or U2382 (N_2382,N_2132,N_2139);
or U2383 (N_2383,N_2202,N_2175);
or U2384 (N_2384,N_2210,N_2230);
nor U2385 (N_2385,N_2165,N_2198);
or U2386 (N_2386,N_2107,N_2212);
or U2387 (N_2387,N_2162,N_2116);
and U2388 (N_2388,N_2209,N_2183);
and U2389 (N_2389,N_2182,N_2165);
and U2390 (N_2390,N_2122,N_2220);
or U2391 (N_2391,N_2196,N_2213);
xnor U2392 (N_2392,N_2219,N_2244);
xnor U2393 (N_2393,N_2220,N_2116);
or U2394 (N_2394,N_2195,N_2210);
nand U2395 (N_2395,N_2177,N_2244);
nand U2396 (N_2396,N_2249,N_2181);
xor U2397 (N_2397,N_2114,N_2199);
and U2398 (N_2398,N_2129,N_2103);
or U2399 (N_2399,N_2243,N_2226);
or U2400 (N_2400,N_2382,N_2338);
and U2401 (N_2401,N_2258,N_2283);
nor U2402 (N_2402,N_2372,N_2345);
xnor U2403 (N_2403,N_2294,N_2321);
or U2404 (N_2404,N_2353,N_2398);
nor U2405 (N_2405,N_2363,N_2328);
and U2406 (N_2406,N_2335,N_2292);
nor U2407 (N_2407,N_2317,N_2354);
or U2408 (N_2408,N_2324,N_2319);
nand U2409 (N_2409,N_2309,N_2323);
and U2410 (N_2410,N_2374,N_2387);
and U2411 (N_2411,N_2355,N_2307);
nand U2412 (N_2412,N_2369,N_2397);
xnor U2413 (N_2413,N_2357,N_2350);
xor U2414 (N_2414,N_2399,N_2266);
and U2415 (N_2415,N_2370,N_2263);
nor U2416 (N_2416,N_2270,N_2305);
or U2417 (N_2417,N_2347,N_2311);
nand U2418 (N_2418,N_2306,N_2389);
xor U2419 (N_2419,N_2272,N_2343);
nor U2420 (N_2420,N_2291,N_2253);
and U2421 (N_2421,N_2348,N_2301);
or U2422 (N_2422,N_2341,N_2379);
nand U2423 (N_2423,N_2349,N_2332);
or U2424 (N_2424,N_2271,N_2286);
and U2425 (N_2425,N_2364,N_2360);
nor U2426 (N_2426,N_2375,N_2386);
nor U2427 (N_2427,N_2388,N_2394);
or U2428 (N_2428,N_2346,N_2279);
xor U2429 (N_2429,N_2289,N_2380);
nand U2430 (N_2430,N_2282,N_2257);
xor U2431 (N_2431,N_2327,N_2390);
xnor U2432 (N_2432,N_2260,N_2318);
xnor U2433 (N_2433,N_2340,N_2320);
xor U2434 (N_2434,N_2269,N_2313);
or U2435 (N_2435,N_2264,N_2250);
nand U2436 (N_2436,N_2381,N_2297);
and U2437 (N_2437,N_2314,N_2310);
xnor U2438 (N_2438,N_2252,N_2367);
nand U2439 (N_2439,N_2396,N_2251);
nand U2440 (N_2440,N_2362,N_2377);
and U2441 (N_2441,N_2392,N_2330);
nor U2442 (N_2442,N_2304,N_2278);
nand U2443 (N_2443,N_2334,N_2322);
and U2444 (N_2444,N_2259,N_2315);
nor U2445 (N_2445,N_2267,N_2261);
xnor U2446 (N_2446,N_2316,N_2290);
nor U2447 (N_2447,N_2277,N_2385);
or U2448 (N_2448,N_2300,N_2276);
nand U2449 (N_2449,N_2352,N_2371);
xor U2450 (N_2450,N_2359,N_2351);
nor U2451 (N_2451,N_2344,N_2395);
and U2452 (N_2452,N_2337,N_2373);
and U2453 (N_2453,N_2384,N_2296);
nor U2454 (N_2454,N_2256,N_2331);
or U2455 (N_2455,N_2299,N_2308);
or U2456 (N_2456,N_2358,N_2287);
nor U2457 (N_2457,N_2339,N_2376);
and U2458 (N_2458,N_2275,N_2333);
or U2459 (N_2459,N_2303,N_2336);
nor U2460 (N_2460,N_2356,N_2295);
nand U2461 (N_2461,N_2293,N_2268);
or U2462 (N_2462,N_2393,N_2273);
nand U2463 (N_2463,N_2281,N_2326);
and U2464 (N_2464,N_2361,N_2284);
nand U2465 (N_2465,N_2366,N_2378);
or U2466 (N_2466,N_2254,N_2265);
xnor U2467 (N_2467,N_2302,N_2383);
nand U2468 (N_2468,N_2342,N_2368);
nor U2469 (N_2469,N_2262,N_2285);
or U2470 (N_2470,N_2312,N_2329);
or U2471 (N_2471,N_2255,N_2365);
nand U2472 (N_2472,N_2298,N_2325);
xor U2473 (N_2473,N_2280,N_2274);
nand U2474 (N_2474,N_2391,N_2288);
xor U2475 (N_2475,N_2345,N_2261);
nor U2476 (N_2476,N_2390,N_2347);
and U2477 (N_2477,N_2350,N_2334);
xor U2478 (N_2478,N_2370,N_2375);
or U2479 (N_2479,N_2258,N_2291);
nor U2480 (N_2480,N_2309,N_2307);
nand U2481 (N_2481,N_2358,N_2375);
or U2482 (N_2482,N_2308,N_2320);
xnor U2483 (N_2483,N_2341,N_2396);
xnor U2484 (N_2484,N_2278,N_2293);
or U2485 (N_2485,N_2329,N_2354);
or U2486 (N_2486,N_2391,N_2254);
xnor U2487 (N_2487,N_2368,N_2353);
nor U2488 (N_2488,N_2371,N_2350);
nor U2489 (N_2489,N_2264,N_2321);
nand U2490 (N_2490,N_2356,N_2370);
nand U2491 (N_2491,N_2307,N_2252);
nor U2492 (N_2492,N_2388,N_2303);
nor U2493 (N_2493,N_2370,N_2270);
xor U2494 (N_2494,N_2398,N_2344);
nor U2495 (N_2495,N_2262,N_2251);
nand U2496 (N_2496,N_2369,N_2254);
xnor U2497 (N_2497,N_2386,N_2344);
xor U2498 (N_2498,N_2351,N_2365);
or U2499 (N_2499,N_2280,N_2256);
nand U2500 (N_2500,N_2296,N_2347);
nor U2501 (N_2501,N_2256,N_2335);
nor U2502 (N_2502,N_2295,N_2349);
nor U2503 (N_2503,N_2383,N_2252);
and U2504 (N_2504,N_2360,N_2317);
xnor U2505 (N_2505,N_2364,N_2367);
nand U2506 (N_2506,N_2307,N_2358);
and U2507 (N_2507,N_2255,N_2278);
or U2508 (N_2508,N_2278,N_2303);
xor U2509 (N_2509,N_2396,N_2331);
and U2510 (N_2510,N_2346,N_2285);
nor U2511 (N_2511,N_2383,N_2258);
xor U2512 (N_2512,N_2340,N_2328);
and U2513 (N_2513,N_2398,N_2393);
xor U2514 (N_2514,N_2252,N_2302);
nand U2515 (N_2515,N_2261,N_2316);
or U2516 (N_2516,N_2284,N_2309);
nand U2517 (N_2517,N_2283,N_2278);
xor U2518 (N_2518,N_2306,N_2262);
and U2519 (N_2519,N_2378,N_2390);
nand U2520 (N_2520,N_2357,N_2312);
or U2521 (N_2521,N_2377,N_2278);
and U2522 (N_2522,N_2287,N_2393);
nand U2523 (N_2523,N_2390,N_2279);
nand U2524 (N_2524,N_2273,N_2299);
nor U2525 (N_2525,N_2342,N_2357);
nor U2526 (N_2526,N_2389,N_2330);
and U2527 (N_2527,N_2294,N_2275);
and U2528 (N_2528,N_2303,N_2391);
xor U2529 (N_2529,N_2369,N_2388);
xnor U2530 (N_2530,N_2290,N_2327);
nor U2531 (N_2531,N_2279,N_2333);
nor U2532 (N_2532,N_2317,N_2397);
xnor U2533 (N_2533,N_2342,N_2352);
xnor U2534 (N_2534,N_2351,N_2386);
or U2535 (N_2535,N_2393,N_2336);
xnor U2536 (N_2536,N_2278,N_2272);
nand U2537 (N_2537,N_2312,N_2386);
or U2538 (N_2538,N_2334,N_2254);
xnor U2539 (N_2539,N_2302,N_2309);
nor U2540 (N_2540,N_2347,N_2303);
nor U2541 (N_2541,N_2311,N_2350);
xnor U2542 (N_2542,N_2268,N_2264);
nor U2543 (N_2543,N_2271,N_2340);
nand U2544 (N_2544,N_2286,N_2299);
nand U2545 (N_2545,N_2395,N_2307);
nor U2546 (N_2546,N_2388,N_2257);
xor U2547 (N_2547,N_2329,N_2372);
nor U2548 (N_2548,N_2316,N_2287);
and U2549 (N_2549,N_2359,N_2272);
or U2550 (N_2550,N_2440,N_2417);
xnor U2551 (N_2551,N_2428,N_2531);
xor U2552 (N_2552,N_2473,N_2480);
and U2553 (N_2553,N_2513,N_2502);
nand U2554 (N_2554,N_2519,N_2477);
or U2555 (N_2555,N_2435,N_2405);
xnor U2556 (N_2556,N_2530,N_2474);
or U2557 (N_2557,N_2490,N_2411);
nand U2558 (N_2558,N_2541,N_2401);
nand U2559 (N_2559,N_2511,N_2548);
xnor U2560 (N_2560,N_2488,N_2445);
xor U2561 (N_2561,N_2497,N_2518);
nor U2562 (N_2562,N_2520,N_2450);
and U2563 (N_2563,N_2458,N_2400);
nor U2564 (N_2564,N_2459,N_2508);
nor U2565 (N_2565,N_2426,N_2489);
nor U2566 (N_2566,N_2464,N_2412);
nor U2567 (N_2567,N_2466,N_2500);
or U2568 (N_2568,N_2421,N_2413);
xor U2569 (N_2569,N_2462,N_2454);
nor U2570 (N_2570,N_2478,N_2501);
or U2571 (N_2571,N_2402,N_2455);
or U2572 (N_2572,N_2496,N_2485);
xor U2573 (N_2573,N_2409,N_2408);
and U2574 (N_2574,N_2546,N_2457);
xnor U2575 (N_2575,N_2536,N_2449);
and U2576 (N_2576,N_2505,N_2448);
or U2577 (N_2577,N_2540,N_2470);
xnor U2578 (N_2578,N_2429,N_2506);
nor U2579 (N_2579,N_2507,N_2503);
or U2580 (N_2580,N_2446,N_2468);
or U2581 (N_2581,N_2492,N_2515);
nand U2582 (N_2582,N_2529,N_2441);
nor U2583 (N_2583,N_2483,N_2527);
xnor U2584 (N_2584,N_2499,N_2542);
nor U2585 (N_2585,N_2410,N_2533);
xnor U2586 (N_2586,N_2420,N_2442);
or U2587 (N_2587,N_2471,N_2437);
or U2588 (N_2588,N_2418,N_2423);
xor U2589 (N_2589,N_2432,N_2427);
nor U2590 (N_2590,N_2539,N_2495);
xor U2591 (N_2591,N_2460,N_2472);
xnor U2592 (N_2592,N_2434,N_2514);
nand U2593 (N_2593,N_2491,N_2532);
nor U2594 (N_2594,N_2461,N_2486);
nor U2595 (N_2595,N_2481,N_2526);
nand U2596 (N_2596,N_2498,N_2444);
xnor U2597 (N_2597,N_2535,N_2494);
nand U2598 (N_2598,N_2537,N_2517);
or U2599 (N_2599,N_2509,N_2414);
nand U2600 (N_2600,N_2504,N_2538);
nand U2601 (N_2601,N_2528,N_2419);
or U2602 (N_2602,N_2453,N_2443);
and U2603 (N_2603,N_2525,N_2415);
and U2604 (N_2604,N_2524,N_2467);
xnor U2605 (N_2605,N_2424,N_2451);
nor U2606 (N_2606,N_2456,N_2493);
nand U2607 (N_2607,N_2487,N_2463);
or U2608 (N_2608,N_2522,N_2403);
xor U2609 (N_2609,N_2447,N_2484);
nor U2610 (N_2610,N_2476,N_2545);
or U2611 (N_2611,N_2475,N_2543);
and U2612 (N_2612,N_2547,N_2406);
xor U2613 (N_2613,N_2510,N_2416);
and U2614 (N_2614,N_2512,N_2479);
nor U2615 (N_2615,N_2404,N_2436);
or U2616 (N_2616,N_2425,N_2438);
nor U2617 (N_2617,N_2549,N_2469);
nor U2618 (N_2618,N_2452,N_2407);
nand U2619 (N_2619,N_2430,N_2482);
nand U2620 (N_2620,N_2523,N_2431);
xor U2621 (N_2621,N_2465,N_2433);
nor U2622 (N_2622,N_2516,N_2521);
xnor U2623 (N_2623,N_2534,N_2422);
or U2624 (N_2624,N_2544,N_2439);
or U2625 (N_2625,N_2437,N_2498);
nor U2626 (N_2626,N_2446,N_2445);
nand U2627 (N_2627,N_2485,N_2503);
nand U2628 (N_2628,N_2457,N_2431);
or U2629 (N_2629,N_2475,N_2412);
nand U2630 (N_2630,N_2537,N_2539);
nor U2631 (N_2631,N_2412,N_2409);
or U2632 (N_2632,N_2504,N_2420);
and U2633 (N_2633,N_2447,N_2419);
nor U2634 (N_2634,N_2445,N_2476);
nor U2635 (N_2635,N_2456,N_2548);
xnor U2636 (N_2636,N_2544,N_2407);
and U2637 (N_2637,N_2534,N_2495);
or U2638 (N_2638,N_2488,N_2437);
xor U2639 (N_2639,N_2405,N_2433);
and U2640 (N_2640,N_2494,N_2407);
nor U2641 (N_2641,N_2512,N_2405);
and U2642 (N_2642,N_2519,N_2548);
nand U2643 (N_2643,N_2405,N_2495);
xnor U2644 (N_2644,N_2402,N_2451);
nor U2645 (N_2645,N_2472,N_2424);
nor U2646 (N_2646,N_2523,N_2400);
nor U2647 (N_2647,N_2481,N_2468);
nor U2648 (N_2648,N_2462,N_2492);
nor U2649 (N_2649,N_2426,N_2524);
xor U2650 (N_2650,N_2475,N_2496);
nor U2651 (N_2651,N_2459,N_2436);
and U2652 (N_2652,N_2516,N_2402);
nor U2653 (N_2653,N_2437,N_2532);
or U2654 (N_2654,N_2522,N_2408);
xor U2655 (N_2655,N_2416,N_2432);
xnor U2656 (N_2656,N_2429,N_2498);
nand U2657 (N_2657,N_2542,N_2432);
or U2658 (N_2658,N_2537,N_2521);
or U2659 (N_2659,N_2442,N_2419);
nor U2660 (N_2660,N_2420,N_2401);
nor U2661 (N_2661,N_2408,N_2476);
or U2662 (N_2662,N_2444,N_2428);
and U2663 (N_2663,N_2468,N_2474);
and U2664 (N_2664,N_2495,N_2436);
xnor U2665 (N_2665,N_2473,N_2410);
nor U2666 (N_2666,N_2460,N_2538);
xor U2667 (N_2667,N_2466,N_2455);
and U2668 (N_2668,N_2480,N_2426);
nor U2669 (N_2669,N_2521,N_2468);
and U2670 (N_2670,N_2429,N_2471);
and U2671 (N_2671,N_2401,N_2514);
xor U2672 (N_2672,N_2522,N_2532);
nand U2673 (N_2673,N_2506,N_2410);
nand U2674 (N_2674,N_2541,N_2438);
nand U2675 (N_2675,N_2455,N_2476);
nor U2676 (N_2676,N_2546,N_2504);
or U2677 (N_2677,N_2435,N_2508);
or U2678 (N_2678,N_2507,N_2492);
xnor U2679 (N_2679,N_2462,N_2458);
or U2680 (N_2680,N_2510,N_2445);
or U2681 (N_2681,N_2402,N_2498);
nand U2682 (N_2682,N_2505,N_2508);
or U2683 (N_2683,N_2466,N_2405);
or U2684 (N_2684,N_2542,N_2486);
xor U2685 (N_2685,N_2515,N_2527);
nand U2686 (N_2686,N_2509,N_2412);
xor U2687 (N_2687,N_2545,N_2506);
nor U2688 (N_2688,N_2480,N_2483);
nor U2689 (N_2689,N_2449,N_2542);
nor U2690 (N_2690,N_2476,N_2493);
xor U2691 (N_2691,N_2514,N_2420);
and U2692 (N_2692,N_2421,N_2477);
nand U2693 (N_2693,N_2506,N_2521);
xnor U2694 (N_2694,N_2500,N_2406);
and U2695 (N_2695,N_2421,N_2521);
or U2696 (N_2696,N_2493,N_2415);
and U2697 (N_2697,N_2504,N_2527);
nor U2698 (N_2698,N_2403,N_2459);
xor U2699 (N_2699,N_2410,N_2420);
or U2700 (N_2700,N_2589,N_2691);
nor U2701 (N_2701,N_2654,N_2588);
xnor U2702 (N_2702,N_2605,N_2582);
nand U2703 (N_2703,N_2623,N_2697);
xor U2704 (N_2704,N_2610,N_2650);
or U2705 (N_2705,N_2642,N_2659);
nand U2706 (N_2706,N_2552,N_2651);
and U2707 (N_2707,N_2551,N_2685);
or U2708 (N_2708,N_2615,N_2566);
or U2709 (N_2709,N_2684,N_2689);
nand U2710 (N_2710,N_2692,N_2641);
and U2711 (N_2711,N_2661,N_2595);
xor U2712 (N_2712,N_2632,N_2590);
nor U2713 (N_2713,N_2672,N_2694);
nand U2714 (N_2714,N_2603,N_2594);
nor U2715 (N_2715,N_2587,N_2624);
xnor U2716 (N_2716,N_2679,N_2686);
nand U2717 (N_2717,N_2565,N_2557);
and U2718 (N_2718,N_2674,N_2563);
xnor U2719 (N_2719,N_2574,N_2673);
nor U2720 (N_2720,N_2611,N_2639);
nor U2721 (N_2721,N_2585,N_2607);
or U2722 (N_2722,N_2627,N_2688);
nor U2723 (N_2723,N_2634,N_2567);
xor U2724 (N_2724,N_2561,N_2581);
xnor U2725 (N_2725,N_2586,N_2649);
or U2726 (N_2726,N_2617,N_2671);
and U2727 (N_2727,N_2643,N_2677);
or U2728 (N_2728,N_2662,N_2644);
nor U2729 (N_2729,N_2690,N_2621);
nand U2730 (N_2730,N_2646,N_2696);
or U2731 (N_2731,N_2616,N_2628);
xor U2732 (N_2732,N_2687,N_2608);
and U2733 (N_2733,N_2602,N_2613);
xor U2734 (N_2734,N_2657,N_2699);
and U2735 (N_2735,N_2667,N_2606);
and U2736 (N_2736,N_2592,N_2575);
xnor U2737 (N_2737,N_2560,N_2577);
and U2738 (N_2738,N_2609,N_2598);
nor U2739 (N_2739,N_2618,N_2625);
xor U2740 (N_2740,N_2555,N_2670);
nand U2741 (N_2741,N_2622,N_2568);
nand U2742 (N_2742,N_2562,N_2573);
and U2743 (N_2743,N_2579,N_2583);
xnor U2744 (N_2744,N_2675,N_2635);
or U2745 (N_2745,N_2653,N_2601);
nor U2746 (N_2746,N_2648,N_2682);
nor U2747 (N_2747,N_2663,N_2550);
and U2748 (N_2748,N_2576,N_2619);
nand U2749 (N_2749,N_2620,N_2669);
nor U2750 (N_2750,N_2570,N_2580);
nand U2751 (N_2751,N_2678,N_2631);
and U2752 (N_2752,N_2665,N_2559);
xnor U2753 (N_2753,N_2614,N_2666);
or U2754 (N_2754,N_2600,N_2640);
or U2755 (N_2755,N_2558,N_2599);
xnor U2756 (N_2756,N_2593,N_2604);
and U2757 (N_2757,N_2578,N_2569);
or U2758 (N_2758,N_2683,N_2668);
nor U2759 (N_2759,N_2591,N_2658);
nand U2760 (N_2760,N_2571,N_2680);
nor U2761 (N_2761,N_2584,N_2693);
and U2762 (N_2762,N_2556,N_2695);
and U2763 (N_2763,N_2664,N_2681);
nand U2764 (N_2764,N_2630,N_2645);
or U2765 (N_2765,N_2655,N_2638);
nor U2766 (N_2766,N_2596,N_2647);
nor U2767 (N_2767,N_2572,N_2564);
xnor U2768 (N_2768,N_2676,N_2553);
or U2769 (N_2769,N_2636,N_2660);
nor U2770 (N_2770,N_2637,N_2554);
nand U2771 (N_2771,N_2626,N_2612);
and U2772 (N_2772,N_2633,N_2652);
nand U2773 (N_2773,N_2597,N_2656);
nand U2774 (N_2774,N_2698,N_2629);
and U2775 (N_2775,N_2695,N_2630);
or U2776 (N_2776,N_2563,N_2557);
xor U2777 (N_2777,N_2688,N_2683);
or U2778 (N_2778,N_2658,N_2575);
nand U2779 (N_2779,N_2582,N_2621);
and U2780 (N_2780,N_2583,N_2668);
and U2781 (N_2781,N_2582,N_2687);
and U2782 (N_2782,N_2669,N_2654);
xnor U2783 (N_2783,N_2641,N_2646);
nor U2784 (N_2784,N_2632,N_2674);
and U2785 (N_2785,N_2576,N_2627);
nor U2786 (N_2786,N_2671,N_2580);
nor U2787 (N_2787,N_2664,N_2606);
nand U2788 (N_2788,N_2622,N_2612);
or U2789 (N_2789,N_2628,N_2675);
or U2790 (N_2790,N_2584,N_2566);
nor U2791 (N_2791,N_2615,N_2605);
xor U2792 (N_2792,N_2688,N_2634);
nor U2793 (N_2793,N_2685,N_2683);
nor U2794 (N_2794,N_2597,N_2689);
nor U2795 (N_2795,N_2576,N_2697);
and U2796 (N_2796,N_2692,N_2604);
nand U2797 (N_2797,N_2647,N_2643);
nand U2798 (N_2798,N_2626,N_2688);
nor U2799 (N_2799,N_2550,N_2677);
and U2800 (N_2800,N_2589,N_2683);
nor U2801 (N_2801,N_2648,N_2693);
xnor U2802 (N_2802,N_2587,N_2670);
or U2803 (N_2803,N_2687,N_2600);
or U2804 (N_2804,N_2646,N_2642);
nor U2805 (N_2805,N_2559,N_2565);
nand U2806 (N_2806,N_2582,N_2644);
and U2807 (N_2807,N_2648,N_2645);
xor U2808 (N_2808,N_2609,N_2676);
nor U2809 (N_2809,N_2633,N_2602);
xnor U2810 (N_2810,N_2647,N_2598);
nand U2811 (N_2811,N_2660,N_2681);
and U2812 (N_2812,N_2588,N_2666);
or U2813 (N_2813,N_2640,N_2594);
and U2814 (N_2814,N_2633,N_2670);
xor U2815 (N_2815,N_2573,N_2588);
xor U2816 (N_2816,N_2565,N_2632);
or U2817 (N_2817,N_2556,N_2674);
xnor U2818 (N_2818,N_2680,N_2575);
nor U2819 (N_2819,N_2605,N_2603);
xor U2820 (N_2820,N_2583,N_2689);
or U2821 (N_2821,N_2598,N_2664);
and U2822 (N_2822,N_2695,N_2552);
and U2823 (N_2823,N_2606,N_2615);
nor U2824 (N_2824,N_2661,N_2690);
and U2825 (N_2825,N_2636,N_2630);
nor U2826 (N_2826,N_2593,N_2632);
nand U2827 (N_2827,N_2694,N_2681);
xnor U2828 (N_2828,N_2663,N_2682);
nand U2829 (N_2829,N_2601,N_2627);
and U2830 (N_2830,N_2675,N_2643);
nand U2831 (N_2831,N_2666,N_2580);
and U2832 (N_2832,N_2679,N_2656);
xnor U2833 (N_2833,N_2588,N_2641);
and U2834 (N_2834,N_2567,N_2646);
nor U2835 (N_2835,N_2599,N_2560);
nand U2836 (N_2836,N_2677,N_2645);
and U2837 (N_2837,N_2591,N_2668);
nand U2838 (N_2838,N_2592,N_2683);
and U2839 (N_2839,N_2558,N_2650);
and U2840 (N_2840,N_2596,N_2573);
xnor U2841 (N_2841,N_2555,N_2658);
or U2842 (N_2842,N_2692,N_2630);
nand U2843 (N_2843,N_2588,N_2590);
nor U2844 (N_2844,N_2683,N_2557);
nand U2845 (N_2845,N_2562,N_2656);
nor U2846 (N_2846,N_2607,N_2697);
xnor U2847 (N_2847,N_2586,N_2553);
or U2848 (N_2848,N_2674,N_2594);
xor U2849 (N_2849,N_2596,N_2604);
nor U2850 (N_2850,N_2805,N_2789);
nand U2851 (N_2851,N_2720,N_2717);
and U2852 (N_2852,N_2806,N_2816);
nor U2853 (N_2853,N_2706,N_2821);
and U2854 (N_2854,N_2739,N_2709);
xnor U2855 (N_2855,N_2741,N_2820);
or U2856 (N_2856,N_2701,N_2813);
nand U2857 (N_2857,N_2800,N_2780);
and U2858 (N_2858,N_2770,N_2817);
or U2859 (N_2859,N_2704,N_2771);
nand U2860 (N_2860,N_2823,N_2812);
nor U2861 (N_2861,N_2788,N_2839);
nand U2862 (N_2862,N_2749,N_2798);
nor U2863 (N_2863,N_2743,N_2795);
or U2864 (N_2864,N_2724,N_2803);
nand U2865 (N_2865,N_2822,N_2744);
xnor U2866 (N_2866,N_2828,N_2792);
or U2867 (N_2867,N_2730,N_2760);
xor U2868 (N_2868,N_2835,N_2745);
nor U2869 (N_2869,N_2759,N_2725);
and U2870 (N_2870,N_2752,N_2735);
nand U2871 (N_2871,N_2818,N_2787);
nor U2872 (N_2872,N_2718,N_2836);
nor U2873 (N_2873,N_2733,N_2826);
or U2874 (N_2874,N_2833,N_2830);
xnor U2875 (N_2875,N_2815,N_2838);
nand U2876 (N_2876,N_2746,N_2827);
or U2877 (N_2877,N_2794,N_2785);
xnor U2878 (N_2878,N_2843,N_2753);
nor U2879 (N_2879,N_2762,N_2778);
or U2880 (N_2880,N_2768,N_2802);
xnor U2881 (N_2881,N_2846,N_2707);
xor U2882 (N_2882,N_2807,N_2829);
nand U2883 (N_2883,N_2755,N_2845);
or U2884 (N_2884,N_2713,N_2723);
nor U2885 (N_2885,N_2775,N_2777);
nor U2886 (N_2886,N_2734,N_2710);
nor U2887 (N_2887,N_2705,N_2757);
nand U2888 (N_2888,N_2832,N_2728);
nand U2889 (N_2889,N_2703,N_2783);
and U2890 (N_2890,N_2808,N_2831);
nand U2891 (N_2891,N_2779,N_2714);
or U2892 (N_2892,N_2736,N_2726);
and U2893 (N_2893,N_2716,N_2715);
nand U2894 (N_2894,N_2748,N_2756);
or U2895 (N_2895,N_2847,N_2731);
or U2896 (N_2896,N_2804,N_2840);
nor U2897 (N_2897,N_2742,N_2786);
or U2898 (N_2898,N_2799,N_2782);
or U2899 (N_2899,N_2824,N_2784);
nor U2900 (N_2900,N_2767,N_2721);
or U2901 (N_2901,N_2740,N_2732);
nor U2902 (N_2902,N_2814,N_2758);
xnor U2903 (N_2903,N_2766,N_2722);
or U2904 (N_2904,N_2708,N_2750);
xor U2905 (N_2905,N_2810,N_2776);
xor U2906 (N_2906,N_2712,N_2774);
nand U2907 (N_2907,N_2773,N_2790);
and U2908 (N_2908,N_2781,N_2765);
nor U2909 (N_2909,N_2737,N_2834);
nand U2910 (N_2910,N_2702,N_2738);
nand U2911 (N_2911,N_2841,N_2769);
xor U2912 (N_2912,N_2729,N_2825);
xnor U2913 (N_2913,N_2791,N_2849);
xor U2914 (N_2914,N_2811,N_2819);
or U2915 (N_2915,N_2809,N_2754);
nor U2916 (N_2916,N_2764,N_2751);
and U2917 (N_2917,N_2842,N_2747);
and U2918 (N_2918,N_2727,N_2711);
and U2919 (N_2919,N_2796,N_2844);
nand U2920 (N_2920,N_2797,N_2837);
or U2921 (N_2921,N_2848,N_2801);
nand U2922 (N_2922,N_2772,N_2719);
or U2923 (N_2923,N_2700,N_2793);
nor U2924 (N_2924,N_2763,N_2761);
or U2925 (N_2925,N_2762,N_2727);
or U2926 (N_2926,N_2766,N_2822);
nor U2927 (N_2927,N_2818,N_2812);
xor U2928 (N_2928,N_2828,N_2830);
or U2929 (N_2929,N_2769,N_2768);
xor U2930 (N_2930,N_2813,N_2783);
or U2931 (N_2931,N_2729,N_2730);
nand U2932 (N_2932,N_2769,N_2711);
xor U2933 (N_2933,N_2763,N_2725);
nor U2934 (N_2934,N_2823,N_2837);
nand U2935 (N_2935,N_2799,N_2795);
or U2936 (N_2936,N_2721,N_2832);
or U2937 (N_2937,N_2836,N_2760);
xor U2938 (N_2938,N_2736,N_2717);
or U2939 (N_2939,N_2770,N_2785);
xnor U2940 (N_2940,N_2827,N_2841);
and U2941 (N_2941,N_2700,N_2727);
nand U2942 (N_2942,N_2779,N_2797);
nand U2943 (N_2943,N_2808,N_2736);
xnor U2944 (N_2944,N_2798,N_2716);
or U2945 (N_2945,N_2807,N_2810);
xnor U2946 (N_2946,N_2762,N_2827);
or U2947 (N_2947,N_2711,N_2786);
nand U2948 (N_2948,N_2790,N_2706);
nor U2949 (N_2949,N_2843,N_2706);
or U2950 (N_2950,N_2738,N_2818);
nor U2951 (N_2951,N_2724,N_2845);
and U2952 (N_2952,N_2846,N_2780);
or U2953 (N_2953,N_2712,N_2763);
nand U2954 (N_2954,N_2764,N_2722);
and U2955 (N_2955,N_2755,N_2821);
xnor U2956 (N_2956,N_2819,N_2846);
nand U2957 (N_2957,N_2822,N_2792);
nor U2958 (N_2958,N_2768,N_2829);
nor U2959 (N_2959,N_2798,N_2755);
or U2960 (N_2960,N_2817,N_2799);
xor U2961 (N_2961,N_2847,N_2730);
nand U2962 (N_2962,N_2829,N_2719);
xor U2963 (N_2963,N_2756,N_2774);
or U2964 (N_2964,N_2833,N_2825);
nand U2965 (N_2965,N_2766,N_2763);
and U2966 (N_2966,N_2840,N_2715);
nor U2967 (N_2967,N_2771,N_2700);
and U2968 (N_2968,N_2839,N_2786);
xnor U2969 (N_2969,N_2812,N_2710);
and U2970 (N_2970,N_2722,N_2825);
or U2971 (N_2971,N_2775,N_2772);
or U2972 (N_2972,N_2714,N_2848);
and U2973 (N_2973,N_2811,N_2773);
nand U2974 (N_2974,N_2745,N_2810);
xor U2975 (N_2975,N_2728,N_2727);
nand U2976 (N_2976,N_2842,N_2838);
nand U2977 (N_2977,N_2846,N_2747);
xor U2978 (N_2978,N_2752,N_2741);
nand U2979 (N_2979,N_2719,N_2760);
or U2980 (N_2980,N_2831,N_2726);
and U2981 (N_2981,N_2816,N_2812);
nand U2982 (N_2982,N_2748,N_2808);
or U2983 (N_2983,N_2811,N_2793);
and U2984 (N_2984,N_2822,N_2745);
nor U2985 (N_2985,N_2752,N_2705);
and U2986 (N_2986,N_2812,N_2761);
nor U2987 (N_2987,N_2804,N_2736);
and U2988 (N_2988,N_2808,N_2762);
nand U2989 (N_2989,N_2806,N_2823);
xnor U2990 (N_2990,N_2794,N_2831);
nor U2991 (N_2991,N_2836,N_2813);
xnor U2992 (N_2992,N_2811,N_2705);
nor U2993 (N_2993,N_2806,N_2796);
nand U2994 (N_2994,N_2804,N_2818);
nor U2995 (N_2995,N_2784,N_2740);
nor U2996 (N_2996,N_2830,N_2835);
or U2997 (N_2997,N_2808,N_2843);
xor U2998 (N_2998,N_2847,N_2708);
xnor U2999 (N_2999,N_2739,N_2716);
nand U3000 (N_3000,N_2917,N_2903);
or U3001 (N_3001,N_2996,N_2891);
or U3002 (N_3002,N_2877,N_2956);
xor U3003 (N_3003,N_2972,N_2985);
and U3004 (N_3004,N_2942,N_2995);
xor U3005 (N_3005,N_2987,N_2909);
nand U3006 (N_3006,N_2912,N_2889);
or U3007 (N_3007,N_2928,N_2870);
and U3008 (N_3008,N_2976,N_2873);
xnor U3009 (N_3009,N_2872,N_2855);
xor U3010 (N_3010,N_2931,N_2863);
xnor U3011 (N_3011,N_2967,N_2990);
or U3012 (N_3012,N_2975,N_2902);
nor U3013 (N_3013,N_2953,N_2957);
nor U3014 (N_3014,N_2858,N_2851);
nand U3015 (N_3015,N_2929,N_2868);
and U3016 (N_3016,N_2983,N_2946);
nor U3017 (N_3017,N_2859,N_2883);
nor U3018 (N_3018,N_2874,N_2962);
and U3019 (N_3019,N_2963,N_2960);
or U3020 (N_3020,N_2939,N_2910);
nor U3021 (N_3021,N_2966,N_2887);
nand U3022 (N_3022,N_2897,N_2854);
or U3023 (N_3023,N_2906,N_2894);
nor U3024 (N_3024,N_2864,N_2878);
or U3025 (N_3025,N_2869,N_2895);
and U3026 (N_3026,N_2850,N_2943);
xor U3027 (N_3027,N_2970,N_2892);
nor U3028 (N_3028,N_2980,N_2937);
or U3029 (N_3029,N_2914,N_2905);
nor U3030 (N_3030,N_2927,N_2979);
or U3031 (N_3031,N_2893,N_2884);
and U3032 (N_3032,N_2926,N_2938);
nand U3033 (N_3033,N_2875,N_2933);
xnor U3034 (N_3034,N_2923,N_2853);
nor U3035 (N_3035,N_2948,N_2860);
and U3036 (N_3036,N_2977,N_2913);
and U3037 (N_3037,N_2919,N_2881);
xnor U3038 (N_3038,N_2888,N_2935);
or U3039 (N_3039,N_2974,N_2982);
nand U3040 (N_3040,N_2994,N_2900);
nor U3041 (N_3041,N_2852,N_2920);
xnor U3042 (N_3042,N_2922,N_2961);
nand U3043 (N_3043,N_2880,N_2867);
and U3044 (N_3044,N_2936,N_2934);
nand U3045 (N_3045,N_2932,N_2861);
xnor U3046 (N_3046,N_2959,N_2930);
and U3047 (N_3047,N_2899,N_2908);
xor U3048 (N_3048,N_2945,N_2882);
and U3049 (N_3049,N_2898,N_2964);
xnor U3050 (N_3050,N_2981,N_2879);
xor U3051 (N_3051,N_2968,N_2904);
nor U3052 (N_3052,N_2997,N_2896);
and U3053 (N_3053,N_2885,N_2984);
and U3054 (N_3054,N_2973,N_2925);
and U3055 (N_3055,N_2971,N_2940);
nor U3056 (N_3056,N_2958,N_2991);
xor U3057 (N_3057,N_2865,N_2857);
or U3058 (N_3058,N_2993,N_2969);
and U3059 (N_3059,N_2921,N_2954);
nand U3060 (N_3060,N_2871,N_2944);
xnor U3061 (N_3061,N_2949,N_2916);
and U3062 (N_3062,N_2915,N_2911);
nand U3063 (N_3063,N_2862,N_2992);
nand U3064 (N_3064,N_2978,N_2856);
and U3065 (N_3065,N_2965,N_2866);
nor U3066 (N_3066,N_2989,N_2988);
nand U3067 (N_3067,N_2950,N_2901);
nand U3068 (N_3068,N_2876,N_2890);
or U3069 (N_3069,N_2955,N_2947);
or U3070 (N_3070,N_2998,N_2907);
nor U3071 (N_3071,N_2918,N_2951);
and U3072 (N_3072,N_2924,N_2886);
and U3073 (N_3073,N_2952,N_2941);
and U3074 (N_3074,N_2986,N_2999);
and U3075 (N_3075,N_2895,N_2997);
nand U3076 (N_3076,N_2942,N_2899);
xor U3077 (N_3077,N_2914,N_2938);
xnor U3078 (N_3078,N_2939,N_2880);
nor U3079 (N_3079,N_2917,N_2991);
nand U3080 (N_3080,N_2902,N_2922);
nand U3081 (N_3081,N_2948,N_2880);
nor U3082 (N_3082,N_2941,N_2901);
nand U3083 (N_3083,N_2941,N_2972);
nor U3084 (N_3084,N_2866,N_2959);
nor U3085 (N_3085,N_2929,N_2903);
nand U3086 (N_3086,N_2900,N_2852);
nor U3087 (N_3087,N_2983,N_2854);
xor U3088 (N_3088,N_2918,N_2926);
or U3089 (N_3089,N_2990,N_2893);
or U3090 (N_3090,N_2883,N_2945);
nand U3091 (N_3091,N_2868,N_2858);
nand U3092 (N_3092,N_2863,N_2985);
nor U3093 (N_3093,N_2983,N_2979);
nand U3094 (N_3094,N_2978,N_2927);
or U3095 (N_3095,N_2933,N_2876);
and U3096 (N_3096,N_2906,N_2943);
and U3097 (N_3097,N_2909,N_2868);
and U3098 (N_3098,N_2889,N_2987);
nand U3099 (N_3099,N_2911,N_2859);
nor U3100 (N_3100,N_2908,N_2906);
nor U3101 (N_3101,N_2877,N_2949);
xor U3102 (N_3102,N_2926,N_2992);
xor U3103 (N_3103,N_2865,N_2855);
nand U3104 (N_3104,N_2919,N_2988);
nor U3105 (N_3105,N_2963,N_2933);
nor U3106 (N_3106,N_2868,N_2885);
and U3107 (N_3107,N_2873,N_2977);
or U3108 (N_3108,N_2934,N_2959);
or U3109 (N_3109,N_2924,N_2932);
nand U3110 (N_3110,N_2973,N_2884);
nand U3111 (N_3111,N_2983,N_2880);
nand U3112 (N_3112,N_2876,N_2888);
or U3113 (N_3113,N_2899,N_2876);
nor U3114 (N_3114,N_2986,N_2985);
nor U3115 (N_3115,N_2869,N_2974);
nand U3116 (N_3116,N_2947,N_2863);
nor U3117 (N_3117,N_2911,N_2987);
and U3118 (N_3118,N_2892,N_2896);
xor U3119 (N_3119,N_2918,N_2963);
xnor U3120 (N_3120,N_2945,N_2855);
nand U3121 (N_3121,N_2973,N_2945);
xnor U3122 (N_3122,N_2994,N_2972);
nor U3123 (N_3123,N_2885,N_2957);
or U3124 (N_3124,N_2875,N_2981);
nand U3125 (N_3125,N_2854,N_2957);
nor U3126 (N_3126,N_2951,N_2870);
and U3127 (N_3127,N_2955,N_2888);
nand U3128 (N_3128,N_2894,N_2910);
or U3129 (N_3129,N_2911,N_2913);
and U3130 (N_3130,N_2937,N_2907);
or U3131 (N_3131,N_2955,N_2880);
nor U3132 (N_3132,N_2972,N_2953);
nor U3133 (N_3133,N_2930,N_2938);
nand U3134 (N_3134,N_2953,N_2866);
nor U3135 (N_3135,N_2944,N_2879);
xnor U3136 (N_3136,N_2934,N_2889);
nor U3137 (N_3137,N_2965,N_2946);
and U3138 (N_3138,N_2967,N_2913);
and U3139 (N_3139,N_2976,N_2876);
nor U3140 (N_3140,N_2973,N_2935);
nor U3141 (N_3141,N_2951,N_2941);
or U3142 (N_3142,N_2975,N_2947);
nand U3143 (N_3143,N_2967,N_2966);
and U3144 (N_3144,N_2978,N_2917);
xor U3145 (N_3145,N_2952,N_2946);
and U3146 (N_3146,N_2885,N_2902);
or U3147 (N_3147,N_2881,N_2988);
xor U3148 (N_3148,N_2889,N_2951);
xnor U3149 (N_3149,N_2910,N_2984);
or U3150 (N_3150,N_3142,N_3104);
or U3151 (N_3151,N_3080,N_3032);
nor U3152 (N_3152,N_3073,N_3018);
nand U3153 (N_3153,N_3108,N_3140);
nand U3154 (N_3154,N_3122,N_3099);
or U3155 (N_3155,N_3047,N_3064);
and U3156 (N_3156,N_3119,N_3051);
xnor U3157 (N_3157,N_3083,N_3093);
xnor U3158 (N_3158,N_3105,N_3075);
nor U3159 (N_3159,N_3026,N_3078);
nor U3160 (N_3160,N_3056,N_3143);
nor U3161 (N_3161,N_3004,N_3035);
and U3162 (N_3162,N_3116,N_3039);
and U3163 (N_3163,N_3081,N_3011);
xor U3164 (N_3164,N_3120,N_3068);
nand U3165 (N_3165,N_3141,N_3144);
nor U3166 (N_3166,N_3028,N_3046);
xor U3167 (N_3167,N_3006,N_3023);
or U3168 (N_3168,N_3045,N_3087);
or U3169 (N_3169,N_3117,N_3054);
and U3170 (N_3170,N_3059,N_3037);
nor U3171 (N_3171,N_3082,N_3149);
nor U3172 (N_3172,N_3049,N_3041);
and U3173 (N_3173,N_3077,N_3000);
xnor U3174 (N_3174,N_3029,N_3094);
or U3175 (N_3175,N_3025,N_3146);
or U3176 (N_3176,N_3020,N_3061);
and U3177 (N_3177,N_3036,N_3015);
nor U3178 (N_3178,N_3050,N_3027);
xor U3179 (N_3179,N_3145,N_3067);
nand U3180 (N_3180,N_3100,N_3113);
nand U3181 (N_3181,N_3024,N_3096);
and U3182 (N_3182,N_3009,N_3103);
xnor U3183 (N_3183,N_3019,N_3044);
xnor U3184 (N_3184,N_3112,N_3005);
nand U3185 (N_3185,N_3069,N_3111);
xor U3186 (N_3186,N_3098,N_3065);
or U3187 (N_3187,N_3127,N_3130);
and U3188 (N_3188,N_3095,N_3126);
nor U3189 (N_3189,N_3106,N_3125);
nor U3190 (N_3190,N_3136,N_3071);
xnor U3191 (N_3191,N_3089,N_3123);
nand U3192 (N_3192,N_3118,N_3090);
nand U3193 (N_3193,N_3086,N_3128);
and U3194 (N_3194,N_3101,N_3102);
nor U3195 (N_3195,N_3129,N_3053);
nand U3196 (N_3196,N_3088,N_3121);
and U3197 (N_3197,N_3042,N_3007);
or U3198 (N_3198,N_3003,N_3002);
nand U3199 (N_3199,N_3135,N_3058);
and U3200 (N_3200,N_3010,N_3017);
or U3201 (N_3201,N_3092,N_3030);
and U3202 (N_3202,N_3132,N_3070);
xnor U3203 (N_3203,N_3016,N_3033);
nor U3204 (N_3204,N_3057,N_3062);
or U3205 (N_3205,N_3079,N_3060);
nand U3206 (N_3206,N_3014,N_3072);
and U3207 (N_3207,N_3031,N_3084);
xnor U3208 (N_3208,N_3133,N_3034);
or U3209 (N_3209,N_3124,N_3063);
xnor U3210 (N_3210,N_3134,N_3137);
or U3211 (N_3211,N_3038,N_3066);
nand U3212 (N_3212,N_3048,N_3110);
and U3213 (N_3213,N_3055,N_3076);
nor U3214 (N_3214,N_3147,N_3091);
nor U3215 (N_3215,N_3040,N_3114);
or U3216 (N_3216,N_3109,N_3107);
nand U3217 (N_3217,N_3085,N_3008);
and U3218 (N_3218,N_3021,N_3148);
nor U3219 (N_3219,N_3013,N_3097);
nor U3220 (N_3220,N_3115,N_3138);
nor U3221 (N_3221,N_3131,N_3139);
nor U3222 (N_3222,N_3001,N_3052);
xor U3223 (N_3223,N_3043,N_3074);
xor U3224 (N_3224,N_3012,N_3022);
and U3225 (N_3225,N_3092,N_3125);
and U3226 (N_3226,N_3052,N_3109);
nand U3227 (N_3227,N_3117,N_3033);
or U3228 (N_3228,N_3070,N_3030);
and U3229 (N_3229,N_3047,N_3032);
or U3230 (N_3230,N_3135,N_3089);
nand U3231 (N_3231,N_3000,N_3137);
and U3232 (N_3232,N_3100,N_3126);
xor U3233 (N_3233,N_3141,N_3005);
or U3234 (N_3234,N_3128,N_3062);
xnor U3235 (N_3235,N_3056,N_3126);
or U3236 (N_3236,N_3142,N_3029);
nand U3237 (N_3237,N_3074,N_3119);
xor U3238 (N_3238,N_3040,N_3025);
nor U3239 (N_3239,N_3116,N_3125);
nor U3240 (N_3240,N_3139,N_3041);
nor U3241 (N_3241,N_3057,N_3142);
nor U3242 (N_3242,N_3014,N_3119);
nand U3243 (N_3243,N_3141,N_3071);
nand U3244 (N_3244,N_3052,N_3027);
or U3245 (N_3245,N_3148,N_3007);
nor U3246 (N_3246,N_3111,N_3135);
xor U3247 (N_3247,N_3109,N_3068);
xor U3248 (N_3248,N_3096,N_3095);
and U3249 (N_3249,N_3113,N_3093);
nor U3250 (N_3250,N_3094,N_3090);
or U3251 (N_3251,N_3002,N_3062);
and U3252 (N_3252,N_3001,N_3051);
nor U3253 (N_3253,N_3097,N_3106);
xor U3254 (N_3254,N_3140,N_3022);
and U3255 (N_3255,N_3113,N_3011);
or U3256 (N_3256,N_3089,N_3126);
nor U3257 (N_3257,N_3053,N_3056);
and U3258 (N_3258,N_3061,N_3080);
nor U3259 (N_3259,N_3021,N_3106);
nor U3260 (N_3260,N_3039,N_3091);
or U3261 (N_3261,N_3144,N_3029);
xnor U3262 (N_3262,N_3072,N_3026);
xnor U3263 (N_3263,N_3053,N_3124);
and U3264 (N_3264,N_3028,N_3048);
and U3265 (N_3265,N_3067,N_3079);
nand U3266 (N_3266,N_3076,N_3140);
and U3267 (N_3267,N_3080,N_3007);
xnor U3268 (N_3268,N_3036,N_3045);
or U3269 (N_3269,N_3098,N_3012);
or U3270 (N_3270,N_3078,N_3145);
xor U3271 (N_3271,N_3065,N_3012);
or U3272 (N_3272,N_3031,N_3018);
nor U3273 (N_3273,N_3105,N_3121);
or U3274 (N_3274,N_3089,N_3139);
or U3275 (N_3275,N_3087,N_3134);
nand U3276 (N_3276,N_3111,N_3056);
xnor U3277 (N_3277,N_3088,N_3066);
or U3278 (N_3278,N_3142,N_3121);
nor U3279 (N_3279,N_3072,N_3092);
nor U3280 (N_3280,N_3014,N_3146);
xor U3281 (N_3281,N_3117,N_3047);
xor U3282 (N_3282,N_3104,N_3087);
xor U3283 (N_3283,N_3116,N_3065);
or U3284 (N_3284,N_3091,N_3094);
and U3285 (N_3285,N_3044,N_3001);
and U3286 (N_3286,N_3128,N_3040);
nor U3287 (N_3287,N_3049,N_3106);
nand U3288 (N_3288,N_3048,N_3149);
xor U3289 (N_3289,N_3070,N_3054);
and U3290 (N_3290,N_3028,N_3066);
and U3291 (N_3291,N_3017,N_3015);
or U3292 (N_3292,N_3010,N_3053);
nor U3293 (N_3293,N_3135,N_3041);
xor U3294 (N_3294,N_3047,N_3120);
or U3295 (N_3295,N_3149,N_3030);
nand U3296 (N_3296,N_3144,N_3065);
xnor U3297 (N_3297,N_3015,N_3002);
nor U3298 (N_3298,N_3116,N_3016);
and U3299 (N_3299,N_3063,N_3100);
xor U3300 (N_3300,N_3297,N_3264);
nand U3301 (N_3301,N_3284,N_3155);
nor U3302 (N_3302,N_3294,N_3181);
nor U3303 (N_3303,N_3208,N_3285);
or U3304 (N_3304,N_3199,N_3157);
nand U3305 (N_3305,N_3267,N_3281);
nor U3306 (N_3306,N_3175,N_3204);
or U3307 (N_3307,N_3184,N_3236);
nand U3308 (N_3308,N_3152,N_3185);
and U3309 (N_3309,N_3273,N_3252);
nand U3310 (N_3310,N_3195,N_3174);
or U3311 (N_3311,N_3156,N_3198);
xnor U3312 (N_3312,N_3235,N_3228);
and U3313 (N_3313,N_3182,N_3286);
nor U3314 (N_3314,N_3176,N_3154);
nor U3315 (N_3315,N_3161,N_3233);
xor U3316 (N_3316,N_3210,N_3200);
nor U3317 (N_3317,N_3205,N_3262);
and U3318 (N_3318,N_3206,N_3258);
and U3319 (N_3319,N_3274,N_3222);
and U3320 (N_3320,N_3295,N_3150);
xnor U3321 (N_3321,N_3272,N_3259);
xnor U3322 (N_3322,N_3250,N_3159);
and U3323 (N_3323,N_3240,N_3291);
nor U3324 (N_3324,N_3194,N_3169);
nor U3325 (N_3325,N_3191,N_3179);
and U3326 (N_3326,N_3217,N_3171);
xor U3327 (N_3327,N_3265,N_3219);
nor U3328 (N_3328,N_3160,N_3266);
nor U3329 (N_3329,N_3153,N_3170);
or U3330 (N_3330,N_3293,N_3212);
and U3331 (N_3331,N_3234,N_3268);
and U3332 (N_3332,N_3213,N_3249);
xnor U3333 (N_3333,N_3244,N_3166);
or U3334 (N_3334,N_3211,N_3231);
nor U3335 (N_3335,N_3237,N_3292);
nor U3336 (N_3336,N_3243,N_3216);
nor U3337 (N_3337,N_3188,N_3271);
nor U3338 (N_3338,N_3256,N_3178);
nand U3339 (N_3339,N_3261,N_3283);
xor U3340 (N_3340,N_3263,N_3203);
and U3341 (N_3341,N_3260,N_3183);
or U3342 (N_3342,N_3289,N_3167);
nor U3343 (N_3343,N_3246,N_3253);
nand U3344 (N_3344,N_3226,N_3296);
or U3345 (N_3345,N_3187,N_3224);
and U3346 (N_3346,N_3248,N_3177);
or U3347 (N_3347,N_3251,N_3270);
nand U3348 (N_3348,N_3280,N_3299);
or U3349 (N_3349,N_3202,N_3232);
nor U3350 (N_3350,N_3201,N_3220);
nand U3351 (N_3351,N_3214,N_3254);
and U3352 (N_3352,N_3290,N_3193);
and U3353 (N_3353,N_3242,N_3239);
and U3354 (N_3354,N_3276,N_3172);
xnor U3355 (N_3355,N_3255,N_3207);
and U3356 (N_3356,N_3238,N_3218);
or U3357 (N_3357,N_3173,N_3278);
nor U3358 (N_3358,N_3215,N_3192);
xor U3359 (N_3359,N_3275,N_3227);
nand U3360 (N_3360,N_3163,N_3282);
or U3361 (N_3361,N_3168,N_3162);
and U3362 (N_3362,N_3196,N_3225);
or U3363 (N_3363,N_3288,N_3245);
nand U3364 (N_3364,N_3223,N_3190);
xnor U3365 (N_3365,N_3180,N_3189);
nor U3366 (N_3366,N_3209,N_3164);
or U3367 (N_3367,N_3165,N_3269);
xnor U3368 (N_3368,N_3151,N_3257);
nand U3369 (N_3369,N_3279,N_3158);
nand U3370 (N_3370,N_3197,N_3287);
and U3371 (N_3371,N_3298,N_3221);
and U3372 (N_3372,N_3230,N_3186);
or U3373 (N_3373,N_3277,N_3247);
and U3374 (N_3374,N_3241,N_3229);
xor U3375 (N_3375,N_3280,N_3225);
and U3376 (N_3376,N_3247,N_3283);
nand U3377 (N_3377,N_3204,N_3211);
nand U3378 (N_3378,N_3253,N_3265);
and U3379 (N_3379,N_3196,N_3195);
nand U3380 (N_3380,N_3279,N_3183);
nand U3381 (N_3381,N_3242,N_3188);
nand U3382 (N_3382,N_3227,N_3248);
nand U3383 (N_3383,N_3255,N_3257);
or U3384 (N_3384,N_3212,N_3196);
nand U3385 (N_3385,N_3179,N_3296);
or U3386 (N_3386,N_3261,N_3282);
nand U3387 (N_3387,N_3157,N_3171);
or U3388 (N_3388,N_3158,N_3196);
and U3389 (N_3389,N_3176,N_3229);
nand U3390 (N_3390,N_3159,N_3217);
nor U3391 (N_3391,N_3172,N_3233);
or U3392 (N_3392,N_3172,N_3197);
or U3393 (N_3393,N_3276,N_3262);
xnor U3394 (N_3394,N_3258,N_3246);
and U3395 (N_3395,N_3277,N_3182);
and U3396 (N_3396,N_3271,N_3210);
xor U3397 (N_3397,N_3258,N_3233);
and U3398 (N_3398,N_3238,N_3158);
xor U3399 (N_3399,N_3167,N_3176);
and U3400 (N_3400,N_3265,N_3258);
xnor U3401 (N_3401,N_3239,N_3171);
nor U3402 (N_3402,N_3264,N_3291);
or U3403 (N_3403,N_3268,N_3292);
nand U3404 (N_3404,N_3155,N_3256);
nand U3405 (N_3405,N_3205,N_3226);
and U3406 (N_3406,N_3216,N_3154);
and U3407 (N_3407,N_3289,N_3245);
nor U3408 (N_3408,N_3259,N_3231);
nor U3409 (N_3409,N_3197,N_3168);
nand U3410 (N_3410,N_3282,N_3210);
nor U3411 (N_3411,N_3227,N_3232);
nand U3412 (N_3412,N_3184,N_3200);
nor U3413 (N_3413,N_3212,N_3166);
and U3414 (N_3414,N_3292,N_3251);
nand U3415 (N_3415,N_3204,N_3299);
xnor U3416 (N_3416,N_3150,N_3224);
or U3417 (N_3417,N_3249,N_3255);
xor U3418 (N_3418,N_3155,N_3262);
nand U3419 (N_3419,N_3291,N_3276);
nor U3420 (N_3420,N_3225,N_3264);
nand U3421 (N_3421,N_3210,N_3156);
nor U3422 (N_3422,N_3160,N_3178);
nor U3423 (N_3423,N_3178,N_3283);
and U3424 (N_3424,N_3193,N_3163);
or U3425 (N_3425,N_3257,N_3192);
nand U3426 (N_3426,N_3161,N_3206);
and U3427 (N_3427,N_3265,N_3200);
nand U3428 (N_3428,N_3168,N_3253);
nor U3429 (N_3429,N_3193,N_3160);
or U3430 (N_3430,N_3299,N_3264);
or U3431 (N_3431,N_3249,N_3266);
nor U3432 (N_3432,N_3254,N_3164);
nor U3433 (N_3433,N_3225,N_3235);
xnor U3434 (N_3434,N_3204,N_3296);
or U3435 (N_3435,N_3299,N_3181);
nor U3436 (N_3436,N_3219,N_3218);
xnor U3437 (N_3437,N_3273,N_3204);
xnor U3438 (N_3438,N_3225,N_3178);
nand U3439 (N_3439,N_3178,N_3220);
and U3440 (N_3440,N_3258,N_3188);
or U3441 (N_3441,N_3283,N_3296);
or U3442 (N_3442,N_3211,N_3283);
nor U3443 (N_3443,N_3264,N_3251);
xor U3444 (N_3444,N_3213,N_3206);
and U3445 (N_3445,N_3179,N_3269);
xnor U3446 (N_3446,N_3267,N_3268);
nand U3447 (N_3447,N_3238,N_3234);
xnor U3448 (N_3448,N_3177,N_3187);
nand U3449 (N_3449,N_3153,N_3207);
nand U3450 (N_3450,N_3314,N_3311);
nor U3451 (N_3451,N_3430,N_3349);
nor U3452 (N_3452,N_3306,N_3360);
nand U3453 (N_3453,N_3307,N_3379);
nor U3454 (N_3454,N_3301,N_3433);
or U3455 (N_3455,N_3352,N_3367);
and U3456 (N_3456,N_3348,N_3309);
nand U3457 (N_3457,N_3401,N_3415);
and U3458 (N_3458,N_3376,N_3381);
or U3459 (N_3459,N_3442,N_3361);
nand U3460 (N_3460,N_3405,N_3357);
xnor U3461 (N_3461,N_3339,N_3341);
or U3462 (N_3462,N_3315,N_3438);
nand U3463 (N_3463,N_3448,N_3305);
nand U3464 (N_3464,N_3300,N_3414);
or U3465 (N_3465,N_3391,N_3358);
or U3466 (N_3466,N_3346,N_3332);
xor U3467 (N_3467,N_3362,N_3343);
nor U3468 (N_3468,N_3388,N_3427);
and U3469 (N_3469,N_3320,N_3340);
and U3470 (N_3470,N_3383,N_3322);
and U3471 (N_3471,N_3359,N_3431);
nand U3472 (N_3472,N_3366,N_3331);
or U3473 (N_3473,N_3390,N_3378);
and U3474 (N_3474,N_3402,N_3373);
nor U3475 (N_3475,N_3428,N_3369);
and U3476 (N_3476,N_3395,N_3308);
nand U3477 (N_3477,N_3344,N_3419);
xor U3478 (N_3478,N_3417,N_3325);
and U3479 (N_3479,N_3304,N_3437);
xnor U3480 (N_3480,N_3434,N_3371);
or U3481 (N_3481,N_3387,N_3432);
nand U3482 (N_3482,N_3412,N_3420);
xnor U3483 (N_3483,N_3338,N_3347);
nand U3484 (N_3484,N_3445,N_3355);
nor U3485 (N_3485,N_3394,N_3404);
xnor U3486 (N_3486,N_3425,N_3345);
and U3487 (N_3487,N_3393,N_3303);
or U3488 (N_3488,N_3422,N_3389);
nand U3489 (N_3489,N_3375,N_3410);
or U3490 (N_3490,N_3319,N_3399);
xnor U3491 (N_3491,N_3374,N_3421);
nor U3492 (N_3492,N_3403,N_3385);
nor U3493 (N_3493,N_3397,N_3372);
or U3494 (N_3494,N_3337,N_3302);
and U3495 (N_3495,N_3313,N_3321);
xor U3496 (N_3496,N_3329,N_3380);
or U3497 (N_3497,N_3416,N_3396);
nor U3498 (N_3498,N_3353,N_3351);
nor U3499 (N_3499,N_3449,N_3446);
and U3500 (N_3500,N_3370,N_3317);
and U3501 (N_3501,N_3409,N_3336);
and U3502 (N_3502,N_3407,N_3368);
xor U3503 (N_3503,N_3333,N_3312);
nor U3504 (N_3504,N_3411,N_3436);
or U3505 (N_3505,N_3310,N_3342);
nand U3506 (N_3506,N_3365,N_3384);
xor U3507 (N_3507,N_3441,N_3350);
and U3508 (N_3508,N_3326,N_3408);
nor U3509 (N_3509,N_3400,N_3382);
and U3510 (N_3510,N_3334,N_3424);
nor U3511 (N_3511,N_3377,N_3327);
nand U3512 (N_3512,N_3318,N_3435);
nor U3513 (N_3513,N_3444,N_3323);
nor U3514 (N_3514,N_3398,N_3413);
and U3515 (N_3515,N_3429,N_3328);
or U3516 (N_3516,N_3363,N_3364);
nor U3517 (N_3517,N_3392,N_3356);
nor U3518 (N_3518,N_3330,N_3335);
or U3519 (N_3519,N_3426,N_3440);
xnor U3520 (N_3520,N_3324,N_3418);
xor U3521 (N_3521,N_3439,N_3447);
xor U3522 (N_3522,N_3316,N_3423);
xor U3523 (N_3523,N_3443,N_3406);
nor U3524 (N_3524,N_3354,N_3386);
or U3525 (N_3525,N_3347,N_3413);
nor U3526 (N_3526,N_3378,N_3339);
nor U3527 (N_3527,N_3405,N_3417);
and U3528 (N_3528,N_3330,N_3411);
nor U3529 (N_3529,N_3381,N_3325);
nor U3530 (N_3530,N_3422,N_3343);
nor U3531 (N_3531,N_3367,N_3312);
xor U3532 (N_3532,N_3383,N_3433);
or U3533 (N_3533,N_3404,N_3351);
and U3534 (N_3534,N_3314,N_3380);
nor U3535 (N_3535,N_3390,N_3415);
xor U3536 (N_3536,N_3363,N_3437);
xor U3537 (N_3537,N_3448,N_3362);
nand U3538 (N_3538,N_3328,N_3369);
and U3539 (N_3539,N_3361,N_3315);
and U3540 (N_3540,N_3340,N_3378);
nor U3541 (N_3541,N_3446,N_3414);
and U3542 (N_3542,N_3323,N_3383);
nor U3543 (N_3543,N_3372,N_3320);
nand U3544 (N_3544,N_3318,N_3409);
and U3545 (N_3545,N_3316,N_3442);
or U3546 (N_3546,N_3441,N_3422);
nand U3547 (N_3547,N_3349,N_3381);
xor U3548 (N_3548,N_3328,N_3446);
xor U3549 (N_3549,N_3362,N_3308);
or U3550 (N_3550,N_3325,N_3330);
xor U3551 (N_3551,N_3338,N_3441);
or U3552 (N_3552,N_3349,N_3427);
or U3553 (N_3553,N_3449,N_3448);
and U3554 (N_3554,N_3395,N_3442);
nor U3555 (N_3555,N_3381,N_3420);
and U3556 (N_3556,N_3320,N_3409);
and U3557 (N_3557,N_3345,N_3361);
xnor U3558 (N_3558,N_3340,N_3408);
or U3559 (N_3559,N_3401,N_3381);
or U3560 (N_3560,N_3318,N_3405);
nor U3561 (N_3561,N_3423,N_3301);
or U3562 (N_3562,N_3323,N_3355);
nor U3563 (N_3563,N_3393,N_3310);
nor U3564 (N_3564,N_3435,N_3391);
or U3565 (N_3565,N_3375,N_3448);
xor U3566 (N_3566,N_3395,N_3413);
and U3567 (N_3567,N_3426,N_3403);
or U3568 (N_3568,N_3341,N_3387);
or U3569 (N_3569,N_3307,N_3337);
nand U3570 (N_3570,N_3321,N_3317);
nand U3571 (N_3571,N_3323,N_3437);
or U3572 (N_3572,N_3322,N_3354);
nand U3573 (N_3573,N_3430,N_3348);
nand U3574 (N_3574,N_3325,N_3427);
and U3575 (N_3575,N_3420,N_3321);
nor U3576 (N_3576,N_3365,N_3330);
and U3577 (N_3577,N_3332,N_3394);
xnor U3578 (N_3578,N_3436,N_3305);
and U3579 (N_3579,N_3369,N_3403);
or U3580 (N_3580,N_3343,N_3384);
nand U3581 (N_3581,N_3338,N_3326);
or U3582 (N_3582,N_3383,N_3329);
nor U3583 (N_3583,N_3326,N_3331);
xor U3584 (N_3584,N_3416,N_3320);
or U3585 (N_3585,N_3346,N_3300);
nor U3586 (N_3586,N_3390,N_3429);
or U3587 (N_3587,N_3418,N_3317);
nand U3588 (N_3588,N_3363,N_3394);
or U3589 (N_3589,N_3448,N_3334);
xor U3590 (N_3590,N_3435,N_3393);
nand U3591 (N_3591,N_3399,N_3356);
and U3592 (N_3592,N_3347,N_3329);
nor U3593 (N_3593,N_3311,N_3402);
xnor U3594 (N_3594,N_3327,N_3368);
nor U3595 (N_3595,N_3430,N_3414);
xnor U3596 (N_3596,N_3346,N_3442);
nor U3597 (N_3597,N_3335,N_3397);
and U3598 (N_3598,N_3353,N_3396);
and U3599 (N_3599,N_3364,N_3419);
and U3600 (N_3600,N_3574,N_3536);
or U3601 (N_3601,N_3455,N_3592);
and U3602 (N_3602,N_3477,N_3544);
nand U3603 (N_3603,N_3462,N_3599);
or U3604 (N_3604,N_3466,N_3553);
xnor U3605 (N_3605,N_3542,N_3469);
or U3606 (N_3606,N_3570,N_3461);
nand U3607 (N_3607,N_3456,N_3509);
or U3608 (N_3608,N_3500,N_3566);
nor U3609 (N_3609,N_3581,N_3525);
xnor U3610 (N_3610,N_3526,N_3593);
nand U3611 (N_3611,N_3490,N_3475);
and U3612 (N_3612,N_3564,N_3559);
and U3613 (N_3613,N_3523,N_3499);
or U3614 (N_3614,N_3585,N_3589);
xnor U3615 (N_3615,N_3545,N_3590);
and U3616 (N_3616,N_3532,N_3598);
or U3617 (N_3617,N_3562,N_3522);
nor U3618 (N_3618,N_3489,N_3549);
xnor U3619 (N_3619,N_3491,N_3494);
and U3620 (N_3620,N_3508,N_3541);
nand U3621 (N_3621,N_3557,N_3463);
nand U3622 (N_3622,N_3534,N_3515);
nor U3623 (N_3623,N_3576,N_3452);
nor U3624 (N_3624,N_3468,N_3498);
or U3625 (N_3625,N_3478,N_3464);
xnor U3626 (N_3626,N_3512,N_3577);
xor U3627 (N_3627,N_3540,N_3529);
or U3628 (N_3628,N_3484,N_3597);
or U3629 (N_3629,N_3516,N_3546);
or U3630 (N_3630,N_3539,N_3483);
nand U3631 (N_3631,N_3518,N_3514);
xor U3632 (N_3632,N_3501,N_3531);
nor U3633 (N_3633,N_3563,N_3521);
or U3634 (N_3634,N_3552,N_3560);
or U3635 (N_3635,N_3450,N_3582);
or U3636 (N_3636,N_3548,N_3485);
nor U3637 (N_3637,N_3473,N_3594);
nor U3638 (N_3638,N_3465,N_3502);
or U3639 (N_3639,N_3480,N_3471);
xor U3640 (N_3640,N_3595,N_3569);
and U3641 (N_3641,N_3535,N_3457);
and U3642 (N_3642,N_3470,N_3556);
nand U3643 (N_3643,N_3504,N_3567);
nand U3644 (N_3644,N_3520,N_3495);
xor U3645 (N_3645,N_3493,N_3558);
xnor U3646 (N_3646,N_3453,N_3481);
and U3647 (N_3647,N_3503,N_3578);
or U3648 (N_3648,N_3474,N_3459);
and U3649 (N_3649,N_3486,N_3505);
or U3650 (N_3650,N_3554,N_3571);
and U3651 (N_3651,N_3555,N_3496);
and U3652 (N_3652,N_3572,N_3507);
and U3653 (N_3653,N_3568,N_3580);
nor U3654 (N_3654,N_3454,N_3561);
xnor U3655 (N_3655,N_3506,N_3487);
nor U3656 (N_3656,N_3467,N_3591);
xnor U3657 (N_3657,N_3583,N_3596);
nand U3658 (N_3658,N_3579,N_3511);
and U3659 (N_3659,N_3530,N_3565);
or U3660 (N_3660,N_3587,N_3588);
nand U3661 (N_3661,N_3458,N_3451);
nor U3662 (N_3662,N_3524,N_3482);
nor U3663 (N_3663,N_3586,N_3492);
xor U3664 (N_3664,N_3460,N_3497);
or U3665 (N_3665,N_3550,N_3547);
and U3666 (N_3666,N_3543,N_3479);
and U3667 (N_3667,N_3573,N_3575);
nand U3668 (N_3668,N_3527,N_3551);
nor U3669 (N_3669,N_3476,N_3510);
nor U3670 (N_3670,N_3519,N_3528);
nor U3671 (N_3671,N_3517,N_3584);
nand U3672 (N_3672,N_3533,N_3538);
nand U3673 (N_3673,N_3537,N_3513);
nor U3674 (N_3674,N_3488,N_3472);
or U3675 (N_3675,N_3461,N_3513);
and U3676 (N_3676,N_3578,N_3552);
xor U3677 (N_3677,N_3590,N_3563);
and U3678 (N_3678,N_3580,N_3523);
xor U3679 (N_3679,N_3498,N_3568);
or U3680 (N_3680,N_3582,N_3585);
and U3681 (N_3681,N_3451,N_3511);
and U3682 (N_3682,N_3527,N_3553);
xnor U3683 (N_3683,N_3480,N_3497);
and U3684 (N_3684,N_3533,N_3475);
xnor U3685 (N_3685,N_3534,N_3557);
nand U3686 (N_3686,N_3508,N_3477);
nand U3687 (N_3687,N_3459,N_3548);
nand U3688 (N_3688,N_3562,N_3538);
and U3689 (N_3689,N_3572,N_3575);
nand U3690 (N_3690,N_3484,N_3518);
xor U3691 (N_3691,N_3580,N_3481);
or U3692 (N_3692,N_3549,N_3518);
nor U3693 (N_3693,N_3552,N_3550);
nand U3694 (N_3694,N_3554,N_3598);
nor U3695 (N_3695,N_3585,N_3495);
nor U3696 (N_3696,N_3554,N_3534);
nand U3697 (N_3697,N_3485,N_3577);
or U3698 (N_3698,N_3507,N_3467);
or U3699 (N_3699,N_3500,N_3549);
and U3700 (N_3700,N_3459,N_3468);
and U3701 (N_3701,N_3521,N_3479);
and U3702 (N_3702,N_3573,N_3461);
nor U3703 (N_3703,N_3580,N_3472);
nand U3704 (N_3704,N_3582,N_3471);
nor U3705 (N_3705,N_3462,N_3499);
nand U3706 (N_3706,N_3484,N_3509);
nand U3707 (N_3707,N_3472,N_3514);
and U3708 (N_3708,N_3517,N_3590);
xnor U3709 (N_3709,N_3572,N_3584);
nor U3710 (N_3710,N_3545,N_3565);
and U3711 (N_3711,N_3510,N_3516);
and U3712 (N_3712,N_3507,N_3544);
xnor U3713 (N_3713,N_3509,N_3531);
and U3714 (N_3714,N_3489,N_3591);
nand U3715 (N_3715,N_3563,N_3537);
nand U3716 (N_3716,N_3463,N_3530);
nand U3717 (N_3717,N_3576,N_3590);
and U3718 (N_3718,N_3452,N_3474);
xor U3719 (N_3719,N_3512,N_3499);
xor U3720 (N_3720,N_3560,N_3571);
nand U3721 (N_3721,N_3466,N_3459);
nand U3722 (N_3722,N_3563,N_3523);
and U3723 (N_3723,N_3585,N_3537);
nor U3724 (N_3724,N_3584,N_3530);
nor U3725 (N_3725,N_3546,N_3470);
xnor U3726 (N_3726,N_3564,N_3562);
or U3727 (N_3727,N_3583,N_3467);
and U3728 (N_3728,N_3450,N_3561);
nor U3729 (N_3729,N_3530,N_3477);
nand U3730 (N_3730,N_3597,N_3483);
nand U3731 (N_3731,N_3487,N_3595);
and U3732 (N_3732,N_3576,N_3534);
or U3733 (N_3733,N_3578,N_3477);
or U3734 (N_3734,N_3549,N_3471);
nand U3735 (N_3735,N_3583,N_3585);
or U3736 (N_3736,N_3591,N_3576);
xnor U3737 (N_3737,N_3567,N_3505);
and U3738 (N_3738,N_3523,N_3487);
or U3739 (N_3739,N_3453,N_3533);
nand U3740 (N_3740,N_3523,N_3502);
or U3741 (N_3741,N_3487,N_3504);
or U3742 (N_3742,N_3521,N_3528);
or U3743 (N_3743,N_3515,N_3485);
or U3744 (N_3744,N_3538,N_3467);
or U3745 (N_3745,N_3510,N_3546);
and U3746 (N_3746,N_3517,N_3567);
or U3747 (N_3747,N_3576,N_3557);
and U3748 (N_3748,N_3586,N_3578);
nor U3749 (N_3749,N_3486,N_3498);
xnor U3750 (N_3750,N_3627,N_3703);
and U3751 (N_3751,N_3678,N_3666);
and U3752 (N_3752,N_3675,N_3652);
and U3753 (N_3753,N_3602,N_3662);
nor U3754 (N_3754,N_3721,N_3713);
nor U3755 (N_3755,N_3746,N_3702);
or U3756 (N_3756,N_3685,N_3710);
nor U3757 (N_3757,N_3735,N_3628);
nand U3758 (N_3758,N_3653,N_3658);
and U3759 (N_3759,N_3711,N_3691);
or U3760 (N_3760,N_3664,N_3733);
nand U3761 (N_3761,N_3625,N_3659);
nand U3762 (N_3762,N_3660,N_3640);
xnor U3763 (N_3763,N_3632,N_3638);
nand U3764 (N_3764,N_3724,N_3695);
or U3765 (N_3765,N_3607,N_3683);
xnor U3766 (N_3766,N_3667,N_3704);
nand U3767 (N_3767,N_3612,N_3737);
xor U3768 (N_3768,N_3604,N_3631);
or U3769 (N_3769,N_3728,N_3620);
xnor U3770 (N_3770,N_3616,N_3749);
nor U3771 (N_3771,N_3633,N_3689);
nor U3772 (N_3772,N_3629,N_3741);
nand U3773 (N_3773,N_3674,N_3693);
nor U3774 (N_3774,N_3697,N_3649);
nand U3775 (N_3775,N_3611,N_3641);
and U3776 (N_3776,N_3606,N_3644);
nand U3777 (N_3777,N_3635,N_3740);
or U3778 (N_3778,N_3643,N_3698);
or U3779 (N_3779,N_3739,N_3670);
nor U3780 (N_3780,N_3731,N_3723);
or U3781 (N_3781,N_3719,N_3716);
nand U3782 (N_3782,N_3679,N_3603);
nor U3783 (N_3783,N_3676,N_3743);
and U3784 (N_3784,N_3673,N_3726);
and U3785 (N_3785,N_3648,N_3677);
nand U3786 (N_3786,N_3617,N_3745);
nand U3787 (N_3787,N_3732,N_3730);
and U3788 (N_3788,N_3655,N_3637);
nand U3789 (N_3789,N_3608,N_3738);
nor U3790 (N_3790,N_3657,N_3729);
nand U3791 (N_3791,N_3684,N_3700);
and U3792 (N_3792,N_3709,N_3610);
or U3793 (N_3793,N_3645,N_3609);
or U3794 (N_3794,N_3720,N_3618);
or U3795 (N_3795,N_3706,N_3601);
nand U3796 (N_3796,N_3682,N_3686);
nand U3797 (N_3797,N_3656,N_3665);
nor U3798 (N_3798,N_3699,N_3651);
and U3799 (N_3799,N_3630,N_3692);
nand U3800 (N_3800,N_3748,N_3680);
and U3801 (N_3801,N_3647,N_3668);
and U3802 (N_3802,N_3661,N_3605);
xnor U3803 (N_3803,N_3623,N_3725);
or U3804 (N_3804,N_3636,N_3744);
xnor U3805 (N_3805,N_3717,N_3654);
and U3806 (N_3806,N_3715,N_3622);
and U3807 (N_3807,N_3615,N_3621);
nor U3808 (N_3808,N_3736,N_3681);
or U3809 (N_3809,N_3600,N_3687);
or U3810 (N_3810,N_3714,N_3626);
xnor U3811 (N_3811,N_3671,N_3747);
xnor U3812 (N_3812,N_3708,N_3694);
nor U3813 (N_3813,N_3624,N_3705);
nand U3814 (N_3814,N_3672,N_3613);
or U3815 (N_3815,N_3669,N_3642);
nand U3816 (N_3816,N_3688,N_3742);
nor U3817 (N_3817,N_3701,N_3634);
xor U3818 (N_3818,N_3639,N_3727);
nand U3819 (N_3819,N_3663,N_3734);
nand U3820 (N_3820,N_3690,N_3712);
nand U3821 (N_3821,N_3696,N_3707);
and U3822 (N_3822,N_3614,N_3619);
and U3823 (N_3823,N_3650,N_3722);
xnor U3824 (N_3824,N_3718,N_3646);
nand U3825 (N_3825,N_3600,N_3698);
nor U3826 (N_3826,N_3615,N_3669);
nand U3827 (N_3827,N_3653,N_3735);
nor U3828 (N_3828,N_3738,N_3707);
nor U3829 (N_3829,N_3693,N_3731);
nor U3830 (N_3830,N_3648,N_3749);
nand U3831 (N_3831,N_3617,N_3635);
and U3832 (N_3832,N_3641,N_3690);
xnor U3833 (N_3833,N_3704,N_3694);
nand U3834 (N_3834,N_3744,N_3749);
xnor U3835 (N_3835,N_3686,N_3610);
and U3836 (N_3836,N_3700,N_3745);
xor U3837 (N_3837,N_3680,N_3685);
nand U3838 (N_3838,N_3691,N_3615);
nor U3839 (N_3839,N_3623,N_3744);
xnor U3840 (N_3840,N_3717,N_3607);
nor U3841 (N_3841,N_3667,N_3690);
or U3842 (N_3842,N_3721,N_3637);
nand U3843 (N_3843,N_3733,N_3735);
and U3844 (N_3844,N_3672,N_3698);
nand U3845 (N_3845,N_3746,N_3638);
or U3846 (N_3846,N_3636,N_3604);
xor U3847 (N_3847,N_3635,N_3706);
xnor U3848 (N_3848,N_3653,N_3667);
and U3849 (N_3849,N_3639,N_3692);
or U3850 (N_3850,N_3717,N_3653);
or U3851 (N_3851,N_3625,N_3603);
and U3852 (N_3852,N_3659,N_3717);
xor U3853 (N_3853,N_3738,N_3652);
xnor U3854 (N_3854,N_3647,N_3703);
nor U3855 (N_3855,N_3720,N_3645);
or U3856 (N_3856,N_3656,N_3689);
and U3857 (N_3857,N_3738,N_3664);
or U3858 (N_3858,N_3601,N_3690);
xnor U3859 (N_3859,N_3669,N_3699);
nand U3860 (N_3860,N_3607,N_3640);
or U3861 (N_3861,N_3616,N_3678);
or U3862 (N_3862,N_3683,N_3652);
nor U3863 (N_3863,N_3629,N_3656);
or U3864 (N_3864,N_3648,N_3747);
xnor U3865 (N_3865,N_3749,N_3738);
nor U3866 (N_3866,N_3678,N_3685);
nand U3867 (N_3867,N_3703,N_3626);
and U3868 (N_3868,N_3606,N_3723);
nor U3869 (N_3869,N_3613,N_3674);
or U3870 (N_3870,N_3644,N_3688);
nor U3871 (N_3871,N_3643,N_3697);
nand U3872 (N_3872,N_3741,N_3648);
or U3873 (N_3873,N_3731,N_3648);
nor U3874 (N_3874,N_3747,N_3635);
nor U3875 (N_3875,N_3736,N_3739);
nor U3876 (N_3876,N_3632,N_3728);
nand U3877 (N_3877,N_3672,N_3734);
xnor U3878 (N_3878,N_3622,N_3685);
xor U3879 (N_3879,N_3709,N_3637);
nor U3880 (N_3880,N_3700,N_3696);
xnor U3881 (N_3881,N_3659,N_3616);
nor U3882 (N_3882,N_3616,N_3655);
or U3883 (N_3883,N_3626,N_3723);
and U3884 (N_3884,N_3636,N_3622);
or U3885 (N_3885,N_3718,N_3711);
xor U3886 (N_3886,N_3641,N_3652);
nand U3887 (N_3887,N_3637,N_3715);
xor U3888 (N_3888,N_3748,N_3695);
or U3889 (N_3889,N_3676,N_3620);
and U3890 (N_3890,N_3601,N_3630);
xor U3891 (N_3891,N_3649,N_3700);
or U3892 (N_3892,N_3724,N_3677);
and U3893 (N_3893,N_3632,N_3697);
nand U3894 (N_3894,N_3654,N_3667);
nor U3895 (N_3895,N_3633,N_3710);
nand U3896 (N_3896,N_3697,N_3641);
nor U3897 (N_3897,N_3705,N_3709);
nand U3898 (N_3898,N_3718,N_3609);
nor U3899 (N_3899,N_3651,N_3629);
and U3900 (N_3900,N_3875,N_3882);
xor U3901 (N_3901,N_3850,N_3791);
nand U3902 (N_3902,N_3832,N_3769);
and U3903 (N_3903,N_3786,N_3780);
nor U3904 (N_3904,N_3838,N_3758);
and U3905 (N_3905,N_3897,N_3873);
xor U3906 (N_3906,N_3849,N_3898);
or U3907 (N_3907,N_3768,N_3864);
xnor U3908 (N_3908,N_3833,N_3896);
nor U3909 (N_3909,N_3868,N_3848);
nor U3910 (N_3910,N_3756,N_3884);
nor U3911 (N_3911,N_3792,N_3829);
xnor U3912 (N_3912,N_3859,N_3798);
nand U3913 (N_3913,N_3801,N_3774);
xor U3914 (N_3914,N_3888,N_3891);
nand U3915 (N_3915,N_3787,N_3809);
and U3916 (N_3916,N_3799,N_3766);
nor U3917 (N_3917,N_3760,N_3824);
xnor U3918 (N_3918,N_3754,N_3821);
and U3919 (N_3919,N_3881,N_3857);
or U3920 (N_3920,N_3861,N_3817);
and U3921 (N_3921,N_3790,N_3851);
xor U3922 (N_3922,N_3810,N_3811);
xnor U3923 (N_3923,N_3759,N_3835);
or U3924 (N_3924,N_3819,N_3797);
nor U3925 (N_3925,N_3842,N_3854);
xor U3926 (N_3926,N_3789,N_3887);
nand U3927 (N_3927,N_3846,N_3852);
or U3928 (N_3928,N_3795,N_3763);
nand U3929 (N_3929,N_3813,N_3834);
or U3930 (N_3930,N_3879,N_3827);
and U3931 (N_3931,N_3755,N_3828);
and U3932 (N_3932,N_3847,N_3820);
xor U3933 (N_3933,N_3867,N_3805);
nand U3934 (N_3934,N_3770,N_3843);
nand U3935 (N_3935,N_3757,N_3767);
and U3936 (N_3936,N_3856,N_3783);
nand U3937 (N_3937,N_3858,N_3812);
or U3938 (N_3938,N_3764,N_3818);
xor U3939 (N_3939,N_3814,N_3836);
or U3940 (N_3940,N_3869,N_3771);
and U3941 (N_3941,N_3753,N_3793);
or U3942 (N_3942,N_3794,N_3830);
xor U3943 (N_3943,N_3895,N_3750);
nand U3944 (N_3944,N_3871,N_3762);
nor U3945 (N_3945,N_3785,N_3822);
and U3946 (N_3946,N_3845,N_3772);
nor U3947 (N_3947,N_3775,N_3800);
or U3948 (N_3948,N_3751,N_3870);
and U3949 (N_3949,N_3781,N_3862);
or U3950 (N_3950,N_3778,N_3885);
nor U3951 (N_3951,N_3782,N_3876);
and U3952 (N_3952,N_3894,N_3806);
nor U3953 (N_3953,N_3807,N_3899);
and U3954 (N_3954,N_3761,N_3866);
or U3955 (N_3955,N_3892,N_3779);
and U3956 (N_3956,N_3825,N_3863);
nor U3957 (N_3957,N_3808,N_3831);
xnor U3958 (N_3958,N_3773,N_3878);
nor U3959 (N_3959,N_3865,N_3880);
and U3960 (N_3960,N_3777,N_3841);
or U3961 (N_3961,N_3860,N_3889);
nor U3962 (N_3962,N_3874,N_3815);
or U3963 (N_3963,N_3776,N_3796);
nand U3964 (N_3964,N_3788,N_3816);
xor U3965 (N_3965,N_3890,N_3886);
xor U3966 (N_3966,N_3844,N_3803);
nand U3967 (N_3967,N_3802,N_3855);
nor U3968 (N_3968,N_3823,N_3853);
nand U3969 (N_3969,N_3893,N_3837);
nor U3970 (N_3970,N_3826,N_3839);
xor U3971 (N_3971,N_3872,N_3877);
xnor U3972 (N_3972,N_3840,N_3752);
and U3973 (N_3973,N_3765,N_3883);
nand U3974 (N_3974,N_3784,N_3804);
nor U3975 (N_3975,N_3808,N_3751);
and U3976 (N_3976,N_3753,N_3804);
xnor U3977 (N_3977,N_3839,N_3764);
or U3978 (N_3978,N_3783,N_3834);
and U3979 (N_3979,N_3834,N_3798);
or U3980 (N_3980,N_3820,N_3779);
and U3981 (N_3981,N_3873,N_3771);
and U3982 (N_3982,N_3828,N_3863);
xnor U3983 (N_3983,N_3893,N_3758);
nor U3984 (N_3984,N_3866,N_3822);
xor U3985 (N_3985,N_3834,N_3800);
nor U3986 (N_3986,N_3853,N_3820);
and U3987 (N_3987,N_3807,N_3872);
xor U3988 (N_3988,N_3830,N_3893);
nor U3989 (N_3989,N_3757,N_3895);
nand U3990 (N_3990,N_3876,N_3783);
nor U3991 (N_3991,N_3834,N_3812);
and U3992 (N_3992,N_3875,N_3806);
and U3993 (N_3993,N_3891,N_3832);
nand U3994 (N_3994,N_3898,N_3861);
xor U3995 (N_3995,N_3856,N_3819);
nand U3996 (N_3996,N_3893,N_3818);
nor U3997 (N_3997,N_3854,N_3864);
or U3998 (N_3998,N_3835,N_3804);
or U3999 (N_3999,N_3885,N_3883);
or U4000 (N_4000,N_3852,N_3751);
nor U4001 (N_4001,N_3868,N_3856);
or U4002 (N_4002,N_3869,N_3846);
nand U4003 (N_4003,N_3772,N_3865);
nand U4004 (N_4004,N_3897,N_3898);
and U4005 (N_4005,N_3879,N_3870);
and U4006 (N_4006,N_3888,N_3845);
or U4007 (N_4007,N_3895,N_3772);
and U4008 (N_4008,N_3891,N_3879);
nor U4009 (N_4009,N_3773,N_3831);
and U4010 (N_4010,N_3762,N_3892);
or U4011 (N_4011,N_3873,N_3814);
nand U4012 (N_4012,N_3775,N_3771);
xor U4013 (N_4013,N_3883,N_3783);
and U4014 (N_4014,N_3870,N_3753);
nor U4015 (N_4015,N_3895,N_3829);
or U4016 (N_4016,N_3807,N_3785);
nor U4017 (N_4017,N_3899,N_3770);
nand U4018 (N_4018,N_3894,N_3780);
nor U4019 (N_4019,N_3830,N_3810);
or U4020 (N_4020,N_3894,N_3838);
nor U4021 (N_4021,N_3829,N_3855);
nor U4022 (N_4022,N_3836,N_3868);
nand U4023 (N_4023,N_3830,N_3799);
nand U4024 (N_4024,N_3763,N_3755);
nor U4025 (N_4025,N_3882,N_3874);
and U4026 (N_4026,N_3812,N_3822);
nor U4027 (N_4027,N_3836,N_3755);
nand U4028 (N_4028,N_3860,N_3830);
or U4029 (N_4029,N_3869,N_3878);
xnor U4030 (N_4030,N_3760,N_3867);
and U4031 (N_4031,N_3795,N_3876);
and U4032 (N_4032,N_3759,N_3866);
nor U4033 (N_4033,N_3877,N_3816);
nor U4034 (N_4034,N_3772,N_3797);
and U4035 (N_4035,N_3771,N_3783);
or U4036 (N_4036,N_3754,N_3880);
nand U4037 (N_4037,N_3817,N_3831);
or U4038 (N_4038,N_3868,N_3892);
nor U4039 (N_4039,N_3782,N_3849);
xor U4040 (N_4040,N_3817,N_3781);
xor U4041 (N_4041,N_3750,N_3894);
and U4042 (N_4042,N_3786,N_3861);
nand U4043 (N_4043,N_3797,N_3892);
nor U4044 (N_4044,N_3827,N_3771);
nand U4045 (N_4045,N_3806,N_3847);
nand U4046 (N_4046,N_3868,N_3776);
or U4047 (N_4047,N_3764,N_3854);
nand U4048 (N_4048,N_3889,N_3878);
or U4049 (N_4049,N_3804,N_3875);
or U4050 (N_4050,N_3902,N_3958);
or U4051 (N_4051,N_3956,N_3974);
and U4052 (N_4052,N_3912,N_3959);
xnor U4053 (N_4053,N_3917,N_3940);
nand U4054 (N_4054,N_3987,N_3947);
and U4055 (N_4055,N_3934,N_4004);
nand U4056 (N_4056,N_4011,N_3997);
and U4057 (N_4057,N_3944,N_4034);
nand U4058 (N_4058,N_3914,N_3968);
nor U4059 (N_4059,N_4024,N_3954);
or U4060 (N_4060,N_4002,N_4031);
or U4061 (N_4061,N_4030,N_4019);
xor U4062 (N_4062,N_3993,N_4035);
or U4063 (N_4063,N_3932,N_3923);
xnor U4064 (N_4064,N_3901,N_3900);
and U4065 (N_4065,N_4027,N_4015);
and U4066 (N_4066,N_4012,N_3936);
nor U4067 (N_4067,N_3965,N_3949);
and U4068 (N_4068,N_3933,N_3913);
or U4069 (N_4069,N_3966,N_3969);
or U4070 (N_4070,N_3942,N_3990);
and U4071 (N_4071,N_4013,N_3938);
and U4072 (N_4072,N_3907,N_3951);
or U4073 (N_4073,N_3941,N_3935);
or U4074 (N_4074,N_4018,N_3928);
nor U4075 (N_4075,N_3962,N_4045);
nand U4076 (N_4076,N_3981,N_3929);
or U4077 (N_4077,N_3989,N_3915);
nand U4078 (N_4078,N_3952,N_3943);
nand U4079 (N_4079,N_3945,N_4026);
or U4080 (N_4080,N_3973,N_3979);
xor U4081 (N_4081,N_3992,N_4016);
nor U4082 (N_4082,N_3995,N_3909);
xnor U4083 (N_4083,N_3994,N_4001);
and U4084 (N_4084,N_3988,N_3980);
and U4085 (N_4085,N_3921,N_3920);
xnor U4086 (N_4086,N_3927,N_4037);
or U4087 (N_4087,N_3955,N_3904);
xnor U4088 (N_4088,N_4032,N_4033);
xor U4089 (N_4089,N_3976,N_3948);
nor U4090 (N_4090,N_4006,N_3975);
nand U4091 (N_4091,N_4042,N_3916);
nand U4092 (N_4092,N_3957,N_4000);
or U4093 (N_4093,N_3905,N_3960);
nor U4094 (N_4094,N_4007,N_4044);
or U4095 (N_4095,N_3939,N_3972);
nor U4096 (N_4096,N_4041,N_3925);
and U4097 (N_4097,N_3906,N_4025);
nand U4098 (N_4098,N_3924,N_3910);
or U4099 (N_4099,N_3986,N_3999);
and U4100 (N_4100,N_4022,N_3937);
nor U4101 (N_4101,N_3996,N_4008);
nand U4102 (N_4102,N_4038,N_3998);
xnor U4103 (N_4103,N_4039,N_4029);
or U4104 (N_4104,N_4020,N_3953);
xor U4105 (N_4105,N_4014,N_3918);
and U4106 (N_4106,N_3978,N_4028);
nand U4107 (N_4107,N_3991,N_3911);
xnor U4108 (N_4108,N_3984,N_3946);
or U4109 (N_4109,N_4021,N_3903);
nand U4110 (N_4110,N_3983,N_3964);
and U4111 (N_4111,N_3982,N_4023);
xnor U4112 (N_4112,N_4046,N_3970);
xnor U4113 (N_4113,N_4040,N_4003);
and U4114 (N_4114,N_3977,N_3950);
or U4115 (N_4115,N_3931,N_3926);
nor U4116 (N_4116,N_3961,N_3930);
nand U4117 (N_4117,N_4036,N_4017);
nor U4118 (N_4118,N_4047,N_4048);
nor U4119 (N_4119,N_3971,N_3963);
xnor U4120 (N_4120,N_3922,N_4005);
nor U4121 (N_4121,N_3985,N_4043);
nor U4122 (N_4122,N_4009,N_3919);
or U4123 (N_4123,N_4049,N_4010);
and U4124 (N_4124,N_3908,N_3967);
or U4125 (N_4125,N_3957,N_3935);
xor U4126 (N_4126,N_3988,N_3937);
nor U4127 (N_4127,N_3938,N_4046);
or U4128 (N_4128,N_3950,N_3933);
or U4129 (N_4129,N_3986,N_3966);
or U4130 (N_4130,N_3964,N_4006);
nand U4131 (N_4131,N_3917,N_3983);
or U4132 (N_4132,N_3996,N_3920);
or U4133 (N_4133,N_3993,N_3921);
or U4134 (N_4134,N_3934,N_3980);
nand U4135 (N_4135,N_3901,N_4029);
nor U4136 (N_4136,N_3972,N_4046);
and U4137 (N_4137,N_3951,N_3953);
or U4138 (N_4138,N_3904,N_3960);
or U4139 (N_4139,N_4047,N_4017);
or U4140 (N_4140,N_3927,N_3905);
or U4141 (N_4141,N_3921,N_4016);
nor U4142 (N_4142,N_3906,N_4039);
nor U4143 (N_4143,N_4037,N_3998);
xor U4144 (N_4144,N_3985,N_4044);
and U4145 (N_4145,N_4002,N_3903);
xor U4146 (N_4146,N_3905,N_3921);
nor U4147 (N_4147,N_3921,N_3945);
or U4148 (N_4148,N_3992,N_3967);
xor U4149 (N_4149,N_4001,N_3927);
nor U4150 (N_4150,N_3950,N_4007);
xor U4151 (N_4151,N_3984,N_3998);
and U4152 (N_4152,N_3949,N_4030);
nor U4153 (N_4153,N_4036,N_3975);
and U4154 (N_4154,N_4027,N_3984);
and U4155 (N_4155,N_3993,N_4044);
nor U4156 (N_4156,N_3920,N_3912);
or U4157 (N_4157,N_4013,N_4033);
nand U4158 (N_4158,N_4029,N_3940);
xnor U4159 (N_4159,N_3985,N_3918);
xor U4160 (N_4160,N_3994,N_3947);
nand U4161 (N_4161,N_3976,N_3917);
nor U4162 (N_4162,N_3934,N_4002);
nand U4163 (N_4163,N_3948,N_4008);
nand U4164 (N_4164,N_3992,N_3927);
xor U4165 (N_4165,N_3985,N_3948);
nor U4166 (N_4166,N_3931,N_3971);
xor U4167 (N_4167,N_3953,N_3965);
xor U4168 (N_4168,N_4004,N_4024);
nand U4169 (N_4169,N_4027,N_3924);
nor U4170 (N_4170,N_3921,N_4043);
or U4171 (N_4171,N_3915,N_3999);
nor U4172 (N_4172,N_4048,N_3969);
and U4173 (N_4173,N_4013,N_3917);
or U4174 (N_4174,N_4034,N_4000);
nand U4175 (N_4175,N_4021,N_3910);
nor U4176 (N_4176,N_4036,N_3955);
xnor U4177 (N_4177,N_3958,N_3907);
nand U4178 (N_4178,N_4009,N_3940);
nor U4179 (N_4179,N_3918,N_3919);
xnor U4180 (N_4180,N_3998,N_4042);
nor U4181 (N_4181,N_4043,N_3904);
nand U4182 (N_4182,N_3954,N_4027);
and U4183 (N_4183,N_4044,N_3913);
and U4184 (N_4184,N_4003,N_4036);
xnor U4185 (N_4185,N_3915,N_3920);
or U4186 (N_4186,N_3928,N_3983);
nor U4187 (N_4187,N_3997,N_3912);
and U4188 (N_4188,N_4041,N_4039);
and U4189 (N_4189,N_3998,N_4015);
nor U4190 (N_4190,N_3972,N_3991);
or U4191 (N_4191,N_3967,N_3927);
nor U4192 (N_4192,N_4027,N_3993);
or U4193 (N_4193,N_4037,N_4019);
nor U4194 (N_4194,N_3977,N_3994);
xnor U4195 (N_4195,N_3966,N_4009);
xnor U4196 (N_4196,N_4030,N_4011);
nor U4197 (N_4197,N_3940,N_3949);
and U4198 (N_4198,N_3954,N_4034);
and U4199 (N_4199,N_4013,N_3900);
nand U4200 (N_4200,N_4156,N_4142);
or U4201 (N_4201,N_4059,N_4159);
and U4202 (N_4202,N_4112,N_4052);
nand U4203 (N_4203,N_4109,N_4095);
or U4204 (N_4204,N_4135,N_4055);
nor U4205 (N_4205,N_4165,N_4153);
nor U4206 (N_4206,N_4140,N_4166);
nand U4207 (N_4207,N_4082,N_4189);
nor U4208 (N_4208,N_4163,N_4193);
xnor U4209 (N_4209,N_4074,N_4057);
and U4210 (N_4210,N_4148,N_4179);
and U4211 (N_4211,N_4102,N_4183);
nor U4212 (N_4212,N_4174,N_4161);
nand U4213 (N_4213,N_4185,N_4155);
and U4214 (N_4214,N_4107,N_4187);
nand U4215 (N_4215,N_4176,N_4113);
and U4216 (N_4216,N_4061,N_4136);
xnor U4217 (N_4217,N_4089,N_4067);
nor U4218 (N_4218,N_4171,N_4103);
nand U4219 (N_4219,N_4180,N_4170);
xor U4220 (N_4220,N_4162,N_4194);
or U4221 (N_4221,N_4118,N_4195);
and U4222 (N_4222,N_4115,N_4092);
xor U4223 (N_4223,N_4110,N_4181);
or U4224 (N_4224,N_4122,N_4128);
or U4225 (N_4225,N_4056,N_4066);
nor U4226 (N_4226,N_4150,N_4152);
and U4227 (N_4227,N_4081,N_4139);
nor U4228 (N_4228,N_4087,N_4063);
nand U4229 (N_4229,N_4116,N_4084);
and U4230 (N_4230,N_4091,N_4164);
and U4231 (N_4231,N_4071,N_4094);
or U4232 (N_4232,N_4132,N_4085);
and U4233 (N_4233,N_4099,N_4121);
nand U4234 (N_4234,N_4124,N_4178);
nand U4235 (N_4235,N_4138,N_4131);
and U4236 (N_4236,N_4098,N_4086);
xor U4237 (N_4237,N_4054,N_4062);
and U4238 (N_4238,N_4114,N_4070);
and U4239 (N_4239,N_4129,N_4111);
nand U4240 (N_4240,N_4072,N_4196);
or U4241 (N_4241,N_4127,N_4119);
nand U4242 (N_4242,N_4173,N_4141);
or U4243 (N_4243,N_4151,N_4053);
and U4244 (N_4244,N_4147,N_4075);
nand U4245 (N_4245,N_4149,N_4058);
xnor U4246 (N_4246,N_4133,N_4096);
and U4247 (N_4247,N_4120,N_4167);
nor U4248 (N_4248,N_4190,N_4175);
xnor U4249 (N_4249,N_4106,N_4100);
xnor U4250 (N_4250,N_4088,N_4146);
nand U4251 (N_4251,N_4199,N_4191);
and U4252 (N_4252,N_4123,N_4064);
and U4253 (N_4253,N_4143,N_4117);
xnor U4254 (N_4254,N_4101,N_4169);
or U4255 (N_4255,N_4080,N_4090);
or U4256 (N_4256,N_4186,N_4078);
and U4257 (N_4257,N_4154,N_4160);
nand U4258 (N_4258,N_4050,N_4126);
nor U4259 (N_4259,N_4083,N_4097);
or U4260 (N_4260,N_4073,N_4198);
or U4261 (N_4261,N_4108,N_4068);
or U4262 (N_4262,N_4184,N_4192);
nor U4263 (N_4263,N_4093,N_4125);
or U4264 (N_4264,N_4158,N_4172);
and U4265 (N_4265,N_4105,N_4197);
and U4266 (N_4266,N_4076,N_4079);
and U4267 (N_4267,N_4182,N_4104);
and U4268 (N_4268,N_4188,N_4051);
nor U4269 (N_4269,N_4137,N_4130);
nand U4270 (N_4270,N_4144,N_4177);
and U4271 (N_4271,N_4157,N_4060);
nand U4272 (N_4272,N_4069,N_4145);
or U4273 (N_4273,N_4065,N_4077);
xor U4274 (N_4274,N_4168,N_4134);
or U4275 (N_4275,N_4091,N_4118);
or U4276 (N_4276,N_4084,N_4130);
nand U4277 (N_4277,N_4126,N_4097);
or U4278 (N_4278,N_4076,N_4132);
xnor U4279 (N_4279,N_4190,N_4127);
nand U4280 (N_4280,N_4098,N_4159);
nor U4281 (N_4281,N_4165,N_4183);
nand U4282 (N_4282,N_4176,N_4189);
or U4283 (N_4283,N_4164,N_4142);
xnor U4284 (N_4284,N_4176,N_4111);
and U4285 (N_4285,N_4126,N_4199);
xnor U4286 (N_4286,N_4130,N_4071);
or U4287 (N_4287,N_4077,N_4153);
nand U4288 (N_4288,N_4127,N_4075);
nand U4289 (N_4289,N_4091,N_4101);
xnor U4290 (N_4290,N_4152,N_4061);
nand U4291 (N_4291,N_4189,N_4129);
xor U4292 (N_4292,N_4151,N_4172);
xor U4293 (N_4293,N_4161,N_4085);
xnor U4294 (N_4294,N_4096,N_4064);
nand U4295 (N_4295,N_4091,N_4085);
nor U4296 (N_4296,N_4054,N_4176);
and U4297 (N_4297,N_4056,N_4119);
or U4298 (N_4298,N_4165,N_4156);
nand U4299 (N_4299,N_4108,N_4054);
or U4300 (N_4300,N_4196,N_4163);
and U4301 (N_4301,N_4104,N_4193);
xnor U4302 (N_4302,N_4117,N_4122);
nand U4303 (N_4303,N_4085,N_4186);
nor U4304 (N_4304,N_4082,N_4166);
or U4305 (N_4305,N_4186,N_4053);
nor U4306 (N_4306,N_4172,N_4070);
nor U4307 (N_4307,N_4058,N_4179);
or U4308 (N_4308,N_4085,N_4090);
nor U4309 (N_4309,N_4181,N_4159);
or U4310 (N_4310,N_4051,N_4072);
nand U4311 (N_4311,N_4199,N_4053);
xor U4312 (N_4312,N_4093,N_4101);
xnor U4313 (N_4313,N_4102,N_4079);
or U4314 (N_4314,N_4091,N_4114);
xnor U4315 (N_4315,N_4137,N_4141);
and U4316 (N_4316,N_4057,N_4120);
xnor U4317 (N_4317,N_4171,N_4141);
and U4318 (N_4318,N_4169,N_4069);
and U4319 (N_4319,N_4176,N_4117);
and U4320 (N_4320,N_4081,N_4105);
or U4321 (N_4321,N_4197,N_4093);
and U4322 (N_4322,N_4065,N_4131);
and U4323 (N_4323,N_4190,N_4126);
xnor U4324 (N_4324,N_4129,N_4101);
nor U4325 (N_4325,N_4091,N_4170);
nand U4326 (N_4326,N_4145,N_4111);
nand U4327 (N_4327,N_4101,N_4088);
or U4328 (N_4328,N_4181,N_4111);
and U4329 (N_4329,N_4133,N_4179);
and U4330 (N_4330,N_4083,N_4085);
or U4331 (N_4331,N_4146,N_4091);
or U4332 (N_4332,N_4170,N_4109);
and U4333 (N_4333,N_4199,N_4109);
nand U4334 (N_4334,N_4137,N_4194);
or U4335 (N_4335,N_4091,N_4128);
nor U4336 (N_4336,N_4197,N_4126);
and U4337 (N_4337,N_4133,N_4102);
xor U4338 (N_4338,N_4079,N_4189);
xnor U4339 (N_4339,N_4073,N_4187);
or U4340 (N_4340,N_4168,N_4091);
nor U4341 (N_4341,N_4099,N_4132);
and U4342 (N_4342,N_4052,N_4187);
and U4343 (N_4343,N_4092,N_4177);
nand U4344 (N_4344,N_4078,N_4160);
and U4345 (N_4345,N_4175,N_4153);
or U4346 (N_4346,N_4124,N_4157);
and U4347 (N_4347,N_4163,N_4148);
nand U4348 (N_4348,N_4139,N_4067);
or U4349 (N_4349,N_4093,N_4162);
nor U4350 (N_4350,N_4349,N_4336);
or U4351 (N_4351,N_4209,N_4322);
nor U4352 (N_4352,N_4248,N_4228);
nand U4353 (N_4353,N_4343,N_4217);
and U4354 (N_4354,N_4263,N_4221);
nand U4355 (N_4355,N_4331,N_4220);
and U4356 (N_4356,N_4272,N_4307);
nor U4357 (N_4357,N_4265,N_4308);
nor U4358 (N_4358,N_4313,N_4269);
xor U4359 (N_4359,N_4235,N_4280);
nand U4360 (N_4360,N_4282,N_4232);
or U4361 (N_4361,N_4320,N_4318);
nand U4362 (N_4362,N_4294,N_4287);
nor U4363 (N_4363,N_4203,N_4296);
nor U4364 (N_4364,N_4305,N_4236);
nand U4365 (N_4365,N_4309,N_4346);
xor U4366 (N_4366,N_4267,N_4335);
or U4367 (N_4367,N_4243,N_4348);
and U4368 (N_4368,N_4241,N_4202);
and U4369 (N_4369,N_4226,N_4326);
nand U4370 (N_4370,N_4225,N_4330);
or U4371 (N_4371,N_4254,N_4339);
or U4372 (N_4372,N_4215,N_4285);
xor U4373 (N_4373,N_4288,N_4275);
or U4374 (N_4374,N_4257,N_4242);
nor U4375 (N_4375,N_4259,N_4207);
nor U4376 (N_4376,N_4312,N_4289);
xor U4377 (N_4377,N_4246,N_4301);
and U4378 (N_4378,N_4344,N_4252);
and U4379 (N_4379,N_4251,N_4237);
nor U4380 (N_4380,N_4214,N_4260);
nor U4381 (N_4381,N_4227,N_4204);
nand U4382 (N_4382,N_4291,N_4321);
nand U4383 (N_4383,N_4333,N_4218);
and U4384 (N_4384,N_4281,N_4276);
and U4385 (N_4385,N_4223,N_4338);
or U4386 (N_4386,N_4270,N_4315);
nand U4387 (N_4387,N_4206,N_4302);
and U4388 (N_4388,N_4304,N_4286);
and U4389 (N_4389,N_4244,N_4211);
nand U4390 (N_4390,N_4323,N_4253);
xor U4391 (N_4391,N_4210,N_4201);
xor U4392 (N_4392,N_4299,N_4306);
nand U4393 (N_4393,N_4311,N_4293);
and U4394 (N_4394,N_4258,N_4222);
nor U4395 (N_4395,N_4324,N_4229);
and U4396 (N_4396,N_4327,N_4250);
xor U4397 (N_4397,N_4239,N_4329);
and U4398 (N_4398,N_4234,N_4310);
nand U4399 (N_4399,N_4255,N_4303);
nor U4400 (N_4400,N_4317,N_4278);
and U4401 (N_4401,N_4231,N_4245);
nor U4402 (N_4402,N_4249,N_4262);
and U4403 (N_4403,N_4297,N_4328);
xnor U4404 (N_4404,N_4298,N_4233);
nor U4405 (N_4405,N_4316,N_4216);
nand U4406 (N_4406,N_4332,N_4342);
xnor U4407 (N_4407,N_4271,N_4224);
nand U4408 (N_4408,N_4238,N_4295);
nand U4409 (N_4409,N_4290,N_4314);
xnor U4410 (N_4410,N_4219,N_4208);
nor U4411 (N_4411,N_4340,N_4261);
and U4412 (N_4412,N_4268,N_4212);
nor U4413 (N_4413,N_4273,N_4337);
xnor U4414 (N_4414,N_4334,N_4300);
nor U4415 (N_4415,N_4283,N_4274);
nor U4416 (N_4416,N_4256,N_4319);
nand U4417 (N_4417,N_4284,N_4345);
xor U4418 (N_4418,N_4266,N_4200);
or U4419 (N_4419,N_4247,N_4213);
and U4420 (N_4420,N_4277,N_4292);
or U4421 (N_4421,N_4264,N_4347);
xnor U4422 (N_4422,N_4240,N_4230);
nor U4423 (N_4423,N_4279,N_4325);
nor U4424 (N_4424,N_4205,N_4341);
nand U4425 (N_4425,N_4277,N_4286);
and U4426 (N_4426,N_4267,N_4244);
or U4427 (N_4427,N_4261,N_4257);
xor U4428 (N_4428,N_4263,N_4226);
and U4429 (N_4429,N_4314,N_4253);
and U4430 (N_4430,N_4307,N_4207);
xor U4431 (N_4431,N_4316,N_4227);
or U4432 (N_4432,N_4272,N_4267);
nand U4433 (N_4433,N_4314,N_4210);
and U4434 (N_4434,N_4248,N_4282);
or U4435 (N_4435,N_4314,N_4332);
xor U4436 (N_4436,N_4320,N_4208);
nand U4437 (N_4437,N_4250,N_4216);
nor U4438 (N_4438,N_4236,N_4315);
nor U4439 (N_4439,N_4328,N_4230);
or U4440 (N_4440,N_4200,N_4214);
and U4441 (N_4441,N_4204,N_4344);
nor U4442 (N_4442,N_4216,N_4238);
xor U4443 (N_4443,N_4231,N_4295);
nand U4444 (N_4444,N_4291,N_4212);
nor U4445 (N_4445,N_4310,N_4259);
xnor U4446 (N_4446,N_4302,N_4254);
or U4447 (N_4447,N_4294,N_4300);
nand U4448 (N_4448,N_4240,N_4347);
and U4449 (N_4449,N_4316,N_4242);
and U4450 (N_4450,N_4202,N_4279);
nand U4451 (N_4451,N_4219,N_4321);
xor U4452 (N_4452,N_4338,N_4349);
xor U4453 (N_4453,N_4263,N_4304);
and U4454 (N_4454,N_4338,N_4239);
nor U4455 (N_4455,N_4267,N_4222);
or U4456 (N_4456,N_4341,N_4236);
and U4457 (N_4457,N_4220,N_4310);
xnor U4458 (N_4458,N_4265,N_4259);
nand U4459 (N_4459,N_4273,N_4221);
or U4460 (N_4460,N_4277,N_4328);
or U4461 (N_4461,N_4284,N_4242);
xor U4462 (N_4462,N_4302,N_4273);
nand U4463 (N_4463,N_4203,N_4202);
nor U4464 (N_4464,N_4274,N_4321);
nand U4465 (N_4465,N_4244,N_4239);
nor U4466 (N_4466,N_4241,N_4283);
nand U4467 (N_4467,N_4285,N_4218);
and U4468 (N_4468,N_4222,N_4245);
and U4469 (N_4469,N_4257,N_4200);
and U4470 (N_4470,N_4287,N_4216);
nor U4471 (N_4471,N_4321,N_4228);
xor U4472 (N_4472,N_4266,N_4282);
and U4473 (N_4473,N_4343,N_4253);
nand U4474 (N_4474,N_4255,N_4290);
nand U4475 (N_4475,N_4243,N_4250);
and U4476 (N_4476,N_4302,N_4259);
xnor U4477 (N_4477,N_4334,N_4337);
nor U4478 (N_4478,N_4215,N_4345);
and U4479 (N_4479,N_4311,N_4245);
and U4480 (N_4480,N_4334,N_4347);
and U4481 (N_4481,N_4276,N_4346);
nor U4482 (N_4482,N_4249,N_4295);
or U4483 (N_4483,N_4230,N_4224);
and U4484 (N_4484,N_4255,N_4262);
and U4485 (N_4485,N_4304,N_4235);
nor U4486 (N_4486,N_4346,N_4313);
and U4487 (N_4487,N_4239,N_4263);
nor U4488 (N_4488,N_4233,N_4334);
nand U4489 (N_4489,N_4335,N_4349);
nand U4490 (N_4490,N_4277,N_4250);
nor U4491 (N_4491,N_4274,N_4239);
nand U4492 (N_4492,N_4338,N_4253);
and U4493 (N_4493,N_4345,N_4332);
xor U4494 (N_4494,N_4328,N_4201);
xor U4495 (N_4495,N_4346,N_4342);
and U4496 (N_4496,N_4252,N_4316);
or U4497 (N_4497,N_4281,N_4347);
nor U4498 (N_4498,N_4205,N_4256);
or U4499 (N_4499,N_4308,N_4258);
nor U4500 (N_4500,N_4414,N_4444);
or U4501 (N_4501,N_4433,N_4431);
nor U4502 (N_4502,N_4432,N_4429);
and U4503 (N_4503,N_4422,N_4360);
nor U4504 (N_4504,N_4495,N_4415);
xor U4505 (N_4505,N_4378,N_4487);
and U4506 (N_4506,N_4483,N_4367);
nor U4507 (N_4507,N_4478,N_4407);
and U4508 (N_4508,N_4498,N_4477);
or U4509 (N_4509,N_4395,N_4370);
nand U4510 (N_4510,N_4399,N_4383);
xnor U4511 (N_4511,N_4352,N_4369);
nand U4512 (N_4512,N_4458,N_4470);
xnor U4513 (N_4513,N_4366,N_4455);
and U4514 (N_4514,N_4394,N_4493);
nand U4515 (N_4515,N_4371,N_4358);
nand U4516 (N_4516,N_4368,N_4488);
nor U4517 (N_4517,N_4476,N_4382);
or U4518 (N_4518,N_4460,N_4441);
nand U4519 (N_4519,N_4452,N_4474);
and U4520 (N_4520,N_4463,N_4428);
nor U4521 (N_4521,N_4438,N_4486);
or U4522 (N_4522,N_4404,N_4381);
and U4523 (N_4523,N_4372,N_4461);
and U4524 (N_4524,N_4393,N_4386);
or U4525 (N_4525,N_4475,N_4396);
or U4526 (N_4526,N_4398,N_4354);
or U4527 (N_4527,N_4436,N_4411);
nand U4528 (N_4528,N_4365,N_4443);
nor U4529 (N_4529,N_4466,N_4362);
or U4530 (N_4530,N_4397,N_4419);
and U4531 (N_4531,N_4388,N_4425);
and U4532 (N_4532,N_4380,N_4359);
and U4533 (N_4533,N_4447,N_4387);
nor U4534 (N_4534,N_4453,N_4465);
xor U4535 (N_4535,N_4364,N_4412);
or U4536 (N_4536,N_4473,N_4405);
and U4537 (N_4537,N_4353,N_4499);
and U4538 (N_4538,N_4408,N_4418);
xor U4539 (N_4539,N_4430,N_4469);
or U4540 (N_4540,N_4435,N_4451);
nand U4541 (N_4541,N_4391,N_4363);
nand U4542 (N_4542,N_4417,N_4472);
nand U4543 (N_4543,N_4491,N_4445);
nor U4544 (N_4544,N_4497,N_4385);
xnor U4545 (N_4545,N_4374,N_4356);
xnor U4546 (N_4546,N_4423,N_4442);
or U4547 (N_4547,N_4457,N_4357);
xnor U4548 (N_4548,N_4492,N_4350);
or U4549 (N_4549,N_4448,N_4454);
nor U4550 (N_4550,N_4390,N_4462);
nand U4551 (N_4551,N_4484,N_4421);
xor U4552 (N_4552,N_4389,N_4379);
nand U4553 (N_4553,N_4489,N_4409);
nand U4554 (N_4554,N_4494,N_4434);
nor U4555 (N_4555,N_4449,N_4424);
nand U4556 (N_4556,N_4361,N_4373);
nand U4557 (N_4557,N_4496,N_4446);
or U4558 (N_4558,N_4490,N_4482);
or U4559 (N_4559,N_4420,N_4402);
nand U4560 (N_4560,N_4376,N_4450);
and U4561 (N_4561,N_4471,N_4355);
nand U4562 (N_4562,N_4427,N_4384);
nand U4563 (N_4563,N_4479,N_4401);
and U4564 (N_4564,N_4400,N_4459);
xnor U4565 (N_4565,N_4406,N_4426);
or U4566 (N_4566,N_4481,N_4456);
or U4567 (N_4567,N_4392,N_4468);
or U4568 (N_4568,N_4485,N_4437);
or U4569 (N_4569,N_4480,N_4467);
or U4570 (N_4570,N_4413,N_4403);
and U4571 (N_4571,N_4375,N_4410);
or U4572 (N_4572,N_4416,N_4351);
nor U4573 (N_4573,N_4439,N_4440);
nand U4574 (N_4574,N_4377,N_4464);
nand U4575 (N_4575,N_4378,N_4477);
nand U4576 (N_4576,N_4361,N_4440);
xor U4577 (N_4577,N_4429,N_4475);
xnor U4578 (N_4578,N_4426,N_4485);
nand U4579 (N_4579,N_4403,N_4371);
or U4580 (N_4580,N_4493,N_4478);
and U4581 (N_4581,N_4386,N_4440);
and U4582 (N_4582,N_4361,N_4471);
xor U4583 (N_4583,N_4395,N_4412);
nand U4584 (N_4584,N_4395,N_4430);
and U4585 (N_4585,N_4437,N_4471);
or U4586 (N_4586,N_4360,N_4432);
nor U4587 (N_4587,N_4483,N_4393);
and U4588 (N_4588,N_4433,N_4495);
or U4589 (N_4589,N_4453,N_4366);
and U4590 (N_4590,N_4388,N_4474);
nor U4591 (N_4591,N_4376,N_4425);
nor U4592 (N_4592,N_4434,N_4378);
and U4593 (N_4593,N_4352,N_4353);
and U4594 (N_4594,N_4447,N_4444);
xor U4595 (N_4595,N_4464,N_4449);
xor U4596 (N_4596,N_4452,N_4472);
and U4597 (N_4597,N_4455,N_4419);
nor U4598 (N_4598,N_4433,N_4483);
or U4599 (N_4599,N_4428,N_4457);
nor U4600 (N_4600,N_4439,N_4488);
xnor U4601 (N_4601,N_4351,N_4393);
nor U4602 (N_4602,N_4407,N_4453);
xor U4603 (N_4603,N_4466,N_4467);
xor U4604 (N_4604,N_4457,N_4473);
nor U4605 (N_4605,N_4400,N_4363);
and U4606 (N_4606,N_4453,N_4481);
nor U4607 (N_4607,N_4490,N_4380);
nor U4608 (N_4608,N_4383,N_4413);
xor U4609 (N_4609,N_4369,N_4435);
or U4610 (N_4610,N_4466,N_4358);
and U4611 (N_4611,N_4359,N_4368);
xnor U4612 (N_4612,N_4429,N_4411);
and U4613 (N_4613,N_4397,N_4449);
nor U4614 (N_4614,N_4403,N_4468);
or U4615 (N_4615,N_4482,N_4421);
xnor U4616 (N_4616,N_4471,N_4466);
and U4617 (N_4617,N_4408,N_4438);
or U4618 (N_4618,N_4401,N_4360);
and U4619 (N_4619,N_4428,N_4365);
or U4620 (N_4620,N_4389,N_4460);
nor U4621 (N_4621,N_4430,N_4490);
and U4622 (N_4622,N_4494,N_4382);
or U4623 (N_4623,N_4456,N_4418);
nand U4624 (N_4624,N_4483,N_4355);
xnor U4625 (N_4625,N_4371,N_4387);
nor U4626 (N_4626,N_4377,N_4403);
nand U4627 (N_4627,N_4401,N_4374);
xor U4628 (N_4628,N_4471,N_4480);
and U4629 (N_4629,N_4392,N_4439);
or U4630 (N_4630,N_4365,N_4488);
and U4631 (N_4631,N_4470,N_4443);
or U4632 (N_4632,N_4394,N_4385);
and U4633 (N_4633,N_4449,N_4452);
and U4634 (N_4634,N_4356,N_4353);
and U4635 (N_4635,N_4468,N_4477);
or U4636 (N_4636,N_4477,N_4458);
and U4637 (N_4637,N_4376,N_4463);
nand U4638 (N_4638,N_4443,N_4361);
nor U4639 (N_4639,N_4478,N_4372);
nor U4640 (N_4640,N_4488,N_4380);
or U4641 (N_4641,N_4462,N_4391);
nor U4642 (N_4642,N_4490,N_4463);
nand U4643 (N_4643,N_4445,N_4466);
nand U4644 (N_4644,N_4410,N_4475);
and U4645 (N_4645,N_4399,N_4438);
nor U4646 (N_4646,N_4415,N_4354);
or U4647 (N_4647,N_4481,N_4411);
and U4648 (N_4648,N_4441,N_4473);
xnor U4649 (N_4649,N_4391,N_4357);
nand U4650 (N_4650,N_4536,N_4538);
or U4651 (N_4651,N_4644,N_4518);
or U4652 (N_4652,N_4539,N_4643);
nor U4653 (N_4653,N_4515,N_4524);
xnor U4654 (N_4654,N_4527,N_4613);
xor U4655 (N_4655,N_4562,N_4555);
xor U4656 (N_4656,N_4566,N_4597);
xor U4657 (N_4657,N_4581,N_4501);
or U4658 (N_4658,N_4530,N_4605);
nor U4659 (N_4659,N_4565,N_4535);
nor U4660 (N_4660,N_4585,N_4507);
or U4661 (N_4661,N_4573,N_4604);
nand U4662 (N_4662,N_4564,N_4598);
or U4663 (N_4663,N_4640,N_4574);
nand U4664 (N_4664,N_4533,N_4624);
nor U4665 (N_4665,N_4645,N_4600);
xnor U4666 (N_4666,N_4607,N_4554);
or U4667 (N_4667,N_4569,N_4578);
xnor U4668 (N_4668,N_4608,N_4638);
or U4669 (N_4669,N_4526,N_4572);
nor U4670 (N_4670,N_4577,N_4513);
nand U4671 (N_4671,N_4519,N_4629);
or U4672 (N_4672,N_4642,N_4571);
nand U4673 (N_4673,N_4529,N_4522);
nor U4674 (N_4674,N_4512,N_4549);
nand U4675 (N_4675,N_4545,N_4619);
nand U4676 (N_4676,N_4556,N_4633);
nand U4677 (N_4677,N_4599,N_4552);
and U4678 (N_4678,N_4550,N_4579);
nor U4679 (N_4679,N_4537,N_4588);
xnor U4680 (N_4680,N_4591,N_4614);
or U4681 (N_4681,N_4531,N_4587);
nand U4682 (N_4682,N_4502,N_4617);
nand U4683 (N_4683,N_4622,N_4632);
xor U4684 (N_4684,N_4611,N_4517);
xor U4685 (N_4685,N_4627,N_4563);
and U4686 (N_4686,N_4557,N_4506);
or U4687 (N_4687,N_4553,N_4561);
xnor U4688 (N_4688,N_4603,N_4635);
xnor U4689 (N_4689,N_4602,N_4543);
nand U4690 (N_4690,N_4631,N_4523);
or U4691 (N_4691,N_4589,N_4510);
xnor U4692 (N_4692,N_4628,N_4504);
nand U4693 (N_4693,N_4647,N_4509);
nor U4694 (N_4694,N_4544,N_4595);
nand U4695 (N_4695,N_4606,N_4596);
and U4696 (N_4696,N_4505,N_4583);
and U4697 (N_4697,N_4639,N_4500);
or U4698 (N_4698,N_4648,N_4503);
nand U4699 (N_4699,N_4516,N_4520);
nor U4700 (N_4700,N_4528,N_4594);
and U4701 (N_4701,N_4586,N_4525);
nor U4702 (N_4702,N_4630,N_4621);
and U4703 (N_4703,N_4612,N_4568);
or U4704 (N_4704,N_4514,N_4576);
and U4705 (N_4705,N_4534,N_4551);
nand U4706 (N_4706,N_4570,N_4626);
nand U4707 (N_4707,N_4615,N_4616);
nor U4708 (N_4708,N_4540,N_4580);
nand U4709 (N_4709,N_4521,N_4637);
nand U4710 (N_4710,N_4623,N_4508);
nor U4711 (N_4711,N_4559,N_4634);
or U4712 (N_4712,N_4582,N_4641);
nand U4713 (N_4713,N_4584,N_4601);
nor U4714 (N_4714,N_4511,N_4532);
nand U4715 (N_4715,N_4542,N_4610);
nor U4716 (N_4716,N_4546,N_4590);
nand U4717 (N_4717,N_4548,N_4547);
or U4718 (N_4718,N_4625,N_4618);
nor U4719 (N_4719,N_4567,N_4649);
or U4720 (N_4720,N_4646,N_4541);
or U4721 (N_4721,N_4609,N_4636);
and U4722 (N_4722,N_4575,N_4592);
nor U4723 (N_4723,N_4558,N_4620);
and U4724 (N_4724,N_4593,N_4560);
and U4725 (N_4725,N_4627,N_4522);
nor U4726 (N_4726,N_4525,N_4523);
and U4727 (N_4727,N_4547,N_4546);
xor U4728 (N_4728,N_4640,N_4644);
or U4729 (N_4729,N_4509,N_4573);
nor U4730 (N_4730,N_4589,N_4514);
and U4731 (N_4731,N_4635,N_4552);
nor U4732 (N_4732,N_4647,N_4576);
nand U4733 (N_4733,N_4544,N_4523);
or U4734 (N_4734,N_4644,N_4610);
and U4735 (N_4735,N_4546,N_4531);
nor U4736 (N_4736,N_4566,N_4628);
xnor U4737 (N_4737,N_4508,N_4603);
xor U4738 (N_4738,N_4548,N_4641);
xor U4739 (N_4739,N_4502,N_4503);
and U4740 (N_4740,N_4518,N_4611);
xor U4741 (N_4741,N_4538,N_4565);
nor U4742 (N_4742,N_4623,N_4522);
xor U4743 (N_4743,N_4525,N_4541);
nor U4744 (N_4744,N_4615,N_4585);
nand U4745 (N_4745,N_4604,N_4521);
nand U4746 (N_4746,N_4537,N_4524);
xnor U4747 (N_4747,N_4599,N_4583);
or U4748 (N_4748,N_4626,N_4521);
nor U4749 (N_4749,N_4502,N_4596);
xor U4750 (N_4750,N_4547,N_4575);
and U4751 (N_4751,N_4542,N_4545);
and U4752 (N_4752,N_4627,N_4611);
nor U4753 (N_4753,N_4610,N_4573);
nor U4754 (N_4754,N_4553,N_4565);
xor U4755 (N_4755,N_4636,N_4537);
nor U4756 (N_4756,N_4597,N_4649);
or U4757 (N_4757,N_4511,N_4519);
and U4758 (N_4758,N_4504,N_4569);
nand U4759 (N_4759,N_4634,N_4501);
and U4760 (N_4760,N_4623,N_4509);
nor U4761 (N_4761,N_4628,N_4538);
xnor U4762 (N_4762,N_4572,N_4603);
nand U4763 (N_4763,N_4578,N_4649);
nor U4764 (N_4764,N_4505,N_4561);
nor U4765 (N_4765,N_4592,N_4522);
or U4766 (N_4766,N_4641,N_4639);
or U4767 (N_4767,N_4561,N_4646);
or U4768 (N_4768,N_4520,N_4630);
or U4769 (N_4769,N_4561,N_4529);
and U4770 (N_4770,N_4539,N_4510);
nor U4771 (N_4771,N_4508,N_4509);
or U4772 (N_4772,N_4628,N_4630);
and U4773 (N_4773,N_4579,N_4507);
nand U4774 (N_4774,N_4543,N_4600);
or U4775 (N_4775,N_4549,N_4628);
and U4776 (N_4776,N_4518,N_4594);
or U4777 (N_4777,N_4574,N_4594);
nor U4778 (N_4778,N_4606,N_4615);
or U4779 (N_4779,N_4514,N_4513);
or U4780 (N_4780,N_4575,N_4603);
or U4781 (N_4781,N_4610,N_4521);
or U4782 (N_4782,N_4621,N_4581);
nand U4783 (N_4783,N_4644,N_4645);
or U4784 (N_4784,N_4584,N_4627);
xor U4785 (N_4785,N_4596,N_4645);
nand U4786 (N_4786,N_4623,N_4527);
xnor U4787 (N_4787,N_4589,N_4530);
and U4788 (N_4788,N_4578,N_4614);
nor U4789 (N_4789,N_4564,N_4612);
nand U4790 (N_4790,N_4600,N_4572);
xor U4791 (N_4791,N_4586,N_4561);
nor U4792 (N_4792,N_4549,N_4585);
xor U4793 (N_4793,N_4599,N_4512);
or U4794 (N_4794,N_4642,N_4566);
nor U4795 (N_4795,N_4591,N_4642);
xnor U4796 (N_4796,N_4611,N_4623);
xnor U4797 (N_4797,N_4523,N_4546);
or U4798 (N_4798,N_4524,N_4561);
xor U4799 (N_4799,N_4616,N_4524);
and U4800 (N_4800,N_4788,N_4660);
and U4801 (N_4801,N_4736,N_4737);
nand U4802 (N_4802,N_4674,N_4652);
nand U4803 (N_4803,N_4794,N_4760);
nand U4804 (N_4804,N_4738,N_4783);
nand U4805 (N_4805,N_4706,N_4779);
xor U4806 (N_4806,N_4755,N_4727);
nand U4807 (N_4807,N_4735,N_4740);
nand U4808 (N_4808,N_4709,N_4792);
or U4809 (N_4809,N_4669,N_4683);
nor U4810 (N_4810,N_4711,N_4656);
and U4811 (N_4811,N_4784,N_4702);
or U4812 (N_4812,N_4797,N_4679);
or U4813 (N_4813,N_4681,N_4745);
xnor U4814 (N_4814,N_4682,N_4742);
xor U4815 (N_4815,N_4690,N_4778);
and U4816 (N_4816,N_4729,N_4724);
nor U4817 (N_4817,N_4734,N_4771);
xnor U4818 (N_4818,N_4657,N_4731);
and U4819 (N_4819,N_4654,N_4667);
nand U4820 (N_4820,N_4758,N_4651);
and U4821 (N_4821,N_4671,N_4685);
nand U4822 (N_4822,N_4746,N_4785);
nand U4823 (N_4823,N_4700,N_4664);
nand U4824 (N_4824,N_4732,N_4678);
nor U4825 (N_4825,N_4789,N_4663);
and U4826 (N_4826,N_4680,N_4676);
xnor U4827 (N_4827,N_4759,N_4790);
nor U4828 (N_4828,N_4672,N_4666);
xnor U4829 (N_4829,N_4753,N_4761);
xnor U4830 (N_4830,N_4775,N_4741);
nor U4831 (N_4831,N_4749,N_4787);
nand U4832 (N_4832,N_4768,N_4744);
and U4833 (N_4833,N_4733,N_4692);
nand U4834 (N_4834,N_4723,N_4747);
xor U4835 (N_4835,N_4714,N_4688);
nand U4836 (N_4836,N_4770,N_4721);
and U4837 (N_4837,N_4748,N_4776);
nand U4838 (N_4838,N_4751,N_4756);
nand U4839 (N_4839,N_4705,N_4754);
nand U4840 (N_4840,N_4693,N_4710);
and U4841 (N_4841,N_4718,N_4726);
or U4842 (N_4842,N_4673,N_4708);
and U4843 (N_4843,N_4655,N_4782);
and U4844 (N_4844,N_4791,N_4798);
or U4845 (N_4845,N_4716,N_4684);
or U4846 (N_4846,N_4717,N_4777);
or U4847 (N_4847,N_4774,N_4765);
xor U4848 (N_4848,N_4668,N_4739);
and U4849 (N_4849,N_4712,N_4725);
or U4850 (N_4850,N_4695,N_4665);
or U4851 (N_4851,N_4764,N_4689);
and U4852 (N_4852,N_4757,N_4769);
nor U4853 (N_4853,N_4661,N_4730);
or U4854 (N_4854,N_4691,N_4767);
and U4855 (N_4855,N_4743,N_4675);
and U4856 (N_4856,N_4658,N_4780);
and U4857 (N_4857,N_4795,N_4686);
and U4858 (N_4858,N_4793,N_4752);
xnor U4859 (N_4859,N_4653,N_4773);
or U4860 (N_4860,N_4694,N_4796);
and U4861 (N_4861,N_4650,N_4670);
nor U4862 (N_4862,N_4719,N_4696);
nand U4863 (N_4863,N_4728,N_4659);
and U4864 (N_4864,N_4699,N_4662);
and U4865 (N_4865,N_4715,N_4677);
or U4866 (N_4866,N_4786,N_4781);
xnor U4867 (N_4867,N_4701,N_4772);
or U4868 (N_4868,N_4707,N_4720);
nor U4869 (N_4869,N_4750,N_4762);
nor U4870 (N_4870,N_4698,N_4704);
or U4871 (N_4871,N_4722,N_4687);
nand U4872 (N_4872,N_4697,N_4766);
and U4873 (N_4873,N_4713,N_4799);
and U4874 (N_4874,N_4763,N_4703);
and U4875 (N_4875,N_4674,N_4758);
and U4876 (N_4876,N_4721,N_4746);
and U4877 (N_4877,N_4733,N_4713);
xor U4878 (N_4878,N_4692,N_4683);
xnor U4879 (N_4879,N_4795,N_4729);
and U4880 (N_4880,N_4752,N_4685);
or U4881 (N_4881,N_4682,N_4792);
nand U4882 (N_4882,N_4735,N_4659);
nor U4883 (N_4883,N_4681,N_4663);
xor U4884 (N_4884,N_4743,N_4730);
and U4885 (N_4885,N_4796,N_4771);
nor U4886 (N_4886,N_4777,N_4738);
and U4887 (N_4887,N_4771,N_4727);
and U4888 (N_4888,N_4761,N_4782);
xnor U4889 (N_4889,N_4693,N_4762);
or U4890 (N_4890,N_4746,N_4790);
nand U4891 (N_4891,N_4798,N_4778);
nand U4892 (N_4892,N_4653,N_4744);
nand U4893 (N_4893,N_4671,N_4657);
nand U4894 (N_4894,N_4664,N_4688);
or U4895 (N_4895,N_4783,N_4768);
xor U4896 (N_4896,N_4705,N_4751);
nand U4897 (N_4897,N_4694,N_4650);
and U4898 (N_4898,N_4683,N_4727);
nor U4899 (N_4899,N_4789,N_4653);
or U4900 (N_4900,N_4781,N_4722);
or U4901 (N_4901,N_4756,N_4701);
and U4902 (N_4902,N_4673,N_4769);
nand U4903 (N_4903,N_4786,N_4716);
xor U4904 (N_4904,N_4761,N_4749);
xor U4905 (N_4905,N_4661,N_4706);
nor U4906 (N_4906,N_4698,N_4778);
nor U4907 (N_4907,N_4790,N_4681);
and U4908 (N_4908,N_4784,N_4747);
and U4909 (N_4909,N_4779,N_4726);
xor U4910 (N_4910,N_4723,N_4734);
nand U4911 (N_4911,N_4725,N_4705);
and U4912 (N_4912,N_4723,N_4770);
nand U4913 (N_4913,N_4791,N_4728);
xnor U4914 (N_4914,N_4747,N_4657);
and U4915 (N_4915,N_4652,N_4730);
and U4916 (N_4916,N_4740,N_4756);
nor U4917 (N_4917,N_4675,N_4693);
nor U4918 (N_4918,N_4762,N_4681);
or U4919 (N_4919,N_4741,N_4759);
nor U4920 (N_4920,N_4677,N_4696);
and U4921 (N_4921,N_4771,N_4797);
or U4922 (N_4922,N_4775,N_4708);
xnor U4923 (N_4923,N_4708,N_4799);
nor U4924 (N_4924,N_4760,N_4739);
and U4925 (N_4925,N_4681,N_4777);
and U4926 (N_4926,N_4690,N_4770);
or U4927 (N_4927,N_4700,N_4695);
nand U4928 (N_4928,N_4726,N_4692);
nand U4929 (N_4929,N_4783,N_4734);
and U4930 (N_4930,N_4687,N_4653);
nor U4931 (N_4931,N_4659,N_4750);
nand U4932 (N_4932,N_4767,N_4695);
or U4933 (N_4933,N_4720,N_4794);
nor U4934 (N_4934,N_4650,N_4692);
nor U4935 (N_4935,N_4771,N_4667);
xor U4936 (N_4936,N_4763,N_4685);
nor U4937 (N_4937,N_4731,N_4720);
and U4938 (N_4938,N_4672,N_4697);
or U4939 (N_4939,N_4710,N_4749);
nand U4940 (N_4940,N_4655,N_4748);
nor U4941 (N_4941,N_4783,N_4701);
or U4942 (N_4942,N_4772,N_4786);
nand U4943 (N_4943,N_4651,N_4679);
or U4944 (N_4944,N_4775,N_4719);
nand U4945 (N_4945,N_4752,N_4733);
xnor U4946 (N_4946,N_4794,N_4709);
or U4947 (N_4947,N_4678,N_4671);
or U4948 (N_4948,N_4773,N_4734);
nor U4949 (N_4949,N_4694,N_4653);
nor U4950 (N_4950,N_4879,N_4920);
and U4951 (N_4951,N_4887,N_4800);
or U4952 (N_4952,N_4845,N_4804);
nand U4953 (N_4953,N_4936,N_4919);
nand U4954 (N_4954,N_4861,N_4940);
xnor U4955 (N_4955,N_4908,N_4906);
xnor U4956 (N_4956,N_4904,N_4889);
or U4957 (N_4957,N_4850,N_4942);
nor U4958 (N_4958,N_4884,N_4941);
nand U4959 (N_4959,N_4905,N_4847);
or U4960 (N_4960,N_4931,N_4860);
xnor U4961 (N_4961,N_4918,N_4934);
nand U4962 (N_4962,N_4807,N_4888);
nor U4963 (N_4963,N_4939,N_4822);
nor U4964 (N_4964,N_4819,N_4829);
or U4965 (N_4965,N_4937,N_4873);
nor U4966 (N_4966,N_4877,N_4897);
nand U4967 (N_4967,N_4870,N_4916);
nor U4968 (N_4968,N_4864,N_4824);
and U4969 (N_4969,N_4945,N_4821);
or U4970 (N_4970,N_4922,N_4869);
xnor U4971 (N_4971,N_4903,N_4896);
nand U4972 (N_4972,N_4849,N_4913);
nand U4973 (N_4973,N_4912,N_4948);
and U4974 (N_4974,N_4833,N_4841);
or U4975 (N_4975,N_4855,N_4909);
nor U4976 (N_4976,N_4932,N_4825);
nand U4977 (N_4977,N_4865,N_4898);
nor U4978 (N_4978,N_4917,N_4823);
xnor U4979 (N_4979,N_4881,N_4843);
and U4980 (N_4980,N_4867,N_4835);
or U4981 (N_4981,N_4911,N_4830);
nor U4982 (N_4982,N_4882,N_4907);
and U4983 (N_4983,N_4885,N_4859);
or U4984 (N_4984,N_4876,N_4811);
or U4985 (N_4985,N_4900,N_4921);
nor U4986 (N_4986,N_4947,N_4828);
or U4987 (N_4987,N_4834,N_4806);
xor U4988 (N_4988,N_4926,N_4915);
or U4989 (N_4989,N_4854,N_4808);
nor U4990 (N_4990,N_4910,N_4868);
nor U4991 (N_4991,N_4928,N_4812);
and U4992 (N_4992,N_4914,N_4944);
nand U4993 (N_4993,N_4815,N_4866);
nand U4994 (N_4994,N_4844,N_4946);
and U4995 (N_4995,N_4878,N_4862);
nor U4996 (N_4996,N_4899,N_4902);
nor U4997 (N_4997,N_4935,N_4943);
nand U4998 (N_4998,N_4933,N_4901);
nor U4999 (N_4999,N_4813,N_4883);
xor U5000 (N_5000,N_4872,N_4927);
or U5001 (N_5001,N_4839,N_4894);
xnor U5002 (N_5002,N_4880,N_4801);
xor U5003 (N_5003,N_4891,N_4851);
and U5004 (N_5004,N_4929,N_4923);
xnor U5005 (N_5005,N_4893,N_4820);
or U5006 (N_5006,N_4837,N_4846);
and U5007 (N_5007,N_4875,N_4842);
xnor U5008 (N_5008,N_4857,N_4805);
and U5009 (N_5009,N_4802,N_4816);
xnor U5010 (N_5010,N_4892,N_4809);
or U5011 (N_5011,N_4852,N_4817);
or U5012 (N_5012,N_4803,N_4871);
or U5013 (N_5013,N_4832,N_4853);
and U5014 (N_5014,N_4826,N_4925);
and U5015 (N_5015,N_4836,N_4938);
xnor U5016 (N_5016,N_4895,N_4856);
nor U5017 (N_5017,N_4831,N_4848);
and U5018 (N_5018,N_4814,N_4840);
nand U5019 (N_5019,N_4863,N_4874);
or U5020 (N_5020,N_4827,N_4949);
or U5021 (N_5021,N_4810,N_4890);
xor U5022 (N_5022,N_4930,N_4924);
and U5023 (N_5023,N_4886,N_4838);
xnor U5024 (N_5024,N_4858,N_4818);
nand U5025 (N_5025,N_4861,N_4850);
and U5026 (N_5026,N_4810,N_4926);
and U5027 (N_5027,N_4945,N_4891);
xnor U5028 (N_5028,N_4834,N_4881);
nor U5029 (N_5029,N_4816,N_4868);
nand U5030 (N_5030,N_4865,N_4820);
nand U5031 (N_5031,N_4941,N_4936);
or U5032 (N_5032,N_4832,N_4899);
nand U5033 (N_5033,N_4901,N_4915);
and U5034 (N_5034,N_4931,N_4899);
nand U5035 (N_5035,N_4934,N_4941);
and U5036 (N_5036,N_4943,N_4934);
and U5037 (N_5037,N_4813,N_4863);
or U5038 (N_5038,N_4934,N_4854);
xor U5039 (N_5039,N_4941,N_4801);
xnor U5040 (N_5040,N_4808,N_4880);
nand U5041 (N_5041,N_4841,N_4801);
nor U5042 (N_5042,N_4859,N_4919);
and U5043 (N_5043,N_4949,N_4811);
nand U5044 (N_5044,N_4802,N_4912);
xor U5045 (N_5045,N_4885,N_4862);
or U5046 (N_5046,N_4927,N_4800);
xnor U5047 (N_5047,N_4888,N_4843);
nor U5048 (N_5048,N_4913,N_4852);
xnor U5049 (N_5049,N_4854,N_4944);
nor U5050 (N_5050,N_4853,N_4947);
nand U5051 (N_5051,N_4942,N_4905);
nand U5052 (N_5052,N_4844,N_4842);
and U5053 (N_5053,N_4908,N_4947);
or U5054 (N_5054,N_4923,N_4874);
and U5055 (N_5055,N_4886,N_4887);
or U5056 (N_5056,N_4892,N_4808);
or U5057 (N_5057,N_4938,N_4850);
and U5058 (N_5058,N_4848,N_4936);
and U5059 (N_5059,N_4857,N_4845);
xor U5060 (N_5060,N_4949,N_4947);
and U5061 (N_5061,N_4876,N_4823);
nand U5062 (N_5062,N_4907,N_4846);
nor U5063 (N_5063,N_4900,N_4826);
nand U5064 (N_5064,N_4894,N_4885);
or U5065 (N_5065,N_4917,N_4872);
nor U5066 (N_5066,N_4831,N_4800);
nor U5067 (N_5067,N_4915,N_4883);
xnor U5068 (N_5068,N_4836,N_4918);
or U5069 (N_5069,N_4808,N_4919);
xnor U5070 (N_5070,N_4829,N_4949);
xor U5071 (N_5071,N_4827,N_4839);
and U5072 (N_5072,N_4874,N_4838);
xor U5073 (N_5073,N_4946,N_4918);
or U5074 (N_5074,N_4902,N_4842);
and U5075 (N_5075,N_4824,N_4848);
nand U5076 (N_5076,N_4895,N_4873);
or U5077 (N_5077,N_4893,N_4833);
nand U5078 (N_5078,N_4871,N_4861);
nand U5079 (N_5079,N_4892,N_4860);
and U5080 (N_5080,N_4919,N_4866);
or U5081 (N_5081,N_4939,N_4876);
and U5082 (N_5082,N_4915,N_4864);
xor U5083 (N_5083,N_4925,N_4823);
and U5084 (N_5084,N_4869,N_4880);
and U5085 (N_5085,N_4892,N_4817);
or U5086 (N_5086,N_4879,N_4802);
nand U5087 (N_5087,N_4941,N_4895);
xor U5088 (N_5088,N_4826,N_4940);
nand U5089 (N_5089,N_4822,N_4870);
or U5090 (N_5090,N_4804,N_4876);
xor U5091 (N_5091,N_4906,N_4813);
xnor U5092 (N_5092,N_4931,N_4888);
and U5093 (N_5093,N_4827,N_4887);
xnor U5094 (N_5094,N_4873,N_4835);
nand U5095 (N_5095,N_4945,N_4829);
and U5096 (N_5096,N_4856,N_4929);
nor U5097 (N_5097,N_4846,N_4801);
and U5098 (N_5098,N_4898,N_4936);
xnor U5099 (N_5099,N_4808,N_4897);
nand U5100 (N_5100,N_5015,N_5030);
nor U5101 (N_5101,N_5006,N_5083);
and U5102 (N_5102,N_4990,N_5093);
nand U5103 (N_5103,N_4968,N_4959);
nand U5104 (N_5104,N_4997,N_5018);
and U5105 (N_5105,N_5053,N_4954);
and U5106 (N_5106,N_5096,N_5028);
nand U5107 (N_5107,N_4975,N_5049);
xnor U5108 (N_5108,N_5062,N_5047);
xnor U5109 (N_5109,N_5034,N_5085);
nor U5110 (N_5110,N_4955,N_4961);
nor U5111 (N_5111,N_4957,N_4981);
xor U5112 (N_5112,N_5029,N_5061);
xor U5113 (N_5113,N_5038,N_4952);
xnor U5114 (N_5114,N_5013,N_5079);
xnor U5115 (N_5115,N_5000,N_4963);
or U5116 (N_5116,N_5005,N_5078);
or U5117 (N_5117,N_4994,N_5050);
nor U5118 (N_5118,N_4982,N_5052);
xnor U5119 (N_5119,N_4970,N_4988);
and U5120 (N_5120,N_5091,N_5039);
or U5121 (N_5121,N_5042,N_4956);
xor U5122 (N_5122,N_4974,N_5023);
and U5123 (N_5123,N_5073,N_5009);
nand U5124 (N_5124,N_4979,N_5011);
nand U5125 (N_5125,N_5003,N_4973);
xor U5126 (N_5126,N_4983,N_5088);
xor U5127 (N_5127,N_4967,N_5066);
nand U5128 (N_5128,N_5097,N_5019);
xnor U5129 (N_5129,N_5072,N_4991);
nand U5130 (N_5130,N_5058,N_5007);
and U5131 (N_5131,N_4984,N_4966);
nand U5132 (N_5132,N_4998,N_5067);
nor U5133 (N_5133,N_5098,N_4960);
and U5134 (N_5134,N_5014,N_4951);
or U5135 (N_5135,N_4962,N_5033);
and U5136 (N_5136,N_5059,N_5046);
and U5137 (N_5137,N_5092,N_5060);
nand U5138 (N_5138,N_4989,N_5032);
nor U5139 (N_5139,N_5081,N_5004);
xnor U5140 (N_5140,N_5041,N_5065);
xnor U5141 (N_5141,N_5087,N_4977);
nand U5142 (N_5142,N_5001,N_5037);
xor U5143 (N_5143,N_5043,N_5063);
or U5144 (N_5144,N_4996,N_5075);
or U5145 (N_5145,N_5054,N_5017);
nand U5146 (N_5146,N_5076,N_5095);
or U5147 (N_5147,N_5055,N_4995);
nor U5148 (N_5148,N_5036,N_4950);
nor U5149 (N_5149,N_5089,N_5031);
or U5150 (N_5150,N_5048,N_5094);
nand U5151 (N_5151,N_5070,N_5040);
or U5152 (N_5152,N_4958,N_5057);
nor U5153 (N_5153,N_5035,N_5024);
or U5154 (N_5154,N_5082,N_5074);
xor U5155 (N_5155,N_4978,N_4999);
xor U5156 (N_5156,N_5077,N_5064);
and U5157 (N_5157,N_4985,N_5051);
and U5158 (N_5158,N_4980,N_5090);
or U5159 (N_5159,N_5071,N_4993);
xor U5160 (N_5160,N_5086,N_5016);
xor U5161 (N_5161,N_4965,N_5020);
nor U5162 (N_5162,N_5084,N_5080);
nor U5163 (N_5163,N_5022,N_5010);
and U5164 (N_5164,N_5002,N_4992);
and U5165 (N_5165,N_4986,N_5068);
nor U5166 (N_5166,N_5008,N_5045);
xor U5167 (N_5167,N_5069,N_5099);
or U5168 (N_5168,N_4976,N_5044);
nand U5169 (N_5169,N_4971,N_5025);
or U5170 (N_5170,N_5026,N_5027);
or U5171 (N_5171,N_4972,N_4987);
or U5172 (N_5172,N_5021,N_4953);
and U5173 (N_5173,N_4964,N_4969);
and U5174 (N_5174,N_5056,N_5012);
xor U5175 (N_5175,N_5089,N_5030);
nor U5176 (N_5176,N_4952,N_4998);
nor U5177 (N_5177,N_5008,N_5033);
nor U5178 (N_5178,N_4956,N_5007);
or U5179 (N_5179,N_5064,N_5012);
or U5180 (N_5180,N_5096,N_5030);
or U5181 (N_5181,N_4993,N_5067);
and U5182 (N_5182,N_5071,N_5006);
and U5183 (N_5183,N_5010,N_5094);
nor U5184 (N_5184,N_5027,N_4999);
or U5185 (N_5185,N_5089,N_5027);
or U5186 (N_5186,N_5012,N_5021);
xor U5187 (N_5187,N_4965,N_4973);
nand U5188 (N_5188,N_4978,N_5009);
nand U5189 (N_5189,N_4962,N_4976);
and U5190 (N_5190,N_5031,N_5069);
nand U5191 (N_5191,N_5030,N_5011);
nor U5192 (N_5192,N_5006,N_4996);
nand U5193 (N_5193,N_5085,N_5007);
or U5194 (N_5194,N_5019,N_5064);
nor U5195 (N_5195,N_5072,N_5032);
xnor U5196 (N_5196,N_4969,N_5020);
nor U5197 (N_5197,N_5042,N_5045);
or U5198 (N_5198,N_5002,N_4998);
and U5199 (N_5199,N_5071,N_5029);
and U5200 (N_5200,N_5041,N_5017);
or U5201 (N_5201,N_4986,N_5008);
nand U5202 (N_5202,N_4994,N_4998);
nand U5203 (N_5203,N_5062,N_5069);
or U5204 (N_5204,N_4958,N_5048);
or U5205 (N_5205,N_5023,N_5062);
or U5206 (N_5206,N_5000,N_5077);
and U5207 (N_5207,N_4973,N_5065);
or U5208 (N_5208,N_5022,N_4977);
or U5209 (N_5209,N_4965,N_5082);
nor U5210 (N_5210,N_5001,N_5006);
nor U5211 (N_5211,N_5009,N_5003);
nor U5212 (N_5212,N_5070,N_4969);
nor U5213 (N_5213,N_5023,N_5079);
nor U5214 (N_5214,N_5078,N_4972);
nor U5215 (N_5215,N_5078,N_4993);
and U5216 (N_5216,N_5018,N_5054);
nor U5217 (N_5217,N_5054,N_5095);
nor U5218 (N_5218,N_5041,N_4958);
nand U5219 (N_5219,N_4956,N_5009);
nor U5220 (N_5220,N_4988,N_5058);
xnor U5221 (N_5221,N_5083,N_4971);
or U5222 (N_5222,N_5008,N_5010);
or U5223 (N_5223,N_4981,N_5006);
xor U5224 (N_5224,N_4962,N_5035);
nor U5225 (N_5225,N_5083,N_5071);
nand U5226 (N_5226,N_5025,N_5009);
xnor U5227 (N_5227,N_5055,N_5044);
nand U5228 (N_5228,N_5030,N_5013);
and U5229 (N_5229,N_5097,N_5047);
nand U5230 (N_5230,N_5040,N_4975);
nor U5231 (N_5231,N_4992,N_4977);
or U5232 (N_5232,N_5075,N_4989);
xnor U5233 (N_5233,N_5033,N_5019);
nand U5234 (N_5234,N_5044,N_4987);
nand U5235 (N_5235,N_5004,N_5037);
nor U5236 (N_5236,N_5063,N_5033);
nand U5237 (N_5237,N_4987,N_5005);
and U5238 (N_5238,N_5087,N_5024);
nor U5239 (N_5239,N_4995,N_5097);
xnor U5240 (N_5240,N_5065,N_5045);
xnor U5241 (N_5241,N_4976,N_4978);
and U5242 (N_5242,N_5084,N_5024);
xnor U5243 (N_5243,N_4965,N_5015);
and U5244 (N_5244,N_5063,N_5066);
xnor U5245 (N_5245,N_5037,N_4999);
nor U5246 (N_5246,N_5032,N_4953);
nor U5247 (N_5247,N_5006,N_5073);
xnor U5248 (N_5248,N_5093,N_4965);
xnor U5249 (N_5249,N_5089,N_5072);
nand U5250 (N_5250,N_5135,N_5165);
nand U5251 (N_5251,N_5191,N_5166);
nand U5252 (N_5252,N_5131,N_5230);
and U5253 (N_5253,N_5163,N_5222);
nand U5254 (N_5254,N_5113,N_5229);
and U5255 (N_5255,N_5245,N_5247);
nor U5256 (N_5256,N_5106,N_5224);
nor U5257 (N_5257,N_5147,N_5182);
nand U5258 (N_5258,N_5204,N_5240);
or U5259 (N_5259,N_5108,N_5136);
and U5260 (N_5260,N_5172,N_5143);
nor U5261 (N_5261,N_5100,N_5128);
nand U5262 (N_5262,N_5155,N_5130);
xnor U5263 (N_5263,N_5110,N_5200);
nor U5264 (N_5264,N_5134,N_5184);
nand U5265 (N_5265,N_5148,N_5176);
xor U5266 (N_5266,N_5209,N_5193);
xnor U5267 (N_5267,N_5178,N_5186);
and U5268 (N_5268,N_5196,N_5208);
or U5269 (N_5269,N_5183,N_5150);
xor U5270 (N_5270,N_5198,N_5239);
nand U5271 (N_5271,N_5149,N_5188);
or U5272 (N_5272,N_5177,N_5158);
nor U5273 (N_5273,N_5132,N_5238);
xnor U5274 (N_5274,N_5161,N_5243);
xor U5275 (N_5275,N_5175,N_5123);
nand U5276 (N_5276,N_5201,N_5151);
and U5277 (N_5277,N_5249,N_5118);
xor U5278 (N_5278,N_5119,N_5212);
nand U5279 (N_5279,N_5223,N_5144);
or U5280 (N_5280,N_5228,N_5107);
nand U5281 (N_5281,N_5174,N_5102);
or U5282 (N_5282,N_5169,N_5237);
nand U5283 (N_5283,N_5211,N_5153);
nand U5284 (N_5284,N_5227,N_5206);
and U5285 (N_5285,N_5111,N_5207);
xnor U5286 (N_5286,N_5127,N_5234);
or U5287 (N_5287,N_5116,N_5197);
nor U5288 (N_5288,N_5125,N_5115);
nand U5289 (N_5289,N_5114,N_5231);
nor U5290 (N_5290,N_5233,N_5202);
nand U5291 (N_5291,N_5164,N_5124);
or U5292 (N_5292,N_5121,N_5242);
nand U5293 (N_5293,N_5225,N_5241);
or U5294 (N_5294,N_5152,N_5146);
nor U5295 (N_5295,N_5112,N_5145);
nand U5296 (N_5296,N_5199,N_5140);
xor U5297 (N_5297,N_5157,N_5101);
xnor U5298 (N_5298,N_5219,N_5194);
or U5299 (N_5299,N_5203,N_5215);
or U5300 (N_5300,N_5120,N_5154);
nor U5301 (N_5301,N_5109,N_5104);
nor U5302 (N_5302,N_5189,N_5179);
nor U5303 (N_5303,N_5137,N_5159);
xnor U5304 (N_5304,N_5213,N_5226);
xor U5305 (N_5305,N_5171,N_5180);
and U5306 (N_5306,N_5192,N_5141);
or U5307 (N_5307,N_5105,N_5216);
and U5308 (N_5308,N_5160,N_5236);
and U5309 (N_5309,N_5217,N_5142);
nand U5310 (N_5310,N_5173,N_5218);
and U5311 (N_5311,N_5181,N_5246);
nor U5312 (N_5312,N_5168,N_5190);
nor U5313 (N_5313,N_5156,N_5117);
xnor U5314 (N_5314,N_5129,N_5210);
nand U5315 (N_5315,N_5220,N_5214);
nor U5316 (N_5316,N_5162,N_5244);
and U5317 (N_5317,N_5185,N_5133);
and U5318 (N_5318,N_5139,N_5103);
and U5319 (N_5319,N_5221,N_5170);
and U5320 (N_5320,N_5235,N_5122);
and U5321 (N_5321,N_5232,N_5187);
xor U5322 (N_5322,N_5138,N_5205);
or U5323 (N_5323,N_5248,N_5195);
nand U5324 (N_5324,N_5126,N_5167);
or U5325 (N_5325,N_5242,N_5102);
nand U5326 (N_5326,N_5191,N_5233);
nor U5327 (N_5327,N_5241,N_5221);
and U5328 (N_5328,N_5248,N_5238);
nand U5329 (N_5329,N_5137,N_5220);
nor U5330 (N_5330,N_5166,N_5141);
and U5331 (N_5331,N_5248,N_5232);
nand U5332 (N_5332,N_5219,N_5118);
or U5333 (N_5333,N_5239,N_5109);
or U5334 (N_5334,N_5187,N_5125);
nor U5335 (N_5335,N_5117,N_5191);
and U5336 (N_5336,N_5224,N_5201);
nor U5337 (N_5337,N_5125,N_5230);
nor U5338 (N_5338,N_5241,N_5111);
nor U5339 (N_5339,N_5144,N_5231);
and U5340 (N_5340,N_5236,N_5185);
and U5341 (N_5341,N_5203,N_5233);
xnor U5342 (N_5342,N_5144,N_5178);
and U5343 (N_5343,N_5208,N_5217);
or U5344 (N_5344,N_5199,N_5223);
or U5345 (N_5345,N_5107,N_5227);
xor U5346 (N_5346,N_5192,N_5220);
nor U5347 (N_5347,N_5208,N_5220);
nor U5348 (N_5348,N_5129,N_5152);
nand U5349 (N_5349,N_5244,N_5215);
xor U5350 (N_5350,N_5140,N_5121);
xnor U5351 (N_5351,N_5179,N_5106);
and U5352 (N_5352,N_5118,N_5115);
nor U5353 (N_5353,N_5203,N_5126);
nand U5354 (N_5354,N_5217,N_5138);
nor U5355 (N_5355,N_5177,N_5153);
and U5356 (N_5356,N_5163,N_5158);
xnor U5357 (N_5357,N_5176,N_5142);
nor U5358 (N_5358,N_5156,N_5247);
nor U5359 (N_5359,N_5110,N_5180);
or U5360 (N_5360,N_5152,N_5182);
nor U5361 (N_5361,N_5188,N_5187);
nand U5362 (N_5362,N_5121,N_5197);
or U5363 (N_5363,N_5186,N_5210);
nand U5364 (N_5364,N_5194,N_5204);
or U5365 (N_5365,N_5203,N_5152);
nand U5366 (N_5366,N_5181,N_5128);
nor U5367 (N_5367,N_5108,N_5247);
and U5368 (N_5368,N_5225,N_5125);
nor U5369 (N_5369,N_5210,N_5242);
xor U5370 (N_5370,N_5153,N_5173);
nor U5371 (N_5371,N_5220,N_5162);
xnor U5372 (N_5372,N_5245,N_5122);
nand U5373 (N_5373,N_5201,N_5236);
nor U5374 (N_5374,N_5144,N_5146);
nand U5375 (N_5375,N_5132,N_5214);
and U5376 (N_5376,N_5144,N_5108);
or U5377 (N_5377,N_5171,N_5225);
and U5378 (N_5378,N_5137,N_5157);
nor U5379 (N_5379,N_5185,N_5206);
and U5380 (N_5380,N_5196,N_5204);
nand U5381 (N_5381,N_5114,N_5132);
or U5382 (N_5382,N_5218,N_5170);
xnor U5383 (N_5383,N_5126,N_5180);
and U5384 (N_5384,N_5143,N_5176);
and U5385 (N_5385,N_5198,N_5114);
or U5386 (N_5386,N_5137,N_5118);
xnor U5387 (N_5387,N_5107,N_5244);
or U5388 (N_5388,N_5241,N_5215);
xnor U5389 (N_5389,N_5128,N_5187);
or U5390 (N_5390,N_5183,N_5153);
and U5391 (N_5391,N_5120,N_5216);
nor U5392 (N_5392,N_5232,N_5199);
or U5393 (N_5393,N_5199,N_5205);
nor U5394 (N_5394,N_5213,N_5183);
xnor U5395 (N_5395,N_5202,N_5154);
nor U5396 (N_5396,N_5117,N_5143);
nor U5397 (N_5397,N_5216,N_5182);
nor U5398 (N_5398,N_5111,N_5104);
and U5399 (N_5399,N_5153,N_5131);
and U5400 (N_5400,N_5278,N_5263);
and U5401 (N_5401,N_5309,N_5381);
nand U5402 (N_5402,N_5299,N_5354);
nor U5403 (N_5403,N_5344,N_5316);
or U5404 (N_5404,N_5269,N_5288);
or U5405 (N_5405,N_5360,N_5320);
or U5406 (N_5406,N_5346,N_5389);
nand U5407 (N_5407,N_5345,N_5370);
nor U5408 (N_5408,N_5347,N_5367);
xnor U5409 (N_5409,N_5268,N_5304);
xor U5410 (N_5410,N_5256,N_5276);
xnor U5411 (N_5411,N_5292,N_5255);
or U5412 (N_5412,N_5379,N_5271);
nand U5413 (N_5413,N_5390,N_5394);
xor U5414 (N_5414,N_5380,N_5369);
or U5415 (N_5415,N_5296,N_5307);
or U5416 (N_5416,N_5387,N_5283);
and U5417 (N_5417,N_5293,N_5374);
or U5418 (N_5418,N_5396,N_5281);
or U5419 (N_5419,N_5253,N_5302);
or U5420 (N_5420,N_5338,N_5393);
xor U5421 (N_5421,N_5258,N_5325);
or U5422 (N_5422,N_5353,N_5286);
nand U5423 (N_5423,N_5371,N_5277);
nand U5424 (N_5424,N_5282,N_5272);
nor U5425 (N_5425,N_5399,N_5388);
nand U5426 (N_5426,N_5359,N_5262);
or U5427 (N_5427,N_5322,N_5358);
nand U5428 (N_5428,N_5334,N_5397);
xor U5429 (N_5429,N_5328,N_5305);
xnor U5430 (N_5430,N_5335,N_5257);
and U5431 (N_5431,N_5294,N_5376);
or U5432 (N_5432,N_5349,N_5364);
and U5433 (N_5433,N_5290,N_5368);
or U5434 (N_5434,N_5297,N_5314);
or U5435 (N_5435,N_5384,N_5264);
and U5436 (N_5436,N_5382,N_5341);
or U5437 (N_5437,N_5357,N_5279);
xnor U5438 (N_5438,N_5348,N_5300);
nor U5439 (N_5439,N_5295,N_5332);
xor U5440 (N_5440,N_5362,N_5356);
nor U5441 (N_5441,N_5267,N_5333);
or U5442 (N_5442,N_5351,N_5339);
nor U5443 (N_5443,N_5327,N_5372);
or U5444 (N_5444,N_5342,N_5317);
nor U5445 (N_5445,N_5323,N_5395);
and U5446 (N_5446,N_5383,N_5251);
and U5447 (N_5447,N_5398,N_5326);
or U5448 (N_5448,N_5385,N_5355);
xor U5449 (N_5449,N_5284,N_5273);
or U5450 (N_5450,N_5291,N_5310);
or U5451 (N_5451,N_5329,N_5319);
nor U5452 (N_5452,N_5254,N_5340);
xor U5453 (N_5453,N_5303,N_5287);
or U5454 (N_5454,N_5361,N_5343);
and U5455 (N_5455,N_5373,N_5306);
and U5456 (N_5456,N_5337,N_5311);
and U5457 (N_5457,N_5391,N_5331);
nor U5458 (N_5458,N_5318,N_5270);
or U5459 (N_5459,N_5261,N_5265);
nor U5460 (N_5460,N_5274,N_5280);
and U5461 (N_5461,N_5392,N_5377);
xnor U5462 (N_5462,N_5285,N_5312);
nor U5463 (N_5463,N_5266,N_5350);
and U5464 (N_5464,N_5298,N_5365);
nand U5465 (N_5465,N_5352,N_5252);
and U5466 (N_5466,N_5386,N_5259);
nand U5467 (N_5467,N_5324,N_5378);
xnor U5468 (N_5468,N_5260,N_5301);
nand U5469 (N_5469,N_5308,N_5313);
xnor U5470 (N_5470,N_5330,N_5315);
and U5471 (N_5471,N_5321,N_5336);
nor U5472 (N_5472,N_5366,N_5250);
and U5473 (N_5473,N_5363,N_5289);
xnor U5474 (N_5474,N_5375,N_5275);
nand U5475 (N_5475,N_5261,N_5292);
nand U5476 (N_5476,N_5272,N_5311);
xor U5477 (N_5477,N_5330,N_5350);
and U5478 (N_5478,N_5308,N_5304);
nor U5479 (N_5479,N_5392,N_5280);
and U5480 (N_5480,N_5362,N_5280);
nand U5481 (N_5481,N_5358,N_5374);
nor U5482 (N_5482,N_5348,N_5380);
or U5483 (N_5483,N_5344,N_5269);
nor U5484 (N_5484,N_5324,N_5341);
xor U5485 (N_5485,N_5332,N_5365);
xnor U5486 (N_5486,N_5355,N_5333);
and U5487 (N_5487,N_5378,N_5290);
nand U5488 (N_5488,N_5332,N_5395);
xor U5489 (N_5489,N_5299,N_5277);
xor U5490 (N_5490,N_5295,N_5304);
xnor U5491 (N_5491,N_5303,N_5263);
xor U5492 (N_5492,N_5259,N_5250);
nand U5493 (N_5493,N_5379,N_5294);
nand U5494 (N_5494,N_5268,N_5289);
and U5495 (N_5495,N_5388,N_5391);
and U5496 (N_5496,N_5287,N_5372);
nand U5497 (N_5497,N_5361,N_5370);
and U5498 (N_5498,N_5371,N_5338);
nand U5499 (N_5499,N_5323,N_5371);
or U5500 (N_5500,N_5360,N_5350);
and U5501 (N_5501,N_5318,N_5269);
nor U5502 (N_5502,N_5331,N_5319);
nor U5503 (N_5503,N_5361,N_5282);
or U5504 (N_5504,N_5270,N_5257);
nor U5505 (N_5505,N_5295,N_5379);
or U5506 (N_5506,N_5264,N_5313);
nor U5507 (N_5507,N_5324,N_5339);
nand U5508 (N_5508,N_5283,N_5318);
xor U5509 (N_5509,N_5273,N_5332);
nand U5510 (N_5510,N_5259,N_5306);
nand U5511 (N_5511,N_5373,N_5314);
nand U5512 (N_5512,N_5327,N_5288);
nor U5513 (N_5513,N_5399,N_5359);
nand U5514 (N_5514,N_5281,N_5364);
or U5515 (N_5515,N_5258,N_5281);
nand U5516 (N_5516,N_5307,N_5347);
or U5517 (N_5517,N_5300,N_5340);
or U5518 (N_5518,N_5334,N_5384);
xor U5519 (N_5519,N_5332,N_5339);
or U5520 (N_5520,N_5395,N_5337);
xnor U5521 (N_5521,N_5295,N_5280);
xnor U5522 (N_5522,N_5254,N_5333);
or U5523 (N_5523,N_5307,N_5321);
nand U5524 (N_5524,N_5273,N_5399);
xnor U5525 (N_5525,N_5358,N_5327);
nor U5526 (N_5526,N_5347,N_5271);
xnor U5527 (N_5527,N_5382,N_5377);
or U5528 (N_5528,N_5384,N_5359);
or U5529 (N_5529,N_5294,N_5363);
or U5530 (N_5530,N_5363,N_5314);
nand U5531 (N_5531,N_5370,N_5289);
or U5532 (N_5532,N_5269,N_5272);
or U5533 (N_5533,N_5258,N_5279);
nor U5534 (N_5534,N_5373,N_5317);
xnor U5535 (N_5535,N_5353,N_5308);
nand U5536 (N_5536,N_5354,N_5348);
xnor U5537 (N_5537,N_5269,N_5371);
xor U5538 (N_5538,N_5316,N_5298);
xor U5539 (N_5539,N_5342,N_5330);
nor U5540 (N_5540,N_5391,N_5272);
nand U5541 (N_5541,N_5345,N_5390);
nand U5542 (N_5542,N_5368,N_5395);
and U5543 (N_5543,N_5329,N_5339);
xnor U5544 (N_5544,N_5360,N_5253);
nand U5545 (N_5545,N_5375,N_5351);
nand U5546 (N_5546,N_5255,N_5358);
nand U5547 (N_5547,N_5304,N_5255);
xor U5548 (N_5548,N_5293,N_5323);
nor U5549 (N_5549,N_5390,N_5365);
nor U5550 (N_5550,N_5426,N_5447);
or U5551 (N_5551,N_5452,N_5542);
nor U5552 (N_5552,N_5470,N_5421);
nor U5553 (N_5553,N_5476,N_5503);
and U5554 (N_5554,N_5514,N_5466);
nand U5555 (N_5555,N_5405,N_5422);
or U5556 (N_5556,N_5533,N_5446);
nand U5557 (N_5557,N_5509,N_5544);
and U5558 (N_5558,N_5454,N_5505);
xor U5559 (N_5559,N_5499,N_5495);
nand U5560 (N_5560,N_5532,N_5529);
and U5561 (N_5561,N_5429,N_5448);
nor U5562 (N_5562,N_5501,N_5545);
nand U5563 (N_5563,N_5469,N_5477);
xor U5564 (N_5564,N_5472,N_5451);
nor U5565 (N_5565,N_5425,N_5481);
nand U5566 (N_5566,N_5415,N_5423);
nor U5567 (N_5567,N_5407,N_5513);
or U5568 (N_5568,N_5468,N_5419);
nor U5569 (N_5569,N_5535,N_5526);
and U5570 (N_5570,N_5504,N_5431);
nand U5571 (N_5571,N_5522,N_5534);
and U5572 (N_5572,N_5546,N_5489);
or U5573 (N_5573,N_5420,N_5538);
or U5574 (N_5574,N_5414,N_5401);
nor U5575 (N_5575,N_5417,N_5443);
and U5576 (N_5576,N_5449,N_5478);
or U5577 (N_5577,N_5536,N_5427);
xnor U5578 (N_5578,N_5496,N_5459);
nor U5579 (N_5579,N_5488,N_5455);
or U5580 (N_5580,N_5528,N_5516);
nand U5581 (N_5581,N_5480,N_5523);
and U5582 (N_5582,N_5436,N_5464);
and U5583 (N_5583,N_5453,N_5402);
nand U5584 (N_5584,N_5530,N_5519);
or U5585 (N_5585,N_5450,N_5465);
xnor U5586 (N_5586,N_5458,N_5457);
or U5587 (N_5587,N_5435,N_5515);
and U5588 (N_5588,N_5487,N_5485);
nand U5589 (N_5589,N_5462,N_5410);
or U5590 (N_5590,N_5537,N_5444);
or U5591 (N_5591,N_5527,N_5441);
nand U5592 (N_5592,N_5437,N_5433);
nor U5593 (N_5593,N_5482,N_5460);
xor U5594 (N_5594,N_5428,N_5409);
xor U5595 (N_5595,N_5467,N_5484);
xor U5596 (N_5596,N_5486,N_5440);
nor U5597 (N_5597,N_5539,N_5524);
and U5598 (N_5598,N_5491,N_5413);
nand U5599 (N_5599,N_5548,N_5434);
nand U5600 (N_5600,N_5461,N_5490);
nor U5601 (N_5601,N_5473,N_5403);
xnor U5602 (N_5602,N_5424,N_5531);
nand U5603 (N_5603,N_5508,N_5521);
xnor U5604 (N_5604,N_5400,N_5525);
or U5605 (N_5605,N_5547,N_5412);
or U5606 (N_5606,N_5549,N_5541);
nand U5607 (N_5607,N_5404,N_5497);
nor U5608 (N_5608,N_5518,N_5411);
nor U5609 (N_5609,N_5498,N_5456);
nor U5610 (N_5610,N_5408,N_5439);
xnor U5611 (N_5611,N_5474,N_5471);
nand U5612 (N_5612,N_5507,N_5479);
and U5613 (N_5613,N_5500,N_5475);
and U5614 (N_5614,N_5442,N_5506);
nand U5615 (N_5615,N_5510,N_5492);
xor U5616 (N_5616,N_5416,N_5483);
nand U5617 (N_5617,N_5430,N_5406);
nor U5618 (N_5618,N_5512,N_5494);
or U5619 (N_5619,N_5493,N_5438);
xor U5620 (N_5620,N_5511,N_5517);
or U5621 (N_5621,N_5540,N_5543);
or U5622 (N_5622,N_5445,N_5418);
nand U5623 (N_5623,N_5432,N_5463);
xnor U5624 (N_5624,N_5502,N_5520);
and U5625 (N_5625,N_5416,N_5505);
nand U5626 (N_5626,N_5493,N_5401);
xor U5627 (N_5627,N_5504,N_5537);
nand U5628 (N_5628,N_5472,N_5431);
nand U5629 (N_5629,N_5431,N_5466);
or U5630 (N_5630,N_5495,N_5502);
nor U5631 (N_5631,N_5439,N_5423);
nand U5632 (N_5632,N_5444,N_5455);
or U5633 (N_5633,N_5458,N_5490);
xnor U5634 (N_5634,N_5407,N_5534);
nor U5635 (N_5635,N_5494,N_5404);
nand U5636 (N_5636,N_5452,N_5494);
xnor U5637 (N_5637,N_5480,N_5509);
nand U5638 (N_5638,N_5432,N_5529);
xor U5639 (N_5639,N_5435,N_5525);
xnor U5640 (N_5640,N_5401,N_5498);
nor U5641 (N_5641,N_5464,N_5444);
xor U5642 (N_5642,N_5454,N_5504);
or U5643 (N_5643,N_5531,N_5455);
and U5644 (N_5644,N_5433,N_5404);
nand U5645 (N_5645,N_5416,N_5437);
xnor U5646 (N_5646,N_5413,N_5527);
nor U5647 (N_5647,N_5446,N_5492);
and U5648 (N_5648,N_5490,N_5405);
and U5649 (N_5649,N_5436,N_5438);
xnor U5650 (N_5650,N_5412,N_5458);
xor U5651 (N_5651,N_5438,N_5458);
nand U5652 (N_5652,N_5538,N_5539);
and U5653 (N_5653,N_5402,N_5475);
nand U5654 (N_5654,N_5425,N_5463);
xnor U5655 (N_5655,N_5432,N_5418);
nor U5656 (N_5656,N_5472,N_5530);
nand U5657 (N_5657,N_5501,N_5487);
xnor U5658 (N_5658,N_5450,N_5441);
or U5659 (N_5659,N_5478,N_5465);
and U5660 (N_5660,N_5474,N_5486);
or U5661 (N_5661,N_5468,N_5533);
nor U5662 (N_5662,N_5536,N_5421);
or U5663 (N_5663,N_5412,N_5407);
and U5664 (N_5664,N_5532,N_5460);
xor U5665 (N_5665,N_5431,N_5447);
nand U5666 (N_5666,N_5503,N_5423);
nor U5667 (N_5667,N_5420,N_5522);
nor U5668 (N_5668,N_5426,N_5466);
nand U5669 (N_5669,N_5532,N_5440);
nand U5670 (N_5670,N_5415,N_5413);
xnor U5671 (N_5671,N_5429,N_5412);
nand U5672 (N_5672,N_5413,N_5495);
nand U5673 (N_5673,N_5515,N_5448);
nor U5674 (N_5674,N_5417,N_5549);
or U5675 (N_5675,N_5459,N_5411);
or U5676 (N_5676,N_5442,N_5420);
nand U5677 (N_5677,N_5444,N_5418);
nor U5678 (N_5678,N_5507,N_5514);
nor U5679 (N_5679,N_5466,N_5438);
xnor U5680 (N_5680,N_5441,N_5459);
or U5681 (N_5681,N_5411,N_5505);
nand U5682 (N_5682,N_5459,N_5517);
and U5683 (N_5683,N_5433,N_5463);
and U5684 (N_5684,N_5416,N_5479);
nand U5685 (N_5685,N_5538,N_5534);
or U5686 (N_5686,N_5490,N_5463);
xnor U5687 (N_5687,N_5433,N_5480);
nor U5688 (N_5688,N_5540,N_5508);
or U5689 (N_5689,N_5532,N_5486);
nand U5690 (N_5690,N_5463,N_5518);
nand U5691 (N_5691,N_5500,N_5483);
xor U5692 (N_5692,N_5488,N_5407);
xnor U5693 (N_5693,N_5528,N_5494);
or U5694 (N_5694,N_5444,N_5469);
nand U5695 (N_5695,N_5479,N_5409);
nor U5696 (N_5696,N_5547,N_5544);
xnor U5697 (N_5697,N_5450,N_5403);
nand U5698 (N_5698,N_5511,N_5482);
nand U5699 (N_5699,N_5411,N_5475);
nand U5700 (N_5700,N_5611,N_5602);
or U5701 (N_5701,N_5635,N_5683);
or U5702 (N_5702,N_5601,N_5637);
nor U5703 (N_5703,N_5674,N_5551);
nand U5704 (N_5704,N_5616,N_5685);
nor U5705 (N_5705,N_5561,N_5647);
nand U5706 (N_5706,N_5628,N_5668);
or U5707 (N_5707,N_5675,N_5580);
and U5708 (N_5708,N_5577,N_5625);
nand U5709 (N_5709,N_5632,N_5665);
xnor U5710 (N_5710,N_5582,N_5688);
nor U5711 (N_5711,N_5680,N_5605);
nand U5712 (N_5712,N_5676,N_5641);
nor U5713 (N_5713,N_5624,N_5699);
xnor U5714 (N_5714,N_5630,N_5642);
nand U5715 (N_5715,N_5644,N_5550);
nand U5716 (N_5716,N_5598,N_5692);
nand U5717 (N_5717,N_5572,N_5650);
or U5718 (N_5718,N_5684,N_5607);
nor U5719 (N_5719,N_5556,N_5571);
nor U5720 (N_5720,N_5640,N_5627);
nand U5721 (N_5721,N_5631,N_5663);
xor U5722 (N_5722,N_5574,N_5664);
nand U5723 (N_5723,N_5660,N_5603);
nand U5724 (N_5724,N_5682,N_5599);
xnor U5725 (N_5725,N_5673,N_5643);
xnor U5726 (N_5726,N_5649,N_5583);
nor U5727 (N_5727,N_5573,N_5587);
nor U5728 (N_5728,N_5648,N_5693);
or U5729 (N_5729,N_5689,N_5557);
or U5730 (N_5730,N_5606,N_5653);
and U5731 (N_5731,N_5698,N_5552);
nand U5732 (N_5732,N_5565,N_5614);
xor U5733 (N_5733,N_5554,N_5652);
or U5734 (N_5734,N_5608,N_5634);
nor U5735 (N_5735,N_5585,N_5618);
nor U5736 (N_5736,N_5656,N_5655);
xnor U5737 (N_5737,N_5591,N_5626);
and U5738 (N_5738,N_5564,N_5669);
xnor U5739 (N_5739,N_5681,N_5622);
nand U5740 (N_5740,N_5687,N_5657);
or U5741 (N_5741,N_5600,N_5579);
nand U5742 (N_5742,N_5570,N_5553);
xor U5743 (N_5743,N_5609,N_5586);
nor U5744 (N_5744,N_5619,N_5612);
and U5745 (N_5745,N_5575,N_5633);
nor U5746 (N_5746,N_5651,N_5679);
or U5747 (N_5747,N_5578,N_5654);
and U5748 (N_5748,N_5666,N_5604);
nor U5749 (N_5749,N_5645,N_5695);
xnor U5750 (N_5750,N_5560,N_5636);
xor U5751 (N_5751,N_5691,N_5596);
xnor U5752 (N_5752,N_5667,N_5590);
nor U5753 (N_5753,N_5610,N_5588);
nor U5754 (N_5754,N_5613,N_5694);
nand U5755 (N_5755,N_5621,N_5697);
xnor U5756 (N_5756,N_5595,N_5672);
nor U5757 (N_5757,N_5562,N_5659);
xnor U5758 (N_5758,N_5563,N_5690);
or U5759 (N_5759,N_5589,N_5638);
xnor U5760 (N_5760,N_5592,N_5566);
xor U5761 (N_5761,N_5558,N_5678);
or U5762 (N_5762,N_5696,N_5568);
nor U5763 (N_5763,N_5661,N_5658);
nor U5764 (N_5764,N_5581,N_5646);
nand U5765 (N_5765,N_5594,N_5623);
nor U5766 (N_5766,N_5593,N_5686);
and U5767 (N_5767,N_5629,N_5670);
nand U5768 (N_5768,N_5615,N_5576);
and U5769 (N_5769,N_5671,N_5559);
or U5770 (N_5770,N_5677,N_5569);
or U5771 (N_5771,N_5617,N_5597);
or U5772 (N_5772,N_5567,N_5555);
xor U5773 (N_5773,N_5620,N_5639);
and U5774 (N_5774,N_5584,N_5662);
or U5775 (N_5775,N_5633,N_5564);
or U5776 (N_5776,N_5567,N_5680);
xor U5777 (N_5777,N_5644,N_5632);
nand U5778 (N_5778,N_5643,N_5682);
or U5779 (N_5779,N_5559,N_5634);
xor U5780 (N_5780,N_5660,N_5685);
xor U5781 (N_5781,N_5683,N_5655);
and U5782 (N_5782,N_5568,N_5624);
or U5783 (N_5783,N_5668,N_5659);
nand U5784 (N_5784,N_5602,N_5558);
and U5785 (N_5785,N_5571,N_5653);
nand U5786 (N_5786,N_5652,N_5635);
nand U5787 (N_5787,N_5613,N_5550);
and U5788 (N_5788,N_5597,N_5676);
or U5789 (N_5789,N_5558,N_5594);
nor U5790 (N_5790,N_5661,N_5617);
or U5791 (N_5791,N_5625,N_5592);
nor U5792 (N_5792,N_5653,N_5649);
nor U5793 (N_5793,N_5555,N_5679);
nand U5794 (N_5794,N_5594,N_5686);
nand U5795 (N_5795,N_5668,N_5685);
or U5796 (N_5796,N_5698,N_5571);
or U5797 (N_5797,N_5584,N_5687);
nand U5798 (N_5798,N_5610,N_5638);
nand U5799 (N_5799,N_5608,N_5564);
nor U5800 (N_5800,N_5674,N_5586);
nand U5801 (N_5801,N_5550,N_5620);
nor U5802 (N_5802,N_5631,N_5616);
and U5803 (N_5803,N_5613,N_5562);
or U5804 (N_5804,N_5647,N_5601);
nand U5805 (N_5805,N_5586,N_5624);
or U5806 (N_5806,N_5669,N_5600);
nand U5807 (N_5807,N_5693,N_5654);
or U5808 (N_5808,N_5579,N_5698);
nand U5809 (N_5809,N_5568,N_5570);
and U5810 (N_5810,N_5671,N_5584);
xnor U5811 (N_5811,N_5676,N_5609);
nand U5812 (N_5812,N_5574,N_5691);
nor U5813 (N_5813,N_5672,N_5662);
nor U5814 (N_5814,N_5593,N_5693);
nand U5815 (N_5815,N_5639,N_5575);
and U5816 (N_5816,N_5623,N_5577);
and U5817 (N_5817,N_5564,N_5651);
nand U5818 (N_5818,N_5622,N_5677);
xnor U5819 (N_5819,N_5665,N_5681);
nor U5820 (N_5820,N_5591,N_5673);
nor U5821 (N_5821,N_5557,N_5653);
nor U5822 (N_5822,N_5559,N_5575);
nand U5823 (N_5823,N_5570,N_5640);
xnor U5824 (N_5824,N_5652,N_5655);
and U5825 (N_5825,N_5673,N_5641);
nor U5826 (N_5826,N_5570,N_5648);
or U5827 (N_5827,N_5673,N_5651);
xor U5828 (N_5828,N_5676,N_5650);
xor U5829 (N_5829,N_5688,N_5637);
or U5830 (N_5830,N_5638,N_5614);
or U5831 (N_5831,N_5634,N_5612);
or U5832 (N_5832,N_5699,N_5580);
and U5833 (N_5833,N_5639,N_5623);
nand U5834 (N_5834,N_5647,N_5609);
nand U5835 (N_5835,N_5635,N_5552);
nand U5836 (N_5836,N_5607,N_5569);
nor U5837 (N_5837,N_5571,N_5595);
xnor U5838 (N_5838,N_5634,N_5661);
xor U5839 (N_5839,N_5670,N_5633);
nand U5840 (N_5840,N_5596,N_5619);
xnor U5841 (N_5841,N_5696,N_5626);
or U5842 (N_5842,N_5644,N_5695);
or U5843 (N_5843,N_5643,N_5626);
xor U5844 (N_5844,N_5628,N_5649);
nor U5845 (N_5845,N_5573,N_5565);
nand U5846 (N_5846,N_5662,N_5560);
or U5847 (N_5847,N_5679,N_5637);
nand U5848 (N_5848,N_5622,N_5636);
xnor U5849 (N_5849,N_5638,N_5626);
xor U5850 (N_5850,N_5754,N_5821);
xor U5851 (N_5851,N_5793,N_5707);
xor U5852 (N_5852,N_5771,N_5764);
nor U5853 (N_5853,N_5768,N_5813);
or U5854 (N_5854,N_5830,N_5752);
and U5855 (N_5855,N_5704,N_5712);
nand U5856 (N_5856,N_5700,N_5790);
or U5857 (N_5857,N_5775,N_5779);
or U5858 (N_5858,N_5806,N_5814);
nand U5859 (N_5859,N_5773,N_5702);
nand U5860 (N_5860,N_5701,N_5737);
nor U5861 (N_5861,N_5747,N_5727);
and U5862 (N_5862,N_5785,N_5759);
nor U5863 (N_5863,N_5834,N_5732);
nand U5864 (N_5864,N_5703,N_5801);
xnor U5865 (N_5865,N_5803,N_5731);
nor U5866 (N_5866,N_5799,N_5817);
and U5867 (N_5867,N_5774,N_5780);
nor U5868 (N_5868,N_5743,N_5825);
xnor U5869 (N_5869,N_5783,N_5789);
xor U5870 (N_5870,N_5820,N_5844);
xnor U5871 (N_5871,N_5812,N_5810);
and U5872 (N_5872,N_5841,N_5787);
xor U5873 (N_5873,N_5795,N_5715);
nor U5874 (N_5874,N_5716,N_5829);
or U5875 (N_5875,N_5815,N_5724);
nand U5876 (N_5876,N_5714,N_5755);
xnor U5877 (N_5877,N_5767,N_5763);
or U5878 (N_5878,N_5746,N_5730);
nand U5879 (N_5879,N_5842,N_5720);
and U5880 (N_5880,N_5710,N_5709);
nand U5881 (N_5881,N_5756,N_5761);
and U5882 (N_5882,N_5753,N_5839);
and U5883 (N_5883,N_5706,N_5765);
nor U5884 (N_5884,N_5837,N_5751);
xor U5885 (N_5885,N_5843,N_5722);
and U5886 (N_5886,N_5729,N_5835);
nand U5887 (N_5887,N_5733,N_5741);
xnor U5888 (N_5888,N_5800,N_5805);
or U5889 (N_5889,N_5705,N_5778);
xnor U5890 (N_5890,N_5723,N_5748);
nand U5891 (N_5891,N_5726,N_5794);
nand U5892 (N_5892,N_5734,N_5827);
and U5893 (N_5893,N_5792,N_5711);
or U5894 (N_5894,N_5848,N_5831);
and U5895 (N_5895,N_5784,N_5725);
nor U5896 (N_5896,N_5760,N_5802);
nor U5897 (N_5897,N_5849,N_5708);
nand U5898 (N_5898,N_5757,N_5797);
and U5899 (N_5899,N_5739,N_5713);
xor U5900 (N_5900,N_5809,N_5736);
or U5901 (N_5901,N_5766,N_5828);
nor U5902 (N_5902,N_5804,N_5788);
nand U5903 (N_5903,N_5798,N_5742);
nor U5904 (N_5904,N_5721,N_5719);
xor U5905 (N_5905,N_5796,N_5777);
and U5906 (N_5906,N_5832,N_5717);
xnor U5907 (N_5907,N_5823,N_5840);
nand U5908 (N_5908,N_5826,N_5818);
nor U5909 (N_5909,N_5847,N_5846);
xor U5910 (N_5910,N_5750,N_5772);
xnor U5911 (N_5911,N_5824,N_5770);
and U5912 (N_5912,N_5776,N_5833);
nand U5913 (N_5913,N_5786,N_5738);
or U5914 (N_5914,N_5745,N_5845);
or U5915 (N_5915,N_5769,N_5740);
nand U5916 (N_5916,N_5735,N_5807);
xor U5917 (N_5917,N_5808,N_5791);
or U5918 (N_5918,N_5811,N_5822);
xor U5919 (N_5919,N_5758,N_5718);
xor U5920 (N_5920,N_5816,N_5728);
or U5921 (N_5921,N_5749,N_5819);
or U5922 (N_5922,N_5838,N_5781);
or U5923 (N_5923,N_5782,N_5744);
and U5924 (N_5924,N_5762,N_5836);
xor U5925 (N_5925,N_5777,N_5845);
or U5926 (N_5926,N_5730,N_5831);
or U5927 (N_5927,N_5772,N_5756);
xnor U5928 (N_5928,N_5824,N_5735);
xor U5929 (N_5929,N_5804,N_5732);
nand U5930 (N_5930,N_5742,N_5760);
and U5931 (N_5931,N_5836,N_5778);
or U5932 (N_5932,N_5845,N_5729);
or U5933 (N_5933,N_5830,N_5700);
and U5934 (N_5934,N_5829,N_5803);
or U5935 (N_5935,N_5708,N_5770);
or U5936 (N_5936,N_5700,N_5763);
and U5937 (N_5937,N_5768,N_5754);
nand U5938 (N_5938,N_5814,N_5834);
xor U5939 (N_5939,N_5779,N_5841);
nor U5940 (N_5940,N_5790,N_5822);
or U5941 (N_5941,N_5828,N_5798);
or U5942 (N_5942,N_5730,N_5719);
and U5943 (N_5943,N_5818,N_5788);
nor U5944 (N_5944,N_5761,N_5813);
or U5945 (N_5945,N_5823,N_5803);
xnor U5946 (N_5946,N_5816,N_5781);
nor U5947 (N_5947,N_5805,N_5806);
nor U5948 (N_5948,N_5771,N_5822);
or U5949 (N_5949,N_5788,N_5731);
nor U5950 (N_5950,N_5778,N_5718);
nand U5951 (N_5951,N_5781,N_5833);
or U5952 (N_5952,N_5717,N_5846);
or U5953 (N_5953,N_5702,N_5737);
or U5954 (N_5954,N_5785,N_5833);
and U5955 (N_5955,N_5747,N_5723);
and U5956 (N_5956,N_5781,N_5819);
xor U5957 (N_5957,N_5764,N_5718);
and U5958 (N_5958,N_5753,N_5760);
or U5959 (N_5959,N_5813,N_5717);
and U5960 (N_5960,N_5742,N_5823);
nand U5961 (N_5961,N_5728,N_5811);
nor U5962 (N_5962,N_5744,N_5730);
xor U5963 (N_5963,N_5781,N_5763);
xnor U5964 (N_5964,N_5777,N_5834);
nand U5965 (N_5965,N_5805,N_5831);
xor U5966 (N_5966,N_5771,N_5818);
or U5967 (N_5967,N_5758,N_5815);
xor U5968 (N_5968,N_5746,N_5787);
or U5969 (N_5969,N_5832,N_5735);
nand U5970 (N_5970,N_5806,N_5837);
nor U5971 (N_5971,N_5748,N_5731);
or U5972 (N_5972,N_5848,N_5837);
nor U5973 (N_5973,N_5768,N_5729);
xnor U5974 (N_5974,N_5825,N_5732);
xnor U5975 (N_5975,N_5823,N_5773);
nor U5976 (N_5976,N_5845,N_5735);
nor U5977 (N_5977,N_5812,N_5712);
xnor U5978 (N_5978,N_5707,N_5723);
nand U5979 (N_5979,N_5707,N_5703);
xor U5980 (N_5980,N_5723,N_5799);
nand U5981 (N_5981,N_5801,N_5812);
xor U5982 (N_5982,N_5750,N_5760);
xnor U5983 (N_5983,N_5815,N_5778);
nand U5984 (N_5984,N_5772,N_5744);
nor U5985 (N_5985,N_5801,N_5775);
nor U5986 (N_5986,N_5808,N_5703);
xor U5987 (N_5987,N_5764,N_5794);
xor U5988 (N_5988,N_5703,N_5813);
nor U5989 (N_5989,N_5727,N_5768);
nor U5990 (N_5990,N_5708,N_5762);
nor U5991 (N_5991,N_5772,N_5791);
nor U5992 (N_5992,N_5847,N_5839);
nor U5993 (N_5993,N_5845,N_5828);
nand U5994 (N_5994,N_5812,N_5732);
nor U5995 (N_5995,N_5803,N_5772);
and U5996 (N_5996,N_5716,N_5824);
xor U5997 (N_5997,N_5752,N_5769);
and U5998 (N_5998,N_5779,N_5734);
or U5999 (N_5999,N_5747,N_5840);
or U6000 (N_6000,N_5857,N_5988);
and U6001 (N_6001,N_5907,N_5903);
and U6002 (N_6002,N_5960,N_5976);
xnor U6003 (N_6003,N_5947,N_5889);
and U6004 (N_6004,N_5860,N_5872);
xnor U6005 (N_6005,N_5906,N_5966);
or U6006 (N_6006,N_5962,N_5929);
nand U6007 (N_6007,N_5922,N_5869);
and U6008 (N_6008,N_5891,N_5924);
or U6009 (N_6009,N_5990,N_5864);
xor U6010 (N_6010,N_5861,N_5865);
nor U6011 (N_6011,N_5913,N_5855);
xnor U6012 (N_6012,N_5925,N_5963);
nor U6013 (N_6013,N_5946,N_5868);
nand U6014 (N_6014,N_5863,N_5854);
and U6015 (N_6015,N_5984,N_5883);
nor U6016 (N_6016,N_5997,N_5888);
and U6017 (N_6017,N_5901,N_5985);
and U6018 (N_6018,N_5916,N_5926);
or U6019 (N_6019,N_5980,N_5944);
nor U6020 (N_6020,N_5853,N_5977);
nor U6021 (N_6021,N_5939,N_5887);
and U6022 (N_6022,N_5996,N_5897);
xor U6023 (N_6023,N_5957,N_5930);
or U6024 (N_6024,N_5974,N_5972);
nor U6025 (N_6025,N_5910,N_5895);
and U6026 (N_6026,N_5904,N_5923);
nand U6027 (N_6027,N_5933,N_5931);
nand U6028 (N_6028,N_5873,N_5870);
nand U6029 (N_6029,N_5973,N_5856);
or U6030 (N_6030,N_5890,N_5880);
or U6031 (N_6031,N_5919,N_5993);
nand U6032 (N_6032,N_5943,N_5859);
nor U6033 (N_6033,N_5852,N_5954);
nand U6034 (N_6034,N_5948,N_5937);
xnor U6035 (N_6035,N_5971,N_5942);
xor U6036 (N_6036,N_5940,N_5884);
or U6037 (N_6037,N_5945,N_5927);
xor U6038 (N_6038,N_5958,N_5979);
xnor U6039 (N_6039,N_5850,N_5885);
xnor U6040 (N_6040,N_5879,N_5967);
nand U6041 (N_6041,N_5982,N_5975);
nor U6042 (N_6042,N_5935,N_5991);
xnor U6043 (N_6043,N_5915,N_5914);
nor U6044 (N_6044,N_5998,N_5871);
and U6045 (N_6045,N_5886,N_5992);
nand U6046 (N_6046,N_5953,N_5983);
xnor U6047 (N_6047,N_5956,N_5858);
nand U6048 (N_6048,N_5909,N_5851);
and U6049 (N_6049,N_5898,N_5866);
nor U6050 (N_6050,N_5874,N_5881);
nor U6051 (N_6051,N_5911,N_5978);
nor U6052 (N_6052,N_5862,N_5892);
or U6053 (N_6053,N_5994,N_5936);
or U6054 (N_6054,N_5900,N_5964);
xnor U6055 (N_6055,N_5917,N_5968);
nor U6056 (N_6056,N_5961,N_5950);
nand U6057 (N_6057,N_5894,N_5918);
or U6058 (N_6058,N_5955,N_5969);
nand U6059 (N_6059,N_5912,N_5965);
nor U6060 (N_6060,N_5986,N_5896);
or U6061 (N_6061,N_5893,N_5920);
xor U6062 (N_6062,N_5949,N_5952);
and U6063 (N_6063,N_5999,N_5989);
and U6064 (N_6064,N_5938,N_5899);
and U6065 (N_6065,N_5867,N_5981);
nor U6066 (N_6066,N_5905,N_5877);
xor U6067 (N_6067,N_5908,N_5902);
nor U6068 (N_6068,N_5878,N_5928);
xor U6069 (N_6069,N_5882,N_5995);
or U6070 (N_6070,N_5959,N_5876);
nor U6071 (N_6071,N_5932,N_5970);
or U6072 (N_6072,N_5951,N_5875);
xnor U6073 (N_6073,N_5921,N_5934);
nor U6074 (N_6074,N_5987,N_5941);
nor U6075 (N_6075,N_5979,N_5850);
or U6076 (N_6076,N_5940,N_5953);
and U6077 (N_6077,N_5962,N_5984);
nand U6078 (N_6078,N_5896,N_5874);
and U6079 (N_6079,N_5853,N_5900);
nand U6080 (N_6080,N_5916,N_5896);
xnor U6081 (N_6081,N_5936,N_5894);
nand U6082 (N_6082,N_5874,N_5972);
nand U6083 (N_6083,N_5902,N_5974);
nand U6084 (N_6084,N_5867,N_5884);
nor U6085 (N_6085,N_5944,N_5914);
nor U6086 (N_6086,N_5922,N_5975);
xor U6087 (N_6087,N_5985,N_5851);
or U6088 (N_6088,N_5864,N_5950);
xnor U6089 (N_6089,N_5979,N_5944);
or U6090 (N_6090,N_5924,N_5887);
or U6091 (N_6091,N_5939,N_5883);
xor U6092 (N_6092,N_5861,N_5903);
xnor U6093 (N_6093,N_5979,N_5861);
xor U6094 (N_6094,N_5988,N_5883);
xnor U6095 (N_6095,N_5954,N_5893);
or U6096 (N_6096,N_5977,N_5917);
and U6097 (N_6097,N_5963,N_5948);
nor U6098 (N_6098,N_5878,N_5933);
nor U6099 (N_6099,N_5861,N_5854);
xnor U6100 (N_6100,N_5943,N_5868);
nor U6101 (N_6101,N_5866,N_5876);
and U6102 (N_6102,N_5853,N_5979);
nor U6103 (N_6103,N_5939,N_5983);
and U6104 (N_6104,N_5915,N_5872);
nor U6105 (N_6105,N_5873,N_5894);
and U6106 (N_6106,N_5977,N_5957);
nand U6107 (N_6107,N_5938,N_5954);
and U6108 (N_6108,N_5906,N_5970);
xnor U6109 (N_6109,N_5911,N_5980);
and U6110 (N_6110,N_5916,N_5972);
xnor U6111 (N_6111,N_5945,N_5982);
or U6112 (N_6112,N_5883,N_5915);
nor U6113 (N_6113,N_5850,N_5995);
xnor U6114 (N_6114,N_5915,N_5977);
or U6115 (N_6115,N_5955,N_5850);
nand U6116 (N_6116,N_5963,N_5926);
xnor U6117 (N_6117,N_5949,N_5947);
xnor U6118 (N_6118,N_5971,N_5950);
and U6119 (N_6119,N_5855,N_5859);
nor U6120 (N_6120,N_5868,N_5956);
and U6121 (N_6121,N_5962,N_5993);
xor U6122 (N_6122,N_5887,N_5880);
xnor U6123 (N_6123,N_5875,N_5974);
nand U6124 (N_6124,N_5873,N_5909);
nor U6125 (N_6125,N_5999,N_5886);
nor U6126 (N_6126,N_5850,N_5877);
or U6127 (N_6127,N_5893,N_5887);
nor U6128 (N_6128,N_5981,N_5889);
xnor U6129 (N_6129,N_5966,N_5984);
xnor U6130 (N_6130,N_5984,N_5854);
nor U6131 (N_6131,N_5941,N_5858);
xnor U6132 (N_6132,N_5961,N_5995);
xor U6133 (N_6133,N_5967,N_5984);
nand U6134 (N_6134,N_5996,N_5882);
and U6135 (N_6135,N_5924,N_5966);
or U6136 (N_6136,N_5953,N_5942);
and U6137 (N_6137,N_5956,N_5856);
and U6138 (N_6138,N_5869,N_5893);
and U6139 (N_6139,N_5979,N_5904);
or U6140 (N_6140,N_5986,N_5868);
xor U6141 (N_6141,N_5980,N_5965);
nor U6142 (N_6142,N_5911,N_5974);
nand U6143 (N_6143,N_5933,N_5873);
or U6144 (N_6144,N_5901,N_5990);
nor U6145 (N_6145,N_5889,N_5942);
nand U6146 (N_6146,N_5956,N_5979);
nor U6147 (N_6147,N_5911,N_5948);
nand U6148 (N_6148,N_5947,N_5930);
nor U6149 (N_6149,N_5851,N_5971);
and U6150 (N_6150,N_6066,N_6026);
nand U6151 (N_6151,N_6079,N_6136);
nand U6152 (N_6152,N_6134,N_6008);
xor U6153 (N_6153,N_6023,N_6055);
nand U6154 (N_6154,N_6046,N_6099);
nand U6155 (N_6155,N_6103,N_6025);
nand U6156 (N_6156,N_6137,N_6140);
and U6157 (N_6157,N_6126,N_6059);
and U6158 (N_6158,N_6132,N_6115);
nand U6159 (N_6159,N_6074,N_6105);
nor U6160 (N_6160,N_6123,N_6147);
nand U6161 (N_6161,N_6083,N_6118);
nor U6162 (N_6162,N_6065,N_6130);
xnor U6163 (N_6163,N_6119,N_6011);
xnor U6164 (N_6164,N_6052,N_6091);
xnor U6165 (N_6165,N_6145,N_6015);
nor U6166 (N_6166,N_6106,N_6019);
xor U6167 (N_6167,N_6043,N_6014);
xnor U6168 (N_6168,N_6100,N_6024);
and U6169 (N_6169,N_6009,N_6050);
xnor U6170 (N_6170,N_6138,N_6064);
nor U6171 (N_6171,N_6040,N_6030);
xor U6172 (N_6172,N_6117,N_6113);
or U6173 (N_6173,N_6000,N_6139);
or U6174 (N_6174,N_6036,N_6054);
and U6175 (N_6175,N_6037,N_6101);
or U6176 (N_6176,N_6095,N_6144);
nand U6177 (N_6177,N_6063,N_6135);
or U6178 (N_6178,N_6068,N_6047);
nand U6179 (N_6179,N_6120,N_6069);
and U6180 (N_6180,N_6114,N_6097);
or U6181 (N_6181,N_6092,N_6041);
nand U6182 (N_6182,N_6027,N_6022);
nand U6183 (N_6183,N_6057,N_6044);
or U6184 (N_6184,N_6004,N_6042);
and U6185 (N_6185,N_6078,N_6010);
or U6186 (N_6186,N_6127,N_6001);
nand U6187 (N_6187,N_6032,N_6107);
and U6188 (N_6188,N_6094,N_6020);
nor U6189 (N_6189,N_6016,N_6072);
xnor U6190 (N_6190,N_6096,N_6076);
nor U6191 (N_6191,N_6141,N_6033);
nor U6192 (N_6192,N_6090,N_6143);
nor U6193 (N_6193,N_6031,N_6039);
nor U6194 (N_6194,N_6070,N_6116);
nand U6195 (N_6195,N_6049,N_6077);
xor U6196 (N_6196,N_6128,N_6111);
and U6197 (N_6197,N_6034,N_6002);
or U6198 (N_6198,N_6075,N_6131);
xnor U6199 (N_6199,N_6082,N_6067);
and U6200 (N_6200,N_6048,N_6029);
or U6201 (N_6201,N_6021,N_6035);
and U6202 (N_6202,N_6003,N_6089);
or U6203 (N_6203,N_6102,N_6084);
xor U6204 (N_6204,N_6017,N_6098);
xor U6205 (N_6205,N_6045,N_6142);
nor U6206 (N_6206,N_6080,N_6129);
xor U6207 (N_6207,N_6088,N_6007);
and U6208 (N_6208,N_6110,N_6028);
or U6209 (N_6209,N_6146,N_6133);
nand U6210 (N_6210,N_6093,N_6018);
or U6211 (N_6211,N_6013,N_6149);
nand U6212 (N_6212,N_6112,N_6053);
and U6213 (N_6213,N_6104,N_6012);
nor U6214 (N_6214,N_6108,N_6058);
nand U6215 (N_6215,N_6086,N_6006);
nand U6216 (N_6216,N_6081,N_6071);
and U6217 (N_6217,N_6056,N_6087);
or U6218 (N_6218,N_6085,N_6148);
xor U6219 (N_6219,N_6062,N_6125);
or U6220 (N_6220,N_6038,N_6051);
xnor U6221 (N_6221,N_6005,N_6124);
nor U6222 (N_6222,N_6109,N_6060);
xnor U6223 (N_6223,N_6122,N_6061);
or U6224 (N_6224,N_6073,N_6121);
and U6225 (N_6225,N_6059,N_6032);
nand U6226 (N_6226,N_6089,N_6052);
and U6227 (N_6227,N_6041,N_6062);
or U6228 (N_6228,N_6033,N_6012);
nor U6229 (N_6229,N_6110,N_6029);
or U6230 (N_6230,N_6109,N_6039);
nand U6231 (N_6231,N_6060,N_6135);
nor U6232 (N_6232,N_6078,N_6134);
nand U6233 (N_6233,N_6123,N_6105);
and U6234 (N_6234,N_6002,N_6041);
and U6235 (N_6235,N_6119,N_6149);
xor U6236 (N_6236,N_6016,N_6083);
xnor U6237 (N_6237,N_6073,N_6052);
nor U6238 (N_6238,N_6132,N_6048);
nor U6239 (N_6239,N_6004,N_6003);
and U6240 (N_6240,N_6143,N_6062);
xor U6241 (N_6241,N_6086,N_6090);
and U6242 (N_6242,N_6023,N_6119);
nand U6243 (N_6243,N_6027,N_6025);
nor U6244 (N_6244,N_6067,N_6004);
nand U6245 (N_6245,N_6062,N_6054);
nand U6246 (N_6246,N_6063,N_6084);
xnor U6247 (N_6247,N_6084,N_6085);
nor U6248 (N_6248,N_6134,N_6143);
and U6249 (N_6249,N_6114,N_6127);
and U6250 (N_6250,N_6099,N_6032);
or U6251 (N_6251,N_6141,N_6121);
nor U6252 (N_6252,N_6053,N_6049);
or U6253 (N_6253,N_6010,N_6022);
nor U6254 (N_6254,N_6006,N_6071);
nor U6255 (N_6255,N_6016,N_6088);
nand U6256 (N_6256,N_6009,N_6041);
nor U6257 (N_6257,N_6071,N_6020);
nor U6258 (N_6258,N_6114,N_6106);
nand U6259 (N_6259,N_6147,N_6115);
and U6260 (N_6260,N_6109,N_6080);
nor U6261 (N_6261,N_6135,N_6082);
xnor U6262 (N_6262,N_6047,N_6053);
or U6263 (N_6263,N_6147,N_6062);
and U6264 (N_6264,N_6148,N_6067);
xnor U6265 (N_6265,N_6018,N_6090);
and U6266 (N_6266,N_6079,N_6142);
xor U6267 (N_6267,N_6044,N_6042);
xor U6268 (N_6268,N_6022,N_6071);
nor U6269 (N_6269,N_6107,N_6069);
nor U6270 (N_6270,N_6000,N_6012);
and U6271 (N_6271,N_6146,N_6119);
and U6272 (N_6272,N_6149,N_6002);
nand U6273 (N_6273,N_6142,N_6086);
or U6274 (N_6274,N_6010,N_6054);
nand U6275 (N_6275,N_6117,N_6034);
or U6276 (N_6276,N_6057,N_6012);
nand U6277 (N_6277,N_6062,N_6059);
nand U6278 (N_6278,N_6075,N_6143);
nand U6279 (N_6279,N_6104,N_6046);
and U6280 (N_6280,N_6124,N_6086);
xor U6281 (N_6281,N_6007,N_6011);
or U6282 (N_6282,N_6041,N_6013);
and U6283 (N_6283,N_6148,N_6001);
or U6284 (N_6284,N_6057,N_6101);
xor U6285 (N_6285,N_6002,N_6032);
xnor U6286 (N_6286,N_6133,N_6051);
nor U6287 (N_6287,N_6083,N_6112);
nor U6288 (N_6288,N_6053,N_6021);
nand U6289 (N_6289,N_6035,N_6080);
nor U6290 (N_6290,N_6105,N_6092);
and U6291 (N_6291,N_6009,N_6028);
and U6292 (N_6292,N_6118,N_6124);
or U6293 (N_6293,N_6130,N_6056);
and U6294 (N_6294,N_6010,N_6113);
or U6295 (N_6295,N_6075,N_6073);
or U6296 (N_6296,N_6051,N_6005);
nand U6297 (N_6297,N_6071,N_6100);
xnor U6298 (N_6298,N_6002,N_6113);
xor U6299 (N_6299,N_6021,N_6114);
or U6300 (N_6300,N_6246,N_6288);
nor U6301 (N_6301,N_6215,N_6290);
and U6302 (N_6302,N_6196,N_6202);
nor U6303 (N_6303,N_6221,N_6199);
xor U6304 (N_6304,N_6225,N_6179);
and U6305 (N_6305,N_6182,N_6240);
and U6306 (N_6306,N_6262,N_6204);
xor U6307 (N_6307,N_6238,N_6211);
nor U6308 (N_6308,N_6227,N_6271);
and U6309 (N_6309,N_6255,N_6224);
or U6310 (N_6310,N_6188,N_6237);
nand U6311 (N_6311,N_6294,N_6181);
nor U6312 (N_6312,N_6287,N_6193);
nand U6313 (N_6313,N_6207,N_6241);
nor U6314 (N_6314,N_6216,N_6169);
nand U6315 (N_6315,N_6158,N_6212);
or U6316 (N_6316,N_6164,N_6279);
or U6317 (N_6317,N_6235,N_6254);
and U6318 (N_6318,N_6257,N_6239);
and U6319 (N_6319,N_6171,N_6285);
xnor U6320 (N_6320,N_6150,N_6208);
xnor U6321 (N_6321,N_6163,N_6242);
or U6322 (N_6322,N_6289,N_6151);
nand U6323 (N_6323,N_6296,N_6186);
nor U6324 (N_6324,N_6190,N_6213);
nand U6325 (N_6325,N_6275,N_6209);
and U6326 (N_6326,N_6201,N_6172);
or U6327 (N_6327,N_6205,N_6286);
and U6328 (N_6328,N_6268,N_6206);
nand U6329 (N_6329,N_6219,N_6234);
nor U6330 (N_6330,N_6230,N_6261);
xor U6331 (N_6331,N_6197,N_6270);
nand U6332 (N_6332,N_6267,N_6249);
or U6333 (N_6333,N_6167,N_6177);
xor U6334 (N_6334,N_6191,N_6168);
xor U6335 (N_6335,N_6252,N_6282);
xor U6336 (N_6336,N_6173,N_6165);
nor U6337 (N_6337,N_6170,N_6272);
nand U6338 (N_6338,N_6217,N_6231);
nor U6339 (N_6339,N_6229,N_6187);
and U6340 (N_6340,N_6274,N_6183);
nand U6341 (N_6341,N_6264,N_6298);
and U6342 (N_6342,N_6218,N_6233);
and U6343 (N_6343,N_6283,N_6281);
nor U6344 (N_6344,N_6260,N_6160);
xor U6345 (N_6345,N_6276,N_6161);
nand U6346 (N_6346,N_6156,N_6266);
and U6347 (N_6347,N_6210,N_6256);
xnor U6348 (N_6348,N_6159,N_6176);
or U6349 (N_6349,N_6189,N_6154);
nand U6350 (N_6350,N_6175,N_6295);
nand U6351 (N_6351,N_6259,N_6299);
xnor U6352 (N_6352,N_6244,N_6198);
xor U6353 (N_6353,N_6245,N_6214);
and U6354 (N_6354,N_6166,N_6152);
nor U6355 (N_6355,N_6155,N_6226);
nand U6356 (N_6356,N_6297,N_6269);
and U6357 (N_6357,N_6280,N_6273);
nor U6358 (N_6358,N_6293,N_6243);
and U6359 (N_6359,N_6153,N_6292);
nand U6360 (N_6360,N_6180,N_6195);
and U6361 (N_6361,N_6185,N_6174);
and U6362 (N_6362,N_6291,N_6162);
nor U6363 (N_6363,N_6248,N_6277);
xor U6364 (N_6364,N_6228,N_6247);
and U6365 (N_6365,N_6192,N_6157);
and U6366 (N_6366,N_6284,N_6278);
and U6367 (N_6367,N_6184,N_6223);
nor U6368 (N_6368,N_6220,N_6236);
nand U6369 (N_6369,N_6253,N_6250);
and U6370 (N_6370,N_6258,N_6200);
xor U6371 (N_6371,N_6194,N_6178);
and U6372 (N_6372,N_6222,N_6232);
nor U6373 (N_6373,N_6263,N_6203);
xor U6374 (N_6374,N_6251,N_6265);
nor U6375 (N_6375,N_6264,N_6268);
or U6376 (N_6376,N_6218,N_6196);
nand U6377 (N_6377,N_6291,N_6278);
nor U6378 (N_6378,N_6220,N_6228);
nor U6379 (N_6379,N_6263,N_6264);
and U6380 (N_6380,N_6263,N_6253);
xor U6381 (N_6381,N_6256,N_6227);
nor U6382 (N_6382,N_6245,N_6150);
and U6383 (N_6383,N_6195,N_6262);
nor U6384 (N_6384,N_6228,N_6198);
and U6385 (N_6385,N_6290,N_6279);
nand U6386 (N_6386,N_6229,N_6151);
xor U6387 (N_6387,N_6223,N_6189);
nor U6388 (N_6388,N_6189,N_6256);
and U6389 (N_6389,N_6224,N_6188);
xor U6390 (N_6390,N_6213,N_6155);
or U6391 (N_6391,N_6287,N_6232);
and U6392 (N_6392,N_6214,N_6297);
xor U6393 (N_6393,N_6178,N_6264);
or U6394 (N_6394,N_6205,N_6190);
or U6395 (N_6395,N_6174,N_6272);
xnor U6396 (N_6396,N_6234,N_6255);
and U6397 (N_6397,N_6185,N_6159);
nand U6398 (N_6398,N_6179,N_6176);
xnor U6399 (N_6399,N_6219,N_6189);
or U6400 (N_6400,N_6234,N_6293);
nor U6401 (N_6401,N_6299,N_6208);
xor U6402 (N_6402,N_6299,N_6297);
or U6403 (N_6403,N_6246,N_6250);
nor U6404 (N_6404,N_6175,N_6183);
and U6405 (N_6405,N_6203,N_6174);
nand U6406 (N_6406,N_6290,N_6294);
nor U6407 (N_6407,N_6272,N_6259);
nand U6408 (N_6408,N_6196,N_6191);
nand U6409 (N_6409,N_6265,N_6157);
nor U6410 (N_6410,N_6297,N_6178);
nand U6411 (N_6411,N_6185,N_6166);
and U6412 (N_6412,N_6152,N_6250);
xor U6413 (N_6413,N_6287,N_6242);
or U6414 (N_6414,N_6253,N_6212);
or U6415 (N_6415,N_6223,N_6222);
nor U6416 (N_6416,N_6161,N_6208);
nand U6417 (N_6417,N_6283,N_6152);
or U6418 (N_6418,N_6155,N_6282);
and U6419 (N_6419,N_6277,N_6280);
and U6420 (N_6420,N_6184,N_6272);
or U6421 (N_6421,N_6277,N_6284);
nand U6422 (N_6422,N_6219,N_6281);
and U6423 (N_6423,N_6204,N_6174);
or U6424 (N_6424,N_6263,N_6208);
or U6425 (N_6425,N_6242,N_6219);
nor U6426 (N_6426,N_6281,N_6254);
or U6427 (N_6427,N_6289,N_6191);
nor U6428 (N_6428,N_6162,N_6219);
nand U6429 (N_6429,N_6220,N_6231);
xor U6430 (N_6430,N_6216,N_6262);
xor U6431 (N_6431,N_6184,N_6192);
nor U6432 (N_6432,N_6260,N_6221);
or U6433 (N_6433,N_6284,N_6219);
and U6434 (N_6434,N_6228,N_6158);
and U6435 (N_6435,N_6274,N_6201);
or U6436 (N_6436,N_6151,N_6203);
nor U6437 (N_6437,N_6263,N_6194);
xnor U6438 (N_6438,N_6182,N_6166);
or U6439 (N_6439,N_6201,N_6288);
xnor U6440 (N_6440,N_6201,N_6234);
nand U6441 (N_6441,N_6262,N_6238);
or U6442 (N_6442,N_6201,N_6179);
nor U6443 (N_6443,N_6277,N_6210);
nor U6444 (N_6444,N_6215,N_6276);
or U6445 (N_6445,N_6151,N_6168);
nand U6446 (N_6446,N_6216,N_6242);
and U6447 (N_6447,N_6193,N_6150);
xnor U6448 (N_6448,N_6165,N_6223);
nor U6449 (N_6449,N_6245,N_6268);
or U6450 (N_6450,N_6392,N_6443);
and U6451 (N_6451,N_6363,N_6368);
and U6452 (N_6452,N_6356,N_6312);
and U6453 (N_6453,N_6409,N_6406);
or U6454 (N_6454,N_6400,N_6426);
xor U6455 (N_6455,N_6313,N_6348);
and U6456 (N_6456,N_6415,N_6387);
nor U6457 (N_6457,N_6414,N_6435);
or U6458 (N_6458,N_6314,N_6413);
nor U6459 (N_6459,N_6304,N_6411);
and U6460 (N_6460,N_6326,N_6359);
xnor U6461 (N_6461,N_6369,N_6315);
and U6462 (N_6462,N_6332,N_6382);
nand U6463 (N_6463,N_6353,N_6333);
xor U6464 (N_6464,N_6378,N_6425);
or U6465 (N_6465,N_6319,N_6335);
or U6466 (N_6466,N_6343,N_6432);
or U6467 (N_6467,N_6419,N_6376);
or U6468 (N_6468,N_6323,N_6385);
nor U6469 (N_6469,N_6324,N_6345);
or U6470 (N_6470,N_6427,N_6441);
xnor U6471 (N_6471,N_6444,N_6377);
nand U6472 (N_6472,N_6311,N_6430);
xnor U6473 (N_6473,N_6307,N_6375);
nor U6474 (N_6474,N_6303,N_6437);
or U6475 (N_6475,N_6418,N_6317);
nor U6476 (N_6476,N_6398,N_6438);
nor U6477 (N_6477,N_6408,N_6320);
nor U6478 (N_6478,N_6397,N_6399);
and U6479 (N_6479,N_6394,N_6349);
nand U6480 (N_6480,N_6440,N_6402);
xor U6481 (N_6481,N_6416,N_6330);
xnor U6482 (N_6482,N_6395,N_6449);
nand U6483 (N_6483,N_6423,N_6322);
nor U6484 (N_6484,N_6391,N_6321);
nor U6485 (N_6485,N_6338,N_6439);
or U6486 (N_6486,N_6355,N_6360);
and U6487 (N_6487,N_6344,N_6352);
nor U6488 (N_6488,N_6421,N_6329);
or U6489 (N_6489,N_6300,N_6340);
nor U6490 (N_6490,N_6350,N_6389);
or U6491 (N_6491,N_6370,N_6366);
nand U6492 (N_6492,N_6401,N_6361);
xor U6493 (N_6493,N_6388,N_6424);
nor U6494 (N_6494,N_6396,N_6405);
or U6495 (N_6495,N_6373,N_6407);
or U6496 (N_6496,N_6364,N_6384);
or U6497 (N_6497,N_6316,N_6433);
nor U6498 (N_6498,N_6337,N_6339);
xnor U6499 (N_6499,N_6417,N_6428);
and U6500 (N_6500,N_6434,N_6346);
or U6501 (N_6501,N_6445,N_6310);
xor U6502 (N_6502,N_6436,N_6442);
nor U6503 (N_6503,N_6420,N_6404);
nand U6504 (N_6504,N_6390,N_6380);
nor U6505 (N_6505,N_6429,N_6393);
nor U6506 (N_6506,N_6306,N_6308);
and U6507 (N_6507,N_6412,N_6302);
and U6508 (N_6508,N_6367,N_6372);
or U6509 (N_6509,N_6357,N_6365);
and U6510 (N_6510,N_6447,N_6328);
or U6511 (N_6511,N_6347,N_6331);
nand U6512 (N_6512,N_6305,N_6422);
or U6513 (N_6513,N_6379,N_6325);
or U6514 (N_6514,N_6358,N_6351);
nor U6515 (N_6515,N_6410,N_6362);
and U6516 (N_6516,N_6383,N_6301);
xnor U6517 (N_6517,N_6341,N_6334);
nor U6518 (N_6518,N_6327,N_6381);
and U6519 (N_6519,N_6448,N_6374);
nor U6520 (N_6520,N_6336,N_6446);
nand U6521 (N_6521,N_6342,N_6318);
xnor U6522 (N_6522,N_6403,N_6431);
xnor U6523 (N_6523,N_6354,N_6386);
and U6524 (N_6524,N_6309,N_6371);
or U6525 (N_6525,N_6348,N_6433);
and U6526 (N_6526,N_6402,N_6344);
nor U6527 (N_6527,N_6301,N_6434);
xor U6528 (N_6528,N_6447,N_6361);
nor U6529 (N_6529,N_6310,N_6391);
and U6530 (N_6530,N_6392,N_6423);
and U6531 (N_6531,N_6432,N_6412);
nor U6532 (N_6532,N_6424,N_6413);
xor U6533 (N_6533,N_6376,N_6380);
xor U6534 (N_6534,N_6414,N_6301);
and U6535 (N_6535,N_6340,N_6368);
xor U6536 (N_6536,N_6302,N_6338);
xor U6537 (N_6537,N_6304,N_6410);
nand U6538 (N_6538,N_6375,N_6347);
xor U6539 (N_6539,N_6338,N_6309);
and U6540 (N_6540,N_6376,N_6375);
nor U6541 (N_6541,N_6364,N_6348);
xnor U6542 (N_6542,N_6406,N_6387);
xnor U6543 (N_6543,N_6358,N_6406);
nor U6544 (N_6544,N_6423,N_6442);
nand U6545 (N_6545,N_6439,N_6372);
and U6546 (N_6546,N_6327,N_6443);
nand U6547 (N_6547,N_6413,N_6312);
xor U6548 (N_6548,N_6305,N_6344);
xor U6549 (N_6549,N_6357,N_6380);
nor U6550 (N_6550,N_6374,N_6443);
nor U6551 (N_6551,N_6360,N_6307);
nand U6552 (N_6552,N_6421,N_6440);
nand U6553 (N_6553,N_6407,N_6329);
or U6554 (N_6554,N_6384,N_6310);
and U6555 (N_6555,N_6416,N_6304);
and U6556 (N_6556,N_6303,N_6434);
and U6557 (N_6557,N_6375,N_6301);
nor U6558 (N_6558,N_6414,N_6316);
or U6559 (N_6559,N_6316,N_6307);
or U6560 (N_6560,N_6332,N_6337);
nor U6561 (N_6561,N_6410,N_6313);
or U6562 (N_6562,N_6402,N_6328);
and U6563 (N_6563,N_6329,N_6403);
xnor U6564 (N_6564,N_6350,N_6368);
and U6565 (N_6565,N_6321,N_6405);
xor U6566 (N_6566,N_6367,N_6346);
xnor U6567 (N_6567,N_6327,N_6305);
nand U6568 (N_6568,N_6403,N_6379);
and U6569 (N_6569,N_6414,N_6359);
nor U6570 (N_6570,N_6446,N_6380);
nand U6571 (N_6571,N_6371,N_6311);
nand U6572 (N_6572,N_6405,N_6410);
xnor U6573 (N_6573,N_6408,N_6328);
xor U6574 (N_6574,N_6390,N_6417);
and U6575 (N_6575,N_6322,N_6309);
xor U6576 (N_6576,N_6388,N_6414);
or U6577 (N_6577,N_6333,N_6370);
xnor U6578 (N_6578,N_6369,N_6375);
and U6579 (N_6579,N_6397,N_6417);
or U6580 (N_6580,N_6357,N_6419);
nor U6581 (N_6581,N_6445,N_6354);
nand U6582 (N_6582,N_6433,N_6304);
or U6583 (N_6583,N_6381,N_6440);
nand U6584 (N_6584,N_6372,N_6423);
nor U6585 (N_6585,N_6315,N_6371);
and U6586 (N_6586,N_6427,N_6340);
nand U6587 (N_6587,N_6377,N_6361);
nor U6588 (N_6588,N_6319,N_6412);
xor U6589 (N_6589,N_6427,N_6356);
nand U6590 (N_6590,N_6448,N_6402);
nand U6591 (N_6591,N_6394,N_6364);
and U6592 (N_6592,N_6442,N_6432);
or U6593 (N_6593,N_6419,N_6439);
and U6594 (N_6594,N_6310,N_6308);
or U6595 (N_6595,N_6433,N_6399);
and U6596 (N_6596,N_6417,N_6355);
nand U6597 (N_6597,N_6432,N_6441);
nand U6598 (N_6598,N_6387,N_6363);
nand U6599 (N_6599,N_6406,N_6335);
nand U6600 (N_6600,N_6555,N_6552);
nand U6601 (N_6601,N_6542,N_6534);
nand U6602 (N_6602,N_6549,N_6509);
nand U6603 (N_6603,N_6516,N_6521);
xnor U6604 (N_6604,N_6452,N_6487);
or U6605 (N_6605,N_6590,N_6491);
nor U6606 (N_6606,N_6507,N_6529);
or U6607 (N_6607,N_6512,N_6515);
xnor U6608 (N_6608,N_6484,N_6556);
xor U6609 (N_6609,N_6559,N_6470);
or U6610 (N_6610,N_6540,N_6458);
nor U6611 (N_6611,N_6535,N_6577);
xnor U6612 (N_6612,N_6573,N_6459);
and U6613 (N_6613,N_6455,N_6465);
and U6614 (N_6614,N_6533,N_6596);
or U6615 (N_6615,N_6494,N_6492);
and U6616 (N_6616,N_6469,N_6499);
or U6617 (N_6617,N_6593,N_6550);
and U6618 (N_6618,N_6576,N_6497);
and U6619 (N_6619,N_6504,N_6500);
nor U6620 (N_6620,N_6514,N_6548);
and U6621 (N_6621,N_6502,N_6486);
and U6622 (N_6622,N_6511,N_6518);
xor U6623 (N_6623,N_6451,N_6572);
nor U6624 (N_6624,N_6546,N_6510);
nor U6625 (N_6625,N_6571,N_6537);
nor U6626 (N_6626,N_6592,N_6583);
nor U6627 (N_6627,N_6508,N_6477);
and U6628 (N_6628,N_6586,N_6489);
xor U6629 (N_6629,N_6581,N_6562);
nand U6630 (N_6630,N_6493,N_6523);
nand U6631 (N_6631,N_6597,N_6563);
and U6632 (N_6632,N_6454,N_6566);
nand U6633 (N_6633,N_6463,N_6575);
and U6634 (N_6634,N_6589,N_6578);
nor U6635 (N_6635,N_6587,N_6560);
nand U6636 (N_6636,N_6564,N_6478);
nor U6637 (N_6637,N_6539,N_6528);
nor U6638 (N_6638,N_6545,N_6482);
nor U6639 (N_6639,N_6517,N_6570);
and U6640 (N_6640,N_6595,N_6591);
and U6641 (N_6641,N_6544,N_6580);
nand U6642 (N_6642,N_6574,N_6468);
nor U6643 (N_6643,N_6488,N_6579);
nor U6644 (N_6644,N_6519,N_6473);
nand U6645 (N_6645,N_6466,N_6490);
xnor U6646 (N_6646,N_6496,N_6485);
xnor U6647 (N_6647,N_6584,N_6457);
xnor U6648 (N_6648,N_6456,N_6503);
xor U6649 (N_6649,N_6464,N_6475);
nand U6650 (N_6650,N_6554,N_6524);
nor U6651 (N_6651,N_6480,N_6495);
or U6652 (N_6652,N_6594,N_6471);
or U6653 (N_6653,N_6526,N_6551);
nand U6654 (N_6654,N_6513,N_6557);
and U6655 (N_6655,N_6476,N_6536);
and U6656 (N_6656,N_6450,N_6585);
xnor U6657 (N_6657,N_6472,N_6527);
nor U6658 (N_6658,N_6474,N_6525);
and U6659 (N_6659,N_6498,N_6479);
and U6660 (N_6660,N_6532,N_6568);
or U6661 (N_6661,N_6553,N_6453);
nand U6662 (N_6662,N_6582,N_6531);
and U6663 (N_6663,N_6561,N_6483);
xnor U6664 (N_6664,N_6467,N_6481);
nand U6665 (N_6665,N_6558,N_6567);
nor U6666 (N_6666,N_6547,N_6520);
xnor U6667 (N_6667,N_6462,N_6538);
or U6668 (N_6668,N_6588,N_6598);
nor U6669 (N_6669,N_6543,N_6565);
or U6670 (N_6670,N_6530,N_6599);
nand U6671 (N_6671,N_6541,N_6460);
nand U6672 (N_6672,N_6569,N_6506);
xnor U6673 (N_6673,N_6505,N_6461);
and U6674 (N_6674,N_6522,N_6501);
or U6675 (N_6675,N_6534,N_6548);
nor U6676 (N_6676,N_6496,N_6507);
and U6677 (N_6677,N_6502,N_6514);
and U6678 (N_6678,N_6529,N_6551);
and U6679 (N_6679,N_6569,N_6510);
or U6680 (N_6680,N_6509,N_6467);
xnor U6681 (N_6681,N_6582,N_6575);
xor U6682 (N_6682,N_6591,N_6526);
nor U6683 (N_6683,N_6588,N_6477);
nand U6684 (N_6684,N_6534,N_6452);
or U6685 (N_6685,N_6451,N_6525);
xnor U6686 (N_6686,N_6469,N_6541);
and U6687 (N_6687,N_6501,N_6519);
and U6688 (N_6688,N_6450,N_6589);
or U6689 (N_6689,N_6560,N_6538);
and U6690 (N_6690,N_6544,N_6585);
and U6691 (N_6691,N_6537,N_6548);
xnor U6692 (N_6692,N_6590,N_6578);
nor U6693 (N_6693,N_6531,N_6512);
nor U6694 (N_6694,N_6596,N_6492);
nand U6695 (N_6695,N_6481,N_6454);
or U6696 (N_6696,N_6568,N_6455);
nand U6697 (N_6697,N_6557,N_6532);
nor U6698 (N_6698,N_6583,N_6562);
or U6699 (N_6699,N_6510,N_6571);
or U6700 (N_6700,N_6559,N_6503);
nand U6701 (N_6701,N_6538,N_6485);
or U6702 (N_6702,N_6582,N_6566);
and U6703 (N_6703,N_6556,N_6462);
nor U6704 (N_6704,N_6454,N_6577);
xnor U6705 (N_6705,N_6511,N_6490);
or U6706 (N_6706,N_6476,N_6565);
nor U6707 (N_6707,N_6554,N_6534);
nor U6708 (N_6708,N_6541,N_6548);
or U6709 (N_6709,N_6538,N_6564);
nor U6710 (N_6710,N_6477,N_6527);
nor U6711 (N_6711,N_6494,N_6498);
and U6712 (N_6712,N_6497,N_6552);
nand U6713 (N_6713,N_6565,N_6475);
nor U6714 (N_6714,N_6484,N_6474);
or U6715 (N_6715,N_6519,N_6514);
and U6716 (N_6716,N_6588,N_6565);
xnor U6717 (N_6717,N_6579,N_6517);
or U6718 (N_6718,N_6468,N_6479);
or U6719 (N_6719,N_6495,N_6469);
xor U6720 (N_6720,N_6550,N_6471);
and U6721 (N_6721,N_6473,N_6578);
and U6722 (N_6722,N_6543,N_6521);
xnor U6723 (N_6723,N_6592,N_6544);
xor U6724 (N_6724,N_6566,N_6515);
or U6725 (N_6725,N_6511,N_6503);
or U6726 (N_6726,N_6484,N_6547);
xor U6727 (N_6727,N_6590,N_6473);
xor U6728 (N_6728,N_6593,N_6561);
and U6729 (N_6729,N_6554,N_6463);
nor U6730 (N_6730,N_6471,N_6470);
and U6731 (N_6731,N_6481,N_6582);
nand U6732 (N_6732,N_6571,N_6548);
nand U6733 (N_6733,N_6486,N_6524);
nand U6734 (N_6734,N_6540,N_6484);
and U6735 (N_6735,N_6579,N_6553);
nor U6736 (N_6736,N_6542,N_6466);
and U6737 (N_6737,N_6499,N_6477);
xor U6738 (N_6738,N_6474,N_6559);
and U6739 (N_6739,N_6596,N_6565);
xnor U6740 (N_6740,N_6576,N_6519);
nor U6741 (N_6741,N_6518,N_6484);
nand U6742 (N_6742,N_6586,N_6594);
or U6743 (N_6743,N_6455,N_6452);
nand U6744 (N_6744,N_6459,N_6507);
nor U6745 (N_6745,N_6571,N_6497);
or U6746 (N_6746,N_6565,N_6467);
or U6747 (N_6747,N_6518,N_6526);
or U6748 (N_6748,N_6462,N_6586);
and U6749 (N_6749,N_6485,N_6511);
and U6750 (N_6750,N_6613,N_6648);
or U6751 (N_6751,N_6611,N_6624);
and U6752 (N_6752,N_6628,N_6688);
xor U6753 (N_6753,N_6627,N_6739);
nor U6754 (N_6754,N_6747,N_6608);
xnor U6755 (N_6755,N_6707,N_6717);
nor U6756 (N_6756,N_6749,N_6643);
nor U6757 (N_6757,N_6649,N_6603);
and U6758 (N_6758,N_6661,N_6697);
nand U6759 (N_6759,N_6715,N_6675);
xnor U6760 (N_6760,N_6635,N_6653);
nor U6761 (N_6761,N_6736,N_6638);
nor U6762 (N_6762,N_6656,N_6623);
and U6763 (N_6763,N_6696,N_6719);
nand U6764 (N_6764,N_6651,N_6704);
xnor U6765 (N_6765,N_6732,N_6742);
or U6766 (N_6766,N_6733,N_6601);
nand U6767 (N_6767,N_6659,N_6657);
nor U6768 (N_6768,N_6668,N_6720);
or U6769 (N_6769,N_6600,N_6722);
and U6770 (N_6770,N_6620,N_6641);
or U6771 (N_6771,N_6701,N_6691);
or U6772 (N_6772,N_6738,N_6626);
and U6773 (N_6773,N_6693,N_6676);
nand U6774 (N_6774,N_6734,N_6702);
nand U6775 (N_6775,N_6618,N_6724);
nor U6776 (N_6776,N_6607,N_6729);
xnor U6777 (N_6777,N_6740,N_6622);
nor U6778 (N_6778,N_6670,N_6714);
nand U6779 (N_6779,N_6671,N_6652);
or U6780 (N_6780,N_6746,N_6687);
and U6781 (N_6781,N_6725,N_6726);
xnor U6782 (N_6782,N_6718,N_6748);
or U6783 (N_6783,N_6713,N_6679);
and U6784 (N_6784,N_6674,N_6602);
or U6785 (N_6785,N_6619,N_6604);
nand U6786 (N_6786,N_6721,N_6728);
or U6787 (N_6787,N_6642,N_6632);
nor U6788 (N_6788,N_6654,N_6612);
and U6789 (N_6789,N_6684,N_6636);
or U6790 (N_6790,N_6686,N_6731);
nor U6791 (N_6791,N_6614,N_6711);
and U6792 (N_6792,N_6699,N_6655);
and U6793 (N_6793,N_6667,N_6700);
xor U6794 (N_6794,N_6744,N_6669);
nor U6795 (N_6795,N_6663,N_6683);
xnor U6796 (N_6796,N_6645,N_6605);
nand U6797 (N_6797,N_6621,N_6616);
and U6798 (N_6798,N_6709,N_6708);
nand U6799 (N_6799,N_6662,N_6609);
and U6800 (N_6800,N_6615,N_6666);
nor U6801 (N_6801,N_6640,N_6658);
nand U6802 (N_6802,N_6617,N_6606);
xor U6803 (N_6803,N_6673,N_6625);
xor U6804 (N_6804,N_6672,N_6639);
or U6805 (N_6805,N_6694,N_6716);
nor U6806 (N_6806,N_6690,N_6650);
or U6807 (N_6807,N_6743,N_6741);
xnor U6808 (N_6808,N_6705,N_6682);
xnor U6809 (N_6809,N_6665,N_6647);
nand U6810 (N_6810,N_6634,N_6727);
xor U6811 (N_6811,N_6629,N_6735);
xor U6812 (N_6812,N_6637,N_6677);
or U6813 (N_6813,N_6664,N_6689);
xnor U6814 (N_6814,N_6698,N_6745);
xnor U6815 (N_6815,N_6723,N_6737);
or U6816 (N_6816,N_6610,N_6630);
or U6817 (N_6817,N_6703,N_6660);
xnor U6818 (N_6818,N_6678,N_6685);
nor U6819 (N_6819,N_6695,N_6712);
xnor U6820 (N_6820,N_6646,N_6644);
nand U6821 (N_6821,N_6680,N_6681);
and U6822 (N_6822,N_6631,N_6706);
xor U6823 (N_6823,N_6710,N_6633);
nand U6824 (N_6824,N_6730,N_6692);
or U6825 (N_6825,N_6695,N_6736);
xnor U6826 (N_6826,N_6622,N_6720);
or U6827 (N_6827,N_6609,N_6624);
and U6828 (N_6828,N_6739,N_6660);
xor U6829 (N_6829,N_6636,N_6661);
and U6830 (N_6830,N_6726,N_6674);
nor U6831 (N_6831,N_6642,N_6687);
nand U6832 (N_6832,N_6681,N_6721);
nand U6833 (N_6833,N_6727,N_6717);
nor U6834 (N_6834,N_6729,N_6700);
or U6835 (N_6835,N_6643,N_6743);
or U6836 (N_6836,N_6705,N_6613);
and U6837 (N_6837,N_6674,N_6625);
nor U6838 (N_6838,N_6648,N_6702);
nand U6839 (N_6839,N_6713,N_6663);
nand U6840 (N_6840,N_6746,N_6638);
nand U6841 (N_6841,N_6708,N_6732);
nor U6842 (N_6842,N_6617,N_6741);
and U6843 (N_6843,N_6648,N_6697);
xor U6844 (N_6844,N_6610,N_6733);
xnor U6845 (N_6845,N_6623,N_6699);
nand U6846 (N_6846,N_6695,N_6669);
nor U6847 (N_6847,N_6682,N_6642);
or U6848 (N_6848,N_6651,N_6740);
nor U6849 (N_6849,N_6723,N_6620);
nand U6850 (N_6850,N_6668,N_6703);
nand U6851 (N_6851,N_6683,N_6738);
xnor U6852 (N_6852,N_6694,N_6707);
xor U6853 (N_6853,N_6626,N_6625);
or U6854 (N_6854,N_6600,N_6628);
or U6855 (N_6855,N_6644,N_6701);
xor U6856 (N_6856,N_6736,N_6611);
xor U6857 (N_6857,N_6655,N_6731);
nor U6858 (N_6858,N_6703,N_6689);
and U6859 (N_6859,N_6706,N_6630);
and U6860 (N_6860,N_6748,N_6662);
xor U6861 (N_6861,N_6720,N_6681);
nand U6862 (N_6862,N_6721,N_6633);
xnor U6863 (N_6863,N_6604,N_6680);
nor U6864 (N_6864,N_6693,N_6670);
nor U6865 (N_6865,N_6715,N_6711);
xnor U6866 (N_6866,N_6615,N_6745);
nor U6867 (N_6867,N_6667,N_6690);
nand U6868 (N_6868,N_6701,N_6611);
nand U6869 (N_6869,N_6722,N_6711);
nor U6870 (N_6870,N_6703,N_6640);
nand U6871 (N_6871,N_6664,N_6698);
nand U6872 (N_6872,N_6681,N_6682);
nor U6873 (N_6873,N_6656,N_6708);
nor U6874 (N_6874,N_6612,N_6717);
nor U6875 (N_6875,N_6682,N_6727);
or U6876 (N_6876,N_6616,N_6605);
or U6877 (N_6877,N_6743,N_6718);
xor U6878 (N_6878,N_6625,N_6710);
or U6879 (N_6879,N_6708,N_6630);
nand U6880 (N_6880,N_6709,N_6692);
xnor U6881 (N_6881,N_6645,N_6631);
nor U6882 (N_6882,N_6706,N_6662);
nor U6883 (N_6883,N_6665,N_6669);
or U6884 (N_6884,N_6703,N_6619);
nor U6885 (N_6885,N_6749,N_6673);
or U6886 (N_6886,N_6711,N_6640);
nor U6887 (N_6887,N_6633,N_6668);
xnor U6888 (N_6888,N_6626,N_6658);
nand U6889 (N_6889,N_6627,N_6690);
nand U6890 (N_6890,N_6699,N_6672);
or U6891 (N_6891,N_6647,N_6680);
xor U6892 (N_6892,N_6640,N_6699);
and U6893 (N_6893,N_6637,N_6642);
xnor U6894 (N_6894,N_6629,N_6699);
xor U6895 (N_6895,N_6623,N_6739);
or U6896 (N_6896,N_6657,N_6647);
and U6897 (N_6897,N_6638,N_6650);
nor U6898 (N_6898,N_6658,N_6613);
nand U6899 (N_6899,N_6617,N_6643);
and U6900 (N_6900,N_6875,N_6810);
or U6901 (N_6901,N_6777,N_6877);
nor U6902 (N_6902,N_6892,N_6831);
xnor U6903 (N_6903,N_6821,N_6899);
nor U6904 (N_6904,N_6890,N_6770);
nor U6905 (N_6905,N_6763,N_6756);
nand U6906 (N_6906,N_6782,N_6797);
and U6907 (N_6907,N_6828,N_6754);
and U6908 (N_6908,N_6768,N_6822);
and U6909 (N_6909,N_6834,N_6854);
nand U6910 (N_6910,N_6765,N_6802);
and U6911 (N_6911,N_6873,N_6848);
xor U6912 (N_6912,N_6863,N_6801);
and U6913 (N_6913,N_6845,N_6889);
xor U6914 (N_6914,N_6851,N_6786);
nand U6915 (N_6915,N_6764,N_6796);
nand U6916 (N_6916,N_6838,N_6852);
nand U6917 (N_6917,N_6776,N_6829);
nand U6918 (N_6918,N_6839,N_6820);
xor U6919 (N_6919,N_6870,N_6826);
xnor U6920 (N_6920,N_6842,N_6879);
nor U6921 (N_6921,N_6806,N_6894);
or U6922 (N_6922,N_6864,N_6751);
xor U6923 (N_6923,N_6823,N_6817);
xnor U6924 (N_6924,N_6862,N_6827);
nand U6925 (N_6925,N_6793,N_6750);
and U6926 (N_6926,N_6783,N_6849);
nor U6927 (N_6927,N_6847,N_6775);
nand U6928 (N_6928,N_6799,N_6830);
or U6929 (N_6929,N_6757,N_6791);
xor U6930 (N_6930,N_6784,N_6853);
or U6931 (N_6931,N_6835,N_6811);
nor U6932 (N_6932,N_6816,N_6798);
nand U6933 (N_6933,N_6787,N_6837);
nand U6934 (N_6934,N_6771,N_6888);
nor U6935 (N_6935,N_6836,N_6790);
nand U6936 (N_6936,N_6878,N_6767);
nand U6937 (N_6937,N_6895,N_6762);
xnor U6938 (N_6938,N_6760,N_6893);
or U6939 (N_6939,N_6865,N_6874);
xor U6940 (N_6940,N_6859,N_6808);
or U6941 (N_6941,N_6841,N_6769);
or U6942 (N_6942,N_6868,N_6833);
xor U6943 (N_6943,N_6881,N_6843);
and U6944 (N_6944,N_6785,N_6887);
nand U6945 (N_6945,N_6860,N_6792);
and U6946 (N_6946,N_6814,N_6759);
or U6947 (N_6947,N_6840,N_6813);
nor U6948 (N_6948,N_6781,N_6804);
nor U6949 (N_6949,N_6773,N_6818);
xor U6950 (N_6950,N_6752,N_6824);
or U6951 (N_6951,N_6891,N_6856);
or U6952 (N_6952,N_6789,N_6815);
nand U6953 (N_6953,N_6898,N_6807);
nand U6954 (N_6954,N_6869,N_6857);
nand U6955 (N_6955,N_6795,N_6780);
nor U6956 (N_6956,N_6755,N_6866);
nand U6957 (N_6957,N_6803,N_6761);
nor U6958 (N_6958,N_6886,N_6880);
nand U6959 (N_6959,N_6819,N_6794);
and U6960 (N_6960,N_6788,N_6861);
or U6961 (N_6961,N_6844,N_6871);
xor U6962 (N_6962,N_6896,N_6884);
xnor U6963 (N_6963,N_6850,N_6858);
nor U6964 (N_6964,N_6897,N_6825);
or U6965 (N_6965,N_6779,N_6758);
nor U6966 (N_6966,N_6778,N_6872);
or U6967 (N_6967,N_6774,N_6876);
nor U6968 (N_6968,N_6846,N_6832);
and U6969 (N_6969,N_6867,N_6766);
and U6970 (N_6970,N_6805,N_6812);
or U6971 (N_6971,N_6883,N_6809);
xor U6972 (N_6972,N_6772,N_6855);
xor U6973 (N_6973,N_6753,N_6885);
nand U6974 (N_6974,N_6800,N_6882);
and U6975 (N_6975,N_6800,N_6818);
and U6976 (N_6976,N_6799,N_6867);
xnor U6977 (N_6977,N_6769,N_6776);
or U6978 (N_6978,N_6882,N_6899);
and U6979 (N_6979,N_6827,N_6829);
and U6980 (N_6980,N_6790,N_6857);
nand U6981 (N_6981,N_6861,N_6867);
and U6982 (N_6982,N_6857,N_6750);
nor U6983 (N_6983,N_6807,N_6832);
xor U6984 (N_6984,N_6890,N_6817);
nor U6985 (N_6985,N_6805,N_6875);
and U6986 (N_6986,N_6773,N_6885);
xnor U6987 (N_6987,N_6813,N_6898);
or U6988 (N_6988,N_6816,N_6877);
nand U6989 (N_6989,N_6856,N_6877);
and U6990 (N_6990,N_6846,N_6863);
and U6991 (N_6991,N_6776,N_6802);
nor U6992 (N_6992,N_6786,N_6787);
nand U6993 (N_6993,N_6839,N_6821);
and U6994 (N_6994,N_6863,N_6869);
xor U6995 (N_6995,N_6767,N_6866);
nand U6996 (N_6996,N_6880,N_6882);
nand U6997 (N_6997,N_6763,N_6808);
xnor U6998 (N_6998,N_6848,N_6843);
xnor U6999 (N_6999,N_6750,N_6794);
or U7000 (N_7000,N_6868,N_6880);
nor U7001 (N_7001,N_6783,N_6780);
nand U7002 (N_7002,N_6855,N_6761);
or U7003 (N_7003,N_6873,N_6830);
or U7004 (N_7004,N_6814,N_6834);
or U7005 (N_7005,N_6881,N_6887);
or U7006 (N_7006,N_6850,N_6837);
xor U7007 (N_7007,N_6825,N_6820);
nand U7008 (N_7008,N_6760,N_6753);
and U7009 (N_7009,N_6866,N_6838);
nand U7010 (N_7010,N_6832,N_6826);
or U7011 (N_7011,N_6810,N_6781);
nand U7012 (N_7012,N_6888,N_6873);
and U7013 (N_7013,N_6777,N_6757);
nor U7014 (N_7014,N_6862,N_6857);
nor U7015 (N_7015,N_6881,N_6837);
or U7016 (N_7016,N_6807,N_6789);
nor U7017 (N_7017,N_6753,N_6839);
nand U7018 (N_7018,N_6875,N_6848);
nor U7019 (N_7019,N_6872,N_6826);
and U7020 (N_7020,N_6876,N_6823);
nor U7021 (N_7021,N_6890,N_6789);
xnor U7022 (N_7022,N_6887,N_6871);
and U7023 (N_7023,N_6781,N_6830);
nor U7024 (N_7024,N_6777,N_6869);
xor U7025 (N_7025,N_6874,N_6831);
and U7026 (N_7026,N_6891,N_6799);
nand U7027 (N_7027,N_6831,N_6763);
or U7028 (N_7028,N_6857,N_6860);
and U7029 (N_7029,N_6824,N_6829);
and U7030 (N_7030,N_6790,N_6870);
xnor U7031 (N_7031,N_6786,N_6845);
or U7032 (N_7032,N_6856,N_6804);
or U7033 (N_7033,N_6848,N_6898);
nand U7034 (N_7034,N_6811,N_6769);
nand U7035 (N_7035,N_6889,N_6760);
and U7036 (N_7036,N_6771,N_6892);
or U7037 (N_7037,N_6782,N_6885);
xnor U7038 (N_7038,N_6888,N_6820);
xnor U7039 (N_7039,N_6885,N_6844);
nor U7040 (N_7040,N_6809,N_6875);
nor U7041 (N_7041,N_6781,N_6788);
nor U7042 (N_7042,N_6791,N_6815);
nor U7043 (N_7043,N_6872,N_6810);
or U7044 (N_7044,N_6899,N_6792);
or U7045 (N_7045,N_6839,N_6798);
nor U7046 (N_7046,N_6809,N_6799);
or U7047 (N_7047,N_6823,N_6782);
nor U7048 (N_7048,N_6758,N_6828);
nand U7049 (N_7049,N_6870,N_6756);
or U7050 (N_7050,N_6903,N_7049);
and U7051 (N_7051,N_6974,N_6944);
xnor U7052 (N_7052,N_6915,N_6910);
xor U7053 (N_7053,N_6962,N_6978);
xor U7054 (N_7054,N_6968,N_6917);
xnor U7055 (N_7055,N_6914,N_6950);
nor U7056 (N_7056,N_6957,N_6926);
nor U7057 (N_7057,N_6925,N_6961);
nor U7058 (N_7058,N_7044,N_6938);
and U7059 (N_7059,N_7036,N_6959);
nand U7060 (N_7060,N_6919,N_6946);
and U7061 (N_7061,N_7038,N_6958);
nand U7062 (N_7062,N_6947,N_7010);
or U7063 (N_7063,N_7006,N_6984);
or U7064 (N_7064,N_6987,N_6969);
nand U7065 (N_7065,N_7033,N_6929);
xor U7066 (N_7066,N_7023,N_7012);
nor U7067 (N_7067,N_6998,N_7030);
nand U7068 (N_7068,N_6912,N_7035);
nor U7069 (N_7069,N_6994,N_6911);
or U7070 (N_7070,N_6918,N_6920);
and U7071 (N_7071,N_6913,N_6993);
nor U7072 (N_7072,N_7034,N_6966);
nor U7073 (N_7073,N_6943,N_7048);
xor U7074 (N_7074,N_7028,N_6953);
xnor U7075 (N_7075,N_6983,N_6949);
nor U7076 (N_7076,N_7020,N_6963);
or U7077 (N_7077,N_6956,N_6934);
xnor U7078 (N_7078,N_7000,N_6922);
xnor U7079 (N_7079,N_6954,N_6916);
or U7080 (N_7080,N_6985,N_6923);
nand U7081 (N_7081,N_6991,N_6928);
nor U7082 (N_7082,N_7003,N_6930);
nand U7083 (N_7083,N_6976,N_6933);
nor U7084 (N_7084,N_7024,N_7026);
nor U7085 (N_7085,N_6960,N_7017);
nor U7086 (N_7086,N_6970,N_6941);
xnor U7087 (N_7087,N_7009,N_6939);
xnor U7088 (N_7088,N_6921,N_6977);
nand U7089 (N_7089,N_6932,N_6997);
or U7090 (N_7090,N_6927,N_6901);
and U7091 (N_7091,N_6945,N_6902);
xnor U7092 (N_7092,N_7007,N_6979);
and U7093 (N_7093,N_6982,N_6904);
or U7094 (N_7094,N_6965,N_6989);
xnor U7095 (N_7095,N_7011,N_7008);
or U7096 (N_7096,N_7018,N_7016);
and U7097 (N_7097,N_6999,N_6952);
xnor U7098 (N_7098,N_7022,N_7046);
or U7099 (N_7099,N_7031,N_7043);
xnor U7100 (N_7100,N_6971,N_6935);
nor U7101 (N_7101,N_6995,N_7029);
nand U7102 (N_7102,N_7005,N_7004);
or U7103 (N_7103,N_6973,N_7032);
or U7104 (N_7104,N_6906,N_6900);
or U7105 (N_7105,N_6964,N_6988);
and U7106 (N_7106,N_7021,N_6948);
xor U7107 (N_7107,N_6905,N_6975);
or U7108 (N_7108,N_6909,N_6907);
xor U7109 (N_7109,N_6967,N_6940);
or U7110 (N_7110,N_7027,N_7037);
xnor U7111 (N_7111,N_7045,N_6924);
xor U7112 (N_7112,N_6908,N_6955);
nand U7113 (N_7113,N_7041,N_6936);
or U7114 (N_7114,N_7019,N_7015);
xnor U7115 (N_7115,N_6951,N_6996);
xor U7116 (N_7116,N_6990,N_7002);
nor U7117 (N_7117,N_6980,N_6981);
nor U7118 (N_7118,N_6992,N_6931);
and U7119 (N_7119,N_6942,N_7001);
or U7120 (N_7120,N_7025,N_6937);
and U7121 (N_7121,N_7042,N_7039);
and U7122 (N_7122,N_6972,N_6986);
nor U7123 (N_7123,N_7014,N_7013);
or U7124 (N_7124,N_7047,N_7040);
xor U7125 (N_7125,N_6938,N_6956);
and U7126 (N_7126,N_6942,N_7037);
nand U7127 (N_7127,N_6969,N_6939);
xor U7128 (N_7128,N_6908,N_7014);
nand U7129 (N_7129,N_6917,N_6971);
and U7130 (N_7130,N_7016,N_6940);
and U7131 (N_7131,N_7035,N_7037);
and U7132 (N_7132,N_7039,N_6902);
nand U7133 (N_7133,N_6963,N_6966);
and U7134 (N_7134,N_6967,N_6969);
or U7135 (N_7135,N_6973,N_7030);
or U7136 (N_7136,N_6996,N_7000);
nand U7137 (N_7137,N_6978,N_7000);
or U7138 (N_7138,N_6976,N_7034);
nor U7139 (N_7139,N_6957,N_7026);
or U7140 (N_7140,N_7049,N_7024);
nand U7141 (N_7141,N_6987,N_6911);
nand U7142 (N_7142,N_7049,N_6991);
or U7143 (N_7143,N_6908,N_7022);
or U7144 (N_7144,N_6956,N_6970);
nor U7145 (N_7145,N_7046,N_7023);
nor U7146 (N_7146,N_6928,N_6957);
and U7147 (N_7147,N_7049,N_7030);
and U7148 (N_7148,N_7039,N_6999);
nand U7149 (N_7149,N_6979,N_7032);
and U7150 (N_7150,N_6958,N_7048);
nand U7151 (N_7151,N_6982,N_7049);
nor U7152 (N_7152,N_6917,N_7019);
nor U7153 (N_7153,N_7019,N_7034);
or U7154 (N_7154,N_6983,N_6960);
nor U7155 (N_7155,N_6984,N_6935);
nand U7156 (N_7156,N_7003,N_7043);
xnor U7157 (N_7157,N_6920,N_6911);
or U7158 (N_7158,N_6929,N_6930);
nand U7159 (N_7159,N_7028,N_7037);
xor U7160 (N_7160,N_6925,N_6969);
nor U7161 (N_7161,N_6980,N_6949);
or U7162 (N_7162,N_6936,N_7002);
nor U7163 (N_7163,N_6962,N_7040);
nand U7164 (N_7164,N_6912,N_6995);
or U7165 (N_7165,N_7005,N_6936);
or U7166 (N_7166,N_6939,N_6965);
xnor U7167 (N_7167,N_6954,N_6962);
and U7168 (N_7168,N_6950,N_6972);
and U7169 (N_7169,N_7039,N_7029);
nor U7170 (N_7170,N_7013,N_6934);
nor U7171 (N_7171,N_7025,N_6962);
xor U7172 (N_7172,N_7042,N_7043);
nand U7173 (N_7173,N_6910,N_6946);
and U7174 (N_7174,N_6970,N_7002);
and U7175 (N_7175,N_6921,N_6923);
nand U7176 (N_7176,N_7031,N_7015);
xor U7177 (N_7177,N_7015,N_6955);
and U7178 (N_7178,N_6906,N_6901);
or U7179 (N_7179,N_6969,N_6940);
and U7180 (N_7180,N_6902,N_6916);
or U7181 (N_7181,N_6967,N_6987);
nand U7182 (N_7182,N_7027,N_7047);
and U7183 (N_7183,N_7017,N_7012);
and U7184 (N_7184,N_7039,N_7009);
nor U7185 (N_7185,N_6910,N_7000);
nand U7186 (N_7186,N_7047,N_7009);
nor U7187 (N_7187,N_6967,N_6913);
nor U7188 (N_7188,N_7045,N_6988);
xor U7189 (N_7189,N_6980,N_6928);
xor U7190 (N_7190,N_7044,N_6929);
and U7191 (N_7191,N_7030,N_6911);
and U7192 (N_7192,N_6974,N_6943);
or U7193 (N_7193,N_6983,N_6910);
and U7194 (N_7194,N_7040,N_6925);
or U7195 (N_7195,N_7045,N_6993);
and U7196 (N_7196,N_6979,N_7036);
xnor U7197 (N_7197,N_6956,N_7018);
or U7198 (N_7198,N_6997,N_6942);
and U7199 (N_7199,N_7012,N_6946);
nand U7200 (N_7200,N_7143,N_7075);
xor U7201 (N_7201,N_7165,N_7114);
nand U7202 (N_7202,N_7066,N_7074);
nor U7203 (N_7203,N_7174,N_7183);
nand U7204 (N_7204,N_7050,N_7090);
and U7205 (N_7205,N_7059,N_7190);
or U7206 (N_7206,N_7067,N_7079);
xnor U7207 (N_7207,N_7142,N_7102);
or U7208 (N_7208,N_7127,N_7122);
nand U7209 (N_7209,N_7149,N_7152);
nand U7210 (N_7210,N_7154,N_7186);
nand U7211 (N_7211,N_7115,N_7105);
xor U7212 (N_7212,N_7130,N_7125);
nor U7213 (N_7213,N_7084,N_7078);
nand U7214 (N_7214,N_7145,N_7129);
nor U7215 (N_7215,N_7099,N_7088);
nor U7216 (N_7216,N_7138,N_7071);
nand U7217 (N_7217,N_7146,N_7182);
and U7218 (N_7218,N_7054,N_7082);
xor U7219 (N_7219,N_7156,N_7060);
nand U7220 (N_7220,N_7180,N_7153);
xor U7221 (N_7221,N_7189,N_7160);
and U7222 (N_7222,N_7052,N_7176);
xnor U7223 (N_7223,N_7140,N_7053);
or U7224 (N_7224,N_7128,N_7135);
and U7225 (N_7225,N_7157,N_7159);
nor U7226 (N_7226,N_7081,N_7167);
nor U7227 (N_7227,N_7070,N_7116);
and U7228 (N_7228,N_7137,N_7080);
xor U7229 (N_7229,N_7057,N_7106);
nand U7230 (N_7230,N_7155,N_7199);
nor U7231 (N_7231,N_7091,N_7136);
xnor U7232 (N_7232,N_7181,N_7178);
nand U7233 (N_7233,N_7147,N_7194);
nor U7234 (N_7234,N_7161,N_7051);
or U7235 (N_7235,N_7092,N_7056);
xnor U7236 (N_7236,N_7058,N_7119);
xnor U7237 (N_7237,N_7134,N_7166);
xnor U7238 (N_7238,N_7192,N_7126);
nand U7239 (N_7239,N_7103,N_7113);
xor U7240 (N_7240,N_7179,N_7132);
nor U7241 (N_7241,N_7120,N_7133);
nand U7242 (N_7242,N_7072,N_7100);
nor U7243 (N_7243,N_7158,N_7170);
or U7244 (N_7244,N_7077,N_7063);
xor U7245 (N_7245,N_7112,N_7089);
xnor U7246 (N_7246,N_7168,N_7188);
or U7247 (N_7247,N_7083,N_7198);
nor U7248 (N_7248,N_7108,N_7148);
xor U7249 (N_7249,N_7191,N_7141);
nand U7250 (N_7250,N_7162,N_7086);
nor U7251 (N_7251,N_7193,N_7110);
xnor U7252 (N_7252,N_7094,N_7096);
and U7253 (N_7253,N_7097,N_7104);
or U7254 (N_7254,N_7123,N_7076);
xnor U7255 (N_7255,N_7195,N_7068);
xnor U7256 (N_7256,N_7069,N_7139);
nor U7257 (N_7257,N_7187,N_7172);
nand U7258 (N_7258,N_7117,N_7109);
nand U7259 (N_7259,N_7064,N_7164);
nand U7260 (N_7260,N_7151,N_7062);
xnor U7261 (N_7261,N_7144,N_7173);
nand U7262 (N_7262,N_7085,N_7185);
xnor U7263 (N_7263,N_7131,N_7197);
xnor U7264 (N_7264,N_7065,N_7163);
and U7265 (N_7265,N_7169,N_7175);
or U7266 (N_7266,N_7171,N_7061);
nor U7267 (N_7267,N_7121,N_7087);
nor U7268 (N_7268,N_7111,N_7093);
and U7269 (N_7269,N_7150,N_7177);
and U7270 (N_7270,N_7124,N_7073);
xor U7271 (N_7271,N_7107,N_7118);
xnor U7272 (N_7272,N_7184,N_7196);
nand U7273 (N_7273,N_7101,N_7095);
xnor U7274 (N_7274,N_7098,N_7055);
nor U7275 (N_7275,N_7174,N_7071);
nand U7276 (N_7276,N_7057,N_7151);
and U7277 (N_7277,N_7157,N_7053);
nor U7278 (N_7278,N_7089,N_7154);
xnor U7279 (N_7279,N_7064,N_7069);
xnor U7280 (N_7280,N_7199,N_7180);
xnor U7281 (N_7281,N_7194,N_7172);
xor U7282 (N_7282,N_7106,N_7130);
nor U7283 (N_7283,N_7129,N_7110);
or U7284 (N_7284,N_7145,N_7191);
nand U7285 (N_7285,N_7068,N_7096);
nor U7286 (N_7286,N_7133,N_7131);
xor U7287 (N_7287,N_7060,N_7052);
nor U7288 (N_7288,N_7072,N_7173);
nor U7289 (N_7289,N_7107,N_7143);
nand U7290 (N_7290,N_7077,N_7152);
xor U7291 (N_7291,N_7062,N_7104);
or U7292 (N_7292,N_7181,N_7136);
and U7293 (N_7293,N_7065,N_7159);
and U7294 (N_7294,N_7073,N_7123);
and U7295 (N_7295,N_7122,N_7197);
nand U7296 (N_7296,N_7103,N_7091);
xor U7297 (N_7297,N_7056,N_7114);
xnor U7298 (N_7298,N_7154,N_7053);
and U7299 (N_7299,N_7079,N_7154);
and U7300 (N_7300,N_7137,N_7057);
nand U7301 (N_7301,N_7164,N_7134);
nand U7302 (N_7302,N_7065,N_7144);
or U7303 (N_7303,N_7181,N_7170);
xor U7304 (N_7304,N_7100,N_7173);
nand U7305 (N_7305,N_7083,N_7069);
xor U7306 (N_7306,N_7170,N_7188);
nor U7307 (N_7307,N_7093,N_7186);
or U7308 (N_7308,N_7104,N_7153);
and U7309 (N_7309,N_7097,N_7065);
nand U7310 (N_7310,N_7067,N_7090);
or U7311 (N_7311,N_7173,N_7162);
nor U7312 (N_7312,N_7167,N_7170);
or U7313 (N_7313,N_7163,N_7072);
and U7314 (N_7314,N_7051,N_7184);
and U7315 (N_7315,N_7197,N_7099);
nor U7316 (N_7316,N_7154,N_7171);
nor U7317 (N_7317,N_7098,N_7146);
nor U7318 (N_7318,N_7068,N_7135);
nand U7319 (N_7319,N_7194,N_7148);
nand U7320 (N_7320,N_7099,N_7050);
nor U7321 (N_7321,N_7115,N_7075);
nor U7322 (N_7322,N_7171,N_7050);
nor U7323 (N_7323,N_7140,N_7050);
xnor U7324 (N_7324,N_7161,N_7191);
and U7325 (N_7325,N_7060,N_7176);
nand U7326 (N_7326,N_7181,N_7123);
nor U7327 (N_7327,N_7078,N_7083);
xor U7328 (N_7328,N_7092,N_7125);
and U7329 (N_7329,N_7060,N_7130);
nand U7330 (N_7330,N_7085,N_7125);
xnor U7331 (N_7331,N_7147,N_7099);
and U7332 (N_7332,N_7197,N_7144);
and U7333 (N_7333,N_7094,N_7079);
xnor U7334 (N_7334,N_7084,N_7125);
nor U7335 (N_7335,N_7153,N_7168);
nor U7336 (N_7336,N_7174,N_7175);
and U7337 (N_7337,N_7146,N_7087);
and U7338 (N_7338,N_7127,N_7051);
nand U7339 (N_7339,N_7126,N_7101);
and U7340 (N_7340,N_7107,N_7134);
or U7341 (N_7341,N_7087,N_7110);
or U7342 (N_7342,N_7117,N_7114);
and U7343 (N_7343,N_7187,N_7059);
nand U7344 (N_7344,N_7079,N_7159);
xnor U7345 (N_7345,N_7118,N_7125);
and U7346 (N_7346,N_7199,N_7119);
and U7347 (N_7347,N_7137,N_7094);
nor U7348 (N_7348,N_7151,N_7197);
nor U7349 (N_7349,N_7151,N_7078);
nor U7350 (N_7350,N_7238,N_7344);
or U7351 (N_7351,N_7201,N_7316);
xnor U7352 (N_7352,N_7273,N_7308);
or U7353 (N_7353,N_7275,N_7317);
xnor U7354 (N_7354,N_7314,N_7286);
or U7355 (N_7355,N_7263,N_7321);
or U7356 (N_7356,N_7300,N_7236);
and U7357 (N_7357,N_7330,N_7265);
and U7358 (N_7358,N_7249,N_7318);
or U7359 (N_7359,N_7328,N_7228);
xnor U7360 (N_7360,N_7223,N_7206);
and U7361 (N_7361,N_7239,N_7205);
xnor U7362 (N_7362,N_7287,N_7209);
nor U7363 (N_7363,N_7227,N_7243);
and U7364 (N_7364,N_7297,N_7242);
nand U7365 (N_7365,N_7241,N_7283);
xor U7366 (N_7366,N_7303,N_7304);
nor U7367 (N_7367,N_7315,N_7302);
nand U7368 (N_7368,N_7234,N_7301);
xor U7369 (N_7369,N_7305,N_7295);
nand U7370 (N_7370,N_7226,N_7310);
nand U7371 (N_7371,N_7222,N_7267);
or U7372 (N_7372,N_7334,N_7340);
nor U7373 (N_7373,N_7341,N_7288);
xor U7374 (N_7374,N_7211,N_7312);
nor U7375 (N_7375,N_7240,N_7285);
and U7376 (N_7376,N_7237,N_7208);
nand U7377 (N_7377,N_7282,N_7327);
nor U7378 (N_7378,N_7233,N_7306);
and U7379 (N_7379,N_7252,N_7232);
nand U7380 (N_7380,N_7218,N_7215);
and U7381 (N_7381,N_7291,N_7214);
or U7382 (N_7382,N_7324,N_7276);
or U7383 (N_7383,N_7348,N_7290);
xor U7384 (N_7384,N_7320,N_7278);
or U7385 (N_7385,N_7202,N_7337);
nor U7386 (N_7386,N_7279,N_7299);
nor U7387 (N_7387,N_7221,N_7212);
xnor U7388 (N_7388,N_7326,N_7210);
nand U7389 (N_7389,N_7246,N_7292);
xor U7390 (N_7390,N_7247,N_7216);
nand U7391 (N_7391,N_7281,N_7270);
xor U7392 (N_7392,N_7333,N_7298);
nor U7393 (N_7393,N_7224,N_7219);
nor U7394 (N_7394,N_7293,N_7229);
nor U7395 (N_7395,N_7280,N_7284);
xor U7396 (N_7396,N_7274,N_7269);
nand U7397 (N_7397,N_7260,N_7335);
or U7398 (N_7398,N_7264,N_7257);
or U7399 (N_7399,N_7261,N_7342);
xor U7400 (N_7400,N_7349,N_7230);
nor U7401 (N_7401,N_7343,N_7323);
nor U7402 (N_7402,N_7254,N_7336);
nor U7403 (N_7403,N_7200,N_7311);
xnor U7404 (N_7404,N_7204,N_7255);
nand U7405 (N_7405,N_7339,N_7313);
nand U7406 (N_7406,N_7268,N_7248);
nand U7407 (N_7407,N_7231,N_7338);
and U7408 (N_7408,N_7235,N_7345);
or U7409 (N_7409,N_7262,N_7258);
and U7410 (N_7410,N_7331,N_7225);
and U7411 (N_7411,N_7256,N_7347);
or U7412 (N_7412,N_7289,N_7203);
nand U7413 (N_7413,N_7319,N_7332);
xor U7414 (N_7414,N_7244,N_7271);
nor U7415 (N_7415,N_7253,N_7294);
xnor U7416 (N_7416,N_7251,N_7207);
xor U7417 (N_7417,N_7329,N_7307);
or U7418 (N_7418,N_7309,N_7266);
and U7419 (N_7419,N_7325,N_7296);
nand U7420 (N_7420,N_7250,N_7259);
and U7421 (N_7421,N_7220,N_7217);
and U7422 (N_7422,N_7213,N_7322);
nand U7423 (N_7423,N_7277,N_7272);
nand U7424 (N_7424,N_7346,N_7245);
nand U7425 (N_7425,N_7329,N_7289);
and U7426 (N_7426,N_7239,N_7291);
xnor U7427 (N_7427,N_7318,N_7237);
xor U7428 (N_7428,N_7256,N_7282);
nor U7429 (N_7429,N_7339,N_7242);
nand U7430 (N_7430,N_7253,N_7265);
or U7431 (N_7431,N_7299,N_7237);
xor U7432 (N_7432,N_7212,N_7340);
nand U7433 (N_7433,N_7268,N_7310);
nor U7434 (N_7434,N_7299,N_7328);
or U7435 (N_7435,N_7204,N_7327);
nor U7436 (N_7436,N_7306,N_7201);
and U7437 (N_7437,N_7204,N_7249);
nand U7438 (N_7438,N_7245,N_7323);
nor U7439 (N_7439,N_7285,N_7295);
and U7440 (N_7440,N_7237,N_7259);
nand U7441 (N_7441,N_7301,N_7207);
xnor U7442 (N_7442,N_7258,N_7290);
nor U7443 (N_7443,N_7334,N_7261);
nand U7444 (N_7444,N_7276,N_7319);
nor U7445 (N_7445,N_7235,N_7347);
and U7446 (N_7446,N_7278,N_7276);
nand U7447 (N_7447,N_7239,N_7344);
nand U7448 (N_7448,N_7201,N_7211);
xor U7449 (N_7449,N_7224,N_7318);
or U7450 (N_7450,N_7301,N_7222);
and U7451 (N_7451,N_7201,N_7251);
nand U7452 (N_7452,N_7223,N_7318);
or U7453 (N_7453,N_7240,N_7269);
nand U7454 (N_7454,N_7214,N_7293);
nor U7455 (N_7455,N_7209,N_7229);
or U7456 (N_7456,N_7238,N_7234);
or U7457 (N_7457,N_7266,N_7202);
nor U7458 (N_7458,N_7270,N_7303);
and U7459 (N_7459,N_7257,N_7338);
or U7460 (N_7460,N_7318,N_7268);
and U7461 (N_7461,N_7302,N_7235);
and U7462 (N_7462,N_7346,N_7259);
xor U7463 (N_7463,N_7250,N_7246);
nand U7464 (N_7464,N_7260,N_7278);
or U7465 (N_7465,N_7260,N_7332);
and U7466 (N_7466,N_7268,N_7277);
or U7467 (N_7467,N_7283,N_7274);
nand U7468 (N_7468,N_7345,N_7297);
xor U7469 (N_7469,N_7343,N_7222);
xnor U7470 (N_7470,N_7281,N_7274);
xnor U7471 (N_7471,N_7223,N_7302);
and U7472 (N_7472,N_7310,N_7346);
nand U7473 (N_7473,N_7231,N_7323);
and U7474 (N_7474,N_7347,N_7250);
and U7475 (N_7475,N_7200,N_7340);
or U7476 (N_7476,N_7311,N_7321);
nor U7477 (N_7477,N_7338,N_7244);
or U7478 (N_7478,N_7308,N_7225);
and U7479 (N_7479,N_7306,N_7331);
xor U7480 (N_7480,N_7250,N_7333);
nand U7481 (N_7481,N_7264,N_7295);
or U7482 (N_7482,N_7204,N_7269);
and U7483 (N_7483,N_7314,N_7299);
or U7484 (N_7484,N_7286,N_7225);
xor U7485 (N_7485,N_7214,N_7288);
xor U7486 (N_7486,N_7286,N_7273);
nand U7487 (N_7487,N_7248,N_7210);
nand U7488 (N_7488,N_7245,N_7343);
xnor U7489 (N_7489,N_7316,N_7338);
xor U7490 (N_7490,N_7316,N_7236);
nand U7491 (N_7491,N_7212,N_7300);
or U7492 (N_7492,N_7289,N_7331);
nor U7493 (N_7493,N_7260,N_7269);
or U7494 (N_7494,N_7332,N_7278);
or U7495 (N_7495,N_7289,N_7295);
and U7496 (N_7496,N_7209,N_7308);
xnor U7497 (N_7497,N_7304,N_7244);
or U7498 (N_7498,N_7257,N_7333);
and U7499 (N_7499,N_7243,N_7282);
or U7500 (N_7500,N_7385,N_7400);
or U7501 (N_7501,N_7387,N_7466);
nor U7502 (N_7502,N_7413,N_7410);
nand U7503 (N_7503,N_7363,N_7352);
nand U7504 (N_7504,N_7493,N_7390);
nor U7505 (N_7505,N_7373,N_7440);
nor U7506 (N_7506,N_7455,N_7388);
nor U7507 (N_7507,N_7483,N_7408);
nand U7508 (N_7508,N_7356,N_7476);
xor U7509 (N_7509,N_7465,N_7470);
nand U7510 (N_7510,N_7454,N_7449);
xor U7511 (N_7511,N_7485,N_7411);
or U7512 (N_7512,N_7362,N_7371);
and U7513 (N_7513,N_7396,N_7372);
nor U7514 (N_7514,N_7488,N_7475);
and U7515 (N_7515,N_7487,N_7361);
nor U7516 (N_7516,N_7486,N_7439);
nor U7517 (N_7517,N_7401,N_7479);
xnor U7518 (N_7518,N_7351,N_7405);
or U7519 (N_7519,N_7393,N_7367);
or U7520 (N_7520,N_7444,N_7350);
and U7521 (N_7521,N_7430,N_7443);
nor U7522 (N_7522,N_7441,N_7419);
and U7523 (N_7523,N_7369,N_7468);
and U7524 (N_7524,N_7417,N_7386);
or U7525 (N_7525,N_7424,N_7459);
xnor U7526 (N_7526,N_7473,N_7482);
nor U7527 (N_7527,N_7433,N_7423);
and U7528 (N_7528,N_7490,N_7447);
nor U7529 (N_7529,N_7404,N_7418);
and U7530 (N_7530,N_7355,N_7354);
and U7531 (N_7531,N_7464,N_7397);
nand U7532 (N_7532,N_7438,N_7406);
or U7533 (N_7533,N_7457,N_7392);
or U7534 (N_7534,N_7415,N_7462);
and U7535 (N_7535,N_7469,N_7420);
or U7536 (N_7536,N_7378,N_7499);
nand U7537 (N_7537,N_7422,N_7357);
xnor U7538 (N_7538,N_7382,N_7414);
nor U7539 (N_7539,N_7365,N_7450);
nand U7540 (N_7540,N_7432,N_7391);
nand U7541 (N_7541,N_7442,N_7460);
nand U7542 (N_7542,N_7384,N_7480);
xor U7543 (N_7543,N_7380,N_7472);
or U7544 (N_7544,N_7495,N_7428);
xor U7545 (N_7545,N_7481,N_7491);
or U7546 (N_7546,N_7467,N_7377);
xor U7547 (N_7547,N_7448,N_7394);
nand U7548 (N_7548,N_7429,N_7403);
xnor U7549 (N_7549,N_7494,N_7395);
and U7550 (N_7550,N_7436,N_7497);
nor U7551 (N_7551,N_7434,N_7478);
and U7552 (N_7552,N_7435,N_7474);
and U7553 (N_7553,N_7402,N_7461);
and U7554 (N_7554,N_7407,N_7452);
nand U7555 (N_7555,N_7409,N_7446);
nor U7556 (N_7556,N_7370,N_7353);
or U7557 (N_7557,N_7453,N_7379);
and U7558 (N_7558,N_7498,N_7456);
or U7559 (N_7559,N_7489,N_7492);
or U7560 (N_7560,N_7364,N_7427);
xor U7561 (N_7561,N_7445,N_7471);
xnor U7562 (N_7562,N_7416,N_7359);
and U7563 (N_7563,N_7360,N_7375);
xnor U7564 (N_7564,N_7431,N_7458);
nor U7565 (N_7565,N_7451,N_7399);
or U7566 (N_7566,N_7496,N_7374);
or U7567 (N_7567,N_7398,N_7383);
nor U7568 (N_7568,N_7381,N_7421);
xor U7569 (N_7569,N_7463,N_7426);
or U7570 (N_7570,N_7477,N_7376);
nand U7571 (N_7571,N_7366,N_7389);
xor U7572 (N_7572,N_7437,N_7425);
or U7573 (N_7573,N_7368,N_7484);
xor U7574 (N_7574,N_7358,N_7412);
xor U7575 (N_7575,N_7351,N_7495);
xnor U7576 (N_7576,N_7422,N_7496);
nand U7577 (N_7577,N_7363,N_7358);
nor U7578 (N_7578,N_7410,N_7456);
xnor U7579 (N_7579,N_7389,N_7400);
nand U7580 (N_7580,N_7455,N_7492);
nand U7581 (N_7581,N_7424,N_7489);
nand U7582 (N_7582,N_7414,N_7436);
and U7583 (N_7583,N_7410,N_7442);
nor U7584 (N_7584,N_7488,N_7453);
nand U7585 (N_7585,N_7393,N_7489);
nor U7586 (N_7586,N_7355,N_7484);
nor U7587 (N_7587,N_7449,N_7351);
or U7588 (N_7588,N_7405,N_7471);
nor U7589 (N_7589,N_7355,N_7391);
nor U7590 (N_7590,N_7388,N_7454);
nor U7591 (N_7591,N_7411,N_7430);
xnor U7592 (N_7592,N_7405,N_7492);
or U7593 (N_7593,N_7493,N_7438);
nor U7594 (N_7594,N_7441,N_7479);
nor U7595 (N_7595,N_7430,N_7438);
xor U7596 (N_7596,N_7448,N_7489);
or U7597 (N_7597,N_7470,N_7455);
and U7598 (N_7598,N_7366,N_7365);
or U7599 (N_7599,N_7380,N_7381);
nand U7600 (N_7600,N_7415,N_7381);
xor U7601 (N_7601,N_7452,N_7375);
nand U7602 (N_7602,N_7406,N_7486);
nor U7603 (N_7603,N_7419,N_7454);
nor U7604 (N_7604,N_7471,N_7474);
and U7605 (N_7605,N_7400,N_7441);
and U7606 (N_7606,N_7374,N_7439);
or U7607 (N_7607,N_7420,N_7446);
and U7608 (N_7608,N_7411,N_7480);
or U7609 (N_7609,N_7388,N_7378);
and U7610 (N_7610,N_7379,N_7368);
or U7611 (N_7611,N_7474,N_7453);
or U7612 (N_7612,N_7416,N_7421);
or U7613 (N_7613,N_7440,N_7407);
xor U7614 (N_7614,N_7445,N_7450);
or U7615 (N_7615,N_7423,N_7476);
or U7616 (N_7616,N_7444,N_7392);
and U7617 (N_7617,N_7439,N_7398);
nor U7618 (N_7618,N_7486,N_7484);
or U7619 (N_7619,N_7453,N_7374);
or U7620 (N_7620,N_7374,N_7396);
and U7621 (N_7621,N_7456,N_7392);
and U7622 (N_7622,N_7360,N_7499);
or U7623 (N_7623,N_7399,N_7359);
nor U7624 (N_7624,N_7409,N_7441);
or U7625 (N_7625,N_7395,N_7495);
and U7626 (N_7626,N_7453,N_7388);
nand U7627 (N_7627,N_7429,N_7487);
and U7628 (N_7628,N_7415,N_7406);
nor U7629 (N_7629,N_7365,N_7397);
or U7630 (N_7630,N_7469,N_7470);
nor U7631 (N_7631,N_7445,N_7356);
nand U7632 (N_7632,N_7370,N_7444);
nand U7633 (N_7633,N_7370,N_7359);
xor U7634 (N_7634,N_7372,N_7350);
nor U7635 (N_7635,N_7460,N_7475);
or U7636 (N_7636,N_7479,N_7445);
nand U7637 (N_7637,N_7456,N_7443);
nor U7638 (N_7638,N_7429,N_7385);
nor U7639 (N_7639,N_7426,N_7425);
and U7640 (N_7640,N_7475,N_7498);
or U7641 (N_7641,N_7382,N_7484);
nor U7642 (N_7642,N_7379,N_7375);
xor U7643 (N_7643,N_7368,N_7383);
xnor U7644 (N_7644,N_7373,N_7418);
or U7645 (N_7645,N_7429,N_7359);
nor U7646 (N_7646,N_7440,N_7470);
and U7647 (N_7647,N_7394,N_7484);
or U7648 (N_7648,N_7394,N_7385);
nor U7649 (N_7649,N_7489,N_7481);
xnor U7650 (N_7650,N_7646,N_7600);
xnor U7651 (N_7651,N_7536,N_7537);
nor U7652 (N_7652,N_7510,N_7581);
nand U7653 (N_7653,N_7596,N_7595);
and U7654 (N_7654,N_7539,N_7629);
nor U7655 (N_7655,N_7647,N_7590);
nor U7656 (N_7656,N_7649,N_7623);
and U7657 (N_7657,N_7565,N_7516);
or U7658 (N_7658,N_7631,N_7507);
nand U7659 (N_7659,N_7558,N_7533);
nor U7660 (N_7660,N_7506,N_7604);
nand U7661 (N_7661,N_7548,N_7622);
xor U7662 (N_7662,N_7619,N_7515);
nor U7663 (N_7663,N_7570,N_7588);
xor U7664 (N_7664,N_7618,N_7645);
or U7665 (N_7665,N_7585,N_7501);
nor U7666 (N_7666,N_7568,N_7643);
xnor U7667 (N_7667,N_7621,N_7566);
nor U7668 (N_7668,N_7526,N_7541);
and U7669 (N_7669,N_7599,N_7626);
or U7670 (N_7670,N_7625,N_7632);
xnor U7671 (N_7671,N_7522,N_7551);
and U7672 (N_7672,N_7577,N_7503);
and U7673 (N_7673,N_7544,N_7606);
or U7674 (N_7674,N_7513,N_7620);
and U7675 (N_7675,N_7628,N_7636);
and U7676 (N_7676,N_7601,N_7584);
or U7677 (N_7677,N_7635,N_7569);
and U7678 (N_7678,N_7564,N_7525);
xnor U7679 (N_7679,N_7500,N_7502);
or U7680 (N_7680,N_7616,N_7561);
or U7681 (N_7681,N_7624,N_7576);
or U7682 (N_7682,N_7614,N_7529);
nand U7683 (N_7683,N_7546,N_7639);
or U7684 (N_7684,N_7598,N_7586);
xor U7685 (N_7685,N_7512,N_7608);
nor U7686 (N_7686,N_7520,N_7610);
nor U7687 (N_7687,N_7572,N_7578);
nor U7688 (N_7688,N_7554,N_7642);
nor U7689 (N_7689,N_7574,N_7550);
nor U7690 (N_7690,N_7607,N_7532);
nand U7691 (N_7691,N_7514,N_7603);
nand U7692 (N_7692,N_7640,N_7555);
or U7693 (N_7693,N_7535,N_7531);
and U7694 (N_7694,N_7509,N_7559);
and U7695 (N_7695,N_7591,N_7644);
and U7696 (N_7696,N_7592,N_7534);
or U7697 (N_7697,N_7567,N_7508);
and U7698 (N_7698,N_7549,N_7580);
and U7699 (N_7699,N_7524,N_7542);
and U7700 (N_7700,N_7527,N_7605);
nand U7701 (N_7701,N_7597,N_7575);
xnor U7702 (N_7702,N_7633,N_7617);
and U7703 (N_7703,N_7517,N_7583);
nand U7704 (N_7704,N_7589,N_7593);
and U7705 (N_7705,N_7530,N_7523);
or U7706 (N_7706,N_7612,N_7521);
nand U7707 (N_7707,N_7602,N_7553);
and U7708 (N_7708,N_7540,N_7638);
or U7709 (N_7709,N_7511,N_7637);
nand U7710 (N_7710,N_7519,N_7563);
xor U7711 (N_7711,N_7594,N_7579);
nor U7712 (N_7712,N_7505,N_7562);
nand U7713 (N_7713,N_7587,N_7648);
nor U7714 (N_7714,N_7543,N_7556);
and U7715 (N_7715,N_7557,N_7518);
nor U7716 (N_7716,N_7615,N_7613);
xnor U7717 (N_7717,N_7547,N_7641);
nor U7718 (N_7718,N_7611,N_7571);
nor U7719 (N_7719,N_7538,N_7560);
nand U7720 (N_7720,N_7634,N_7528);
nand U7721 (N_7721,N_7630,N_7552);
nor U7722 (N_7722,N_7627,N_7504);
xor U7723 (N_7723,N_7609,N_7573);
xor U7724 (N_7724,N_7582,N_7545);
nand U7725 (N_7725,N_7646,N_7503);
xnor U7726 (N_7726,N_7621,N_7539);
xor U7727 (N_7727,N_7542,N_7522);
or U7728 (N_7728,N_7584,N_7506);
xnor U7729 (N_7729,N_7522,N_7517);
and U7730 (N_7730,N_7605,N_7564);
xnor U7731 (N_7731,N_7546,N_7649);
xnor U7732 (N_7732,N_7539,N_7524);
and U7733 (N_7733,N_7592,N_7565);
and U7734 (N_7734,N_7617,N_7529);
nand U7735 (N_7735,N_7614,N_7583);
or U7736 (N_7736,N_7599,N_7555);
nor U7737 (N_7737,N_7571,N_7602);
and U7738 (N_7738,N_7633,N_7601);
and U7739 (N_7739,N_7607,N_7621);
and U7740 (N_7740,N_7609,N_7627);
nor U7741 (N_7741,N_7611,N_7586);
nand U7742 (N_7742,N_7518,N_7519);
nor U7743 (N_7743,N_7522,N_7587);
or U7744 (N_7744,N_7649,N_7613);
xor U7745 (N_7745,N_7544,N_7511);
nand U7746 (N_7746,N_7595,N_7610);
nand U7747 (N_7747,N_7615,N_7557);
and U7748 (N_7748,N_7541,N_7615);
or U7749 (N_7749,N_7606,N_7510);
nor U7750 (N_7750,N_7590,N_7526);
and U7751 (N_7751,N_7635,N_7559);
nand U7752 (N_7752,N_7606,N_7576);
nor U7753 (N_7753,N_7516,N_7582);
nor U7754 (N_7754,N_7565,N_7544);
and U7755 (N_7755,N_7534,N_7589);
nor U7756 (N_7756,N_7540,N_7589);
xor U7757 (N_7757,N_7508,N_7631);
nor U7758 (N_7758,N_7605,N_7525);
or U7759 (N_7759,N_7623,N_7622);
or U7760 (N_7760,N_7521,N_7510);
nor U7761 (N_7761,N_7630,N_7553);
xnor U7762 (N_7762,N_7546,N_7593);
or U7763 (N_7763,N_7632,N_7591);
nor U7764 (N_7764,N_7603,N_7576);
xnor U7765 (N_7765,N_7542,N_7584);
and U7766 (N_7766,N_7561,N_7623);
xor U7767 (N_7767,N_7615,N_7528);
nor U7768 (N_7768,N_7647,N_7501);
nor U7769 (N_7769,N_7530,N_7604);
or U7770 (N_7770,N_7569,N_7648);
xnor U7771 (N_7771,N_7525,N_7544);
nor U7772 (N_7772,N_7606,N_7608);
or U7773 (N_7773,N_7550,N_7561);
xor U7774 (N_7774,N_7597,N_7538);
xnor U7775 (N_7775,N_7564,N_7610);
nand U7776 (N_7776,N_7543,N_7627);
or U7777 (N_7777,N_7506,N_7634);
xnor U7778 (N_7778,N_7501,N_7638);
and U7779 (N_7779,N_7584,N_7573);
and U7780 (N_7780,N_7519,N_7520);
and U7781 (N_7781,N_7541,N_7511);
or U7782 (N_7782,N_7618,N_7530);
and U7783 (N_7783,N_7591,N_7534);
xor U7784 (N_7784,N_7540,N_7577);
and U7785 (N_7785,N_7530,N_7553);
nor U7786 (N_7786,N_7549,N_7597);
nand U7787 (N_7787,N_7570,N_7595);
or U7788 (N_7788,N_7630,N_7591);
nor U7789 (N_7789,N_7504,N_7539);
or U7790 (N_7790,N_7579,N_7503);
and U7791 (N_7791,N_7565,N_7642);
nor U7792 (N_7792,N_7572,N_7564);
xnor U7793 (N_7793,N_7597,N_7516);
xnor U7794 (N_7794,N_7564,N_7645);
or U7795 (N_7795,N_7515,N_7556);
xor U7796 (N_7796,N_7521,N_7619);
or U7797 (N_7797,N_7509,N_7580);
or U7798 (N_7798,N_7542,N_7578);
nand U7799 (N_7799,N_7643,N_7614);
nor U7800 (N_7800,N_7746,N_7683);
nand U7801 (N_7801,N_7795,N_7673);
nor U7802 (N_7802,N_7679,N_7655);
or U7803 (N_7803,N_7704,N_7786);
or U7804 (N_7804,N_7656,N_7799);
or U7805 (N_7805,N_7792,N_7692);
or U7806 (N_7806,N_7740,N_7775);
nor U7807 (N_7807,N_7712,N_7744);
nor U7808 (N_7808,N_7785,N_7757);
and U7809 (N_7809,N_7690,N_7768);
xor U7810 (N_7810,N_7791,N_7688);
or U7811 (N_7811,N_7670,N_7695);
or U7812 (N_7812,N_7748,N_7666);
or U7813 (N_7813,N_7675,N_7715);
nand U7814 (N_7814,N_7796,N_7742);
xnor U7815 (N_7815,N_7677,N_7662);
or U7816 (N_7816,N_7671,N_7797);
nand U7817 (N_7817,N_7723,N_7722);
nor U7818 (N_7818,N_7706,N_7778);
or U7819 (N_7819,N_7769,N_7794);
nor U7820 (N_7820,N_7729,N_7650);
nand U7821 (N_7821,N_7686,N_7784);
nand U7822 (N_7822,N_7698,N_7709);
and U7823 (N_7823,N_7682,N_7703);
or U7824 (N_7824,N_7667,N_7759);
or U7825 (N_7825,N_7788,N_7754);
nor U7826 (N_7826,N_7750,N_7770);
and U7827 (N_7827,N_7763,N_7745);
or U7828 (N_7828,N_7730,N_7718);
nor U7829 (N_7829,N_7669,N_7705);
nor U7830 (N_7830,N_7762,N_7687);
xnor U7831 (N_7831,N_7774,N_7761);
nand U7832 (N_7832,N_7676,N_7689);
and U7833 (N_7833,N_7772,N_7760);
xor U7834 (N_7834,N_7732,N_7674);
nor U7835 (N_7835,N_7766,N_7776);
nor U7836 (N_7836,N_7696,N_7659);
and U7837 (N_7837,N_7779,N_7678);
nand U7838 (N_7838,N_7664,N_7777);
and U7839 (N_7839,N_7665,N_7658);
or U7840 (N_7840,N_7739,N_7681);
nand U7841 (N_7841,N_7780,N_7652);
xor U7842 (N_7842,N_7700,N_7691);
or U7843 (N_7843,N_7771,N_7728);
xor U7844 (N_7844,N_7767,N_7790);
nand U7845 (N_7845,N_7753,N_7793);
nor U7846 (N_7846,N_7716,N_7756);
nor U7847 (N_7847,N_7708,N_7720);
or U7848 (N_7848,N_7765,N_7694);
and U7849 (N_7849,N_7651,N_7713);
or U7850 (N_7850,N_7755,N_7782);
xor U7851 (N_7851,N_7725,N_7680);
nand U7852 (N_7852,N_7734,N_7714);
or U7853 (N_7853,N_7727,N_7668);
or U7854 (N_7854,N_7781,N_7653);
xnor U7855 (N_7855,N_7697,N_7654);
or U7856 (N_7856,N_7693,N_7657);
or U7857 (N_7857,N_7751,N_7661);
xnor U7858 (N_7858,N_7733,N_7738);
nand U7859 (N_7859,N_7717,N_7702);
xor U7860 (N_7860,N_7749,N_7731);
nand U7861 (N_7861,N_7672,N_7660);
and U7862 (N_7862,N_7726,N_7707);
nor U7863 (N_7863,N_7741,N_7736);
xor U7864 (N_7864,N_7758,N_7719);
nor U7865 (N_7865,N_7685,N_7721);
nor U7866 (N_7866,N_7699,N_7737);
nand U7867 (N_7867,N_7787,N_7711);
and U7868 (N_7868,N_7783,N_7724);
nor U7869 (N_7869,N_7701,N_7798);
and U7870 (N_7870,N_7752,N_7743);
xor U7871 (N_7871,N_7747,N_7710);
or U7872 (N_7872,N_7789,N_7684);
xnor U7873 (N_7873,N_7773,N_7764);
nand U7874 (N_7874,N_7663,N_7735);
and U7875 (N_7875,N_7702,N_7672);
xor U7876 (N_7876,N_7674,N_7684);
nand U7877 (N_7877,N_7668,N_7666);
nor U7878 (N_7878,N_7792,N_7776);
xnor U7879 (N_7879,N_7770,N_7722);
xnor U7880 (N_7880,N_7797,N_7733);
xnor U7881 (N_7881,N_7782,N_7692);
and U7882 (N_7882,N_7703,N_7773);
or U7883 (N_7883,N_7741,N_7786);
nor U7884 (N_7884,N_7758,N_7774);
or U7885 (N_7885,N_7748,N_7722);
nor U7886 (N_7886,N_7653,N_7686);
or U7887 (N_7887,N_7668,N_7735);
nor U7888 (N_7888,N_7700,N_7690);
nand U7889 (N_7889,N_7793,N_7667);
and U7890 (N_7890,N_7718,N_7680);
nor U7891 (N_7891,N_7719,N_7683);
or U7892 (N_7892,N_7703,N_7731);
xor U7893 (N_7893,N_7682,N_7755);
xnor U7894 (N_7894,N_7653,N_7651);
or U7895 (N_7895,N_7761,N_7773);
and U7896 (N_7896,N_7777,N_7706);
xor U7897 (N_7897,N_7695,N_7714);
and U7898 (N_7898,N_7715,N_7655);
nor U7899 (N_7899,N_7713,N_7799);
and U7900 (N_7900,N_7760,N_7749);
nor U7901 (N_7901,N_7706,N_7669);
xor U7902 (N_7902,N_7732,N_7767);
nand U7903 (N_7903,N_7784,N_7723);
or U7904 (N_7904,N_7657,N_7686);
xor U7905 (N_7905,N_7750,N_7756);
and U7906 (N_7906,N_7745,N_7796);
nand U7907 (N_7907,N_7747,N_7672);
nand U7908 (N_7908,N_7678,N_7694);
or U7909 (N_7909,N_7761,N_7676);
and U7910 (N_7910,N_7747,N_7741);
nor U7911 (N_7911,N_7772,N_7780);
or U7912 (N_7912,N_7664,N_7775);
nor U7913 (N_7913,N_7714,N_7670);
nor U7914 (N_7914,N_7740,N_7788);
xnor U7915 (N_7915,N_7727,N_7670);
nor U7916 (N_7916,N_7789,N_7696);
nand U7917 (N_7917,N_7762,N_7767);
nand U7918 (N_7918,N_7797,N_7652);
xor U7919 (N_7919,N_7671,N_7740);
nand U7920 (N_7920,N_7780,N_7718);
xor U7921 (N_7921,N_7754,N_7797);
nor U7922 (N_7922,N_7722,N_7701);
nand U7923 (N_7923,N_7658,N_7785);
or U7924 (N_7924,N_7724,N_7680);
and U7925 (N_7925,N_7673,N_7794);
nor U7926 (N_7926,N_7765,N_7788);
or U7927 (N_7927,N_7770,N_7656);
nand U7928 (N_7928,N_7659,N_7791);
nand U7929 (N_7929,N_7767,N_7734);
or U7930 (N_7930,N_7767,N_7794);
or U7931 (N_7931,N_7692,N_7774);
nor U7932 (N_7932,N_7714,N_7787);
nor U7933 (N_7933,N_7686,N_7676);
nand U7934 (N_7934,N_7723,N_7799);
nand U7935 (N_7935,N_7719,N_7734);
and U7936 (N_7936,N_7714,N_7685);
nor U7937 (N_7937,N_7794,N_7650);
and U7938 (N_7938,N_7721,N_7698);
nor U7939 (N_7939,N_7770,N_7779);
nand U7940 (N_7940,N_7788,N_7692);
nor U7941 (N_7941,N_7758,N_7760);
xnor U7942 (N_7942,N_7759,N_7762);
and U7943 (N_7943,N_7694,N_7699);
and U7944 (N_7944,N_7784,N_7735);
nor U7945 (N_7945,N_7793,N_7727);
nor U7946 (N_7946,N_7774,N_7791);
nor U7947 (N_7947,N_7748,N_7699);
or U7948 (N_7948,N_7794,N_7729);
nand U7949 (N_7949,N_7771,N_7720);
and U7950 (N_7950,N_7917,N_7872);
nand U7951 (N_7951,N_7805,N_7845);
or U7952 (N_7952,N_7842,N_7819);
and U7953 (N_7953,N_7939,N_7924);
or U7954 (N_7954,N_7887,N_7889);
and U7955 (N_7955,N_7854,N_7847);
nand U7956 (N_7956,N_7945,N_7828);
nand U7957 (N_7957,N_7808,N_7803);
or U7958 (N_7958,N_7886,N_7859);
or U7959 (N_7959,N_7885,N_7850);
or U7960 (N_7960,N_7841,N_7949);
and U7961 (N_7961,N_7915,N_7825);
and U7962 (N_7962,N_7895,N_7912);
or U7963 (N_7963,N_7944,N_7906);
nor U7964 (N_7964,N_7946,N_7880);
or U7965 (N_7965,N_7925,N_7849);
and U7966 (N_7966,N_7879,N_7883);
xor U7967 (N_7967,N_7901,N_7827);
and U7968 (N_7968,N_7856,N_7852);
or U7969 (N_7969,N_7903,N_7869);
and U7970 (N_7970,N_7812,N_7826);
or U7971 (N_7971,N_7862,N_7909);
and U7972 (N_7972,N_7908,N_7913);
xor U7973 (N_7973,N_7898,N_7824);
xnor U7974 (N_7974,N_7848,N_7911);
and U7975 (N_7975,N_7907,N_7882);
or U7976 (N_7976,N_7834,N_7910);
and U7977 (N_7977,N_7840,N_7864);
xnor U7978 (N_7978,N_7890,N_7893);
xor U7979 (N_7979,N_7936,N_7846);
nand U7980 (N_7980,N_7838,N_7873);
nand U7981 (N_7981,N_7875,N_7918);
nor U7982 (N_7982,N_7916,N_7823);
nor U7983 (N_7983,N_7837,N_7899);
and U7984 (N_7984,N_7802,N_7855);
nand U7985 (N_7985,N_7923,N_7931);
and U7986 (N_7986,N_7930,N_7919);
nand U7987 (N_7987,N_7858,N_7804);
xor U7988 (N_7988,N_7822,N_7932);
nand U7989 (N_7989,N_7868,N_7843);
xnor U7990 (N_7990,N_7829,N_7857);
nor U7991 (N_7991,N_7806,N_7947);
or U7992 (N_7992,N_7820,N_7920);
or U7993 (N_7993,N_7897,N_7814);
nand U7994 (N_7994,N_7813,N_7884);
nand U7995 (N_7995,N_7877,N_7940);
or U7996 (N_7996,N_7874,N_7891);
nor U7997 (N_7997,N_7922,N_7800);
and U7998 (N_7998,N_7832,N_7836);
nor U7999 (N_7999,N_7948,N_7863);
or U8000 (N_8000,N_7810,N_7926);
xor U8001 (N_8001,N_7928,N_7815);
xnor U8002 (N_8002,N_7878,N_7833);
nor U8003 (N_8003,N_7943,N_7865);
nand U8004 (N_8004,N_7807,N_7902);
and U8005 (N_8005,N_7938,N_7892);
or U8006 (N_8006,N_7830,N_7817);
nor U8007 (N_8007,N_7835,N_7937);
nor U8008 (N_8008,N_7941,N_7881);
and U8009 (N_8009,N_7853,N_7818);
nand U8010 (N_8010,N_7866,N_7929);
or U8011 (N_8011,N_7811,N_7809);
nor U8012 (N_8012,N_7851,N_7844);
and U8013 (N_8013,N_7921,N_7870);
or U8014 (N_8014,N_7867,N_7876);
nor U8015 (N_8015,N_7914,N_7927);
nor U8016 (N_8016,N_7831,N_7861);
nand U8017 (N_8017,N_7905,N_7934);
or U8018 (N_8018,N_7816,N_7801);
or U8019 (N_8019,N_7839,N_7904);
xor U8020 (N_8020,N_7933,N_7888);
or U8021 (N_8021,N_7821,N_7896);
nor U8022 (N_8022,N_7871,N_7860);
or U8023 (N_8023,N_7894,N_7900);
nor U8024 (N_8024,N_7935,N_7942);
nor U8025 (N_8025,N_7916,N_7933);
xor U8026 (N_8026,N_7897,N_7869);
xnor U8027 (N_8027,N_7894,N_7801);
and U8028 (N_8028,N_7931,N_7910);
or U8029 (N_8029,N_7832,N_7949);
or U8030 (N_8030,N_7903,N_7824);
nand U8031 (N_8031,N_7822,N_7852);
nor U8032 (N_8032,N_7907,N_7922);
xor U8033 (N_8033,N_7870,N_7895);
or U8034 (N_8034,N_7918,N_7820);
and U8035 (N_8035,N_7919,N_7944);
and U8036 (N_8036,N_7890,N_7927);
or U8037 (N_8037,N_7811,N_7900);
nand U8038 (N_8038,N_7945,N_7821);
and U8039 (N_8039,N_7804,N_7851);
nor U8040 (N_8040,N_7901,N_7867);
or U8041 (N_8041,N_7907,N_7901);
nand U8042 (N_8042,N_7896,N_7944);
nand U8043 (N_8043,N_7941,N_7882);
or U8044 (N_8044,N_7911,N_7818);
nor U8045 (N_8045,N_7889,N_7816);
nor U8046 (N_8046,N_7894,N_7880);
or U8047 (N_8047,N_7845,N_7881);
or U8048 (N_8048,N_7891,N_7838);
and U8049 (N_8049,N_7818,N_7928);
nor U8050 (N_8050,N_7900,N_7853);
or U8051 (N_8051,N_7827,N_7833);
xor U8052 (N_8052,N_7873,N_7923);
nand U8053 (N_8053,N_7815,N_7897);
xnor U8054 (N_8054,N_7897,N_7827);
nor U8055 (N_8055,N_7840,N_7865);
or U8056 (N_8056,N_7941,N_7923);
and U8057 (N_8057,N_7928,N_7887);
or U8058 (N_8058,N_7836,N_7948);
nor U8059 (N_8059,N_7915,N_7947);
and U8060 (N_8060,N_7921,N_7839);
xnor U8061 (N_8061,N_7869,N_7940);
or U8062 (N_8062,N_7818,N_7832);
or U8063 (N_8063,N_7824,N_7895);
nand U8064 (N_8064,N_7806,N_7929);
and U8065 (N_8065,N_7898,N_7859);
xnor U8066 (N_8066,N_7848,N_7910);
nor U8067 (N_8067,N_7879,N_7937);
xor U8068 (N_8068,N_7868,N_7894);
xnor U8069 (N_8069,N_7807,N_7945);
nand U8070 (N_8070,N_7879,N_7839);
xnor U8071 (N_8071,N_7851,N_7873);
xnor U8072 (N_8072,N_7824,N_7915);
xor U8073 (N_8073,N_7813,N_7886);
xnor U8074 (N_8074,N_7907,N_7906);
and U8075 (N_8075,N_7806,N_7855);
nand U8076 (N_8076,N_7838,N_7830);
nand U8077 (N_8077,N_7804,N_7923);
nor U8078 (N_8078,N_7888,N_7817);
or U8079 (N_8079,N_7916,N_7811);
nor U8080 (N_8080,N_7870,N_7939);
xnor U8081 (N_8081,N_7859,N_7889);
nand U8082 (N_8082,N_7925,N_7946);
xor U8083 (N_8083,N_7891,N_7920);
nand U8084 (N_8084,N_7858,N_7812);
nor U8085 (N_8085,N_7838,N_7836);
and U8086 (N_8086,N_7814,N_7874);
or U8087 (N_8087,N_7847,N_7818);
xnor U8088 (N_8088,N_7934,N_7863);
and U8089 (N_8089,N_7863,N_7946);
nand U8090 (N_8090,N_7942,N_7872);
or U8091 (N_8091,N_7882,N_7827);
nand U8092 (N_8092,N_7859,N_7857);
or U8093 (N_8093,N_7935,N_7931);
or U8094 (N_8094,N_7903,N_7884);
or U8095 (N_8095,N_7876,N_7934);
and U8096 (N_8096,N_7837,N_7818);
nand U8097 (N_8097,N_7836,N_7822);
nor U8098 (N_8098,N_7810,N_7918);
nand U8099 (N_8099,N_7857,N_7910);
nor U8100 (N_8100,N_8047,N_7967);
xnor U8101 (N_8101,N_8044,N_8032);
or U8102 (N_8102,N_8010,N_8082);
nor U8103 (N_8103,N_8056,N_8094);
or U8104 (N_8104,N_8012,N_7955);
and U8105 (N_8105,N_7960,N_7972);
or U8106 (N_8106,N_8051,N_8045);
xnor U8107 (N_8107,N_8035,N_8055);
nor U8108 (N_8108,N_8089,N_8039);
xor U8109 (N_8109,N_7973,N_8066);
and U8110 (N_8110,N_8067,N_8096);
nor U8111 (N_8111,N_8093,N_8073);
or U8112 (N_8112,N_8088,N_8018);
or U8113 (N_8113,N_7968,N_7999);
xnor U8114 (N_8114,N_8024,N_8098);
and U8115 (N_8115,N_8091,N_8041);
or U8116 (N_8116,N_8075,N_7989);
nand U8117 (N_8117,N_8011,N_8020);
or U8118 (N_8118,N_8050,N_8009);
and U8119 (N_8119,N_8076,N_7977);
or U8120 (N_8120,N_8037,N_8092);
or U8121 (N_8121,N_8071,N_8061);
or U8122 (N_8122,N_7959,N_8030);
or U8123 (N_8123,N_7954,N_8084);
nor U8124 (N_8124,N_7971,N_8079);
xnor U8125 (N_8125,N_8033,N_8019);
nor U8126 (N_8126,N_8048,N_7975);
nand U8127 (N_8127,N_7965,N_8074);
and U8128 (N_8128,N_8028,N_8002);
and U8129 (N_8129,N_7987,N_8078);
nand U8130 (N_8130,N_7982,N_8099);
nor U8131 (N_8131,N_8008,N_7962);
or U8132 (N_8132,N_8046,N_8022);
xor U8133 (N_8133,N_7956,N_8081);
and U8134 (N_8134,N_8083,N_8053);
xnor U8135 (N_8135,N_8001,N_7952);
nor U8136 (N_8136,N_8031,N_7953);
nand U8137 (N_8137,N_8080,N_8023);
or U8138 (N_8138,N_8043,N_8027);
and U8139 (N_8139,N_7983,N_8049);
nand U8140 (N_8140,N_8070,N_8007);
or U8141 (N_8141,N_7992,N_7958);
or U8142 (N_8142,N_8059,N_8064);
or U8143 (N_8143,N_7961,N_7964);
or U8144 (N_8144,N_8054,N_7981);
and U8145 (N_8145,N_8085,N_8077);
and U8146 (N_8146,N_7957,N_7998);
and U8147 (N_8147,N_7995,N_8097);
and U8148 (N_8148,N_8000,N_8052);
xor U8149 (N_8149,N_8060,N_8014);
and U8150 (N_8150,N_7994,N_8038);
nand U8151 (N_8151,N_7980,N_7985);
nor U8152 (N_8152,N_8040,N_8029);
xor U8153 (N_8153,N_8026,N_8063);
xor U8154 (N_8154,N_7993,N_8072);
xor U8155 (N_8155,N_8034,N_8062);
nor U8156 (N_8156,N_7976,N_8015);
or U8157 (N_8157,N_7951,N_7988);
xor U8158 (N_8158,N_8087,N_8006);
or U8159 (N_8159,N_8003,N_7969);
nand U8160 (N_8160,N_8013,N_8058);
and U8161 (N_8161,N_7996,N_7978);
nor U8162 (N_8162,N_8005,N_8025);
nor U8163 (N_8163,N_8068,N_8090);
xnor U8164 (N_8164,N_8086,N_8017);
nand U8165 (N_8165,N_8021,N_7974);
nand U8166 (N_8166,N_8065,N_7966);
xnor U8167 (N_8167,N_8057,N_8036);
xor U8168 (N_8168,N_8016,N_7991);
nor U8169 (N_8169,N_7986,N_7997);
nor U8170 (N_8170,N_7963,N_8042);
and U8171 (N_8171,N_7984,N_8004);
nor U8172 (N_8172,N_7970,N_8095);
nand U8173 (N_8173,N_7950,N_7990);
nor U8174 (N_8174,N_8069,N_7979);
xnor U8175 (N_8175,N_8048,N_8033);
nor U8176 (N_8176,N_8018,N_7974);
or U8177 (N_8177,N_8067,N_7951);
or U8178 (N_8178,N_8027,N_7998);
nor U8179 (N_8179,N_8040,N_8001);
nand U8180 (N_8180,N_7981,N_8096);
nor U8181 (N_8181,N_8007,N_7999);
xor U8182 (N_8182,N_8049,N_7974);
xor U8183 (N_8183,N_7950,N_8059);
nor U8184 (N_8184,N_7971,N_7977);
nor U8185 (N_8185,N_8039,N_8063);
xor U8186 (N_8186,N_7970,N_8074);
or U8187 (N_8187,N_8034,N_7974);
nand U8188 (N_8188,N_7969,N_7990);
xor U8189 (N_8189,N_8069,N_8056);
xor U8190 (N_8190,N_8016,N_7965);
xnor U8191 (N_8191,N_8051,N_7988);
xnor U8192 (N_8192,N_8095,N_7955);
or U8193 (N_8193,N_8081,N_7967);
and U8194 (N_8194,N_8059,N_8000);
xnor U8195 (N_8195,N_7988,N_7958);
nor U8196 (N_8196,N_8090,N_7996);
nand U8197 (N_8197,N_7963,N_8071);
xor U8198 (N_8198,N_7986,N_8011);
nor U8199 (N_8199,N_7992,N_8073);
xor U8200 (N_8200,N_8035,N_8066);
and U8201 (N_8201,N_8013,N_7954);
or U8202 (N_8202,N_8010,N_8020);
xor U8203 (N_8203,N_8087,N_8009);
nand U8204 (N_8204,N_8082,N_7984);
or U8205 (N_8205,N_7961,N_8071);
and U8206 (N_8206,N_7982,N_8042);
and U8207 (N_8207,N_7962,N_7979);
nor U8208 (N_8208,N_7996,N_8019);
xnor U8209 (N_8209,N_8062,N_7977);
xnor U8210 (N_8210,N_7989,N_8039);
nor U8211 (N_8211,N_8023,N_8092);
and U8212 (N_8212,N_7961,N_8072);
or U8213 (N_8213,N_8032,N_7999);
xor U8214 (N_8214,N_8080,N_7987);
and U8215 (N_8215,N_7973,N_8030);
and U8216 (N_8216,N_7987,N_7960);
nand U8217 (N_8217,N_8018,N_7953);
or U8218 (N_8218,N_7957,N_8025);
nand U8219 (N_8219,N_8091,N_8049);
nand U8220 (N_8220,N_7955,N_8089);
or U8221 (N_8221,N_7967,N_8083);
and U8222 (N_8222,N_7974,N_8022);
or U8223 (N_8223,N_8079,N_8090);
nor U8224 (N_8224,N_7984,N_8009);
xnor U8225 (N_8225,N_8058,N_8029);
nor U8226 (N_8226,N_8004,N_8081);
nand U8227 (N_8227,N_8090,N_8098);
or U8228 (N_8228,N_8058,N_8035);
or U8229 (N_8229,N_8078,N_8011);
xnor U8230 (N_8230,N_7952,N_8066);
nor U8231 (N_8231,N_7999,N_8080);
and U8232 (N_8232,N_8096,N_8007);
xor U8233 (N_8233,N_7962,N_8049);
nor U8234 (N_8234,N_8062,N_8043);
and U8235 (N_8235,N_7988,N_8062);
and U8236 (N_8236,N_8010,N_8003);
xnor U8237 (N_8237,N_8075,N_7977);
xnor U8238 (N_8238,N_8059,N_7955);
xnor U8239 (N_8239,N_8035,N_8037);
nor U8240 (N_8240,N_8010,N_8057);
nor U8241 (N_8241,N_7988,N_8029);
nor U8242 (N_8242,N_8055,N_8093);
and U8243 (N_8243,N_8051,N_8046);
or U8244 (N_8244,N_7950,N_8096);
and U8245 (N_8245,N_7980,N_8097);
nor U8246 (N_8246,N_8002,N_8043);
nand U8247 (N_8247,N_8096,N_8052);
and U8248 (N_8248,N_7997,N_8021);
nor U8249 (N_8249,N_7980,N_8002);
nor U8250 (N_8250,N_8132,N_8206);
and U8251 (N_8251,N_8177,N_8139);
or U8252 (N_8252,N_8209,N_8110);
and U8253 (N_8253,N_8238,N_8242);
or U8254 (N_8254,N_8223,N_8166);
nor U8255 (N_8255,N_8131,N_8228);
nand U8256 (N_8256,N_8195,N_8170);
nand U8257 (N_8257,N_8126,N_8106);
nor U8258 (N_8258,N_8232,N_8130);
nand U8259 (N_8259,N_8158,N_8247);
xor U8260 (N_8260,N_8118,N_8148);
nor U8261 (N_8261,N_8113,N_8154);
and U8262 (N_8262,N_8194,N_8101);
or U8263 (N_8263,N_8171,N_8202);
and U8264 (N_8264,N_8155,N_8161);
nand U8265 (N_8265,N_8122,N_8236);
or U8266 (N_8266,N_8229,N_8150);
xnor U8267 (N_8267,N_8149,N_8203);
and U8268 (N_8268,N_8127,N_8117);
xnor U8269 (N_8269,N_8239,N_8102);
nand U8270 (N_8270,N_8215,N_8124);
or U8271 (N_8271,N_8186,N_8189);
and U8272 (N_8272,N_8157,N_8164);
nand U8273 (N_8273,N_8241,N_8199);
and U8274 (N_8274,N_8167,N_8190);
nor U8275 (N_8275,N_8141,N_8196);
or U8276 (N_8276,N_8244,N_8147);
nor U8277 (N_8277,N_8192,N_8140);
or U8278 (N_8278,N_8103,N_8128);
nor U8279 (N_8279,N_8152,N_8129);
xnor U8280 (N_8280,N_8248,N_8144);
nor U8281 (N_8281,N_8201,N_8153);
nor U8282 (N_8282,N_8207,N_8225);
or U8283 (N_8283,N_8137,N_8208);
xnor U8284 (N_8284,N_8226,N_8125);
xor U8285 (N_8285,N_8178,N_8221);
or U8286 (N_8286,N_8135,N_8114);
nand U8287 (N_8287,N_8172,N_8134);
and U8288 (N_8288,N_8151,N_8197);
xor U8289 (N_8289,N_8214,N_8174);
or U8290 (N_8290,N_8185,N_8200);
or U8291 (N_8291,N_8224,N_8187);
nand U8292 (N_8292,N_8100,N_8159);
or U8293 (N_8293,N_8240,N_8182);
or U8294 (N_8294,N_8218,N_8175);
or U8295 (N_8295,N_8145,N_8179);
xnor U8296 (N_8296,N_8181,N_8249);
nand U8297 (N_8297,N_8243,N_8191);
nor U8298 (N_8298,N_8142,N_8235);
nor U8299 (N_8299,N_8233,N_8212);
nor U8300 (N_8300,N_8205,N_8213);
and U8301 (N_8301,N_8176,N_8245);
nor U8302 (N_8302,N_8133,N_8237);
nand U8303 (N_8303,N_8246,N_8111);
xor U8304 (N_8304,N_8146,N_8227);
nor U8305 (N_8305,N_8234,N_8230);
or U8306 (N_8306,N_8165,N_8112);
or U8307 (N_8307,N_8123,N_8169);
nand U8308 (N_8308,N_8168,N_8198);
nor U8309 (N_8309,N_8211,N_8184);
nor U8310 (N_8310,N_8108,N_8162);
and U8311 (N_8311,N_8217,N_8121);
or U8312 (N_8312,N_8193,N_8138);
nand U8313 (N_8313,N_8180,N_8204);
xor U8314 (N_8314,N_8104,N_8107);
nand U8315 (N_8315,N_8210,N_8143);
xor U8316 (N_8316,N_8183,N_8105);
nor U8317 (N_8317,N_8231,N_8160);
xor U8318 (N_8318,N_8216,N_8156);
xnor U8319 (N_8319,N_8119,N_8222);
nor U8320 (N_8320,N_8163,N_8219);
and U8321 (N_8321,N_8115,N_8120);
xnor U8322 (N_8322,N_8220,N_8188);
nor U8323 (N_8323,N_8116,N_8136);
nor U8324 (N_8324,N_8109,N_8173);
nand U8325 (N_8325,N_8220,N_8177);
or U8326 (N_8326,N_8150,N_8137);
xnor U8327 (N_8327,N_8106,N_8238);
or U8328 (N_8328,N_8238,N_8143);
xor U8329 (N_8329,N_8231,N_8188);
xnor U8330 (N_8330,N_8233,N_8120);
xor U8331 (N_8331,N_8141,N_8161);
nand U8332 (N_8332,N_8121,N_8124);
and U8333 (N_8333,N_8199,N_8230);
nor U8334 (N_8334,N_8134,N_8137);
xor U8335 (N_8335,N_8217,N_8231);
nor U8336 (N_8336,N_8215,N_8152);
or U8337 (N_8337,N_8247,N_8227);
nor U8338 (N_8338,N_8161,N_8239);
and U8339 (N_8339,N_8183,N_8237);
nand U8340 (N_8340,N_8211,N_8246);
or U8341 (N_8341,N_8197,N_8244);
or U8342 (N_8342,N_8227,N_8148);
nand U8343 (N_8343,N_8231,N_8247);
and U8344 (N_8344,N_8213,N_8118);
and U8345 (N_8345,N_8241,N_8137);
nand U8346 (N_8346,N_8226,N_8161);
nand U8347 (N_8347,N_8118,N_8194);
nor U8348 (N_8348,N_8147,N_8182);
xor U8349 (N_8349,N_8139,N_8183);
nor U8350 (N_8350,N_8196,N_8206);
nor U8351 (N_8351,N_8231,N_8128);
or U8352 (N_8352,N_8180,N_8114);
or U8353 (N_8353,N_8128,N_8234);
or U8354 (N_8354,N_8146,N_8181);
and U8355 (N_8355,N_8173,N_8242);
nor U8356 (N_8356,N_8225,N_8218);
xor U8357 (N_8357,N_8123,N_8128);
xnor U8358 (N_8358,N_8241,N_8218);
nor U8359 (N_8359,N_8231,N_8138);
and U8360 (N_8360,N_8102,N_8182);
xnor U8361 (N_8361,N_8245,N_8146);
nor U8362 (N_8362,N_8208,N_8178);
or U8363 (N_8363,N_8206,N_8171);
nand U8364 (N_8364,N_8226,N_8238);
nand U8365 (N_8365,N_8139,N_8124);
xor U8366 (N_8366,N_8114,N_8171);
xnor U8367 (N_8367,N_8195,N_8166);
or U8368 (N_8368,N_8187,N_8164);
or U8369 (N_8369,N_8234,N_8213);
or U8370 (N_8370,N_8201,N_8228);
xnor U8371 (N_8371,N_8188,N_8138);
nand U8372 (N_8372,N_8209,N_8141);
xor U8373 (N_8373,N_8215,N_8224);
and U8374 (N_8374,N_8189,N_8210);
or U8375 (N_8375,N_8212,N_8138);
and U8376 (N_8376,N_8117,N_8142);
and U8377 (N_8377,N_8222,N_8211);
nor U8378 (N_8378,N_8164,N_8194);
and U8379 (N_8379,N_8162,N_8188);
or U8380 (N_8380,N_8240,N_8125);
xnor U8381 (N_8381,N_8206,N_8129);
and U8382 (N_8382,N_8215,N_8233);
nor U8383 (N_8383,N_8106,N_8183);
xnor U8384 (N_8384,N_8118,N_8119);
and U8385 (N_8385,N_8119,N_8206);
xnor U8386 (N_8386,N_8156,N_8185);
nand U8387 (N_8387,N_8228,N_8173);
nand U8388 (N_8388,N_8210,N_8209);
or U8389 (N_8389,N_8161,N_8139);
xor U8390 (N_8390,N_8178,N_8197);
or U8391 (N_8391,N_8241,N_8151);
nor U8392 (N_8392,N_8206,N_8243);
or U8393 (N_8393,N_8133,N_8208);
xnor U8394 (N_8394,N_8156,N_8108);
or U8395 (N_8395,N_8125,N_8231);
nand U8396 (N_8396,N_8197,N_8184);
nand U8397 (N_8397,N_8219,N_8234);
and U8398 (N_8398,N_8189,N_8143);
nand U8399 (N_8399,N_8195,N_8202);
and U8400 (N_8400,N_8372,N_8361);
xor U8401 (N_8401,N_8260,N_8269);
nor U8402 (N_8402,N_8395,N_8398);
nand U8403 (N_8403,N_8265,N_8326);
or U8404 (N_8404,N_8349,N_8351);
xnor U8405 (N_8405,N_8280,N_8320);
nand U8406 (N_8406,N_8263,N_8368);
or U8407 (N_8407,N_8381,N_8303);
xnor U8408 (N_8408,N_8360,N_8331);
or U8409 (N_8409,N_8370,N_8250);
nor U8410 (N_8410,N_8310,N_8386);
and U8411 (N_8411,N_8282,N_8288);
or U8412 (N_8412,N_8252,N_8287);
or U8413 (N_8413,N_8325,N_8311);
and U8414 (N_8414,N_8305,N_8391);
xnor U8415 (N_8415,N_8394,N_8388);
nor U8416 (N_8416,N_8307,N_8332);
and U8417 (N_8417,N_8369,N_8354);
or U8418 (N_8418,N_8261,N_8299);
or U8419 (N_8419,N_8383,N_8290);
nor U8420 (N_8420,N_8297,N_8306);
nand U8421 (N_8421,N_8289,N_8379);
nand U8422 (N_8422,N_8367,N_8266);
nor U8423 (N_8423,N_8251,N_8316);
nor U8424 (N_8424,N_8276,N_8301);
and U8425 (N_8425,N_8359,N_8283);
or U8426 (N_8426,N_8302,N_8323);
or U8427 (N_8427,N_8380,N_8258);
nand U8428 (N_8428,N_8279,N_8378);
or U8429 (N_8429,N_8340,N_8322);
and U8430 (N_8430,N_8376,N_8335);
or U8431 (N_8431,N_8382,N_8371);
nand U8432 (N_8432,N_8362,N_8344);
nor U8433 (N_8433,N_8339,N_8374);
nand U8434 (N_8434,N_8328,N_8313);
nor U8435 (N_8435,N_8356,N_8273);
nor U8436 (N_8436,N_8365,N_8385);
xnor U8437 (N_8437,N_8314,N_8304);
nand U8438 (N_8438,N_8284,N_8286);
nand U8439 (N_8439,N_8377,N_8342);
nand U8440 (N_8440,N_8330,N_8281);
nand U8441 (N_8441,N_8327,N_8318);
nand U8442 (N_8442,N_8357,N_8384);
nor U8443 (N_8443,N_8393,N_8271);
or U8444 (N_8444,N_8253,N_8338);
nand U8445 (N_8445,N_8262,N_8294);
nand U8446 (N_8446,N_8300,N_8272);
xor U8447 (N_8447,N_8312,N_8355);
nor U8448 (N_8448,N_8268,N_8348);
nand U8449 (N_8449,N_8324,N_8392);
and U8450 (N_8450,N_8256,N_8347);
nand U8451 (N_8451,N_8295,N_8350);
and U8452 (N_8452,N_8277,N_8317);
and U8453 (N_8453,N_8373,N_8399);
xnor U8454 (N_8454,N_8363,N_8343);
xor U8455 (N_8455,N_8333,N_8285);
and U8456 (N_8456,N_8396,N_8387);
and U8457 (N_8457,N_8308,N_8275);
nand U8458 (N_8458,N_8257,N_8352);
or U8459 (N_8459,N_8296,N_8254);
nand U8460 (N_8460,N_8390,N_8375);
xor U8461 (N_8461,N_8292,N_8291);
nor U8462 (N_8462,N_8315,N_8293);
and U8463 (N_8463,N_8397,N_8329);
nor U8464 (N_8464,N_8364,N_8259);
and U8465 (N_8465,N_8334,N_8278);
nand U8466 (N_8466,N_8341,N_8321);
nand U8467 (N_8467,N_8274,N_8353);
nor U8468 (N_8468,N_8309,N_8267);
nor U8469 (N_8469,N_8336,N_8319);
nand U8470 (N_8470,N_8264,N_8389);
xor U8471 (N_8471,N_8255,N_8366);
nor U8472 (N_8472,N_8345,N_8270);
or U8473 (N_8473,N_8358,N_8337);
nor U8474 (N_8474,N_8346,N_8298);
xor U8475 (N_8475,N_8257,N_8369);
nand U8476 (N_8476,N_8259,N_8260);
nor U8477 (N_8477,N_8260,N_8317);
and U8478 (N_8478,N_8340,N_8352);
or U8479 (N_8479,N_8297,N_8271);
and U8480 (N_8480,N_8325,N_8260);
and U8481 (N_8481,N_8392,N_8251);
nand U8482 (N_8482,N_8348,N_8358);
xor U8483 (N_8483,N_8300,N_8355);
nor U8484 (N_8484,N_8351,N_8386);
or U8485 (N_8485,N_8263,N_8286);
nand U8486 (N_8486,N_8324,N_8269);
xor U8487 (N_8487,N_8338,N_8267);
or U8488 (N_8488,N_8377,N_8272);
and U8489 (N_8489,N_8294,N_8386);
or U8490 (N_8490,N_8372,N_8289);
xor U8491 (N_8491,N_8313,N_8341);
or U8492 (N_8492,N_8295,N_8395);
and U8493 (N_8493,N_8284,N_8279);
or U8494 (N_8494,N_8396,N_8302);
or U8495 (N_8495,N_8253,N_8281);
xnor U8496 (N_8496,N_8266,N_8349);
and U8497 (N_8497,N_8318,N_8303);
nand U8498 (N_8498,N_8263,N_8359);
nor U8499 (N_8499,N_8363,N_8362);
nor U8500 (N_8500,N_8358,N_8317);
nand U8501 (N_8501,N_8276,N_8271);
nand U8502 (N_8502,N_8263,N_8366);
nand U8503 (N_8503,N_8339,N_8326);
xnor U8504 (N_8504,N_8359,N_8305);
or U8505 (N_8505,N_8257,N_8374);
nand U8506 (N_8506,N_8365,N_8391);
nor U8507 (N_8507,N_8390,N_8289);
nand U8508 (N_8508,N_8387,N_8397);
xnor U8509 (N_8509,N_8331,N_8324);
nand U8510 (N_8510,N_8273,N_8396);
xnor U8511 (N_8511,N_8282,N_8295);
nand U8512 (N_8512,N_8277,N_8373);
nand U8513 (N_8513,N_8277,N_8334);
and U8514 (N_8514,N_8326,N_8288);
and U8515 (N_8515,N_8353,N_8348);
nor U8516 (N_8516,N_8387,N_8334);
and U8517 (N_8517,N_8383,N_8267);
or U8518 (N_8518,N_8335,N_8328);
or U8519 (N_8519,N_8353,N_8276);
nand U8520 (N_8520,N_8309,N_8366);
nand U8521 (N_8521,N_8307,N_8396);
and U8522 (N_8522,N_8342,N_8354);
or U8523 (N_8523,N_8348,N_8332);
nor U8524 (N_8524,N_8350,N_8261);
or U8525 (N_8525,N_8325,N_8282);
nand U8526 (N_8526,N_8391,N_8293);
nor U8527 (N_8527,N_8344,N_8322);
nand U8528 (N_8528,N_8318,N_8373);
nand U8529 (N_8529,N_8271,N_8377);
nor U8530 (N_8530,N_8397,N_8296);
nand U8531 (N_8531,N_8271,N_8339);
and U8532 (N_8532,N_8357,N_8288);
nor U8533 (N_8533,N_8271,N_8272);
and U8534 (N_8534,N_8273,N_8275);
and U8535 (N_8535,N_8363,N_8339);
xor U8536 (N_8536,N_8343,N_8351);
nand U8537 (N_8537,N_8346,N_8310);
or U8538 (N_8538,N_8272,N_8372);
and U8539 (N_8539,N_8340,N_8362);
and U8540 (N_8540,N_8337,N_8320);
and U8541 (N_8541,N_8365,N_8253);
or U8542 (N_8542,N_8339,N_8365);
nand U8543 (N_8543,N_8367,N_8296);
nand U8544 (N_8544,N_8266,N_8360);
xnor U8545 (N_8545,N_8374,N_8274);
or U8546 (N_8546,N_8312,N_8381);
or U8547 (N_8547,N_8355,N_8277);
xnor U8548 (N_8548,N_8331,N_8362);
nor U8549 (N_8549,N_8388,N_8348);
xnor U8550 (N_8550,N_8434,N_8435);
or U8551 (N_8551,N_8464,N_8401);
or U8552 (N_8552,N_8541,N_8408);
nand U8553 (N_8553,N_8505,N_8500);
nand U8554 (N_8554,N_8511,N_8446);
and U8555 (N_8555,N_8473,N_8415);
and U8556 (N_8556,N_8516,N_8439);
or U8557 (N_8557,N_8403,N_8444);
xnor U8558 (N_8558,N_8449,N_8529);
nand U8559 (N_8559,N_8432,N_8538);
or U8560 (N_8560,N_8427,N_8531);
nor U8561 (N_8561,N_8419,N_8466);
or U8562 (N_8562,N_8527,N_8518);
xnor U8563 (N_8563,N_8496,N_8507);
nor U8564 (N_8564,N_8440,N_8478);
or U8565 (N_8565,N_8503,N_8498);
xnor U8566 (N_8566,N_8521,N_8520);
xor U8567 (N_8567,N_8429,N_8479);
nand U8568 (N_8568,N_8407,N_8420);
nor U8569 (N_8569,N_8418,N_8459);
nor U8570 (N_8570,N_8467,N_8471);
or U8571 (N_8571,N_8542,N_8412);
and U8572 (N_8572,N_8512,N_8448);
xnor U8573 (N_8573,N_8442,N_8428);
nor U8574 (N_8574,N_8411,N_8499);
nand U8575 (N_8575,N_8438,N_8400);
xor U8576 (N_8576,N_8447,N_8517);
nor U8577 (N_8577,N_8483,N_8453);
nand U8578 (N_8578,N_8534,N_8417);
and U8579 (N_8579,N_8470,N_8406);
nor U8580 (N_8580,N_8508,N_8480);
or U8581 (N_8581,N_8457,N_8533);
and U8582 (N_8582,N_8497,N_8509);
nor U8583 (N_8583,N_8515,N_8477);
nand U8584 (N_8584,N_8425,N_8528);
nand U8585 (N_8585,N_8426,N_8422);
and U8586 (N_8586,N_8548,N_8460);
and U8587 (N_8587,N_8539,N_8445);
xnor U8588 (N_8588,N_8482,N_8532);
xor U8589 (N_8589,N_8476,N_8462);
or U8590 (N_8590,N_8540,N_8535);
xor U8591 (N_8591,N_8547,N_8524);
xnor U8592 (N_8592,N_8495,N_8404);
nand U8593 (N_8593,N_8485,N_8486);
nand U8594 (N_8594,N_8488,N_8506);
or U8595 (N_8595,N_8484,N_8546);
nand U8596 (N_8596,N_8409,N_8443);
and U8597 (N_8597,N_8431,N_8530);
or U8598 (N_8598,N_8414,N_8514);
or U8599 (N_8599,N_8452,N_8504);
nand U8600 (N_8600,N_8469,N_8455);
nand U8601 (N_8601,N_8549,N_8502);
or U8602 (N_8602,N_8490,N_8410);
nand U8603 (N_8603,N_8436,N_8522);
xor U8604 (N_8604,N_8492,N_8402);
and U8605 (N_8605,N_8474,N_8454);
or U8606 (N_8606,N_8433,N_8416);
nor U8607 (N_8607,N_8501,N_8487);
or U8608 (N_8608,N_8489,N_8405);
xor U8609 (N_8609,N_8481,N_8441);
nor U8610 (N_8610,N_8450,N_8475);
xnor U8611 (N_8611,N_8430,N_8526);
nor U8612 (N_8612,N_8465,N_8413);
and U8613 (N_8613,N_8491,N_8423);
nor U8614 (N_8614,N_8437,N_8458);
nor U8615 (N_8615,N_8510,N_8463);
nand U8616 (N_8616,N_8525,N_8472);
nor U8617 (N_8617,N_8537,N_8513);
nor U8618 (N_8618,N_8523,N_8545);
xor U8619 (N_8619,N_8461,N_8536);
nor U8620 (N_8620,N_8494,N_8421);
nand U8621 (N_8621,N_8456,N_8543);
nand U8622 (N_8622,N_8424,N_8468);
xor U8623 (N_8623,N_8519,N_8493);
nor U8624 (N_8624,N_8451,N_8544);
xnor U8625 (N_8625,N_8482,N_8406);
and U8626 (N_8626,N_8479,N_8401);
nand U8627 (N_8627,N_8535,N_8523);
or U8628 (N_8628,N_8497,N_8444);
nand U8629 (N_8629,N_8542,N_8435);
xnor U8630 (N_8630,N_8474,N_8445);
nand U8631 (N_8631,N_8457,N_8512);
and U8632 (N_8632,N_8452,N_8526);
and U8633 (N_8633,N_8535,N_8512);
nand U8634 (N_8634,N_8548,N_8439);
nor U8635 (N_8635,N_8417,N_8538);
and U8636 (N_8636,N_8513,N_8505);
or U8637 (N_8637,N_8498,N_8404);
nor U8638 (N_8638,N_8521,N_8485);
or U8639 (N_8639,N_8423,N_8457);
nor U8640 (N_8640,N_8505,N_8482);
or U8641 (N_8641,N_8423,N_8434);
or U8642 (N_8642,N_8425,N_8414);
or U8643 (N_8643,N_8432,N_8478);
and U8644 (N_8644,N_8546,N_8508);
and U8645 (N_8645,N_8533,N_8549);
nor U8646 (N_8646,N_8541,N_8476);
xnor U8647 (N_8647,N_8468,N_8532);
and U8648 (N_8648,N_8510,N_8418);
nor U8649 (N_8649,N_8477,N_8473);
and U8650 (N_8650,N_8441,N_8454);
nor U8651 (N_8651,N_8462,N_8527);
nor U8652 (N_8652,N_8419,N_8461);
nand U8653 (N_8653,N_8547,N_8458);
xnor U8654 (N_8654,N_8522,N_8544);
nor U8655 (N_8655,N_8450,N_8492);
xor U8656 (N_8656,N_8499,N_8544);
and U8657 (N_8657,N_8535,N_8463);
nor U8658 (N_8658,N_8454,N_8546);
nor U8659 (N_8659,N_8513,N_8481);
and U8660 (N_8660,N_8500,N_8510);
nor U8661 (N_8661,N_8456,N_8488);
nand U8662 (N_8662,N_8504,N_8508);
xor U8663 (N_8663,N_8534,N_8473);
xnor U8664 (N_8664,N_8433,N_8409);
nand U8665 (N_8665,N_8508,N_8519);
and U8666 (N_8666,N_8504,N_8526);
or U8667 (N_8667,N_8533,N_8480);
or U8668 (N_8668,N_8538,N_8406);
xor U8669 (N_8669,N_8506,N_8543);
xnor U8670 (N_8670,N_8548,N_8451);
and U8671 (N_8671,N_8548,N_8424);
or U8672 (N_8672,N_8480,N_8458);
nand U8673 (N_8673,N_8465,N_8545);
or U8674 (N_8674,N_8502,N_8542);
and U8675 (N_8675,N_8547,N_8456);
or U8676 (N_8676,N_8447,N_8523);
xor U8677 (N_8677,N_8437,N_8419);
or U8678 (N_8678,N_8507,N_8457);
nor U8679 (N_8679,N_8532,N_8400);
xnor U8680 (N_8680,N_8505,N_8412);
or U8681 (N_8681,N_8411,N_8446);
and U8682 (N_8682,N_8473,N_8528);
xnor U8683 (N_8683,N_8528,N_8536);
or U8684 (N_8684,N_8487,N_8401);
or U8685 (N_8685,N_8442,N_8433);
xnor U8686 (N_8686,N_8536,N_8472);
nand U8687 (N_8687,N_8486,N_8448);
nand U8688 (N_8688,N_8408,N_8472);
nor U8689 (N_8689,N_8536,N_8458);
and U8690 (N_8690,N_8534,N_8522);
and U8691 (N_8691,N_8543,N_8441);
and U8692 (N_8692,N_8525,N_8464);
nor U8693 (N_8693,N_8520,N_8435);
nand U8694 (N_8694,N_8476,N_8427);
or U8695 (N_8695,N_8421,N_8471);
xor U8696 (N_8696,N_8483,N_8488);
nand U8697 (N_8697,N_8490,N_8512);
nor U8698 (N_8698,N_8441,N_8537);
and U8699 (N_8699,N_8545,N_8522);
xor U8700 (N_8700,N_8567,N_8677);
nand U8701 (N_8701,N_8644,N_8608);
nand U8702 (N_8702,N_8666,N_8591);
and U8703 (N_8703,N_8635,N_8667);
and U8704 (N_8704,N_8647,N_8616);
nor U8705 (N_8705,N_8585,N_8695);
nor U8706 (N_8706,N_8682,N_8562);
and U8707 (N_8707,N_8661,N_8606);
xnor U8708 (N_8708,N_8602,N_8638);
and U8709 (N_8709,N_8684,N_8654);
nor U8710 (N_8710,N_8651,N_8561);
nand U8711 (N_8711,N_8572,N_8577);
nand U8712 (N_8712,N_8587,N_8565);
or U8713 (N_8713,N_8680,N_8632);
xnor U8714 (N_8714,N_8552,N_8629);
nor U8715 (N_8715,N_8662,N_8653);
nor U8716 (N_8716,N_8576,N_8643);
nor U8717 (N_8717,N_8641,N_8683);
nor U8718 (N_8718,N_8622,N_8696);
nand U8719 (N_8719,N_8551,N_8697);
xor U8720 (N_8720,N_8580,N_8681);
or U8721 (N_8721,N_8627,N_8672);
or U8722 (N_8722,N_8573,N_8671);
nand U8723 (N_8723,N_8659,N_8615);
nor U8724 (N_8724,N_8694,N_8612);
or U8725 (N_8725,N_8636,N_8620);
and U8726 (N_8726,N_8621,N_8673);
xor U8727 (N_8727,N_8613,N_8578);
nand U8728 (N_8728,N_8554,N_8656);
nor U8729 (N_8729,N_8639,N_8588);
or U8730 (N_8730,N_8664,N_8598);
xnor U8731 (N_8731,N_8586,N_8571);
nor U8732 (N_8732,N_8600,N_8560);
nor U8733 (N_8733,N_8611,N_8557);
and U8734 (N_8734,N_8698,N_8678);
and U8735 (N_8735,N_8556,N_8569);
and U8736 (N_8736,N_8607,N_8626);
nor U8737 (N_8737,N_8592,N_8674);
xnor U8738 (N_8738,N_8633,N_8668);
nand U8739 (N_8739,N_8687,N_8583);
or U8740 (N_8740,N_8614,N_8564);
nor U8741 (N_8741,N_8589,N_8693);
nand U8742 (N_8742,N_8652,N_8566);
and U8743 (N_8743,N_8675,N_8679);
xnor U8744 (N_8744,N_8563,N_8686);
xor U8745 (N_8745,N_8555,N_8619);
nand U8746 (N_8746,N_8550,N_8649);
and U8747 (N_8747,N_8581,N_8558);
or U8748 (N_8748,N_8692,N_8574);
and U8749 (N_8749,N_8665,N_8603);
xnor U8750 (N_8750,N_8630,N_8658);
or U8751 (N_8751,N_8669,N_8594);
nand U8752 (N_8752,N_8690,N_8617);
nand U8753 (N_8753,N_8624,N_8648);
xor U8754 (N_8754,N_8568,N_8590);
or U8755 (N_8755,N_8605,N_8559);
and U8756 (N_8756,N_8642,N_8640);
xor U8757 (N_8757,N_8609,N_8655);
nor U8758 (N_8758,N_8645,N_8610);
nand U8759 (N_8759,N_8618,N_8553);
or U8760 (N_8760,N_8593,N_8646);
nand U8761 (N_8761,N_8604,N_8685);
nor U8762 (N_8762,N_8579,N_8570);
nand U8763 (N_8763,N_8582,N_8628);
nand U8764 (N_8764,N_8595,N_8596);
and U8765 (N_8765,N_8637,N_8689);
xor U8766 (N_8766,N_8699,N_8625);
nor U8767 (N_8767,N_8634,N_8599);
and U8768 (N_8768,N_8663,N_8676);
nand U8769 (N_8769,N_8688,N_8575);
nand U8770 (N_8770,N_8650,N_8660);
xnor U8771 (N_8771,N_8601,N_8623);
or U8772 (N_8772,N_8691,N_8597);
and U8773 (N_8773,N_8584,N_8670);
and U8774 (N_8774,N_8631,N_8657);
nand U8775 (N_8775,N_8698,N_8636);
or U8776 (N_8776,N_8665,N_8623);
and U8777 (N_8777,N_8590,N_8610);
nand U8778 (N_8778,N_8695,N_8604);
or U8779 (N_8779,N_8679,N_8691);
or U8780 (N_8780,N_8631,N_8569);
nor U8781 (N_8781,N_8632,N_8670);
nor U8782 (N_8782,N_8600,N_8680);
nor U8783 (N_8783,N_8651,N_8662);
nand U8784 (N_8784,N_8690,N_8673);
xor U8785 (N_8785,N_8690,N_8685);
nor U8786 (N_8786,N_8696,N_8566);
or U8787 (N_8787,N_8639,N_8559);
nor U8788 (N_8788,N_8677,N_8579);
nor U8789 (N_8789,N_8553,N_8650);
and U8790 (N_8790,N_8659,N_8550);
xnor U8791 (N_8791,N_8696,N_8685);
nor U8792 (N_8792,N_8601,N_8660);
or U8793 (N_8793,N_8584,N_8550);
or U8794 (N_8794,N_8557,N_8698);
and U8795 (N_8795,N_8577,N_8690);
or U8796 (N_8796,N_8631,N_8675);
nor U8797 (N_8797,N_8695,N_8615);
or U8798 (N_8798,N_8564,N_8590);
or U8799 (N_8799,N_8608,N_8671);
and U8800 (N_8800,N_8629,N_8587);
nor U8801 (N_8801,N_8631,N_8656);
nand U8802 (N_8802,N_8694,N_8685);
and U8803 (N_8803,N_8603,N_8682);
or U8804 (N_8804,N_8572,N_8584);
xor U8805 (N_8805,N_8638,N_8599);
nand U8806 (N_8806,N_8613,N_8696);
xor U8807 (N_8807,N_8602,N_8609);
xor U8808 (N_8808,N_8561,N_8635);
and U8809 (N_8809,N_8688,N_8623);
and U8810 (N_8810,N_8683,N_8668);
nand U8811 (N_8811,N_8617,N_8693);
or U8812 (N_8812,N_8576,N_8561);
or U8813 (N_8813,N_8627,N_8639);
xnor U8814 (N_8814,N_8610,N_8594);
xnor U8815 (N_8815,N_8599,N_8612);
nor U8816 (N_8816,N_8649,N_8590);
nand U8817 (N_8817,N_8550,N_8681);
nand U8818 (N_8818,N_8633,N_8604);
xor U8819 (N_8819,N_8566,N_8657);
nand U8820 (N_8820,N_8671,N_8625);
xnor U8821 (N_8821,N_8611,N_8631);
nand U8822 (N_8822,N_8604,N_8664);
nand U8823 (N_8823,N_8699,N_8664);
nor U8824 (N_8824,N_8554,N_8695);
xnor U8825 (N_8825,N_8625,N_8690);
or U8826 (N_8826,N_8684,N_8638);
nor U8827 (N_8827,N_8667,N_8684);
nor U8828 (N_8828,N_8590,N_8653);
nand U8829 (N_8829,N_8589,N_8670);
or U8830 (N_8830,N_8602,N_8657);
xnor U8831 (N_8831,N_8664,N_8634);
xor U8832 (N_8832,N_8687,N_8557);
nand U8833 (N_8833,N_8580,N_8677);
nor U8834 (N_8834,N_8622,N_8629);
nand U8835 (N_8835,N_8627,N_8593);
nor U8836 (N_8836,N_8574,N_8671);
nand U8837 (N_8837,N_8690,N_8576);
or U8838 (N_8838,N_8573,N_8690);
xor U8839 (N_8839,N_8629,N_8599);
nor U8840 (N_8840,N_8553,N_8566);
nand U8841 (N_8841,N_8660,N_8557);
or U8842 (N_8842,N_8602,N_8601);
nand U8843 (N_8843,N_8675,N_8643);
or U8844 (N_8844,N_8666,N_8679);
nand U8845 (N_8845,N_8557,N_8559);
and U8846 (N_8846,N_8560,N_8615);
and U8847 (N_8847,N_8577,N_8648);
or U8848 (N_8848,N_8623,N_8644);
xor U8849 (N_8849,N_8605,N_8617);
and U8850 (N_8850,N_8822,N_8847);
nor U8851 (N_8851,N_8708,N_8802);
nor U8852 (N_8852,N_8761,N_8746);
nor U8853 (N_8853,N_8739,N_8801);
nor U8854 (N_8854,N_8831,N_8724);
xnor U8855 (N_8855,N_8799,N_8743);
nand U8856 (N_8856,N_8737,N_8808);
or U8857 (N_8857,N_8753,N_8702);
xnor U8858 (N_8858,N_8738,N_8744);
and U8859 (N_8859,N_8717,N_8778);
nor U8860 (N_8860,N_8712,N_8757);
xnor U8861 (N_8861,N_8843,N_8760);
and U8862 (N_8862,N_8785,N_8789);
nand U8863 (N_8863,N_8833,N_8770);
nand U8864 (N_8864,N_8820,N_8787);
and U8865 (N_8865,N_8707,N_8837);
or U8866 (N_8866,N_8719,N_8741);
or U8867 (N_8867,N_8726,N_8705);
nand U8868 (N_8868,N_8764,N_8797);
or U8869 (N_8869,N_8735,N_8718);
nor U8870 (N_8870,N_8790,N_8756);
and U8871 (N_8871,N_8765,N_8767);
xnor U8872 (N_8872,N_8710,N_8824);
nor U8873 (N_8873,N_8723,N_8832);
nand U8874 (N_8874,N_8751,N_8821);
nand U8875 (N_8875,N_8734,N_8749);
nand U8876 (N_8876,N_8836,N_8810);
or U8877 (N_8877,N_8758,N_8781);
and U8878 (N_8878,N_8812,N_8748);
and U8879 (N_8879,N_8809,N_8828);
xnor U8880 (N_8880,N_8774,N_8716);
nor U8881 (N_8881,N_8816,N_8700);
xnor U8882 (N_8882,N_8784,N_8732);
xor U8883 (N_8883,N_8762,N_8701);
and U8884 (N_8884,N_8793,N_8763);
and U8885 (N_8885,N_8792,N_8834);
and U8886 (N_8886,N_8750,N_8829);
and U8887 (N_8887,N_8840,N_8706);
or U8888 (N_8888,N_8703,N_8807);
and U8889 (N_8889,N_8733,N_8827);
or U8890 (N_8890,N_8742,N_8715);
or U8891 (N_8891,N_8804,N_8740);
xnor U8892 (N_8892,N_8817,N_8846);
and U8893 (N_8893,N_8704,N_8768);
and U8894 (N_8894,N_8796,N_8711);
nor U8895 (N_8895,N_8783,N_8800);
or U8896 (N_8896,N_8811,N_8813);
and U8897 (N_8897,N_8776,N_8754);
xor U8898 (N_8898,N_8771,N_8835);
xor U8899 (N_8899,N_8798,N_8721);
xor U8900 (N_8900,N_8780,N_8806);
xor U8901 (N_8901,N_8823,N_8775);
nor U8902 (N_8902,N_8745,N_8839);
or U8903 (N_8903,N_8842,N_8730);
nand U8904 (N_8904,N_8729,N_8814);
nand U8905 (N_8905,N_8845,N_8747);
xnor U8906 (N_8906,N_8803,N_8825);
nor U8907 (N_8907,N_8727,N_8819);
or U8908 (N_8908,N_8728,N_8722);
xnor U8909 (N_8909,N_8791,N_8759);
xor U8910 (N_8910,N_8755,N_8725);
nand U8911 (N_8911,N_8713,N_8795);
and U8912 (N_8912,N_8815,N_8779);
and U8913 (N_8913,N_8782,N_8752);
and U8914 (N_8914,N_8772,N_8736);
or U8915 (N_8915,N_8769,N_8794);
and U8916 (N_8916,N_8830,N_8714);
and U8917 (N_8917,N_8838,N_8848);
or U8918 (N_8918,N_8841,N_8805);
nand U8919 (N_8919,N_8773,N_8777);
nand U8920 (N_8920,N_8731,N_8849);
and U8921 (N_8921,N_8709,N_8786);
xnor U8922 (N_8922,N_8818,N_8826);
xnor U8923 (N_8923,N_8766,N_8844);
xor U8924 (N_8924,N_8788,N_8720);
nand U8925 (N_8925,N_8775,N_8733);
nand U8926 (N_8926,N_8753,N_8705);
nor U8927 (N_8927,N_8840,N_8755);
xor U8928 (N_8928,N_8783,N_8716);
and U8929 (N_8929,N_8732,N_8777);
and U8930 (N_8930,N_8823,N_8839);
nor U8931 (N_8931,N_8816,N_8702);
nor U8932 (N_8932,N_8833,N_8701);
xnor U8933 (N_8933,N_8775,N_8842);
nor U8934 (N_8934,N_8840,N_8805);
nor U8935 (N_8935,N_8714,N_8783);
and U8936 (N_8936,N_8728,N_8760);
nand U8937 (N_8937,N_8735,N_8817);
nand U8938 (N_8938,N_8823,N_8731);
nor U8939 (N_8939,N_8749,N_8778);
xnor U8940 (N_8940,N_8789,N_8732);
or U8941 (N_8941,N_8820,N_8759);
nor U8942 (N_8942,N_8833,N_8842);
nor U8943 (N_8943,N_8828,N_8753);
and U8944 (N_8944,N_8767,N_8807);
and U8945 (N_8945,N_8828,N_8780);
nand U8946 (N_8946,N_8828,N_8778);
or U8947 (N_8947,N_8828,N_8837);
and U8948 (N_8948,N_8770,N_8725);
nor U8949 (N_8949,N_8731,N_8818);
or U8950 (N_8950,N_8759,N_8708);
and U8951 (N_8951,N_8820,N_8812);
nor U8952 (N_8952,N_8730,N_8748);
nand U8953 (N_8953,N_8734,N_8837);
xnor U8954 (N_8954,N_8830,N_8752);
nor U8955 (N_8955,N_8837,N_8787);
or U8956 (N_8956,N_8798,N_8814);
and U8957 (N_8957,N_8818,N_8767);
and U8958 (N_8958,N_8839,N_8805);
and U8959 (N_8959,N_8777,N_8728);
nor U8960 (N_8960,N_8756,N_8728);
and U8961 (N_8961,N_8845,N_8728);
xnor U8962 (N_8962,N_8788,N_8819);
nand U8963 (N_8963,N_8792,N_8785);
or U8964 (N_8964,N_8733,N_8738);
nor U8965 (N_8965,N_8779,N_8823);
and U8966 (N_8966,N_8795,N_8803);
and U8967 (N_8967,N_8808,N_8756);
nor U8968 (N_8968,N_8784,N_8735);
xor U8969 (N_8969,N_8775,N_8758);
or U8970 (N_8970,N_8796,N_8813);
or U8971 (N_8971,N_8757,N_8734);
nand U8972 (N_8972,N_8805,N_8798);
or U8973 (N_8973,N_8739,N_8842);
xnor U8974 (N_8974,N_8831,N_8718);
xnor U8975 (N_8975,N_8791,N_8746);
nor U8976 (N_8976,N_8789,N_8773);
xor U8977 (N_8977,N_8822,N_8715);
nor U8978 (N_8978,N_8840,N_8712);
xnor U8979 (N_8979,N_8809,N_8762);
or U8980 (N_8980,N_8811,N_8812);
nor U8981 (N_8981,N_8799,N_8840);
xor U8982 (N_8982,N_8732,N_8797);
nand U8983 (N_8983,N_8737,N_8756);
and U8984 (N_8984,N_8827,N_8811);
and U8985 (N_8985,N_8764,N_8803);
xor U8986 (N_8986,N_8774,N_8835);
nor U8987 (N_8987,N_8737,N_8782);
nor U8988 (N_8988,N_8735,N_8800);
nor U8989 (N_8989,N_8784,N_8773);
or U8990 (N_8990,N_8723,N_8724);
nand U8991 (N_8991,N_8829,N_8749);
nor U8992 (N_8992,N_8731,N_8811);
or U8993 (N_8993,N_8765,N_8788);
and U8994 (N_8994,N_8750,N_8746);
or U8995 (N_8995,N_8831,N_8799);
nand U8996 (N_8996,N_8818,N_8795);
nand U8997 (N_8997,N_8838,N_8804);
and U8998 (N_8998,N_8817,N_8763);
and U8999 (N_8999,N_8799,N_8766);
xnor U9000 (N_9000,N_8853,N_8911);
nor U9001 (N_9001,N_8936,N_8869);
xor U9002 (N_9002,N_8897,N_8862);
nand U9003 (N_9003,N_8874,N_8992);
or U9004 (N_9004,N_8993,N_8888);
xnor U9005 (N_9005,N_8918,N_8925);
and U9006 (N_9006,N_8931,N_8904);
xnor U9007 (N_9007,N_8948,N_8863);
nand U9008 (N_9008,N_8946,N_8972);
xor U9009 (N_9009,N_8951,N_8937);
or U9010 (N_9010,N_8980,N_8908);
or U9011 (N_9011,N_8933,N_8958);
or U9012 (N_9012,N_8995,N_8916);
and U9013 (N_9013,N_8967,N_8921);
or U9014 (N_9014,N_8883,N_8989);
nand U9015 (N_9015,N_8867,N_8943);
nor U9016 (N_9016,N_8930,N_8978);
xnor U9017 (N_9017,N_8985,N_8945);
nor U9018 (N_9018,N_8969,N_8947);
or U9019 (N_9019,N_8968,N_8927);
or U9020 (N_9020,N_8857,N_8878);
or U9021 (N_9021,N_8966,N_8971);
and U9022 (N_9022,N_8917,N_8890);
xor U9023 (N_9023,N_8892,N_8942);
or U9024 (N_9024,N_8975,N_8919);
nand U9025 (N_9025,N_8962,N_8981);
nand U9026 (N_9026,N_8898,N_8987);
or U9027 (N_9027,N_8858,N_8870);
nor U9028 (N_9028,N_8938,N_8896);
nor U9029 (N_9029,N_8868,N_8952);
xor U9030 (N_9030,N_8889,N_8865);
nor U9031 (N_9031,N_8950,N_8965);
nor U9032 (N_9032,N_8997,N_8913);
nor U9033 (N_9033,N_8949,N_8875);
or U9034 (N_9034,N_8902,N_8986);
and U9035 (N_9035,N_8994,N_8998);
and U9036 (N_9036,N_8929,N_8923);
or U9037 (N_9037,N_8999,N_8909);
or U9038 (N_9038,N_8934,N_8852);
or U9039 (N_9039,N_8871,N_8982);
nand U9040 (N_9040,N_8940,N_8895);
nand U9041 (N_9041,N_8922,N_8939);
nor U9042 (N_9042,N_8899,N_8864);
nand U9043 (N_9043,N_8894,N_8963);
and U9044 (N_9044,N_8988,N_8944);
nand U9045 (N_9045,N_8906,N_8970);
nor U9046 (N_9046,N_8915,N_8920);
nor U9047 (N_9047,N_8880,N_8861);
nand U9048 (N_9048,N_8910,N_8854);
xor U9049 (N_9049,N_8905,N_8856);
or U9050 (N_9050,N_8964,N_8996);
xor U9051 (N_9051,N_8876,N_8957);
nand U9052 (N_9052,N_8907,N_8961);
or U9053 (N_9053,N_8873,N_8954);
or U9054 (N_9054,N_8860,N_8991);
xor U9055 (N_9055,N_8872,N_8900);
nand U9056 (N_9056,N_8983,N_8941);
and U9057 (N_9057,N_8974,N_8886);
or U9058 (N_9058,N_8851,N_8914);
nor U9059 (N_9059,N_8879,N_8887);
xor U9060 (N_9060,N_8893,N_8932);
or U9061 (N_9061,N_8990,N_8912);
xnor U9062 (N_9062,N_8855,N_8960);
or U9063 (N_9063,N_8928,N_8901);
and U9064 (N_9064,N_8953,N_8973);
and U9065 (N_9065,N_8955,N_8956);
nand U9066 (N_9066,N_8926,N_8903);
nor U9067 (N_9067,N_8977,N_8959);
and U9068 (N_9068,N_8976,N_8850);
nand U9069 (N_9069,N_8859,N_8866);
nor U9070 (N_9070,N_8924,N_8881);
nand U9071 (N_9071,N_8877,N_8935);
nor U9072 (N_9072,N_8979,N_8885);
and U9073 (N_9073,N_8882,N_8984);
nor U9074 (N_9074,N_8891,N_8884);
xnor U9075 (N_9075,N_8859,N_8875);
nand U9076 (N_9076,N_8877,N_8851);
or U9077 (N_9077,N_8859,N_8955);
or U9078 (N_9078,N_8959,N_8919);
nor U9079 (N_9079,N_8972,N_8906);
xnor U9080 (N_9080,N_8983,N_8981);
nor U9081 (N_9081,N_8899,N_8892);
nand U9082 (N_9082,N_8857,N_8946);
or U9083 (N_9083,N_8969,N_8906);
nand U9084 (N_9084,N_8893,N_8870);
nand U9085 (N_9085,N_8915,N_8997);
and U9086 (N_9086,N_8992,N_8927);
or U9087 (N_9087,N_8981,N_8912);
nand U9088 (N_9088,N_8932,N_8925);
xnor U9089 (N_9089,N_8898,N_8951);
or U9090 (N_9090,N_8930,N_8982);
nand U9091 (N_9091,N_8984,N_8919);
nor U9092 (N_9092,N_8902,N_8959);
nor U9093 (N_9093,N_8972,N_8930);
and U9094 (N_9094,N_8951,N_8917);
nor U9095 (N_9095,N_8984,N_8955);
nand U9096 (N_9096,N_8918,N_8877);
xnor U9097 (N_9097,N_8998,N_8905);
and U9098 (N_9098,N_8884,N_8979);
nand U9099 (N_9099,N_8859,N_8998);
and U9100 (N_9100,N_8995,N_8863);
nor U9101 (N_9101,N_8855,N_8922);
xor U9102 (N_9102,N_8965,N_8986);
or U9103 (N_9103,N_8874,N_8872);
xor U9104 (N_9104,N_8885,N_8960);
or U9105 (N_9105,N_8945,N_8865);
xor U9106 (N_9106,N_8924,N_8853);
nor U9107 (N_9107,N_8859,N_8991);
nor U9108 (N_9108,N_8946,N_8886);
nand U9109 (N_9109,N_8993,N_8936);
or U9110 (N_9110,N_8985,N_8976);
or U9111 (N_9111,N_8968,N_8856);
and U9112 (N_9112,N_8927,N_8886);
nor U9113 (N_9113,N_8868,N_8959);
and U9114 (N_9114,N_8881,N_8932);
or U9115 (N_9115,N_8995,N_8991);
nand U9116 (N_9116,N_8898,N_8879);
nand U9117 (N_9117,N_8859,N_8905);
and U9118 (N_9118,N_8988,N_8935);
nor U9119 (N_9119,N_8914,N_8925);
and U9120 (N_9120,N_8863,N_8902);
or U9121 (N_9121,N_8969,N_8996);
nand U9122 (N_9122,N_8905,N_8855);
nor U9123 (N_9123,N_8940,N_8865);
nor U9124 (N_9124,N_8970,N_8936);
xnor U9125 (N_9125,N_8911,N_8964);
or U9126 (N_9126,N_8949,N_8922);
nor U9127 (N_9127,N_8879,N_8942);
nor U9128 (N_9128,N_8992,N_8938);
nand U9129 (N_9129,N_8965,N_8977);
nor U9130 (N_9130,N_8950,N_8879);
nand U9131 (N_9131,N_8960,N_8952);
or U9132 (N_9132,N_8909,N_8955);
nor U9133 (N_9133,N_8952,N_8895);
nor U9134 (N_9134,N_8896,N_8996);
and U9135 (N_9135,N_8943,N_8936);
or U9136 (N_9136,N_8933,N_8962);
xnor U9137 (N_9137,N_8948,N_8851);
xnor U9138 (N_9138,N_8858,N_8885);
nor U9139 (N_9139,N_8949,N_8899);
nor U9140 (N_9140,N_8927,N_8947);
nor U9141 (N_9141,N_8901,N_8906);
and U9142 (N_9142,N_8868,N_8940);
nor U9143 (N_9143,N_8899,N_8919);
nor U9144 (N_9144,N_8941,N_8863);
xnor U9145 (N_9145,N_8856,N_8999);
nand U9146 (N_9146,N_8899,N_8875);
or U9147 (N_9147,N_8976,N_8981);
nor U9148 (N_9148,N_8950,N_8880);
and U9149 (N_9149,N_8925,N_8967);
and U9150 (N_9150,N_9094,N_9060);
or U9151 (N_9151,N_9118,N_9048);
xnor U9152 (N_9152,N_9076,N_9037);
and U9153 (N_9153,N_9080,N_9050);
or U9154 (N_9154,N_9003,N_9126);
nand U9155 (N_9155,N_9063,N_9082);
xor U9156 (N_9156,N_9128,N_9091);
xor U9157 (N_9157,N_9135,N_9131);
nand U9158 (N_9158,N_9001,N_9140);
nand U9159 (N_9159,N_9083,N_9054);
nand U9160 (N_9160,N_9115,N_9088);
nand U9161 (N_9161,N_9109,N_9134);
nor U9162 (N_9162,N_9071,N_9033);
xor U9163 (N_9163,N_9043,N_9129);
xor U9164 (N_9164,N_9046,N_9078);
or U9165 (N_9165,N_9018,N_9072);
or U9166 (N_9166,N_9102,N_9123);
nor U9167 (N_9167,N_9004,N_9002);
or U9168 (N_9168,N_9007,N_9005);
nand U9169 (N_9169,N_9064,N_9111);
or U9170 (N_9170,N_9144,N_9055);
nand U9171 (N_9171,N_9119,N_9014);
and U9172 (N_9172,N_9039,N_9034);
and U9173 (N_9173,N_9085,N_9139);
or U9174 (N_9174,N_9106,N_9056);
and U9175 (N_9175,N_9010,N_9125);
nand U9176 (N_9176,N_9017,N_9022);
xnor U9177 (N_9177,N_9121,N_9124);
nor U9178 (N_9178,N_9012,N_9027);
and U9179 (N_9179,N_9141,N_9073);
nand U9180 (N_9180,N_9104,N_9137);
or U9181 (N_9181,N_9113,N_9036);
nor U9182 (N_9182,N_9000,N_9024);
nor U9183 (N_9183,N_9103,N_9026);
or U9184 (N_9184,N_9074,N_9108);
and U9185 (N_9185,N_9136,N_9040);
nand U9186 (N_9186,N_9011,N_9021);
or U9187 (N_9187,N_9122,N_9120);
or U9188 (N_9188,N_9016,N_9093);
and U9189 (N_9189,N_9029,N_9051);
nor U9190 (N_9190,N_9112,N_9077);
xor U9191 (N_9191,N_9032,N_9075);
nand U9192 (N_9192,N_9035,N_9068);
and U9193 (N_9193,N_9028,N_9052);
or U9194 (N_9194,N_9110,N_9096);
nand U9195 (N_9195,N_9066,N_9081);
xnor U9196 (N_9196,N_9042,N_9101);
and U9197 (N_9197,N_9138,N_9053);
and U9198 (N_9198,N_9009,N_9069);
xor U9199 (N_9199,N_9067,N_9130);
or U9200 (N_9200,N_9019,N_9105);
xor U9201 (N_9201,N_9058,N_9147);
or U9202 (N_9202,N_9107,N_9038);
xor U9203 (N_9203,N_9062,N_9097);
nor U9204 (N_9204,N_9057,N_9133);
xor U9205 (N_9205,N_9116,N_9070);
and U9206 (N_9206,N_9099,N_9020);
or U9207 (N_9207,N_9030,N_9098);
nor U9208 (N_9208,N_9008,N_9145);
xnor U9209 (N_9209,N_9095,N_9006);
nand U9210 (N_9210,N_9059,N_9065);
and U9211 (N_9211,N_9092,N_9047);
nor U9212 (N_9212,N_9087,N_9114);
and U9213 (N_9213,N_9132,N_9013);
or U9214 (N_9214,N_9031,N_9090);
or U9215 (N_9215,N_9045,N_9041);
or U9216 (N_9216,N_9117,N_9084);
or U9217 (N_9217,N_9100,N_9061);
nor U9218 (N_9218,N_9015,N_9127);
nand U9219 (N_9219,N_9049,N_9142);
nand U9220 (N_9220,N_9044,N_9148);
and U9221 (N_9221,N_9089,N_9025);
xnor U9222 (N_9222,N_9143,N_9086);
or U9223 (N_9223,N_9079,N_9149);
nor U9224 (N_9224,N_9023,N_9146);
nand U9225 (N_9225,N_9148,N_9119);
xnor U9226 (N_9226,N_9006,N_9126);
xor U9227 (N_9227,N_9130,N_9035);
and U9228 (N_9228,N_9109,N_9078);
or U9229 (N_9229,N_9073,N_9054);
or U9230 (N_9230,N_9037,N_9144);
xnor U9231 (N_9231,N_9010,N_9036);
or U9232 (N_9232,N_9050,N_9110);
nand U9233 (N_9233,N_9114,N_9105);
nor U9234 (N_9234,N_9033,N_9005);
or U9235 (N_9235,N_9053,N_9020);
or U9236 (N_9236,N_9048,N_9094);
nand U9237 (N_9237,N_9070,N_9138);
nor U9238 (N_9238,N_9121,N_9014);
or U9239 (N_9239,N_9055,N_9082);
or U9240 (N_9240,N_9034,N_9059);
and U9241 (N_9241,N_9089,N_9124);
and U9242 (N_9242,N_9035,N_9143);
or U9243 (N_9243,N_9021,N_9106);
and U9244 (N_9244,N_9038,N_9138);
nand U9245 (N_9245,N_9074,N_9130);
nand U9246 (N_9246,N_9127,N_9134);
xor U9247 (N_9247,N_9049,N_9118);
xnor U9248 (N_9248,N_9024,N_9014);
nand U9249 (N_9249,N_9114,N_9028);
nand U9250 (N_9250,N_9143,N_9126);
xnor U9251 (N_9251,N_9098,N_9081);
nor U9252 (N_9252,N_9023,N_9098);
or U9253 (N_9253,N_9125,N_9002);
nor U9254 (N_9254,N_9100,N_9092);
and U9255 (N_9255,N_9137,N_9126);
xor U9256 (N_9256,N_9034,N_9064);
xnor U9257 (N_9257,N_9051,N_9090);
and U9258 (N_9258,N_9144,N_9019);
nand U9259 (N_9259,N_9083,N_9070);
nand U9260 (N_9260,N_9132,N_9121);
nor U9261 (N_9261,N_9000,N_9130);
nand U9262 (N_9262,N_9102,N_9040);
or U9263 (N_9263,N_9149,N_9092);
nor U9264 (N_9264,N_9141,N_9097);
or U9265 (N_9265,N_9044,N_9074);
and U9266 (N_9266,N_9069,N_9128);
xnor U9267 (N_9267,N_9049,N_9093);
or U9268 (N_9268,N_9093,N_9067);
nand U9269 (N_9269,N_9068,N_9124);
xor U9270 (N_9270,N_9051,N_9019);
or U9271 (N_9271,N_9104,N_9073);
nor U9272 (N_9272,N_9136,N_9147);
nand U9273 (N_9273,N_9054,N_9114);
or U9274 (N_9274,N_9003,N_9143);
xor U9275 (N_9275,N_9139,N_9147);
xnor U9276 (N_9276,N_9059,N_9085);
and U9277 (N_9277,N_9084,N_9120);
nor U9278 (N_9278,N_9128,N_9120);
or U9279 (N_9279,N_9047,N_9079);
or U9280 (N_9280,N_9073,N_9143);
nor U9281 (N_9281,N_9031,N_9143);
nor U9282 (N_9282,N_9125,N_9036);
or U9283 (N_9283,N_9096,N_9008);
nand U9284 (N_9284,N_9149,N_9048);
and U9285 (N_9285,N_9004,N_9053);
nand U9286 (N_9286,N_9030,N_9034);
nor U9287 (N_9287,N_9014,N_9000);
nor U9288 (N_9288,N_9021,N_9120);
xnor U9289 (N_9289,N_9006,N_9125);
and U9290 (N_9290,N_9027,N_9128);
and U9291 (N_9291,N_9048,N_9084);
nor U9292 (N_9292,N_9008,N_9022);
nor U9293 (N_9293,N_9026,N_9015);
nor U9294 (N_9294,N_9019,N_9049);
and U9295 (N_9295,N_9143,N_9142);
and U9296 (N_9296,N_9090,N_9079);
and U9297 (N_9297,N_9030,N_9084);
or U9298 (N_9298,N_9096,N_9050);
nand U9299 (N_9299,N_9082,N_9127);
and U9300 (N_9300,N_9255,N_9264);
and U9301 (N_9301,N_9180,N_9279);
nand U9302 (N_9302,N_9245,N_9265);
nor U9303 (N_9303,N_9184,N_9178);
and U9304 (N_9304,N_9167,N_9215);
and U9305 (N_9305,N_9291,N_9155);
or U9306 (N_9306,N_9203,N_9223);
xnor U9307 (N_9307,N_9290,N_9213);
nand U9308 (N_9308,N_9277,N_9270);
or U9309 (N_9309,N_9217,N_9278);
xor U9310 (N_9310,N_9182,N_9285);
xor U9311 (N_9311,N_9162,N_9282);
nor U9312 (N_9312,N_9229,N_9170);
nand U9313 (N_9313,N_9226,N_9189);
xnor U9314 (N_9314,N_9160,N_9153);
and U9315 (N_9315,N_9274,N_9201);
xnor U9316 (N_9316,N_9241,N_9159);
and U9317 (N_9317,N_9262,N_9283);
or U9318 (N_9318,N_9251,N_9200);
nand U9319 (N_9319,N_9267,N_9295);
nor U9320 (N_9320,N_9192,N_9284);
nor U9321 (N_9321,N_9219,N_9176);
nand U9322 (N_9322,N_9294,N_9296);
nor U9323 (N_9323,N_9227,N_9280);
nand U9324 (N_9324,N_9190,N_9173);
xor U9325 (N_9325,N_9187,N_9286);
nor U9326 (N_9326,N_9234,N_9156);
nand U9327 (N_9327,N_9263,N_9287);
and U9328 (N_9328,N_9150,N_9161);
or U9329 (N_9329,N_9289,N_9194);
or U9330 (N_9330,N_9211,N_9233);
nor U9331 (N_9331,N_9236,N_9166);
xnor U9332 (N_9332,N_9158,N_9185);
or U9333 (N_9333,N_9232,N_9240);
or U9334 (N_9334,N_9222,N_9253);
nor U9335 (N_9335,N_9181,N_9216);
or U9336 (N_9336,N_9244,N_9206);
xor U9337 (N_9337,N_9183,N_9258);
and U9338 (N_9338,N_9247,N_9250);
or U9339 (N_9339,N_9218,N_9193);
or U9340 (N_9340,N_9157,N_9179);
and U9341 (N_9341,N_9174,N_9202);
nand U9342 (N_9342,N_9273,N_9186);
and U9343 (N_9343,N_9220,N_9242);
nand U9344 (N_9344,N_9249,N_9259);
or U9345 (N_9345,N_9172,N_9195);
and U9346 (N_9346,N_9297,N_9152);
xor U9347 (N_9347,N_9171,N_9246);
or U9348 (N_9348,N_9210,N_9238);
xnor U9349 (N_9349,N_9230,N_9235);
nand U9350 (N_9350,N_9256,N_9243);
xor U9351 (N_9351,N_9224,N_9299);
nor U9352 (N_9352,N_9168,N_9151);
and U9353 (N_9353,N_9288,N_9239);
xnor U9354 (N_9354,N_9272,N_9221);
or U9355 (N_9355,N_9298,N_9204);
nand U9356 (N_9356,N_9254,N_9197);
or U9357 (N_9357,N_9163,N_9252);
and U9358 (N_9358,N_9268,N_9209);
nand U9359 (N_9359,N_9281,N_9196);
or U9360 (N_9360,N_9165,N_9293);
or U9361 (N_9361,N_9257,N_9271);
or U9362 (N_9362,N_9261,N_9225);
xnor U9363 (N_9363,N_9177,N_9208);
nand U9364 (N_9364,N_9228,N_9275);
or U9365 (N_9365,N_9231,N_9266);
xnor U9366 (N_9366,N_9205,N_9212);
and U9367 (N_9367,N_9169,N_9269);
or U9368 (N_9368,N_9199,N_9248);
or U9369 (N_9369,N_9175,N_9276);
or U9370 (N_9370,N_9260,N_9191);
xnor U9371 (N_9371,N_9207,N_9198);
nand U9372 (N_9372,N_9154,N_9214);
or U9373 (N_9373,N_9292,N_9237);
and U9374 (N_9374,N_9188,N_9164);
nor U9375 (N_9375,N_9194,N_9215);
nor U9376 (N_9376,N_9173,N_9159);
nor U9377 (N_9377,N_9187,N_9252);
or U9378 (N_9378,N_9220,N_9229);
or U9379 (N_9379,N_9154,N_9249);
or U9380 (N_9380,N_9164,N_9201);
and U9381 (N_9381,N_9299,N_9150);
nand U9382 (N_9382,N_9292,N_9179);
and U9383 (N_9383,N_9197,N_9268);
and U9384 (N_9384,N_9277,N_9210);
nand U9385 (N_9385,N_9261,N_9151);
nor U9386 (N_9386,N_9274,N_9222);
or U9387 (N_9387,N_9254,N_9190);
xnor U9388 (N_9388,N_9258,N_9151);
nor U9389 (N_9389,N_9199,N_9193);
xnor U9390 (N_9390,N_9212,N_9221);
xor U9391 (N_9391,N_9228,N_9234);
nor U9392 (N_9392,N_9272,N_9248);
nand U9393 (N_9393,N_9274,N_9266);
nor U9394 (N_9394,N_9279,N_9201);
and U9395 (N_9395,N_9290,N_9237);
nand U9396 (N_9396,N_9195,N_9270);
or U9397 (N_9397,N_9292,N_9164);
and U9398 (N_9398,N_9181,N_9199);
and U9399 (N_9399,N_9264,N_9217);
nor U9400 (N_9400,N_9213,N_9187);
and U9401 (N_9401,N_9294,N_9226);
nand U9402 (N_9402,N_9259,N_9212);
nor U9403 (N_9403,N_9199,N_9240);
or U9404 (N_9404,N_9293,N_9151);
xnor U9405 (N_9405,N_9167,N_9216);
or U9406 (N_9406,N_9157,N_9229);
nor U9407 (N_9407,N_9176,N_9205);
xnor U9408 (N_9408,N_9285,N_9283);
nor U9409 (N_9409,N_9267,N_9233);
nor U9410 (N_9410,N_9197,N_9252);
nor U9411 (N_9411,N_9219,N_9252);
or U9412 (N_9412,N_9184,N_9190);
or U9413 (N_9413,N_9251,N_9159);
nor U9414 (N_9414,N_9256,N_9197);
xor U9415 (N_9415,N_9213,N_9263);
nor U9416 (N_9416,N_9225,N_9168);
and U9417 (N_9417,N_9214,N_9188);
nor U9418 (N_9418,N_9289,N_9250);
nor U9419 (N_9419,N_9217,N_9166);
and U9420 (N_9420,N_9221,N_9173);
nand U9421 (N_9421,N_9242,N_9244);
nor U9422 (N_9422,N_9277,N_9227);
nor U9423 (N_9423,N_9176,N_9183);
nor U9424 (N_9424,N_9153,N_9217);
and U9425 (N_9425,N_9206,N_9258);
or U9426 (N_9426,N_9174,N_9161);
nand U9427 (N_9427,N_9257,N_9261);
and U9428 (N_9428,N_9277,N_9175);
nor U9429 (N_9429,N_9263,N_9246);
xnor U9430 (N_9430,N_9235,N_9259);
xnor U9431 (N_9431,N_9246,N_9288);
nand U9432 (N_9432,N_9268,N_9156);
or U9433 (N_9433,N_9184,N_9162);
or U9434 (N_9434,N_9242,N_9228);
nor U9435 (N_9435,N_9189,N_9271);
nor U9436 (N_9436,N_9192,N_9201);
and U9437 (N_9437,N_9299,N_9242);
nor U9438 (N_9438,N_9176,N_9238);
nor U9439 (N_9439,N_9220,N_9180);
and U9440 (N_9440,N_9268,N_9159);
or U9441 (N_9441,N_9240,N_9287);
xnor U9442 (N_9442,N_9248,N_9162);
nand U9443 (N_9443,N_9156,N_9208);
or U9444 (N_9444,N_9220,N_9198);
nand U9445 (N_9445,N_9284,N_9262);
nand U9446 (N_9446,N_9265,N_9274);
nand U9447 (N_9447,N_9246,N_9293);
nand U9448 (N_9448,N_9206,N_9186);
and U9449 (N_9449,N_9210,N_9269);
and U9450 (N_9450,N_9311,N_9416);
and U9451 (N_9451,N_9413,N_9309);
nand U9452 (N_9452,N_9382,N_9369);
nor U9453 (N_9453,N_9390,N_9410);
nand U9454 (N_9454,N_9415,N_9327);
nor U9455 (N_9455,N_9337,N_9372);
or U9456 (N_9456,N_9300,N_9322);
or U9457 (N_9457,N_9374,N_9354);
xnor U9458 (N_9458,N_9446,N_9345);
or U9459 (N_9459,N_9329,N_9396);
xor U9460 (N_9460,N_9306,N_9417);
nand U9461 (N_9461,N_9428,N_9394);
xnor U9462 (N_9462,N_9328,N_9380);
xnor U9463 (N_9463,N_9378,N_9356);
nand U9464 (N_9464,N_9365,N_9397);
nand U9465 (N_9465,N_9408,N_9422);
or U9466 (N_9466,N_9319,N_9436);
or U9467 (N_9467,N_9331,N_9404);
and U9468 (N_9468,N_9373,N_9320);
nand U9469 (N_9469,N_9425,N_9370);
nand U9470 (N_9470,N_9400,N_9430);
and U9471 (N_9471,N_9305,N_9350);
or U9472 (N_9472,N_9437,N_9363);
xnor U9473 (N_9473,N_9401,N_9387);
nand U9474 (N_9474,N_9351,N_9332);
xnor U9475 (N_9475,N_9395,N_9432);
nand U9476 (N_9476,N_9448,N_9323);
nor U9477 (N_9477,N_9355,N_9386);
or U9478 (N_9478,N_9317,N_9335);
and U9479 (N_9479,N_9358,N_9407);
or U9480 (N_9480,N_9409,N_9301);
xnor U9481 (N_9481,N_9418,N_9344);
and U9482 (N_9482,N_9375,N_9393);
and U9483 (N_9483,N_9315,N_9403);
nand U9484 (N_9484,N_9352,N_9441);
nor U9485 (N_9485,N_9307,N_9316);
nor U9486 (N_9486,N_9312,N_9349);
nand U9487 (N_9487,N_9427,N_9357);
nand U9488 (N_9488,N_9444,N_9353);
xnor U9489 (N_9489,N_9445,N_9381);
or U9490 (N_9490,N_9421,N_9367);
or U9491 (N_9491,N_9442,N_9389);
xnor U9492 (N_9492,N_9334,N_9359);
or U9493 (N_9493,N_9330,N_9377);
and U9494 (N_9494,N_9399,N_9429);
and U9495 (N_9495,N_9426,N_9412);
or U9496 (N_9496,N_9440,N_9447);
and U9497 (N_9497,N_9325,N_9385);
nor U9498 (N_9498,N_9434,N_9342);
or U9499 (N_9499,N_9392,N_9423);
nand U9500 (N_9500,N_9414,N_9420);
xor U9501 (N_9501,N_9398,N_9366);
or U9502 (N_9502,N_9435,N_9361);
nor U9503 (N_9503,N_9364,N_9303);
nand U9504 (N_9504,N_9371,N_9348);
or U9505 (N_9505,N_9368,N_9324);
and U9506 (N_9506,N_9449,N_9439);
and U9507 (N_9507,N_9424,N_9419);
or U9508 (N_9508,N_9321,N_9443);
or U9509 (N_9509,N_9341,N_9379);
and U9510 (N_9510,N_9346,N_9402);
xnor U9511 (N_9511,N_9406,N_9383);
nand U9512 (N_9512,N_9339,N_9433);
and U9513 (N_9513,N_9340,N_9302);
nand U9514 (N_9514,N_9338,N_9308);
nor U9515 (N_9515,N_9310,N_9343);
or U9516 (N_9516,N_9336,N_9360);
nand U9517 (N_9517,N_9362,N_9314);
nor U9518 (N_9518,N_9313,N_9391);
and U9519 (N_9519,N_9438,N_9347);
nor U9520 (N_9520,N_9411,N_9388);
nor U9521 (N_9521,N_9384,N_9376);
nand U9522 (N_9522,N_9326,N_9318);
nand U9523 (N_9523,N_9405,N_9431);
and U9524 (N_9524,N_9333,N_9304);
nand U9525 (N_9525,N_9340,N_9312);
and U9526 (N_9526,N_9400,N_9412);
nand U9527 (N_9527,N_9448,N_9400);
xor U9528 (N_9528,N_9334,N_9430);
or U9529 (N_9529,N_9319,N_9361);
nand U9530 (N_9530,N_9384,N_9345);
nor U9531 (N_9531,N_9310,N_9387);
nor U9532 (N_9532,N_9414,N_9394);
and U9533 (N_9533,N_9424,N_9410);
nand U9534 (N_9534,N_9445,N_9354);
nand U9535 (N_9535,N_9316,N_9339);
nand U9536 (N_9536,N_9404,N_9419);
nand U9537 (N_9537,N_9426,N_9402);
nand U9538 (N_9538,N_9392,N_9399);
xnor U9539 (N_9539,N_9307,N_9362);
nor U9540 (N_9540,N_9371,N_9333);
and U9541 (N_9541,N_9388,N_9395);
nor U9542 (N_9542,N_9333,N_9375);
xnor U9543 (N_9543,N_9398,N_9309);
nor U9544 (N_9544,N_9425,N_9376);
xor U9545 (N_9545,N_9422,N_9376);
nor U9546 (N_9546,N_9439,N_9333);
nor U9547 (N_9547,N_9310,N_9319);
nand U9548 (N_9548,N_9380,N_9403);
xnor U9549 (N_9549,N_9431,N_9331);
nand U9550 (N_9550,N_9335,N_9411);
and U9551 (N_9551,N_9423,N_9313);
and U9552 (N_9552,N_9319,N_9399);
and U9553 (N_9553,N_9396,N_9431);
nor U9554 (N_9554,N_9438,N_9341);
and U9555 (N_9555,N_9400,N_9348);
nor U9556 (N_9556,N_9345,N_9448);
xnor U9557 (N_9557,N_9443,N_9318);
nand U9558 (N_9558,N_9338,N_9365);
or U9559 (N_9559,N_9346,N_9376);
or U9560 (N_9560,N_9417,N_9320);
nand U9561 (N_9561,N_9341,N_9371);
nand U9562 (N_9562,N_9398,N_9399);
and U9563 (N_9563,N_9426,N_9392);
and U9564 (N_9564,N_9370,N_9405);
nand U9565 (N_9565,N_9410,N_9341);
and U9566 (N_9566,N_9363,N_9409);
xor U9567 (N_9567,N_9373,N_9389);
or U9568 (N_9568,N_9405,N_9379);
nor U9569 (N_9569,N_9312,N_9348);
nor U9570 (N_9570,N_9405,N_9320);
or U9571 (N_9571,N_9385,N_9434);
xor U9572 (N_9572,N_9379,N_9443);
nand U9573 (N_9573,N_9348,N_9406);
nor U9574 (N_9574,N_9343,N_9389);
nor U9575 (N_9575,N_9434,N_9396);
xnor U9576 (N_9576,N_9328,N_9352);
nand U9577 (N_9577,N_9353,N_9437);
nand U9578 (N_9578,N_9403,N_9360);
nand U9579 (N_9579,N_9324,N_9379);
nand U9580 (N_9580,N_9383,N_9309);
nor U9581 (N_9581,N_9357,N_9337);
nor U9582 (N_9582,N_9344,N_9422);
and U9583 (N_9583,N_9419,N_9374);
and U9584 (N_9584,N_9366,N_9410);
nor U9585 (N_9585,N_9414,N_9407);
nand U9586 (N_9586,N_9432,N_9422);
and U9587 (N_9587,N_9392,N_9362);
and U9588 (N_9588,N_9406,N_9332);
nand U9589 (N_9589,N_9427,N_9382);
xnor U9590 (N_9590,N_9441,N_9367);
xnor U9591 (N_9591,N_9325,N_9429);
and U9592 (N_9592,N_9338,N_9301);
or U9593 (N_9593,N_9309,N_9340);
nand U9594 (N_9594,N_9440,N_9352);
and U9595 (N_9595,N_9410,N_9312);
xnor U9596 (N_9596,N_9349,N_9301);
or U9597 (N_9597,N_9380,N_9417);
xor U9598 (N_9598,N_9301,N_9336);
and U9599 (N_9599,N_9300,N_9372);
or U9600 (N_9600,N_9517,N_9568);
or U9601 (N_9601,N_9550,N_9532);
and U9602 (N_9602,N_9530,N_9475);
xnor U9603 (N_9603,N_9597,N_9471);
or U9604 (N_9604,N_9587,N_9505);
xnor U9605 (N_9605,N_9519,N_9548);
xnor U9606 (N_9606,N_9545,N_9466);
nand U9607 (N_9607,N_9483,N_9467);
nand U9608 (N_9608,N_9491,N_9584);
xor U9609 (N_9609,N_9513,N_9539);
nor U9610 (N_9610,N_9509,N_9525);
nor U9611 (N_9611,N_9486,N_9575);
nor U9612 (N_9612,N_9591,N_9592);
nor U9613 (N_9613,N_9463,N_9520);
nand U9614 (N_9614,N_9533,N_9534);
nor U9615 (N_9615,N_9543,N_9456);
nand U9616 (N_9616,N_9565,N_9537);
nor U9617 (N_9617,N_9468,N_9572);
nor U9618 (N_9618,N_9457,N_9502);
or U9619 (N_9619,N_9510,N_9454);
nor U9620 (N_9620,N_9485,N_9526);
xor U9621 (N_9621,N_9585,N_9582);
nor U9622 (N_9622,N_9474,N_9559);
nor U9623 (N_9623,N_9590,N_9498);
or U9624 (N_9624,N_9594,N_9561);
or U9625 (N_9625,N_9544,N_9560);
nor U9626 (N_9626,N_9451,N_9493);
or U9627 (N_9627,N_9599,N_9556);
nand U9628 (N_9628,N_9479,N_9464);
xnor U9629 (N_9629,N_9484,N_9518);
nand U9630 (N_9630,N_9508,N_9573);
and U9631 (N_9631,N_9527,N_9583);
or U9632 (N_9632,N_9566,N_9492);
nand U9633 (N_9633,N_9487,N_9542);
and U9634 (N_9634,N_9558,N_9563);
and U9635 (N_9635,N_9529,N_9453);
xnor U9636 (N_9636,N_9586,N_9528);
and U9637 (N_9637,N_9553,N_9535);
xor U9638 (N_9638,N_9450,N_9452);
xnor U9639 (N_9639,N_9465,N_9579);
nor U9640 (N_9640,N_9596,N_9554);
and U9641 (N_9641,N_9576,N_9562);
nand U9642 (N_9642,N_9469,N_9551);
nor U9643 (N_9643,N_9460,N_9462);
nor U9644 (N_9644,N_9488,N_9495);
and U9645 (N_9645,N_9477,N_9459);
nand U9646 (N_9646,N_9557,N_9473);
or U9647 (N_9647,N_9489,N_9580);
nor U9648 (N_9648,N_9514,N_9541);
or U9649 (N_9649,N_9564,N_9507);
nor U9650 (N_9650,N_9536,N_9490);
nor U9651 (N_9651,N_9555,N_9506);
nand U9652 (N_9652,N_9540,N_9516);
or U9653 (N_9653,N_9588,N_9458);
nand U9654 (N_9654,N_9515,N_9503);
nor U9655 (N_9655,N_9598,N_9511);
and U9656 (N_9656,N_9523,N_9470);
and U9657 (N_9657,N_9497,N_9499);
and U9658 (N_9658,N_9593,N_9481);
xor U9659 (N_9659,N_9549,N_9478);
or U9660 (N_9660,N_9570,N_9504);
and U9661 (N_9661,N_9531,N_9480);
xor U9662 (N_9662,N_9496,N_9574);
nand U9663 (N_9663,N_9482,N_9546);
nand U9664 (N_9664,N_9455,N_9577);
or U9665 (N_9665,N_9567,N_9547);
xnor U9666 (N_9666,N_9501,N_9571);
and U9667 (N_9667,N_9521,N_9578);
xor U9668 (N_9668,N_9500,N_9512);
or U9669 (N_9669,N_9524,N_9522);
nand U9670 (N_9670,N_9589,N_9552);
nor U9671 (N_9671,N_9472,N_9476);
xnor U9672 (N_9672,N_9569,N_9595);
nand U9673 (N_9673,N_9494,N_9461);
or U9674 (N_9674,N_9581,N_9538);
xnor U9675 (N_9675,N_9468,N_9537);
xor U9676 (N_9676,N_9510,N_9585);
and U9677 (N_9677,N_9543,N_9574);
or U9678 (N_9678,N_9482,N_9572);
nand U9679 (N_9679,N_9529,N_9565);
or U9680 (N_9680,N_9534,N_9530);
nor U9681 (N_9681,N_9469,N_9495);
or U9682 (N_9682,N_9587,N_9548);
nor U9683 (N_9683,N_9585,N_9453);
xnor U9684 (N_9684,N_9593,N_9485);
or U9685 (N_9685,N_9481,N_9517);
and U9686 (N_9686,N_9593,N_9544);
nor U9687 (N_9687,N_9452,N_9490);
nand U9688 (N_9688,N_9574,N_9478);
nor U9689 (N_9689,N_9500,N_9572);
or U9690 (N_9690,N_9548,N_9540);
nand U9691 (N_9691,N_9508,N_9521);
and U9692 (N_9692,N_9522,N_9532);
or U9693 (N_9693,N_9541,N_9469);
xnor U9694 (N_9694,N_9563,N_9480);
or U9695 (N_9695,N_9493,N_9542);
xor U9696 (N_9696,N_9475,N_9456);
nand U9697 (N_9697,N_9552,N_9475);
or U9698 (N_9698,N_9454,N_9549);
or U9699 (N_9699,N_9495,N_9517);
nor U9700 (N_9700,N_9566,N_9595);
or U9701 (N_9701,N_9475,N_9452);
or U9702 (N_9702,N_9591,N_9470);
and U9703 (N_9703,N_9570,N_9533);
or U9704 (N_9704,N_9473,N_9502);
or U9705 (N_9705,N_9529,N_9479);
xor U9706 (N_9706,N_9477,N_9508);
or U9707 (N_9707,N_9450,N_9575);
nand U9708 (N_9708,N_9455,N_9459);
nand U9709 (N_9709,N_9598,N_9553);
or U9710 (N_9710,N_9544,N_9570);
xnor U9711 (N_9711,N_9546,N_9591);
nor U9712 (N_9712,N_9454,N_9557);
or U9713 (N_9713,N_9458,N_9511);
or U9714 (N_9714,N_9486,N_9515);
and U9715 (N_9715,N_9454,N_9498);
and U9716 (N_9716,N_9575,N_9504);
nor U9717 (N_9717,N_9514,N_9512);
xnor U9718 (N_9718,N_9545,N_9548);
xnor U9719 (N_9719,N_9575,N_9532);
or U9720 (N_9720,N_9523,N_9484);
or U9721 (N_9721,N_9484,N_9590);
xnor U9722 (N_9722,N_9496,N_9462);
nand U9723 (N_9723,N_9542,N_9464);
nand U9724 (N_9724,N_9566,N_9527);
nor U9725 (N_9725,N_9464,N_9546);
nand U9726 (N_9726,N_9479,N_9506);
or U9727 (N_9727,N_9498,N_9596);
and U9728 (N_9728,N_9473,N_9567);
and U9729 (N_9729,N_9456,N_9532);
xnor U9730 (N_9730,N_9568,N_9557);
nor U9731 (N_9731,N_9490,N_9470);
or U9732 (N_9732,N_9450,N_9559);
xor U9733 (N_9733,N_9521,N_9556);
xnor U9734 (N_9734,N_9554,N_9589);
nand U9735 (N_9735,N_9583,N_9581);
xor U9736 (N_9736,N_9556,N_9514);
or U9737 (N_9737,N_9484,N_9470);
or U9738 (N_9738,N_9480,N_9533);
nand U9739 (N_9739,N_9580,N_9499);
or U9740 (N_9740,N_9590,N_9491);
and U9741 (N_9741,N_9487,N_9544);
nor U9742 (N_9742,N_9464,N_9525);
xnor U9743 (N_9743,N_9487,N_9564);
nor U9744 (N_9744,N_9584,N_9481);
and U9745 (N_9745,N_9590,N_9466);
nor U9746 (N_9746,N_9567,N_9512);
nand U9747 (N_9747,N_9453,N_9524);
xor U9748 (N_9748,N_9598,N_9483);
xnor U9749 (N_9749,N_9490,N_9595);
or U9750 (N_9750,N_9658,N_9619);
and U9751 (N_9751,N_9742,N_9672);
nand U9752 (N_9752,N_9737,N_9671);
nor U9753 (N_9753,N_9673,N_9633);
xnor U9754 (N_9754,N_9662,N_9724);
xor U9755 (N_9755,N_9725,N_9601);
and U9756 (N_9756,N_9684,N_9629);
nor U9757 (N_9757,N_9636,N_9704);
nand U9758 (N_9758,N_9606,N_9697);
nand U9759 (N_9759,N_9749,N_9650);
or U9760 (N_9760,N_9678,N_9748);
or U9761 (N_9761,N_9693,N_9634);
xnor U9762 (N_9762,N_9615,N_9628);
and U9763 (N_9763,N_9746,N_9632);
xnor U9764 (N_9764,N_9705,N_9626);
and U9765 (N_9765,N_9679,N_9608);
nand U9766 (N_9766,N_9713,N_9676);
or U9767 (N_9767,N_9730,N_9701);
or U9768 (N_9768,N_9702,N_9641);
nand U9769 (N_9769,N_9734,N_9717);
and U9770 (N_9770,N_9689,N_9692);
and U9771 (N_9771,N_9647,N_9613);
and U9772 (N_9772,N_9674,N_9667);
and U9773 (N_9773,N_9708,N_9740);
or U9774 (N_9774,N_9733,N_9660);
and U9775 (N_9775,N_9683,N_9700);
xnor U9776 (N_9776,N_9745,N_9719);
and U9777 (N_9777,N_9666,N_9621);
nor U9778 (N_9778,N_9723,N_9682);
nand U9779 (N_9779,N_9670,N_9685);
nor U9780 (N_9780,N_9649,N_9696);
and U9781 (N_9781,N_9744,N_9698);
nand U9782 (N_9782,N_9681,N_9677);
nand U9783 (N_9783,N_9664,N_9642);
xnor U9784 (N_9784,N_9653,N_9656);
nand U9785 (N_9785,N_9669,N_9688);
and U9786 (N_9786,N_9602,N_9651);
xnor U9787 (N_9787,N_9741,N_9635);
xor U9788 (N_9788,N_9646,N_9707);
nand U9789 (N_9789,N_9703,N_9645);
xor U9790 (N_9790,N_9699,N_9610);
nor U9791 (N_9791,N_9729,N_9739);
nand U9792 (N_9792,N_9747,N_9735);
nor U9793 (N_9793,N_9712,N_9668);
nand U9794 (N_9794,N_9600,N_9675);
nand U9795 (N_9795,N_9612,N_9652);
nand U9796 (N_9796,N_9625,N_9715);
and U9797 (N_9797,N_9630,N_9623);
or U9798 (N_9798,N_9631,N_9640);
or U9799 (N_9799,N_9663,N_9611);
and U9800 (N_9800,N_9620,N_9607);
xnor U9801 (N_9801,N_9654,N_9694);
nor U9802 (N_9802,N_9637,N_9680);
nand U9803 (N_9803,N_9617,N_9661);
nor U9804 (N_9804,N_9686,N_9639);
nand U9805 (N_9805,N_9718,N_9691);
nand U9806 (N_9806,N_9727,N_9690);
and U9807 (N_9807,N_9618,N_9603);
xor U9808 (N_9808,N_9604,N_9711);
and U9809 (N_9809,N_9687,N_9657);
nand U9810 (N_9810,N_9722,N_9643);
or U9811 (N_9811,N_9695,N_9720);
and U9812 (N_9812,N_9732,N_9665);
xor U9813 (N_9813,N_9716,N_9721);
nand U9814 (N_9814,N_9616,N_9648);
nor U9815 (N_9815,N_9644,N_9743);
xor U9816 (N_9816,N_9710,N_9736);
nor U9817 (N_9817,N_9609,N_9706);
nand U9818 (N_9818,N_9714,N_9605);
or U9819 (N_9819,N_9638,N_9655);
or U9820 (N_9820,N_9709,N_9738);
nor U9821 (N_9821,N_9731,N_9726);
or U9822 (N_9822,N_9728,N_9622);
nand U9823 (N_9823,N_9659,N_9627);
or U9824 (N_9824,N_9624,N_9614);
nand U9825 (N_9825,N_9604,N_9643);
and U9826 (N_9826,N_9711,N_9715);
nor U9827 (N_9827,N_9602,N_9740);
or U9828 (N_9828,N_9614,N_9610);
nand U9829 (N_9829,N_9640,N_9612);
nor U9830 (N_9830,N_9733,N_9723);
nor U9831 (N_9831,N_9615,N_9694);
nor U9832 (N_9832,N_9690,N_9654);
or U9833 (N_9833,N_9727,N_9614);
nand U9834 (N_9834,N_9610,N_9640);
nand U9835 (N_9835,N_9637,N_9728);
xnor U9836 (N_9836,N_9604,N_9737);
xnor U9837 (N_9837,N_9723,N_9709);
xor U9838 (N_9838,N_9727,N_9684);
and U9839 (N_9839,N_9620,N_9733);
nor U9840 (N_9840,N_9601,N_9624);
and U9841 (N_9841,N_9669,N_9672);
nor U9842 (N_9842,N_9655,N_9649);
xor U9843 (N_9843,N_9625,N_9653);
or U9844 (N_9844,N_9694,N_9604);
nand U9845 (N_9845,N_9712,N_9623);
nor U9846 (N_9846,N_9672,N_9666);
nand U9847 (N_9847,N_9660,N_9658);
and U9848 (N_9848,N_9723,N_9713);
nor U9849 (N_9849,N_9627,N_9733);
xor U9850 (N_9850,N_9716,N_9655);
or U9851 (N_9851,N_9658,N_9621);
and U9852 (N_9852,N_9602,N_9699);
or U9853 (N_9853,N_9704,N_9728);
nand U9854 (N_9854,N_9675,N_9720);
xor U9855 (N_9855,N_9748,N_9602);
xnor U9856 (N_9856,N_9679,N_9725);
nor U9857 (N_9857,N_9656,N_9693);
or U9858 (N_9858,N_9603,N_9730);
nor U9859 (N_9859,N_9608,N_9676);
xnor U9860 (N_9860,N_9682,N_9744);
and U9861 (N_9861,N_9604,N_9645);
and U9862 (N_9862,N_9702,N_9685);
or U9863 (N_9863,N_9695,N_9740);
and U9864 (N_9864,N_9656,N_9679);
nand U9865 (N_9865,N_9656,N_9721);
or U9866 (N_9866,N_9743,N_9639);
xnor U9867 (N_9867,N_9644,N_9731);
nand U9868 (N_9868,N_9629,N_9687);
nor U9869 (N_9869,N_9706,N_9645);
xnor U9870 (N_9870,N_9662,N_9731);
or U9871 (N_9871,N_9682,N_9636);
and U9872 (N_9872,N_9637,N_9727);
and U9873 (N_9873,N_9640,N_9728);
xor U9874 (N_9874,N_9713,N_9620);
and U9875 (N_9875,N_9644,N_9637);
or U9876 (N_9876,N_9711,N_9613);
nand U9877 (N_9877,N_9692,N_9611);
xor U9878 (N_9878,N_9667,N_9606);
xor U9879 (N_9879,N_9681,N_9658);
nand U9880 (N_9880,N_9699,N_9637);
and U9881 (N_9881,N_9627,N_9745);
and U9882 (N_9882,N_9603,N_9625);
xnor U9883 (N_9883,N_9640,N_9626);
or U9884 (N_9884,N_9708,N_9735);
nor U9885 (N_9885,N_9726,N_9686);
and U9886 (N_9886,N_9742,N_9744);
xor U9887 (N_9887,N_9623,N_9650);
xnor U9888 (N_9888,N_9686,N_9683);
and U9889 (N_9889,N_9600,N_9693);
nand U9890 (N_9890,N_9658,N_9728);
nand U9891 (N_9891,N_9673,N_9607);
and U9892 (N_9892,N_9717,N_9676);
nand U9893 (N_9893,N_9680,N_9713);
and U9894 (N_9894,N_9676,N_9747);
xnor U9895 (N_9895,N_9614,N_9618);
and U9896 (N_9896,N_9626,N_9736);
and U9897 (N_9897,N_9613,N_9619);
nand U9898 (N_9898,N_9606,N_9626);
xor U9899 (N_9899,N_9715,N_9709);
or U9900 (N_9900,N_9778,N_9752);
xnor U9901 (N_9901,N_9780,N_9814);
xor U9902 (N_9902,N_9758,N_9790);
nor U9903 (N_9903,N_9786,N_9757);
and U9904 (N_9904,N_9879,N_9803);
and U9905 (N_9905,N_9840,N_9865);
or U9906 (N_9906,N_9796,N_9772);
and U9907 (N_9907,N_9877,N_9891);
and U9908 (N_9908,N_9872,N_9751);
nand U9909 (N_9909,N_9851,N_9806);
xor U9910 (N_9910,N_9876,N_9855);
nor U9911 (N_9911,N_9767,N_9871);
nand U9912 (N_9912,N_9849,N_9889);
or U9913 (N_9913,N_9784,N_9843);
or U9914 (N_9914,N_9863,N_9848);
and U9915 (N_9915,N_9774,N_9844);
and U9916 (N_9916,N_9789,N_9823);
nand U9917 (N_9917,N_9811,N_9856);
nand U9918 (N_9918,N_9777,N_9787);
and U9919 (N_9919,N_9792,N_9883);
nand U9920 (N_9920,N_9887,N_9832);
xnor U9921 (N_9921,N_9853,N_9776);
xnor U9922 (N_9922,N_9818,N_9866);
and U9923 (N_9923,N_9797,N_9847);
and U9924 (N_9924,N_9799,N_9765);
xor U9925 (N_9925,N_9886,N_9756);
xor U9926 (N_9926,N_9822,N_9770);
or U9927 (N_9927,N_9852,N_9804);
nor U9928 (N_9928,N_9816,N_9807);
nor U9929 (N_9929,N_9858,N_9861);
and U9930 (N_9930,N_9753,N_9766);
xor U9931 (N_9931,N_9895,N_9817);
xnor U9932 (N_9932,N_9763,N_9859);
xor U9933 (N_9933,N_9831,N_9845);
nand U9934 (N_9934,N_9826,N_9841);
xor U9935 (N_9935,N_9829,N_9870);
nand U9936 (N_9936,N_9836,N_9830);
nand U9937 (N_9937,N_9890,N_9802);
and U9938 (N_9938,N_9825,N_9898);
or U9939 (N_9939,N_9838,N_9782);
or U9940 (N_9940,N_9769,N_9893);
nand U9941 (N_9941,N_9771,N_9800);
nand U9942 (N_9942,N_9795,N_9762);
nand U9943 (N_9943,N_9827,N_9812);
nand U9944 (N_9944,N_9839,N_9768);
nor U9945 (N_9945,N_9834,N_9750);
nand U9946 (N_9946,N_9791,N_9835);
nand U9947 (N_9947,N_9899,N_9779);
or U9948 (N_9948,N_9819,N_9788);
nor U9949 (N_9949,N_9837,N_9781);
and U9950 (N_9950,N_9760,N_9793);
and U9951 (N_9951,N_9821,N_9878);
nor U9952 (N_9952,N_9828,N_9755);
nand U9953 (N_9953,N_9894,N_9860);
nand U9954 (N_9954,N_9761,N_9850);
or U9955 (N_9955,N_9809,N_9764);
xnor U9956 (N_9956,N_9846,N_9754);
xnor U9957 (N_9957,N_9773,N_9884);
nor U9958 (N_9958,N_9815,N_9775);
and U9959 (N_9959,N_9874,N_9897);
xor U9960 (N_9960,N_9867,N_9869);
and U9961 (N_9961,N_9813,N_9820);
or U9962 (N_9962,N_9896,N_9785);
xor U9963 (N_9963,N_9888,N_9842);
nand U9964 (N_9964,N_9892,N_9798);
xnor U9965 (N_9965,N_9759,N_9885);
xnor U9966 (N_9966,N_9881,N_9873);
nor U9967 (N_9967,N_9783,N_9864);
nand U9968 (N_9968,N_9808,N_9805);
xor U9969 (N_9969,N_9882,N_9833);
xor U9970 (N_9970,N_9880,N_9824);
or U9971 (N_9971,N_9875,N_9857);
or U9972 (N_9972,N_9862,N_9810);
and U9973 (N_9973,N_9868,N_9854);
nor U9974 (N_9974,N_9801,N_9794);
nor U9975 (N_9975,N_9789,N_9862);
or U9976 (N_9976,N_9823,N_9796);
xor U9977 (N_9977,N_9817,N_9866);
and U9978 (N_9978,N_9762,N_9773);
or U9979 (N_9979,N_9811,N_9834);
or U9980 (N_9980,N_9816,N_9892);
nor U9981 (N_9981,N_9859,N_9886);
nand U9982 (N_9982,N_9753,N_9897);
nand U9983 (N_9983,N_9808,N_9777);
and U9984 (N_9984,N_9875,N_9790);
or U9985 (N_9985,N_9828,N_9822);
nand U9986 (N_9986,N_9760,N_9806);
and U9987 (N_9987,N_9834,N_9793);
or U9988 (N_9988,N_9840,N_9775);
nand U9989 (N_9989,N_9773,N_9769);
or U9990 (N_9990,N_9806,N_9765);
nor U9991 (N_9991,N_9869,N_9761);
nor U9992 (N_9992,N_9896,N_9761);
nor U9993 (N_9993,N_9883,N_9815);
nor U9994 (N_9994,N_9829,N_9850);
or U9995 (N_9995,N_9842,N_9750);
nor U9996 (N_9996,N_9873,N_9835);
xnor U9997 (N_9997,N_9888,N_9755);
nand U9998 (N_9998,N_9884,N_9890);
and U9999 (N_9999,N_9895,N_9772);
nor U10000 (N_10000,N_9819,N_9859);
or U10001 (N_10001,N_9874,N_9849);
xor U10002 (N_10002,N_9841,N_9800);
and U10003 (N_10003,N_9899,N_9807);
xor U10004 (N_10004,N_9813,N_9835);
and U10005 (N_10005,N_9779,N_9803);
nor U10006 (N_10006,N_9775,N_9800);
and U10007 (N_10007,N_9829,N_9867);
xor U10008 (N_10008,N_9847,N_9845);
nand U10009 (N_10009,N_9837,N_9882);
xor U10010 (N_10010,N_9861,N_9782);
xnor U10011 (N_10011,N_9844,N_9818);
and U10012 (N_10012,N_9807,N_9856);
and U10013 (N_10013,N_9799,N_9768);
and U10014 (N_10014,N_9846,N_9878);
or U10015 (N_10015,N_9771,N_9799);
xor U10016 (N_10016,N_9824,N_9849);
and U10017 (N_10017,N_9753,N_9760);
xor U10018 (N_10018,N_9863,N_9840);
nor U10019 (N_10019,N_9893,N_9805);
nor U10020 (N_10020,N_9849,N_9764);
or U10021 (N_10021,N_9789,N_9863);
or U10022 (N_10022,N_9833,N_9809);
and U10023 (N_10023,N_9865,N_9866);
or U10024 (N_10024,N_9899,N_9776);
xnor U10025 (N_10025,N_9777,N_9811);
nor U10026 (N_10026,N_9824,N_9751);
nor U10027 (N_10027,N_9797,N_9837);
nor U10028 (N_10028,N_9799,N_9801);
nor U10029 (N_10029,N_9799,N_9879);
xor U10030 (N_10030,N_9778,N_9761);
nand U10031 (N_10031,N_9833,N_9889);
or U10032 (N_10032,N_9829,N_9806);
or U10033 (N_10033,N_9771,N_9857);
nand U10034 (N_10034,N_9784,N_9867);
or U10035 (N_10035,N_9863,N_9877);
and U10036 (N_10036,N_9856,N_9794);
and U10037 (N_10037,N_9786,N_9778);
nor U10038 (N_10038,N_9793,N_9890);
nor U10039 (N_10039,N_9849,N_9899);
nand U10040 (N_10040,N_9804,N_9896);
nand U10041 (N_10041,N_9833,N_9860);
and U10042 (N_10042,N_9789,N_9794);
or U10043 (N_10043,N_9819,N_9839);
nor U10044 (N_10044,N_9824,N_9819);
or U10045 (N_10045,N_9870,N_9888);
nor U10046 (N_10046,N_9837,N_9859);
nand U10047 (N_10047,N_9799,N_9845);
and U10048 (N_10048,N_9874,N_9770);
xor U10049 (N_10049,N_9779,N_9774);
xnor U10050 (N_10050,N_10041,N_9986);
or U10051 (N_10051,N_9975,N_9994);
nor U10052 (N_10052,N_10001,N_10047);
nand U10053 (N_10053,N_9928,N_10022);
and U10054 (N_10054,N_10014,N_9990);
and U10055 (N_10055,N_10005,N_10002);
nor U10056 (N_10056,N_10042,N_9919);
nor U10057 (N_10057,N_9909,N_9944);
xnor U10058 (N_10058,N_9992,N_9934);
nor U10059 (N_10059,N_9958,N_9966);
nor U10060 (N_10060,N_9955,N_9991);
xor U10061 (N_10061,N_9937,N_9925);
and U10062 (N_10062,N_9930,N_9961);
nor U10063 (N_10063,N_9912,N_10039);
and U10064 (N_10064,N_9964,N_9924);
xor U10065 (N_10065,N_10049,N_10025);
xor U10066 (N_10066,N_9939,N_9979);
or U10067 (N_10067,N_9922,N_10016);
xnor U10068 (N_10068,N_10031,N_9945);
or U10069 (N_10069,N_9926,N_10003);
nor U10070 (N_10070,N_9936,N_9910);
xor U10071 (N_10071,N_9987,N_9977);
nor U10072 (N_10072,N_9943,N_10045);
nand U10073 (N_10073,N_10043,N_9941);
nor U10074 (N_10074,N_9971,N_10019);
xor U10075 (N_10075,N_9938,N_9962);
or U10076 (N_10076,N_10000,N_9931);
xnor U10077 (N_10077,N_9996,N_9963);
xnor U10078 (N_10078,N_9969,N_9970);
xor U10079 (N_10079,N_9956,N_9976);
nor U10080 (N_10080,N_9983,N_10021);
nand U10081 (N_10081,N_9918,N_9940);
and U10082 (N_10082,N_10009,N_10018);
and U10083 (N_10083,N_9998,N_9968);
nor U10084 (N_10084,N_10011,N_10032);
nand U10085 (N_10085,N_10024,N_10037);
xnor U10086 (N_10086,N_9920,N_10035);
and U10087 (N_10087,N_9985,N_9916);
or U10088 (N_10088,N_10030,N_9917);
nor U10089 (N_10089,N_9914,N_9960);
and U10090 (N_10090,N_9953,N_9905);
nand U10091 (N_10091,N_9906,N_9974);
and U10092 (N_10092,N_9942,N_9957);
and U10093 (N_10093,N_10046,N_9932);
xnor U10094 (N_10094,N_9935,N_9967);
nand U10095 (N_10095,N_9921,N_10029);
or U10096 (N_10096,N_9959,N_10026);
or U10097 (N_10097,N_9965,N_9923);
nor U10098 (N_10098,N_9927,N_10027);
and U10099 (N_10099,N_10007,N_9915);
or U10100 (N_10100,N_10033,N_9993);
nand U10101 (N_10101,N_9981,N_9997);
xor U10102 (N_10102,N_10036,N_9933);
and U10103 (N_10103,N_10044,N_9952);
nor U10104 (N_10104,N_9950,N_9972);
xnor U10105 (N_10105,N_9984,N_9900);
or U10106 (N_10106,N_10015,N_9954);
xnor U10107 (N_10107,N_9901,N_10006);
or U10108 (N_10108,N_9982,N_9988);
or U10109 (N_10109,N_9946,N_10028);
xnor U10110 (N_10110,N_10004,N_10048);
xnor U10111 (N_10111,N_9949,N_9947);
or U10112 (N_10112,N_10013,N_9907);
or U10113 (N_10113,N_9913,N_9995);
nor U10114 (N_10114,N_9903,N_10020);
nand U10115 (N_10115,N_9904,N_9951);
xor U10116 (N_10116,N_10010,N_9989);
nor U10117 (N_10117,N_10040,N_9999);
or U10118 (N_10118,N_10038,N_9948);
xor U10119 (N_10119,N_9973,N_9929);
xnor U10120 (N_10120,N_9978,N_10012);
xor U10121 (N_10121,N_10034,N_10008);
nor U10122 (N_10122,N_9908,N_9911);
and U10123 (N_10123,N_9980,N_10023);
xor U10124 (N_10124,N_10017,N_9902);
nand U10125 (N_10125,N_9937,N_9933);
nand U10126 (N_10126,N_9987,N_10041);
nand U10127 (N_10127,N_10013,N_10008);
nand U10128 (N_10128,N_9989,N_9908);
and U10129 (N_10129,N_9989,N_10046);
xnor U10130 (N_10130,N_9940,N_9967);
or U10131 (N_10131,N_9950,N_9980);
nand U10132 (N_10132,N_10029,N_9936);
and U10133 (N_10133,N_9929,N_10013);
nand U10134 (N_10134,N_9963,N_10034);
xnor U10135 (N_10135,N_9983,N_9994);
nand U10136 (N_10136,N_9965,N_9909);
xor U10137 (N_10137,N_9938,N_9988);
and U10138 (N_10138,N_9964,N_9958);
xnor U10139 (N_10139,N_10040,N_10038);
or U10140 (N_10140,N_9914,N_10022);
xnor U10141 (N_10141,N_9936,N_9931);
nand U10142 (N_10142,N_9907,N_9987);
nor U10143 (N_10143,N_10004,N_9968);
and U10144 (N_10144,N_10005,N_9915);
or U10145 (N_10145,N_9965,N_10006);
xnor U10146 (N_10146,N_9919,N_9964);
nor U10147 (N_10147,N_9921,N_9935);
nand U10148 (N_10148,N_9959,N_10042);
and U10149 (N_10149,N_9978,N_10040);
or U10150 (N_10150,N_10017,N_10041);
and U10151 (N_10151,N_9919,N_9942);
nor U10152 (N_10152,N_9938,N_10038);
xor U10153 (N_10153,N_9950,N_9952);
and U10154 (N_10154,N_10024,N_9966);
nand U10155 (N_10155,N_9917,N_9942);
nor U10156 (N_10156,N_9936,N_9914);
or U10157 (N_10157,N_10045,N_9951);
xor U10158 (N_10158,N_10028,N_10033);
nor U10159 (N_10159,N_9997,N_9967);
or U10160 (N_10160,N_10039,N_10018);
and U10161 (N_10161,N_9974,N_9987);
xor U10162 (N_10162,N_9947,N_10034);
nand U10163 (N_10163,N_9900,N_10004);
nand U10164 (N_10164,N_9912,N_9999);
xnor U10165 (N_10165,N_9955,N_9936);
or U10166 (N_10166,N_9971,N_10026);
xnor U10167 (N_10167,N_9984,N_10020);
nor U10168 (N_10168,N_9963,N_9955);
and U10169 (N_10169,N_9992,N_9988);
and U10170 (N_10170,N_9908,N_10033);
nand U10171 (N_10171,N_10016,N_9997);
nand U10172 (N_10172,N_10037,N_10001);
xnor U10173 (N_10173,N_10006,N_10001);
or U10174 (N_10174,N_9914,N_9975);
and U10175 (N_10175,N_9968,N_9976);
and U10176 (N_10176,N_9996,N_9903);
nor U10177 (N_10177,N_9917,N_10024);
nor U10178 (N_10178,N_10013,N_9939);
or U10179 (N_10179,N_9950,N_10027);
nand U10180 (N_10180,N_9975,N_10030);
and U10181 (N_10181,N_9930,N_9938);
or U10182 (N_10182,N_9935,N_9926);
or U10183 (N_10183,N_9959,N_9997);
xor U10184 (N_10184,N_9906,N_9967);
and U10185 (N_10185,N_9967,N_9977);
xor U10186 (N_10186,N_9995,N_9911);
and U10187 (N_10187,N_9922,N_10031);
nand U10188 (N_10188,N_9918,N_10015);
and U10189 (N_10189,N_9963,N_9919);
xor U10190 (N_10190,N_9900,N_9948);
or U10191 (N_10191,N_9908,N_9971);
and U10192 (N_10192,N_9982,N_10034);
nand U10193 (N_10193,N_9995,N_9958);
or U10194 (N_10194,N_9940,N_9987);
and U10195 (N_10195,N_9933,N_9990);
nor U10196 (N_10196,N_9971,N_10039);
and U10197 (N_10197,N_9942,N_9953);
xnor U10198 (N_10198,N_9909,N_9914);
and U10199 (N_10199,N_9927,N_9928);
nor U10200 (N_10200,N_10199,N_10075);
nand U10201 (N_10201,N_10096,N_10115);
nand U10202 (N_10202,N_10184,N_10080);
and U10203 (N_10203,N_10167,N_10169);
nand U10204 (N_10204,N_10114,N_10142);
and U10205 (N_10205,N_10143,N_10174);
or U10206 (N_10206,N_10178,N_10062);
nand U10207 (N_10207,N_10188,N_10104);
nor U10208 (N_10208,N_10088,N_10098);
nand U10209 (N_10209,N_10158,N_10120);
nor U10210 (N_10210,N_10086,N_10113);
nand U10211 (N_10211,N_10166,N_10112);
xor U10212 (N_10212,N_10194,N_10129);
and U10213 (N_10213,N_10138,N_10177);
or U10214 (N_10214,N_10157,N_10121);
xor U10215 (N_10215,N_10050,N_10068);
nand U10216 (N_10216,N_10066,N_10141);
nor U10217 (N_10217,N_10124,N_10052);
nand U10218 (N_10218,N_10134,N_10160);
and U10219 (N_10219,N_10172,N_10144);
xnor U10220 (N_10220,N_10084,N_10180);
nor U10221 (N_10221,N_10196,N_10065);
xor U10222 (N_10222,N_10101,N_10153);
and U10223 (N_10223,N_10155,N_10181);
nand U10224 (N_10224,N_10074,N_10179);
or U10225 (N_10225,N_10097,N_10132);
and U10226 (N_10226,N_10130,N_10067);
or U10227 (N_10227,N_10136,N_10054);
and U10228 (N_10228,N_10145,N_10056);
and U10229 (N_10229,N_10140,N_10061);
xnor U10230 (N_10230,N_10150,N_10105);
xor U10231 (N_10231,N_10090,N_10070);
nor U10232 (N_10232,N_10182,N_10118);
xnor U10233 (N_10233,N_10058,N_10135);
or U10234 (N_10234,N_10116,N_10192);
xnor U10235 (N_10235,N_10149,N_10064);
nor U10236 (N_10236,N_10091,N_10102);
and U10237 (N_10237,N_10103,N_10082);
or U10238 (N_10238,N_10193,N_10165);
or U10239 (N_10239,N_10173,N_10077);
and U10240 (N_10240,N_10139,N_10108);
and U10241 (N_10241,N_10163,N_10133);
xnor U10242 (N_10242,N_10175,N_10146);
nand U10243 (N_10243,N_10176,N_10151);
and U10244 (N_10244,N_10126,N_10161);
nor U10245 (N_10245,N_10168,N_10100);
xnor U10246 (N_10246,N_10131,N_10164);
nor U10247 (N_10247,N_10076,N_10189);
nor U10248 (N_10248,N_10128,N_10187);
or U10249 (N_10249,N_10081,N_10190);
and U10250 (N_10250,N_10198,N_10060);
nor U10251 (N_10251,N_10093,N_10170);
nor U10252 (N_10252,N_10117,N_10183);
nand U10253 (N_10253,N_10125,N_10071);
xnor U10254 (N_10254,N_10085,N_10099);
nor U10255 (N_10255,N_10057,N_10094);
nor U10256 (N_10256,N_10195,N_10059);
or U10257 (N_10257,N_10156,N_10092);
or U10258 (N_10258,N_10111,N_10191);
or U10259 (N_10259,N_10197,N_10185);
and U10260 (N_10260,N_10069,N_10110);
nor U10261 (N_10261,N_10087,N_10083);
nor U10262 (N_10262,N_10148,N_10122);
and U10263 (N_10263,N_10137,N_10162);
xor U10264 (N_10264,N_10079,N_10152);
xor U10265 (N_10265,N_10123,N_10051);
nor U10266 (N_10266,N_10154,N_10053);
and U10267 (N_10267,N_10109,N_10107);
and U10268 (N_10268,N_10072,N_10073);
or U10269 (N_10269,N_10147,N_10078);
and U10270 (N_10270,N_10106,N_10089);
or U10271 (N_10271,N_10095,N_10186);
or U10272 (N_10272,N_10063,N_10055);
nand U10273 (N_10273,N_10127,N_10159);
or U10274 (N_10274,N_10171,N_10119);
and U10275 (N_10275,N_10124,N_10100);
xnor U10276 (N_10276,N_10173,N_10184);
nand U10277 (N_10277,N_10124,N_10064);
or U10278 (N_10278,N_10090,N_10076);
and U10279 (N_10279,N_10103,N_10183);
xnor U10280 (N_10280,N_10162,N_10123);
nand U10281 (N_10281,N_10073,N_10114);
xnor U10282 (N_10282,N_10122,N_10184);
and U10283 (N_10283,N_10088,N_10138);
or U10284 (N_10284,N_10101,N_10190);
and U10285 (N_10285,N_10097,N_10120);
nand U10286 (N_10286,N_10068,N_10194);
or U10287 (N_10287,N_10197,N_10198);
and U10288 (N_10288,N_10194,N_10105);
nand U10289 (N_10289,N_10164,N_10062);
xor U10290 (N_10290,N_10064,N_10144);
nand U10291 (N_10291,N_10157,N_10129);
nor U10292 (N_10292,N_10063,N_10093);
xnor U10293 (N_10293,N_10188,N_10138);
or U10294 (N_10294,N_10113,N_10128);
nor U10295 (N_10295,N_10116,N_10175);
and U10296 (N_10296,N_10141,N_10122);
nor U10297 (N_10297,N_10053,N_10197);
and U10298 (N_10298,N_10187,N_10175);
or U10299 (N_10299,N_10066,N_10099);
xnor U10300 (N_10300,N_10096,N_10160);
xor U10301 (N_10301,N_10131,N_10154);
nand U10302 (N_10302,N_10062,N_10179);
and U10303 (N_10303,N_10169,N_10059);
xor U10304 (N_10304,N_10144,N_10161);
and U10305 (N_10305,N_10131,N_10155);
nor U10306 (N_10306,N_10081,N_10076);
or U10307 (N_10307,N_10124,N_10188);
nor U10308 (N_10308,N_10161,N_10092);
nand U10309 (N_10309,N_10098,N_10147);
and U10310 (N_10310,N_10134,N_10192);
nand U10311 (N_10311,N_10066,N_10090);
or U10312 (N_10312,N_10186,N_10129);
nor U10313 (N_10313,N_10113,N_10080);
xor U10314 (N_10314,N_10087,N_10141);
and U10315 (N_10315,N_10120,N_10125);
xnor U10316 (N_10316,N_10162,N_10110);
and U10317 (N_10317,N_10166,N_10095);
or U10318 (N_10318,N_10093,N_10055);
and U10319 (N_10319,N_10190,N_10168);
nor U10320 (N_10320,N_10099,N_10104);
xor U10321 (N_10321,N_10112,N_10051);
or U10322 (N_10322,N_10172,N_10146);
nor U10323 (N_10323,N_10055,N_10154);
or U10324 (N_10324,N_10195,N_10109);
and U10325 (N_10325,N_10054,N_10053);
nand U10326 (N_10326,N_10174,N_10178);
or U10327 (N_10327,N_10145,N_10139);
nand U10328 (N_10328,N_10151,N_10130);
and U10329 (N_10329,N_10166,N_10076);
nor U10330 (N_10330,N_10104,N_10080);
or U10331 (N_10331,N_10059,N_10100);
nand U10332 (N_10332,N_10076,N_10100);
and U10333 (N_10333,N_10185,N_10136);
and U10334 (N_10334,N_10079,N_10092);
nand U10335 (N_10335,N_10179,N_10139);
and U10336 (N_10336,N_10130,N_10150);
nand U10337 (N_10337,N_10173,N_10159);
nor U10338 (N_10338,N_10097,N_10103);
or U10339 (N_10339,N_10068,N_10139);
and U10340 (N_10340,N_10158,N_10093);
and U10341 (N_10341,N_10108,N_10135);
nand U10342 (N_10342,N_10101,N_10174);
nor U10343 (N_10343,N_10092,N_10130);
and U10344 (N_10344,N_10091,N_10100);
xnor U10345 (N_10345,N_10068,N_10147);
and U10346 (N_10346,N_10113,N_10117);
or U10347 (N_10347,N_10199,N_10182);
or U10348 (N_10348,N_10088,N_10116);
or U10349 (N_10349,N_10171,N_10179);
xnor U10350 (N_10350,N_10211,N_10237);
nand U10351 (N_10351,N_10296,N_10309);
nor U10352 (N_10352,N_10231,N_10249);
xnor U10353 (N_10353,N_10256,N_10252);
and U10354 (N_10354,N_10315,N_10325);
nand U10355 (N_10355,N_10208,N_10205);
and U10356 (N_10356,N_10333,N_10348);
and U10357 (N_10357,N_10234,N_10220);
xor U10358 (N_10358,N_10340,N_10259);
and U10359 (N_10359,N_10204,N_10241);
and U10360 (N_10360,N_10213,N_10347);
and U10361 (N_10361,N_10219,N_10297);
nor U10362 (N_10362,N_10304,N_10308);
nor U10363 (N_10363,N_10262,N_10223);
xnor U10364 (N_10364,N_10332,N_10277);
and U10365 (N_10365,N_10286,N_10287);
or U10366 (N_10366,N_10268,N_10320);
and U10367 (N_10367,N_10246,N_10322);
xor U10368 (N_10368,N_10225,N_10214);
or U10369 (N_10369,N_10337,N_10294);
or U10370 (N_10370,N_10215,N_10218);
nor U10371 (N_10371,N_10321,N_10284);
xnor U10372 (N_10372,N_10282,N_10257);
nand U10373 (N_10373,N_10221,N_10289);
xor U10374 (N_10374,N_10343,N_10317);
xor U10375 (N_10375,N_10318,N_10226);
and U10376 (N_10376,N_10349,N_10310);
nor U10377 (N_10377,N_10291,N_10207);
and U10378 (N_10378,N_10327,N_10244);
xor U10379 (N_10379,N_10316,N_10261);
or U10380 (N_10380,N_10224,N_10243);
and U10381 (N_10381,N_10341,N_10295);
and U10382 (N_10382,N_10330,N_10279);
nand U10383 (N_10383,N_10212,N_10278);
and U10384 (N_10384,N_10344,N_10245);
xnor U10385 (N_10385,N_10339,N_10281);
or U10386 (N_10386,N_10273,N_10301);
and U10387 (N_10387,N_10331,N_10326);
nand U10388 (N_10388,N_10306,N_10222);
or U10389 (N_10389,N_10323,N_10230);
nand U10390 (N_10390,N_10227,N_10233);
nor U10391 (N_10391,N_10255,N_10209);
and U10392 (N_10392,N_10258,N_10229);
nand U10393 (N_10393,N_10283,N_10239);
nand U10394 (N_10394,N_10314,N_10298);
nor U10395 (N_10395,N_10250,N_10248);
and U10396 (N_10396,N_10345,N_10200);
xor U10397 (N_10397,N_10238,N_10276);
or U10398 (N_10398,N_10311,N_10251);
nand U10399 (N_10399,N_10293,N_10299);
or U10400 (N_10400,N_10236,N_10232);
or U10401 (N_10401,N_10280,N_10267);
nor U10402 (N_10402,N_10285,N_10324);
nor U10403 (N_10403,N_10206,N_10272);
and U10404 (N_10404,N_10263,N_10292);
or U10405 (N_10405,N_10228,N_10240);
nand U10406 (N_10406,N_10307,N_10329);
and U10407 (N_10407,N_10203,N_10328);
and U10408 (N_10408,N_10201,N_10217);
and U10409 (N_10409,N_10290,N_10335);
and U10410 (N_10410,N_10346,N_10247);
or U10411 (N_10411,N_10271,N_10313);
nor U10412 (N_10412,N_10303,N_10242);
nor U10413 (N_10413,N_10338,N_10275);
nand U10414 (N_10414,N_10288,N_10270);
and U10415 (N_10415,N_10312,N_10269);
xnor U10416 (N_10416,N_10302,N_10260);
or U10417 (N_10417,N_10253,N_10264);
xor U10418 (N_10418,N_10254,N_10266);
nor U10419 (N_10419,N_10305,N_10336);
or U10420 (N_10420,N_10342,N_10300);
and U10421 (N_10421,N_10265,N_10210);
and U10422 (N_10422,N_10274,N_10235);
or U10423 (N_10423,N_10216,N_10319);
nor U10424 (N_10424,N_10334,N_10202);
nand U10425 (N_10425,N_10292,N_10306);
or U10426 (N_10426,N_10342,N_10231);
nand U10427 (N_10427,N_10220,N_10325);
or U10428 (N_10428,N_10337,N_10233);
nor U10429 (N_10429,N_10209,N_10330);
xnor U10430 (N_10430,N_10270,N_10215);
and U10431 (N_10431,N_10249,N_10346);
nand U10432 (N_10432,N_10331,N_10330);
or U10433 (N_10433,N_10218,N_10323);
or U10434 (N_10434,N_10303,N_10250);
or U10435 (N_10435,N_10281,N_10258);
or U10436 (N_10436,N_10202,N_10284);
or U10437 (N_10437,N_10251,N_10341);
nand U10438 (N_10438,N_10297,N_10336);
xnor U10439 (N_10439,N_10203,N_10245);
or U10440 (N_10440,N_10242,N_10316);
nand U10441 (N_10441,N_10268,N_10293);
or U10442 (N_10442,N_10227,N_10202);
nor U10443 (N_10443,N_10348,N_10239);
or U10444 (N_10444,N_10238,N_10273);
or U10445 (N_10445,N_10201,N_10232);
or U10446 (N_10446,N_10247,N_10325);
nor U10447 (N_10447,N_10238,N_10257);
and U10448 (N_10448,N_10342,N_10272);
or U10449 (N_10449,N_10347,N_10277);
nand U10450 (N_10450,N_10242,N_10229);
or U10451 (N_10451,N_10329,N_10260);
or U10452 (N_10452,N_10280,N_10330);
and U10453 (N_10453,N_10310,N_10327);
and U10454 (N_10454,N_10315,N_10200);
nand U10455 (N_10455,N_10316,N_10235);
or U10456 (N_10456,N_10243,N_10210);
and U10457 (N_10457,N_10346,N_10289);
nor U10458 (N_10458,N_10321,N_10307);
or U10459 (N_10459,N_10294,N_10347);
xnor U10460 (N_10460,N_10346,N_10310);
and U10461 (N_10461,N_10208,N_10292);
xor U10462 (N_10462,N_10276,N_10278);
nor U10463 (N_10463,N_10317,N_10287);
nor U10464 (N_10464,N_10246,N_10235);
nand U10465 (N_10465,N_10316,N_10210);
nor U10466 (N_10466,N_10213,N_10303);
and U10467 (N_10467,N_10230,N_10286);
nor U10468 (N_10468,N_10335,N_10252);
or U10469 (N_10469,N_10208,N_10347);
and U10470 (N_10470,N_10223,N_10290);
nor U10471 (N_10471,N_10313,N_10220);
xnor U10472 (N_10472,N_10322,N_10287);
xnor U10473 (N_10473,N_10345,N_10264);
and U10474 (N_10474,N_10228,N_10243);
xnor U10475 (N_10475,N_10233,N_10309);
nor U10476 (N_10476,N_10336,N_10300);
or U10477 (N_10477,N_10227,N_10205);
and U10478 (N_10478,N_10255,N_10337);
xor U10479 (N_10479,N_10305,N_10307);
nand U10480 (N_10480,N_10247,N_10215);
or U10481 (N_10481,N_10218,N_10313);
xor U10482 (N_10482,N_10333,N_10317);
nor U10483 (N_10483,N_10212,N_10330);
xnor U10484 (N_10484,N_10233,N_10253);
xor U10485 (N_10485,N_10283,N_10326);
nand U10486 (N_10486,N_10255,N_10298);
xor U10487 (N_10487,N_10299,N_10215);
and U10488 (N_10488,N_10232,N_10251);
or U10489 (N_10489,N_10231,N_10301);
or U10490 (N_10490,N_10338,N_10310);
or U10491 (N_10491,N_10255,N_10309);
xor U10492 (N_10492,N_10298,N_10336);
nor U10493 (N_10493,N_10212,N_10283);
or U10494 (N_10494,N_10291,N_10267);
nand U10495 (N_10495,N_10267,N_10271);
nor U10496 (N_10496,N_10315,N_10322);
nand U10497 (N_10497,N_10311,N_10284);
xor U10498 (N_10498,N_10260,N_10228);
nand U10499 (N_10499,N_10346,N_10307);
and U10500 (N_10500,N_10356,N_10428);
nand U10501 (N_10501,N_10360,N_10371);
nand U10502 (N_10502,N_10495,N_10430);
nand U10503 (N_10503,N_10449,N_10413);
and U10504 (N_10504,N_10433,N_10374);
nand U10505 (N_10505,N_10411,N_10405);
nor U10506 (N_10506,N_10358,N_10440);
nor U10507 (N_10507,N_10462,N_10456);
or U10508 (N_10508,N_10441,N_10499);
nand U10509 (N_10509,N_10385,N_10444);
nor U10510 (N_10510,N_10412,N_10457);
or U10511 (N_10511,N_10453,N_10437);
xnor U10512 (N_10512,N_10459,N_10467);
xnor U10513 (N_10513,N_10410,N_10447);
and U10514 (N_10514,N_10471,N_10470);
nor U10515 (N_10515,N_10469,N_10364);
xnor U10516 (N_10516,N_10480,N_10435);
xor U10517 (N_10517,N_10481,N_10479);
nand U10518 (N_10518,N_10420,N_10376);
nand U10519 (N_10519,N_10366,N_10357);
and U10520 (N_10520,N_10386,N_10373);
nor U10521 (N_10521,N_10372,N_10363);
xor U10522 (N_10522,N_10391,N_10408);
nand U10523 (N_10523,N_10354,N_10416);
and U10524 (N_10524,N_10370,N_10443);
and U10525 (N_10525,N_10406,N_10442);
xnor U10526 (N_10526,N_10380,N_10432);
or U10527 (N_10527,N_10446,N_10384);
or U10528 (N_10528,N_10421,N_10427);
and U10529 (N_10529,N_10353,N_10492);
and U10530 (N_10530,N_10468,N_10483);
or U10531 (N_10531,N_10445,N_10450);
or U10532 (N_10532,N_10381,N_10389);
and U10533 (N_10533,N_10403,N_10418);
and U10534 (N_10534,N_10434,N_10489);
xnor U10535 (N_10535,N_10491,N_10362);
nor U10536 (N_10536,N_10390,N_10448);
nor U10537 (N_10537,N_10394,N_10439);
nand U10538 (N_10538,N_10407,N_10458);
xor U10539 (N_10539,N_10388,N_10397);
nand U10540 (N_10540,N_10415,N_10367);
nand U10541 (N_10541,N_10361,N_10350);
nor U10542 (N_10542,N_10478,N_10438);
nor U10543 (N_10543,N_10486,N_10369);
and U10544 (N_10544,N_10429,N_10375);
xnor U10545 (N_10545,N_10378,N_10383);
nand U10546 (N_10546,N_10393,N_10417);
and U10547 (N_10547,N_10498,N_10382);
nor U10548 (N_10548,N_10454,N_10436);
or U10549 (N_10549,N_10404,N_10493);
xnor U10550 (N_10550,N_10475,N_10422);
or U10551 (N_10551,N_10401,N_10472);
or U10552 (N_10552,N_10423,N_10482);
or U10553 (N_10553,N_10368,N_10365);
xnor U10554 (N_10554,N_10451,N_10351);
and U10555 (N_10555,N_10359,N_10485);
or U10556 (N_10556,N_10496,N_10488);
xnor U10557 (N_10557,N_10398,N_10352);
xnor U10558 (N_10558,N_10490,N_10419);
xnor U10559 (N_10559,N_10477,N_10402);
and U10560 (N_10560,N_10377,N_10395);
xnor U10561 (N_10561,N_10399,N_10466);
or U10562 (N_10562,N_10476,N_10461);
and U10563 (N_10563,N_10473,N_10464);
nor U10564 (N_10564,N_10487,N_10424);
nand U10565 (N_10565,N_10431,N_10452);
xor U10566 (N_10566,N_10474,N_10425);
nor U10567 (N_10567,N_10460,N_10494);
xor U10568 (N_10568,N_10484,N_10379);
nand U10569 (N_10569,N_10396,N_10463);
and U10570 (N_10570,N_10409,N_10400);
nor U10571 (N_10571,N_10387,N_10455);
or U10572 (N_10572,N_10414,N_10426);
and U10573 (N_10573,N_10392,N_10355);
xnor U10574 (N_10574,N_10465,N_10497);
nor U10575 (N_10575,N_10482,N_10489);
and U10576 (N_10576,N_10427,N_10422);
nand U10577 (N_10577,N_10437,N_10430);
or U10578 (N_10578,N_10448,N_10399);
or U10579 (N_10579,N_10476,N_10380);
xnor U10580 (N_10580,N_10413,N_10415);
or U10581 (N_10581,N_10458,N_10424);
xnor U10582 (N_10582,N_10414,N_10498);
or U10583 (N_10583,N_10474,N_10398);
or U10584 (N_10584,N_10378,N_10482);
or U10585 (N_10585,N_10375,N_10470);
nor U10586 (N_10586,N_10432,N_10369);
xor U10587 (N_10587,N_10469,N_10431);
xnor U10588 (N_10588,N_10455,N_10400);
nand U10589 (N_10589,N_10499,N_10398);
or U10590 (N_10590,N_10419,N_10455);
nand U10591 (N_10591,N_10360,N_10405);
nor U10592 (N_10592,N_10374,N_10416);
and U10593 (N_10593,N_10490,N_10486);
nand U10594 (N_10594,N_10487,N_10449);
nand U10595 (N_10595,N_10490,N_10480);
and U10596 (N_10596,N_10466,N_10430);
nor U10597 (N_10597,N_10354,N_10357);
xnor U10598 (N_10598,N_10378,N_10449);
nand U10599 (N_10599,N_10403,N_10434);
nor U10600 (N_10600,N_10353,N_10437);
nor U10601 (N_10601,N_10427,N_10461);
or U10602 (N_10602,N_10398,N_10394);
nand U10603 (N_10603,N_10369,N_10385);
and U10604 (N_10604,N_10439,N_10428);
nor U10605 (N_10605,N_10479,N_10394);
nor U10606 (N_10606,N_10466,N_10435);
nand U10607 (N_10607,N_10494,N_10375);
or U10608 (N_10608,N_10404,N_10496);
nand U10609 (N_10609,N_10403,N_10382);
or U10610 (N_10610,N_10363,N_10378);
and U10611 (N_10611,N_10392,N_10413);
or U10612 (N_10612,N_10465,N_10442);
nand U10613 (N_10613,N_10409,N_10393);
xor U10614 (N_10614,N_10392,N_10466);
and U10615 (N_10615,N_10370,N_10368);
or U10616 (N_10616,N_10498,N_10486);
or U10617 (N_10617,N_10354,N_10418);
xor U10618 (N_10618,N_10416,N_10373);
or U10619 (N_10619,N_10380,N_10477);
or U10620 (N_10620,N_10401,N_10384);
or U10621 (N_10621,N_10488,N_10364);
or U10622 (N_10622,N_10470,N_10478);
and U10623 (N_10623,N_10359,N_10417);
or U10624 (N_10624,N_10386,N_10385);
and U10625 (N_10625,N_10426,N_10369);
nand U10626 (N_10626,N_10492,N_10354);
or U10627 (N_10627,N_10482,N_10412);
and U10628 (N_10628,N_10477,N_10379);
or U10629 (N_10629,N_10366,N_10413);
and U10630 (N_10630,N_10457,N_10468);
and U10631 (N_10631,N_10449,N_10383);
xnor U10632 (N_10632,N_10369,N_10441);
xor U10633 (N_10633,N_10493,N_10367);
xor U10634 (N_10634,N_10363,N_10448);
and U10635 (N_10635,N_10498,N_10351);
and U10636 (N_10636,N_10376,N_10451);
nor U10637 (N_10637,N_10498,N_10422);
or U10638 (N_10638,N_10379,N_10496);
xor U10639 (N_10639,N_10452,N_10466);
and U10640 (N_10640,N_10454,N_10496);
xnor U10641 (N_10641,N_10404,N_10489);
nand U10642 (N_10642,N_10379,N_10372);
or U10643 (N_10643,N_10376,N_10497);
nand U10644 (N_10644,N_10356,N_10412);
nand U10645 (N_10645,N_10409,N_10456);
and U10646 (N_10646,N_10366,N_10472);
nand U10647 (N_10647,N_10393,N_10489);
and U10648 (N_10648,N_10417,N_10442);
xnor U10649 (N_10649,N_10411,N_10472);
or U10650 (N_10650,N_10603,N_10568);
nand U10651 (N_10651,N_10633,N_10619);
nor U10652 (N_10652,N_10548,N_10615);
or U10653 (N_10653,N_10599,N_10592);
xnor U10654 (N_10654,N_10639,N_10546);
nor U10655 (N_10655,N_10503,N_10635);
nor U10656 (N_10656,N_10521,N_10628);
or U10657 (N_10657,N_10645,N_10544);
and U10658 (N_10658,N_10528,N_10648);
and U10659 (N_10659,N_10508,N_10573);
xor U10660 (N_10660,N_10579,N_10595);
or U10661 (N_10661,N_10514,N_10609);
xnor U10662 (N_10662,N_10625,N_10640);
nor U10663 (N_10663,N_10598,N_10551);
nand U10664 (N_10664,N_10578,N_10506);
xor U10665 (N_10665,N_10560,N_10563);
nor U10666 (N_10666,N_10618,N_10602);
and U10667 (N_10667,N_10580,N_10583);
xnor U10668 (N_10668,N_10525,N_10536);
or U10669 (N_10669,N_10574,N_10561);
xor U10670 (N_10670,N_10611,N_10638);
or U10671 (N_10671,N_10559,N_10509);
and U10672 (N_10672,N_10636,N_10620);
nor U10673 (N_10673,N_10555,N_10607);
and U10674 (N_10674,N_10532,N_10564);
and U10675 (N_10675,N_10537,N_10637);
and U10676 (N_10676,N_10549,N_10629);
xor U10677 (N_10677,N_10566,N_10510);
xnor U10678 (N_10678,N_10647,N_10591);
xnor U10679 (N_10679,N_10502,N_10540);
nand U10680 (N_10680,N_10535,N_10505);
xnor U10681 (N_10681,N_10501,N_10558);
or U10682 (N_10682,N_10569,N_10634);
nand U10683 (N_10683,N_10538,N_10530);
nor U10684 (N_10684,N_10621,N_10588);
nand U10685 (N_10685,N_10557,N_10526);
or U10686 (N_10686,N_10614,N_10570);
xnor U10687 (N_10687,N_10594,N_10527);
or U10688 (N_10688,N_10512,N_10523);
xnor U10689 (N_10689,N_10584,N_10642);
and U10690 (N_10690,N_10517,N_10518);
nor U10691 (N_10691,N_10507,N_10575);
or U10692 (N_10692,N_10533,N_10643);
and U10693 (N_10693,N_10612,N_10622);
xnor U10694 (N_10694,N_10596,N_10547);
and U10695 (N_10695,N_10605,N_10606);
nor U10696 (N_10696,N_10554,N_10562);
nor U10697 (N_10697,N_10577,N_10631);
nor U10698 (N_10698,N_10520,N_10627);
xor U10699 (N_10699,N_10593,N_10597);
and U10700 (N_10700,N_10610,N_10511);
xnor U10701 (N_10701,N_10617,N_10531);
nor U10702 (N_10702,N_10600,N_10542);
or U10703 (N_10703,N_10582,N_10571);
nor U10704 (N_10704,N_10587,N_10589);
xor U10705 (N_10705,N_10601,N_10604);
nand U10706 (N_10706,N_10646,N_10541);
xnor U10707 (N_10707,N_10626,N_10556);
xnor U10708 (N_10708,N_10641,N_10552);
xnor U10709 (N_10709,N_10567,N_10504);
nor U10710 (N_10710,N_10545,N_10515);
and U10711 (N_10711,N_10529,N_10585);
and U10712 (N_10712,N_10616,N_10590);
xor U10713 (N_10713,N_10581,N_10623);
and U10714 (N_10714,N_10500,N_10649);
xor U10715 (N_10715,N_10553,N_10519);
xnor U10716 (N_10716,N_10516,N_10613);
xnor U10717 (N_10717,N_10608,N_10543);
or U10718 (N_10718,N_10550,N_10565);
and U10719 (N_10719,N_10644,N_10513);
nor U10720 (N_10720,N_10522,N_10630);
or U10721 (N_10721,N_10534,N_10524);
nor U10722 (N_10722,N_10576,N_10586);
and U10723 (N_10723,N_10624,N_10539);
xor U10724 (N_10724,N_10632,N_10572);
or U10725 (N_10725,N_10584,N_10618);
or U10726 (N_10726,N_10539,N_10531);
nor U10727 (N_10727,N_10503,N_10522);
or U10728 (N_10728,N_10546,N_10535);
xor U10729 (N_10729,N_10566,N_10571);
and U10730 (N_10730,N_10559,N_10501);
nor U10731 (N_10731,N_10646,N_10559);
xnor U10732 (N_10732,N_10513,N_10562);
xor U10733 (N_10733,N_10566,N_10533);
nor U10734 (N_10734,N_10607,N_10554);
and U10735 (N_10735,N_10524,N_10540);
or U10736 (N_10736,N_10556,N_10514);
nand U10737 (N_10737,N_10625,N_10577);
nand U10738 (N_10738,N_10636,N_10616);
nand U10739 (N_10739,N_10554,N_10620);
xnor U10740 (N_10740,N_10594,N_10644);
or U10741 (N_10741,N_10627,N_10555);
xnor U10742 (N_10742,N_10528,N_10587);
nor U10743 (N_10743,N_10579,N_10539);
or U10744 (N_10744,N_10598,N_10501);
xnor U10745 (N_10745,N_10552,N_10615);
or U10746 (N_10746,N_10631,N_10530);
xor U10747 (N_10747,N_10561,N_10636);
xnor U10748 (N_10748,N_10541,N_10567);
or U10749 (N_10749,N_10583,N_10516);
xor U10750 (N_10750,N_10536,N_10618);
xnor U10751 (N_10751,N_10602,N_10500);
and U10752 (N_10752,N_10550,N_10646);
or U10753 (N_10753,N_10555,N_10578);
or U10754 (N_10754,N_10626,N_10583);
nand U10755 (N_10755,N_10620,N_10593);
xor U10756 (N_10756,N_10624,N_10557);
nor U10757 (N_10757,N_10520,N_10576);
nand U10758 (N_10758,N_10648,N_10513);
nor U10759 (N_10759,N_10593,N_10592);
or U10760 (N_10760,N_10610,N_10632);
or U10761 (N_10761,N_10599,N_10612);
or U10762 (N_10762,N_10605,N_10635);
and U10763 (N_10763,N_10532,N_10581);
nor U10764 (N_10764,N_10633,N_10500);
or U10765 (N_10765,N_10590,N_10579);
nand U10766 (N_10766,N_10562,N_10551);
nand U10767 (N_10767,N_10611,N_10603);
nor U10768 (N_10768,N_10511,N_10517);
or U10769 (N_10769,N_10573,N_10645);
nor U10770 (N_10770,N_10500,N_10515);
nand U10771 (N_10771,N_10634,N_10510);
nor U10772 (N_10772,N_10601,N_10611);
or U10773 (N_10773,N_10625,N_10570);
xor U10774 (N_10774,N_10645,N_10558);
or U10775 (N_10775,N_10598,N_10555);
xnor U10776 (N_10776,N_10615,N_10622);
and U10777 (N_10777,N_10561,N_10638);
xor U10778 (N_10778,N_10642,N_10623);
xnor U10779 (N_10779,N_10550,N_10636);
and U10780 (N_10780,N_10613,N_10612);
xnor U10781 (N_10781,N_10548,N_10566);
nand U10782 (N_10782,N_10561,N_10626);
nand U10783 (N_10783,N_10534,N_10611);
and U10784 (N_10784,N_10625,N_10518);
and U10785 (N_10785,N_10597,N_10569);
nor U10786 (N_10786,N_10501,N_10538);
and U10787 (N_10787,N_10547,N_10522);
nand U10788 (N_10788,N_10523,N_10617);
and U10789 (N_10789,N_10503,N_10647);
nor U10790 (N_10790,N_10644,N_10581);
xnor U10791 (N_10791,N_10638,N_10612);
and U10792 (N_10792,N_10608,N_10633);
xnor U10793 (N_10793,N_10550,N_10511);
and U10794 (N_10794,N_10607,N_10615);
or U10795 (N_10795,N_10624,N_10545);
nand U10796 (N_10796,N_10629,N_10553);
or U10797 (N_10797,N_10616,N_10574);
and U10798 (N_10798,N_10555,N_10537);
xnor U10799 (N_10799,N_10638,N_10596);
or U10800 (N_10800,N_10685,N_10711);
xor U10801 (N_10801,N_10656,N_10770);
nand U10802 (N_10802,N_10679,N_10767);
nor U10803 (N_10803,N_10762,N_10728);
nor U10804 (N_10804,N_10778,N_10664);
nor U10805 (N_10805,N_10673,N_10743);
nand U10806 (N_10806,N_10694,N_10666);
nand U10807 (N_10807,N_10742,N_10697);
nand U10808 (N_10808,N_10713,N_10754);
nor U10809 (N_10809,N_10796,N_10683);
xnor U10810 (N_10810,N_10702,N_10750);
nor U10811 (N_10811,N_10721,N_10655);
nand U10812 (N_10812,N_10791,N_10689);
and U10813 (N_10813,N_10756,N_10717);
nand U10814 (N_10814,N_10797,N_10736);
xnor U10815 (N_10815,N_10744,N_10708);
nor U10816 (N_10816,N_10723,N_10740);
and U10817 (N_10817,N_10735,N_10775);
nor U10818 (N_10818,N_10786,N_10653);
and U10819 (N_10819,N_10782,N_10672);
nand U10820 (N_10820,N_10651,N_10752);
and U10821 (N_10821,N_10707,N_10729);
or U10822 (N_10822,N_10719,N_10773);
nand U10823 (N_10823,N_10692,N_10709);
xor U10824 (N_10824,N_10706,N_10737);
nand U10825 (N_10825,N_10678,N_10720);
and U10826 (N_10826,N_10712,N_10789);
or U10827 (N_10827,N_10691,N_10768);
nand U10828 (N_10828,N_10670,N_10659);
and U10829 (N_10829,N_10686,N_10682);
nor U10830 (N_10830,N_10765,N_10671);
nand U10831 (N_10831,N_10779,N_10718);
and U10832 (N_10832,N_10746,N_10763);
and U10833 (N_10833,N_10792,N_10663);
and U10834 (N_10834,N_10677,N_10668);
xnor U10835 (N_10835,N_10755,N_10784);
xor U10836 (N_10836,N_10724,N_10794);
and U10837 (N_10837,N_10722,N_10738);
and U10838 (N_10838,N_10681,N_10688);
and U10839 (N_10839,N_10795,N_10799);
xnor U10840 (N_10840,N_10714,N_10667);
nor U10841 (N_10841,N_10749,N_10731);
nor U10842 (N_10842,N_10696,N_10758);
nand U10843 (N_10843,N_10761,N_10725);
xnor U10844 (N_10844,N_10751,N_10662);
or U10845 (N_10845,N_10787,N_10780);
and U10846 (N_10846,N_10734,N_10650);
xor U10847 (N_10847,N_10716,N_10699);
and U10848 (N_10848,N_10747,N_10698);
and U10849 (N_10849,N_10703,N_10652);
or U10850 (N_10850,N_10772,N_10766);
and U10851 (N_10851,N_10785,N_10764);
nand U10852 (N_10852,N_10730,N_10657);
and U10853 (N_10853,N_10661,N_10654);
nand U10854 (N_10854,N_10669,N_10675);
or U10855 (N_10855,N_10790,N_10660);
nor U10856 (N_10856,N_10704,N_10769);
or U10857 (N_10857,N_10788,N_10753);
nor U10858 (N_10858,N_10727,N_10760);
nand U10859 (N_10859,N_10690,N_10715);
or U10860 (N_10860,N_10684,N_10798);
or U10861 (N_10861,N_10732,N_10674);
nand U10862 (N_10862,N_10774,N_10726);
nor U10863 (N_10863,N_10759,N_10695);
nand U10864 (N_10864,N_10700,N_10777);
nand U10865 (N_10865,N_10741,N_10676);
and U10866 (N_10866,N_10757,N_10771);
nand U10867 (N_10867,N_10710,N_10793);
or U10868 (N_10868,N_10680,N_10745);
and U10869 (N_10869,N_10733,N_10687);
nand U10870 (N_10870,N_10658,N_10748);
xor U10871 (N_10871,N_10739,N_10783);
xnor U10872 (N_10872,N_10781,N_10701);
nor U10873 (N_10873,N_10776,N_10705);
nor U10874 (N_10874,N_10665,N_10693);
or U10875 (N_10875,N_10672,N_10775);
xnor U10876 (N_10876,N_10743,N_10667);
nor U10877 (N_10877,N_10790,N_10733);
xnor U10878 (N_10878,N_10797,N_10796);
nand U10879 (N_10879,N_10707,N_10663);
xnor U10880 (N_10880,N_10678,N_10797);
nand U10881 (N_10881,N_10701,N_10798);
xor U10882 (N_10882,N_10732,N_10686);
nand U10883 (N_10883,N_10701,N_10795);
and U10884 (N_10884,N_10654,N_10702);
or U10885 (N_10885,N_10731,N_10654);
or U10886 (N_10886,N_10668,N_10697);
and U10887 (N_10887,N_10722,N_10753);
xnor U10888 (N_10888,N_10701,N_10664);
or U10889 (N_10889,N_10793,N_10707);
and U10890 (N_10890,N_10763,N_10773);
nor U10891 (N_10891,N_10693,N_10750);
nand U10892 (N_10892,N_10706,N_10670);
or U10893 (N_10893,N_10661,N_10752);
xor U10894 (N_10894,N_10656,N_10736);
xor U10895 (N_10895,N_10781,N_10754);
xor U10896 (N_10896,N_10737,N_10681);
and U10897 (N_10897,N_10672,N_10703);
nand U10898 (N_10898,N_10739,N_10737);
or U10899 (N_10899,N_10668,N_10769);
xnor U10900 (N_10900,N_10794,N_10743);
or U10901 (N_10901,N_10659,N_10761);
xnor U10902 (N_10902,N_10761,N_10696);
or U10903 (N_10903,N_10774,N_10763);
and U10904 (N_10904,N_10652,N_10685);
or U10905 (N_10905,N_10779,N_10696);
and U10906 (N_10906,N_10655,N_10702);
nor U10907 (N_10907,N_10779,N_10772);
nor U10908 (N_10908,N_10796,N_10653);
nor U10909 (N_10909,N_10743,N_10727);
nand U10910 (N_10910,N_10794,N_10736);
or U10911 (N_10911,N_10793,N_10720);
or U10912 (N_10912,N_10744,N_10694);
nand U10913 (N_10913,N_10765,N_10688);
or U10914 (N_10914,N_10693,N_10748);
xor U10915 (N_10915,N_10663,N_10716);
and U10916 (N_10916,N_10732,N_10754);
and U10917 (N_10917,N_10704,N_10732);
and U10918 (N_10918,N_10776,N_10790);
xnor U10919 (N_10919,N_10730,N_10694);
xor U10920 (N_10920,N_10662,N_10793);
and U10921 (N_10921,N_10708,N_10766);
xnor U10922 (N_10922,N_10756,N_10746);
xnor U10923 (N_10923,N_10715,N_10726);
nor U10924 (N_10924,N_10672,N_10669);
nand U10925 (N_10925,N_10708,N_10785);
nand U10926 (N_10926,N_10764,N_10696);
xor U10927 (N_10927,N_10744,N_10670);
and U10928 (N_10928,N_10661,N_10737);
nor U10929 (N_10929,N_10723,N_10677);
nor U10930 (N_10930,N_10748,N_10768);
or U10931 (N_10931,N_10777,N_10753);
nor U10932 (N_10932,N_10716,N_10741);
xor U10933 (N_10933,N_10684,N_10704);
or U10934 (N_10934,N_10726,N_10745);
nand U10935 (N_10935,N_10719,N_10790);
nor U10936 (N_10936,N_10749,N_10796);
nand U10937 (N_10937,N_10681,N_10729);
nor U10938 (N_10938,N_10667,N_10710);
or U10939 (N_10939,N_10717,N_10689);
or U10940 (N_10940,N_10733,N_10650);
and U10941 (N_10941,N_10748,N_10696);
nand U10942 (N_10942,N_10704,N_10658);
or U10943 (N_10943,N_10750,N_10731);
nand U10944 (N_10944,N_10662,N_10721);
nor U10945 (N_10945,N_10681,N_10771);
nor U10946 (N_10946,N_10712,N_10711);
nor U10947 (N_10947,N_10695,N_10736);
or U10948 (N_10948,N_10771,N_10744);
xor U10949 (N_10949,N_10782,N_10721);
and U10950 (N_10950,N_10827,N_10826);
and U10951 (N_10951,N_10808,N_10840);
xnor U10952 (N_10952,N_10922,N_10888);
xor U10953 (N_10953,N_10835,N_10897);
nor U10954 (N_10954,N_10871,N_10830);
xnor U10955 (N_10955,N_10834,N_10884);
nand U10956 (N_10956,N_10866,N_10880);
xor U10957 (N_10957,N_10921,N_10806);
xor U10958 (N_10958,N_10890,N_10900);
xnor U10959 (N_10959,N_10839,N_10849);
nand U10960 (N_10960,N_10882,N_10885);
and U10961 (N_10961,N_10813,N_10899);
xnor U10962 (N_10962,N_10910,N_10877);
and U10963 (N_10963,N_10847,N_10829);
and U10964 (N_10964,N_10843,N_10929);
nor U10965 (N_10965,N_10824,N_10889);
nand U10966 (N_10966,N_10886,N_10821);
xor U10967 (N_10967,N_10935,N_10944);
and U10968 (N_10968,N_10836,N_10807);
xor U10969 (N_10969,N_10855,N_10859);
and U10970 (N_10970,N_10869,N_10862);
nand U10971 (N_10971,N_10918,N_10802);
or U10972 (N_10972,N_10924,N_10898);
and U10973 (N_10973,N_10915,N_10810);
nor U10974 (N_10974,N_10861,N_10865);
or U10975 (N_10975,N_10872,N_10928);
nand U10976 (N_10976,N_10833,N_10901);
nand U10977 (N_10977,N_10853,N_10914);
nor U10978 (N_10978,N_10870,N_10907);
nor U10979 (N_10979,N_10815,N_10819);
or U10980 (N_10980,N_10863,N_10904);
xor U10981 (N_10981,N_10868,N_10945);
nor U10982 (N_10982,N_10818,N_10800);
xor U10983 (N_10983,N_10801,N_10822);
xnor U10984 (N_10984,N_10892,N_10857);
and U10985 (N_10985,N_10947,N_10940);
nor U10986 (N_10986,N_10905,N_10903);
nand U10987 (N_10987,N_10939,N_10923);
nand U10988 (N_10988,N_10932,N_10842);
nor U10989 (N_10989,N_10906,N_10883);
nand U10990 (N_10990,N_10841,N_10876);
and U10991 (N_10991,N_10850,N_10858);
nor U10992 (N_10992,N_10874,N_10817);
and U10993 (N_10993,N_10948,N_10902);
nand U10994 (N_10994,N_10927,N_10887);
nand U10995 (N_10995,N_10933,N_10930);
or U10996 (N_10996,N_10891,N_10846);
nor U10997 (N_10997,N_10941,N_10912);
or U10998 (N_10998,N_10804,N_10828);
nand U10999 (N_10999,N_10943,N_10864);
and U11000 (N_11000,N_10832,N_10931);
and U11001 (N_11001,N_10820,N_10831);
nor U11002 (N_11002,N_10937,N_10925);
xnor U11003 (N_11003,N_10805,N_10875);
or U11004 (N_11004,N_10938,N_10934);
and U11005 (N_11005,N_10881,N_10844);
and U11006 (N_11006,N_10809,N_10845);
or U11007 (N_11007,N_10811,N_10867);
and U11008 (N_11008,N_10946,N_10926);
nor U11009 (N_11009,N_10949,N_10816);
nor U11010 (N_11010,N_10852,N_10856);
nor U11011 (N_11011,N_10854,N_10908);
or U11012 (N_11012,N_10936,N_10860);
nand U11013 (N_11013,N_10942,N_10838);
or U11014 (N_11014,N_10919,N_10837);
and U11015 (N_11015,N_10917,N_10916);
or U11016 (N_11016,N_10879,N_10896);
xnor U11017 (N_11017,N_10851,N_10920);
nand U11018 (N_11018,N_10913,N_10825);
nor U11019 (N_11019,N_10893,N_10823);
nor U11020 (N_11020,N_10873,N_10894);
nor U11021 (N_11021,N_10848,N_10911);
and U11022 (N_11022,N_10909,N_10814);
and U11023 (N_11023,N_10895,N_10812);
and U11024 (N_11024,N_10878,N_10803);
xnor U11025 (N_11025,N_10878,N_10949);
or U11026 (N_11026,N_10874,N_10847);
nor U11027 (N_11027,N_10932,N_10944);
nand U11028 (N_11028,N_10898,N_10834);
or U11029 (N_11029,N_10805,N_10913);
or U11030 (N_11030,N_10926,N_10845);
nor U11031 (N_11031,N_10814,N_10927);
xor U11032 (N_11032,N_10839,N_10887);
or U11033 (N_11033,N_10820,N_10930);
or U11034 (N_11034,N_10925,N_10874);
and U11035 (N_11035,N_10912,N_10934);
nor U11036 (N_11036,N_10851,N_10921);
or U11037 (N_11037,N_10908,N_10884);
nand U11038 (N_11038,N_10852,N_10864);
nand U11039 (N_11039,N_10931,N_10945);
and U11040 (N_11040,N_10850,N_10861);
nand U11041 (N_11041,N_10840,N_10903);
or U11042 (N_11042,N_10893,N_10947);
xnor U11043 (N_11043,N_10904,N_10919);
nor U11044 (N_11044,N_10899,N_10875);
nand U11045 (N_11045,N_10938,N_10931);
nor U11046 (N_11046,N_10880,N_10846);
and U11047 (N_11047,N_10900,N_10932);
or U11048 (N_11048,N_10932,N_10917);
xor U11049 (N_11049,N_10918,N_10908);
or U11050 (N_11050,N_10890,N_10940);
or U11051 (N_11051,N_10828,N_10807);
nor U11052 (N_11052,N_10890,N_10903);
nand U11053 (N_11053,N_10933,N_10818);
and U11054 (N_11054,N_10934,N_10821);
nor U11055 (N_11055,N_10943,N_10811);
and U11056 (N_11056,N_10821,N_10883);
or U11057 (N_11057,N_10926,N_10901);
and U11058 (N_11058,N_10909,N_10945);
nor U11059 (N_11059,N_10913,N_10921);
or U11060 (N_11060,N_10858,N_10938);
nand U11061 (N_11061,N_10874,N_10936);
and U11062 (N_11062,N_10929,N_10922);
or U11063 (N_11063,N_10847,N_10843);
or U11064 (N_11064,N_10903,N_10832);
nand U11065 (N_11065,N_10907,N_10890);
and U11066 (N_11066,N_10931,N_10923);
xnor U11067 (N_11067,N_10832,N_10932);
or U11068 (N_11068,N_10831,N_10814);
or U11069 (N_11069,N_10874,N_10944);
xnor U11070 (N_11070,N_10838,N_10880);
and U11071 (N_11071,N_10944,N_10820);
nand U11072 (N_11072,N_10815,N_10900);
or U11073 (N_11073,N_10800,N_10828);
or U11074 (N_11074,N_10900,N_10883);
nand U11075 (N_11075,N_10872,N_10828);
or U11076 (N_11076,N_10941,N_10837);
or U11077 (N_11077,N_10928,N_10800);
or U11078 (N_11078,N_10810,N_10830);
xor U11079 (N_11079,N_10818,N_10826);
or U11080 (N_11080,N_10882,N_10917);
nand U11081 (N_11081,N_10895,N_10902);
nand U11082 (N_11082,N_10832,N_10804);
nor U11083 (N_11083,N_10906,N_10826);
or U11084 (N_11084,N_10832,N_10901);
xnor U11085 (N_11085,N_10848,N_10925);
nand U11086 (N_11086,N_10843,N_10860);
or U11087 (N_11087,N_10935,N_10877);
nor U11088 (N_11088,N_10935,N_10868);
or U11089 (N_11089,N_10826,N_10832);
and U11090 (N_11090,N_10917,N_10809);
and U11091 (N_11091,N_10945,N_10827);
or U11092 (N_11092,N_10871,N_10806);
xnor U11093 (N_11093,N_10827,N_10936);
nand U11094 (N_11094,N_10906,N_10804);
and U11095 (N_11095,N_10817,N_10881);
and U11096 (N_11096,N_10923,N_10849);
and U11097 (N_11097,N_10918,N_10882);
or U11098 (N_11098,N_10889,N_10830);
nand U11099 (N_11099,N_10896,N_10876);
or U11100 (N_11100,N_11076,N_11034);
and U11101 (N_11101,N_10964,N_11029);
nand U11102 (N_11102,N_11097,N_11014);
xor U11103 (N_11103,N_11015,N_11046);
xor U11104 (N_11104,N_11004,N_11081);
or U11105 (N_11105,N_11016,N_10992);
nor U11106 (N_11106,N_11091,N_11098);
or U11107 (N_11107,N_10985,N_11033);
nand U11108 (N_11108,N_11042,N_11041);
or U11109 (N_11109,N_11008,N_10999);
xnor U11110 (N_11110,N_11073,N_11053);
xnor U11111 (N_11111,N_11071,N_11082);
and U11112 (N_11112,N_11013,N_11026);
xor U11113 (N_11113,N_11035,N_10995);
or U11114 (N_11114,N_11025,N_11017);
xnor U11115 (N_11115,N_10967,N_10953);
nand U11116 (N_11116,N_11020,N_10994);
xor U11117 (N_11117,N_11022,N_11010);
nor U11118 (N_11118,N_10971,N_11093);
nand U11119 (N_11119,N_11051,N_10974);
nand U11120 (N_11120,N_10965,N_11018);
nand U11121 (N_11121,N_10989,N_10952);
nor U11122 (N_11122,N_11024,N_11021);
and U11123 (N_11123,N_11011,N_11040);
or U11124 (N_11124,N_11000,N_10986);
xor U11125 (N_11125,N_10957,N_10960);
nand U11126 (N_11126,N_11087,N_11095);
nor U11127 (N_11127,N_11030,N_11031);
xor U11128 (N_11128,N_11055,N_11074);
nand U11129 (N_11129,N_11059,N_10990);
nand U11130 (N_11130,N_10972,N_11079);
xor U11131 (N_11131,N_10961,N_10956);
nand U11132 (N_11132,N_10978,N_10996);
nand U11133 (N_11133,N_10997,N_10977);
nor U11134 (N_11134,N_11047,N_11067);
and U11135 (N_11135,N_11088,N_11065);
or U11136 (N_11136,N_11089,N_11023);
and U11137 (N_11137,N_11039,N_11069);
and U11138 (N_11138,N_11058,N_11057);
and U11139 (N_11139,N_10991,N_10951);
and U11140 (N_11140,N_10988,N_10955);
and U11141 (N_11141,N_11019,N_11012);
and U11142 (N_11142,N_10973,N_11070);
nand U11143 (N_11143,N_10954,N_11045);
nand U11144 (N_11144,N_11077,N_11038);
or U11145 (N_11145,N_11092,N_10987);
or U11146 (N_11146,N_11099,N_10976);
or U11147 (N_11147,N_10969,N_11064);
xor U11148 (N_11148,N_10982,N_10984);
and U11149 (N_11149,N_11062,N_11009);
nand U11150 (N_11150,N_11007,N_11027);
nand U11151 (N_11151,N_10993,N_11060);
or U11152 (N_11152,N_11085,N_11003);
or U11153 (N_11153,N_11005,N_11090);
and U11154 (N_11154,N_10983,N_10979);
xnor U11155 (N_11155,N_11072,N_11037);
or U11156 (N_11156,N_11054,N_11043);
nor U11157 (N_11157,N_10959,N_11052);
nand U11158 (N_11158,N_10962,N_11056);
nor U11159 (N_11159,N_11078,N_11044);
or U11160 (N_11160,N_10998,N_10968);
nand U11161 (N_11161,N_10975,N_11083);
xor U11162 (N_11162,N_10958,N_11028);
and U11163 (N_11163,N_11061,N_10980);
xnor U11164 (N_11164,N_10981,N_11096);
and U11165 (N_11165,N_11066,N_11094);
nor U11166 (N_11166,N_11006,N_11049);
xnor U11167 (N_11167,N_10966,N_10963);
xnor U11168 (N_11168,N_11036,N_11032);
xnor U11169 (N_11169,N_11048,N_10950);
nand U11170 (N_11170,N_10970,N_11075);
or U11171 (N_11171,N_11050,N_11063);
xor U11172 (N_11172,N_11080,N_11086);
nor U11173 (N_11173,N_11084,N_11002);
and U11174 (N_11174,N_11068,N_11001);
xnor U11175 (N_11175,N_11078,N_11077);
nand U11176 (N_11176,N_11081,N_11096);
nor U11177 (N_11177,N_10984,N_11091);
or U11178 (N_11178,N_10987,N_10981);
nand U11179 (N_11179,N_10991,N_11040);
xor U11180 (N_11180,N_11098,N_10987);
nand U11181 (N_11181,N_11078,N_10962);
xnor U11182 (N_11182,N_11051,N_11018);
or U11183 (N_11183,N_11068,N_11040);
and U11184 (N_11184,N_11044,N_11003);
nor U11185 (N_11185,N_11050,N_11089);
and U11186 (N_11186,N_11034,N_11056);
nor U11187 (N_11187,N_11008,N_11073);
and U11188 (N_11188,N_11057,N_11013);
xnor U11189 (N_11189,N_11007,N_11044);
nand U11190 (N_11190,N_10969,N_11022);
xnor U11191 (N_11191,N_11041,N_11016);
nor U11192 (N_11192,N_11014,N_11019);
nor U11193 (N_11193,N_11078,N_11095);
and U11194 (N_11194,N_11051,N_11010);
xnor U11195 (N_11195,N_11010,N_11001);
nand U11196 (N_11196,N_11001,N_10962);
xor U11197 (N_11197,N_11003,N_10970);
and U11198 (N_11198,N_11072,N_11078);
or U11199 (N_11199,N_10996,N_11071);
or U11200 (N_11200,N_10984,N_11010);
nand U11201 (N_11201,N_10951,N_10980);
nand U11202 (N_11202,N_10986,N_10957);
xnor U11203 (N_11203,N_10957,N_11063);
nand U11204 (N_11204,N_11080,N_11091);
nor U11205 (N_11205,N_11005,N_10970);
nand U11206 (N_11206,N_11039,N_11038);
and U11207 (N_11207,N_10957,N_11090);
xnor U11208 (N_11208,N_11080,N_11075);
and U11209 (N_11209,N_11088,N_11056);
or U11210 (N_11210,N_10958,N_11076);
and U11211 (N_11211,N_11046,N_11055);
nand U11212 (N_11212,N_10988,N_10978);
or U11213 (N_11213,N_11099,N_11088);
nand U11214 (N_11214,N_11066,N_11039);
and U11215 (N_11215,N_11057,N_10991);
or U11216 (N_11216,N_10976,N_11090);
nand U11217 (N_11217,N_11006,N_11089);
and U11218 (N_11218,N_11086,N_11062);
nand U11219 (N_11219,N_11068,N_11034);
nor U11220 (N_11220,N_11023,N_11015);
or U11221 (N_11221,N_11020,N_11068);
nor U11222 (N_11222,N_11047,N_11040);
or U11223 (N_11223,N_11046,N_11093);
or U11224 (N_11224,N_11058,N_11027);
xor U11225 (N_11225,N_10961,N_11097);
and U11226 (N_11226,N_10977,N_10953);
xor U11227 (N_11227,N_11067,N_11092);
xor U11228 (N_11228,N_11070,N_10975);
or U11229 (N_11229,N_10997,N_11066);
or U11230 (N_11230,N_10997,N_11047);
xor U11231 (N_11231,N_11057,N_11014);
xnor U11232 (N_11232,N_11060,N_10974);
nand U11233 (N_11233,N_11053,N_11007);
nor U11234 (N_11234,N_11064,N_10994);
xor U11235 (N_11235,N_10997,N_10969);
nand U11236 (N_11236,N_11020,N_11024);
or U11237 (N_11237,N_11065,N_11083);
nand U11238 (N_11238,N_11039,N_11084);
xnor U11239 (N_11239,N_11078,N_11035);
and U11240 (N_11240,N_11042,N_10981);
nor U11241 (N_11241,N_10990,N_11015);
nand U11242 (N_11242,N_11029,N_11015);
or U11243 (N_11243,N_11003,N_11067);
nand U11244 (N_11244,N_10990,N_11008);
and U11245 (N_11245,N_10961,N_11028);
or U11246 (N_11246,N_11081,N_11019);
nand U11247 (N_11247,N_11089,N_11012);
nor U11248 (N_11248,N_10980,N_11005);
xnor U11249 (N_11249,N_11015,N_11054);
xor U11250 (N_11250,N_11218,N_11228);
xor U11251 (N_11251,N_11115,N_11199);
xnor U11252 (N_11252,N_11201,N_11108);
and U11253 (N_11253,N_11198,N_11157);
or U11254 (N_11254,N_11196,N_11154);
xor U11255 (N_11255,N_11131,N_11122);
and U11256 (N_11256,N_11224,N_11104);
or U11257 (N_11257,N_11112,N_11232);
nor U11258 (N_11258,N_11239,N_11103);
or U11259 (N_11259,N_11139,N_11133);
xor U11260 (N_11260,N_11185,N_11138);
and U11261 (N_11261,N_11181,N_11222);
nand U11262 (N_11262,N_11136,N_11163);
nand U11263 (N_11263,N_11164,N_11182);
nand U11264 (N_11264,N_11178,N_11145);
and U11265 (N_11265,N_11223,N_11177);
nor U11266 (N_11266,N_11137,N_11221);
nand U11267 (N_11267,N_11105,N_11100);
or U11268 (N_11268,N_11158,N_11226);
nor U11269 (N_11269,N_11188,N_11209);
xor U11270 (N_11270,N_11118,N_11202);
and U11271 (N_11271,N_11121,N_11244);
nand U11272 (N_11272,N_11146,N_11159);
nand U11273 (N_11273,N_11195,N_11143);
xor U11274 (N_11274,N_11134,N_11106);
and U11275 (N_11275,N_11109,N_11200);
nand U11276 (N_11276,N_11194,N_11243);
or U11277 (N_11277,N_11191,N_11160);
xnor U11278 (N_11278,N_11183,N_11124);
or U11279 (N_11279,N_11149,N_11208);
and U11280 (N_11280,N_11150,N_11231);
and U11281 (N_11281,N_11190,N_11207);
and U11282 (N_11282,N_11173,N_11176);
and U11283 (N_11283,N_11170,N_11229);
nor U11284 (N_11284,N_11249,N_11210);
xnor U11285 (N_11285,N_11135,N_11203);
nand U11286 (N_11286,N_11125,N_11197);
and U11287 (N_11287,N_11225,N_11107);
nor U11288 (N_11288,N_11171,N_11240);
nand U11289 (N_11289,N_11227,N_11237);
xnor U11290 (N_11290,N_11248,N_11175);
nor U11291 (N_11291,N_11230,N_11167);
or U11292 (N_11292,N_11241,N_11162);
or U11293 (N_11293,N_11238,N_11233);
and U11294 (N_11294,N_11142,N_11214);
nor U11295 (N_11295,N_11219,N_11102);
xor U11296 (N_11296,N_11111,N_11245);
or U11297 (N_11297,N_11168,N_11206);
nand U11298 (N_11298,N_11165,N_11130);
xor U11299 (N_11299,N_11161,N_11129);
or U11300 (N_11300,N_11235,N_11117);
or U11301 (N_11301,N_11216,N_11189);
nor U11302 (N_11302,N_11147,N_11152);
nor U11303 (N_11303,N_11242,N_11141);
xnor U11304 (N_11304,N_11110,N_11174);
nor U11305 (N_11305,N_11234,N_11128);
nand U11306 (N_11306,N_11236,N_11186);
or U11307 (N_11307,N_11155,N_11113);
nand U11308 (N_11308,N_11169,N_11184);
or U11309 (N_11309,N_11114,N_11192);
xnor U11310 (N_11310,N_11247,N_11215);
and U11311 (N_11311,N_11156,N_11120);
xor U11312 (N_11312,N_11153,N_11151);
xnor U11313 (N_11313,N_11213,N_11132);
nor U11314 (N_11314,N_11123,N_11205);
or U11315 (N_11315,N_11211,N_11172);
nand U11316 (N_11316,N_11144,N_11140);
and U11317 (N_11317,N_11193,N_11166);
or U11318 (N_11318,N_11217,N_11179);
nand U11319 (N_11319,N_11119,N_11116);
xor U11320 (N_11320,N_11204,N_11126);
nor U11321 (N_11321,N_11180,N_11127);
nor U11322 (N_11322,N_11187,N_11101);
nor U11323 (N_11323,N_11212,N_11220);
xor U11324 (N_11324,N_11246,N_11148);
nor U11325 (N_11325,N_11121,N_11103);
nor U11326 (N_11326,N_11242,N_11136);
nand U11327 (N_11327,N_11162,N_11170);
nand U11328 (N_11328,N_11129,N_11186);
xnor U11329 (N_11329,N_11239,N_11245);
and U11330 (N_11330,N_11115,N_11238);
or U11331 (N_11331,N_11199,N_11150);
nor U11332 (N_11332,N_11156,N_11105);
nor U11333 (N_11333,N_11171,N_11243);
and U11334 (N_11334,N_11247,N_11222);
nor U11335 (N_11335,N_11100,N_11190);
nand U11336 (N_11336,N_11178,N_11113);
xnor U11337 (N_11337,N_11141,N_11144);
nor U11338 (N_11338,N_11246,N_11108);
xnor U11339 (N_11339,N_11209,N_11201);
nand U11340 (N_11340,N_11187,N_11154);
and U11341 (N_11341,N_11160,N_11243);
or U11342 (N_11342,N_11206,N_11120);
xnor U11343 (N_11343,N_11205,N_11162);
and U11344 (N_11344,N_11137,N_11160);
nor U11345 (N_11345,N_11177,N_11129);
or U11346 (N_11346,N_11234,N_11197);
and U11347 (N_11347,N_11188,N_11201);
xnor U11348 (N_11348,N_11227,N_11112);
and U11349 (N_11349,N_11149,N_11190);
or U11350 (N_11350,N_11140,N_11220);
xor U11351 (N_11351,N_11216,N_11246);
nand U11352 (N_11352,N_11105,N_11235);
or U11353 (N_11353,N_11158,N_11171);
nand U11354 (N_11354,N_11215,N_11224);
and U11355 (N_11355,N_11109,N_11233);
or U11356 (N_11356,N_11196,N_11167);
nor U11357 (N_11357,N_11103,N_11129);
and U11358 (N_11358,N_11130,N_11198);
xnor U11359 (N_11359,N_11146,N_11247);
xor U11360 (N_11360,N_11165,N_11205);
and U11361 (N_11361,N_11106,N_11219);
nand U11362 (N_11362,N_11111,N_11143);
and U11363 (N_11363,N_11179,N_11140);
nand U11364 (N_11364,N_11164,N_11214);
or U11365 (N_11365,N_11125,N_11101);
nor U11366 (N_11366,N_11106,N_11177);
nand U11367 (N_11367,N_11179,N_11184);
nand U11368 (N_11368,N_11227,N_11129);
or U11369 (N_11369,N_11204,N_11158);
or U11370 (N_11370,N_11142,N_11115);
nand U11371 (N_11371,N_11123,N_11214);
nand U11372 (N_11372,N_11222,N_11183);
nor U11373 (N_11373,N_11219,N_11119);
or U11374 (N_11374,N_11193,N_11142);
or U11375 (N_11375,N_11153,N_11207);
and U11376 (N_11376,N_11108,N_11142);
nand U11377 (N_11377,N_11140,N_11142);
nor U11378 (N_11378,N_11193,N_11245);
and U11379 (N_11379,N_11218,N_11124);
or U11380 (N_11380,N_11148,N_11243);
xor U11381 (N_11381,N_11126,N_11246);
or U11382 (N_11382,N_11211,N_11231);
xor U11383 (N_11383,N_11145,N_11114);
nor U11384 (N_11384,N_11172,N_11150);
xor U11385 (N_11385,N_11202,N_11141);
and U11386 (N_11386,N_11132,N_11166);
xnor U11387 (N_11387,N_11158,N_11183);
xnor U11388 (N_11388,N_11123,N_11126);
and U11389 (N_11389,N_11196,N_11143);
nand U11390 (N_11390,N_11240,N_11153);
or U11391 (N_11391,N_11102,N_11135);
nand U11392 (N_11392,N_11228,N_11244);
xor U11393 (N_11393,N_11134,N_11244);
or U11394 (N_11394,N_11124,N_11171);
nor U11395 (N_11395,N_11194,N_11246);
nor U11396 (N_11396,N_11156,N_11113);
and U11397 (N_11397,N_11247,N_11156);
nor U11398 (N_11398,N_11125,N_11182);
nor U11399 (N_11399,N_11225,N_11116);
and U11400 (N_11400,N_11295,N_11359);
and U11401 (N_11401,N_11390,N_11259);
nand U11402 (N_11402,N_11364,N_11363);
xnor U11403 (N_11403,N_11285,N_11288);
xor U11404 (N_11404,N_11383,N_11251);
or U11405 (N_11405,N_11371,N_11277);
or U11406 (N_11406,N_11339,N_11312);
and U11407 (N_11407,N_11276,N_11348);
xor U11408 (N_11408,N_11310,N_11264);
and U11409 (N_11409,N_11340,N_11337);
and U11410 (N_11410,N_11283,N_11303);
or U11411 (N_11411,N_11279,N_11373);
nand U11412 (N_11412,N_11356,N_11378);
or U11413 (N_11413,N_11326,N_11381);
nand U11414 (N_11414,N_11270,N_11307);
and U11415 (N_11415,N_11389,N_11306);
xor U11416 (N_11416,N_11395,N_11369);
or U11417 (N_11417,N_11281,N_11282);
nor U11418 (N_11418,N_11380,N_11302);
nor U11419 (N_11419,N_11260,N_11304);
nor U11420 (N_11420,N_11316,N_11372);
or U11421 (N_11421,N_11313,N_11322);
and U11422 (N_11422,N_11323,N_11328);
xor U11423 (N_11423,N_11366,N_11342);
nand U11424 (N_11424,N_11387,N_11351);
or U11425 (N_11425,N_11346,N_11257);
nor U11426 (N_11426,N_11382,N_11355);
nor U11427 (N_11427,N_11334,N_11278);
and U11428 (N_11428,N_11273,N_11375);
nor U11429 (N_11429,N_11286,N_11290);
nor U11430 (N_11430,N_11358,N_11311);
xnor U11431 (N_11431,N_11338,N_11268);
and U11432 (N_11432,N_11396,N_11391);
nand U11433 (N_11433,N_11350,N_11393);
nor U11434 (N_11434,N_11319,N_11291);
nor U11435 (N_11435,N_11284,N_11333);
nor U11436 (N_11436,N_11332,N_11392);
and U11437 (N_11437,N_11292,N_11398);
or U11438 (N_11438,N_11388,N_11309);
or U11439 (N_11439,N_11379,N_11308);
and U11440 (N_11440,N_11327,N_11377);
or U11441 (N_11441,N_11343,N_11321);
nand U11442 (N_11442,N_11258,N_11301);
and U11443 (N_11443,N_11280,N_11266);
or U11444 (N_11444,N_11275,N_11265);
xor U11445 (N_11445,N_11385,N_11252);
and U11446 (N_11446,N_11324,N_11360);
nor U11447 (N_11447,N_11330,N_11271);
or U11448 (N_11448,N_11294,N_11354);
nand U11449 (N_11449,N_11329,N_11298);
or U11450 (N_11450,N_11344,N_11386);
xor U11451 (N_11451,N_11345,N_11255);
nor U11452 (N_11452,N_11315,N_11331);
nor U11453 (N_11453,N_11297,N_11341);
and U11454 (N_11454,N_11335,N_11370);
and U11455 (N_11455,N_11293,N_11254);
xnor U11456 (N_11456,N_11325,N_11274);
or U11457 (N_11457,N_11374,N_11394);
or U11458 (N_11458,N_11314,N_11317);
xnor U11459 (N_11459,N_11361,N_11368);
nor U11460 (N_11460,N_11376,N_11253);
or U11461 (N_11461,N_11287,N_11256);
and U11462 (N_11462,N_11399,N_11289);
xnor U11463 (N_11463,N_11262,N_11299);
nor U11464 (N_11464,N_11261,N_11353);
nand U11465 (N_11465,N_11263,N_11362);
nor U11466 (N_11466,N_11357,N_11272);
xor U11467 (N_11467,N_11318,N_11397);
xor U11468 (N_11468,N_11352,N_11367);
xnor U11469 (N_11469,N_11250,N_11300);
xor U11470 (N_11470,N_11347,N_11349);
nor U11471 (N_11471,N_11305,N_11269);
nor U11472 (N_11472,N_11296,N_11267);
xor U11473 (N_11473,N_11365,N_11384);
nor U11474 (N_11474,N_11336,N_11320);
xnor U11475 (N_11475,N_11351,N_11344);
nand U11476 (N_11476,N_11398,N_11281);
xnor U11477 (N_11477,N_11259,N_11286);
and U11478 (N_11478,N_11363,N_11376);
xor U11479 (N_11479,N_11274,N_11397);
xor U11480 (N_11480,N_11385,N_11357);
xor U11481 (N_11481,N_11364,N_11382);
and U11482 (N_11482,N_11269,N_11349);
or U11483 (N_11483,N_11361,N_11280);
nand U11484 (N_11484,N_11266,N_11366);
xnor U11485 (N_11485,N_11385,N_11381);
or U11486 (N_11486,N_11331,N_11318);
or U11487 (N_11487,N_11371,N_11384);
or U11488 (N_11488,N_11382,N_11387);
nand U11489 (N_11489,N_11320,N_11377);
xor U11490 (N_11490,N_11257,N_11263);
or U11491 (N_11491,N_11341,N_11251);
nor U11492 (N_11492,N_11379,N_11280);
nand U11493 (N_11493,N_11308,N_11385);
xor U11494 (N_11494,N_11291,N_11356);
xnor U11495 (N_11495,N_11325,N_11379);
xnor U11496 (N_11496,N_11278,N_11291);
nor U11497 (N_11497,N_11284,N_11339);
xnor U11498 (N_11498,N_11308,N_11392);
and U11499 (N_11499,N_11271,N_11290);
nor U11500 (N_11500,N_11299,N_11328);
and U11501 (N_11501,N_11354,N_11385);
or U11502 (N_11502,N_11336,N_11345);
nor U11503 (N_11503,N_11254,N_11378);
nor U11504 (N_11504,N_11271,N_11259);
and U11505 (N_11505,N_11342,N_11311);
nor U11506 (N_11506,N_11327,N_11360);
or U11507 (N_11507,N_11355,N_11359);
or U11508 (N_11508,N_11388,N_11354);
nor U11509 (N_11509,N_11365,N_11393);
nand U11510 (N_11510,N_11389,N_11332);
or U11511 (N_11511,N_11355,N_11366);
nand U11512 (N_11512,N_11358,N_11296);
and U11513 (N_11513,N_11391,N_11336);
or U11514 (N_11514,N_11384,N_11392);
xnor U11515 (N_11515,N_11299,N_11327);
and U11516 (N_11516,N_11257,N_11289);
or U11517 (N_11517,N_11272,N_11348);
nand U11518 (N_11518,N_11302,N_11288);
xor U11519 (N_11519,N_11276,N_11320);
nor U11520 (N_11520,N_11329,N_11312);
nor U11521 (N_11521,N_11305,N_11260);
nand U11522 (N_11522,N_11272,N_11337);
and U11523 (N_11523,N_11274,N_11254);
nor U11524 (N_11524,N_11251,N_11332);
or U11525 (N_11525,N_11258,N_11383);
or U11526 (N_11526,N_11339,N_11332);
xor U11527 (N_11527,N_11341,N_11354);
or U11528 (N_11528,N_11348,N_11354);
nor U11529 (N_11529,N_11373,N_11337);
and U11530 (N_11530,N_11343,N_11347);
xnor U11531 (N_11531,N_11369,N_11254);
or U11532 (N_11532,N_11355,N_11348);
nand U11533 (N_11533,N_11378,N_11342);
nand U11534 (N_11534,N_11397,N_11264);
and U11535 (N_11535,N_11280,N_11343);
nand U11536 (N_11536,N_11361,N_11279);
nand U11537 (N_11537,N_11382,N_11294);
nor U11538 (N_11538,N_11373,N_11372);
nand U11539 (N_11539,N_11386,N_11352);
nand U11540 (N_11540,N_11304,N_11379);
or U11541 (N_11541,N_11313,N_11319);
or U11542 (N_11542,N_11255,N_11348);
xnor U11543 (N_11543,N_11263,N_11258);
and U11544 (N_11544,N_11315,N_11339);
and U11545 (N_11545,N_11279,N_11308);
or U11546 (N_11546,N_11398,N_11348);
and U11547 (N_11547,N_11312,N_11364);
and U11548 (N_11548,N_11380,N_11326);
or U11549 (N_11549,N_11399,N_11311);
nand U11550 (N_11550,N_11476,N_11520);
or U11551 (N_11551,N_11452,N_11437);
xnor U11552 (N_11552,N_11433,N_11513);
nor U11553 (N_11553,N_11465,N_11500);
nor U11554 (N_11554,N_11431,N_11538);
xor U11555 (N_11555,N_11470,N_11473);
nor U11556 (N_11556,N_11480,N_11472);
or U11557 (N_11557,N_11469,N_11421);
or U11558 (N_11558,N_11474,N_11406);
and U11559 (N_11559,N_11468,N_11478);
nor U11560 (N_11560,N_11403,N_11549);
nand U11561 (N_11561,N_11455,N_11507);
and U11562 (N_11562,N_11442,N_11453);
and U11563 (N_11563,N_11541,N_11435);
nand U11564 (N_11564,N_11451,N_11488);
and U11565 (N_11565,N_11492,N_11545);
nand U11566 (N_11566,N_11425,N_11511);
nor U11567 (N_11567,N_11445,N_11432);
xnor U11568 (N_11568,N_11461,N_11544);
nand U11569 (N_11569,N_11439,N_11503);
nor U11570 (N_11570,N_11547,N_11493);
and U11571 (N_11571,N_11510,N_11517);
nor U11572 (N_11572,N_11426,N_11419);
nor U11573 (N_11573,N_11423,N_11477);
or U11574 (N_11574,N_11402,N_11463);
nand U11575 (N_11575,N_11514,N_11416);
xor U11576 (N_11576,N_11498,N_11515);
nor U11577 (N_11577,N_11428,N_11429);
and U11578 (N_11578,N_11494,N_11519);
nor U11579 (N_11579,N_11530,N_11524);
nor U11580 (N_11580,N_11427,N_11489);
nand U11581 (N_11581,N_11518,N_11546);
xnor U11582 (N_11582,N_11438,N_11504);
or U11583 (N_11583,N_11525,N_11440);
or U11584 (N_11584,N_11490,N_11516);
nand U11585 (N_11585,N_11505,N_11526);
or U11586 (N_11586,N_11506,N_11449);
nand U11587 (N_11587,N_11482,N_11412);
nand U11588 (N_11588,N_11537,N_11418);
xnor U11589 (N_11589,N_11434,N_11430);
nand U11590 (N_11590,N_11415,N_11499);
and U11591 (N_11591,N_11496,N_11441);
and U11592 (N_11592,N_11481,N_11529);
or U11593 (N_11593,N_11467,N_11475);
and U11594 (N_11594,N_11527,N_11422);
and U11595 (N_11595,N_11409,N_11533);
nand U11596 (N_11596,N_11497,N_11444);
or U11597 (N_11597,N_11456,N_11491);
nand U11598 (N_11598,N_11443,N_11531);
nor U11599 (N_11599,N_11466,N_11447);
and U11600 (N_11600,N_11414,N_11548);
or U11601 (N_11601,N_11407,N_11532);
nor U11602 (N_11602,N_11509,N_11522);
or U11603 (N_11603,N_11471,N_11408);
and U11604 (N_11604,N_11436,N_11521);
nand U11605 (N_11605,N_11424,N_11523);
and U11606 (N_11606,N_11457,N_11536);
or U11607 (N_11607,N_11512,N_11485);
nand U11608 (N_11608,N_11405,N_11450);
xor U11609 (N_11609,N_11417,N_11454);
xor U11610 (N_11610,N_11486,N_11535);
or U11611 (N_11611,N_11534,N_11410);
and U11612 (N_11612,N_11479,N_11459);
xnor U11613 (N_11613,N_11464,N_11400);
nand U11614 (N_11614,N_11411,N_11404);
nor U11615 (N_11615,N_11542,N_11462);
nor U11616 (N_11616,N_11413,N_11528);
and U11617 (N_11617,N_11540,N_11501);
nor U11618 (N_11618,N_11458,N_11539);
xnor U11619 (N_11619,N_11483,N_11448);
xor U11620 (N_11620,N_11420,N_11446);
xnor U11621 (N_11621,N_11460,N_11487);
xnor U11622 (N_11622,N_11401,N_11502);
or U11623 (N_11623,N_11495,N_11543);
nor U11624 (N_11624,N_11484,N_11508);
nand U11625 (N_11625,N_11423,N_11470);
nand U11626 (N_11626,N_11462,N_11504);
nand U11627 (N_11627,N_11486,N_11529);
xnor U11628 (N_11628,N_11530,N_11427);
xnor U11629 (N_11629,N_11501,N_11479);
xnor U11630 (N_11630,N_11523,N_11529);
or U11631 (N_11631,N_11518,N_11500);
xnor U11632 (N_11632,N_11491,N_11477);
and U11633 (N_11633,N_11428,N_11520);
nor U11634 (N_11634,N_11540,N_11471);
nor U11635 (N_11635,N_11490,N_11548);
xor U11636 (N_11636,N_11499,N_11543);
and U11637 (N_11637,N_11482,N_11522);
or U11638 (N_11638,N_11471,N_11443);
nor U11639 (N_11639,N_11521,N_11419);
xor U11640 (N_11640,N_11490,N_11466);
or U11641 (N_11641,N_11476,N_11430);
nand U11642 (N_11642,N_11455,N_11514);
and U11643 (N_11643,N_11453,N_11448);
or U11644 (N_11644,N_11481,N_11425);
xor U11645 (N_11645,N_11533,N_11412);
nand U11646 (N_11646,N_11549,N_11488);
and U11647 (N_11647,N_11431,N_11412);
and U11648 (N_11648,N_11548,N_11435);
nand U11649 (N_11649,N_11474,N_11481);
and U11650 (N_11650,N_11414,N_11426);
xnor U11651 (N_11651,N_11451,N_11535);
and U11652 (N_11652,N_11481,N_11542);
or U11653 (N_11653,N_11411,N_11519);
or U11654 (N_11654,N_11470,N_11524);
nand U11655 (N_11655,N_11438,N_11496);
or U11656 (N_11656,N_11533,N_11516);
and U11657 (N_11657,N_11417,N_11428);
or U11658 (N_11658,N_11476,N_11490);
nor U11659 (N_11659,N_11528,N_11478);
nand U11660 (N_11660,N_11492,N_11424);
or U11661 (N_11661,N_11400,N_11449);
xnor U11662 (N_11662,N_11498,N_11466);
and U11663 (N_11663,N_11457,N_11472);
nand U11664 (N_11664,N_11433,N_11518);
nand U11665 (N_11665,N_11469,N_11459);
xor U11666 (N_11666,N_11411,N_11505);
nand U11667 (N_11667,N_11410,N_11474);
xnor U11668 (N_11668,N_11451,N_11507);
nand U11669 (N_11669,N_11430,N_11420);
and U11670 (N_11670,N_11511,N_11483);
nor U11671 (N_11671,N_11411,N_11522);
xnor U11672 (N_11672,N_11423,N_11400);
nand U11673 (N_11673,N_11414,N_11481);
nor U11674 (N_11674,N_11415,N_11437);
and U11675 (N_11675,N_11505,N_11496);
or U11676 (N_11676,N_11530,N_11509);
nand U11677 (N_11677,N_11540,N_11449);
nor U11678 (N_11678,N_11473,N_11508);
or U11679 (N_11679,N_11524,N_11413);
nor U11680 (N_11680,N_11461,N_11501);
xnor U11681 (N_11681,N_11512,N_11414);
nor U11682 (N_11682,N_11462,N_11545);
nor U11683 (N_11683,N_11526,N_11473);
nor U11684 (N_11684,N_11441,N_11543);
nand U11685 (N_11685,N_11544,N_11522);
or U11686 (N_11686,N_11409,N_11541);
nand U11687 (N_11687,N_11493,N_11548);
nand U11688 (N_11688,N_11449,N_11493);
or U11689 (N_11689,N_11509,N_11440);
and U11690 (N_11690,N_11465,N_11459);
or U11691 (N_11691,N_11488,N_11415);
nand U11692 (N_11692,N_11470,N_11498);
or U11693 (N_11693,N_11532,N_11516);
or U11694 (N_11694,N_11458,N_11517);
nor U11695 (N_11695,N_11451,N_11410);
xnor U11696 (N_11696,N_11438,N_11549);
or U11697 (N_11697,N_11538,N_11518);
nand U11698 (N_11698,N_11513,N_11468);
xor U11699 (N_11699,N_11474,N_11507);
nor U11700 (N_11700,N_11587,N_11589);
and U11701 (N_11701,N_11657,N_11683);
xnor U11702 (N_11702,N_11573,N_11583);
and U11703 (N_11703,N_11682,N_11640);
or U11704 (N_11704,N_11679,N_11699);
or U11705 (N_11705,N_11665,N_11588);
nand U11706 (N_11706,N_11580,N_11693);
xor U11707 (N_11707,N_11664,N_11570);
or U11708 (N_11708,N_11565,N_11610);
and U11709 (N_11709,N_11681,N_11658);
and U11710 (N_11710,N_11666,N_11619);
nor U11711 (N_11711,N_11590,N_11551);
xor U11712 (N_11712,N_11661,N_11611);
nand U11713 (N_11713,N_11566,N_11642);
xnor U11714 (N_11714,N_11595,N_11596);
or U11715 (N_11715,N_11585,N_11689);
nand U11716 (N_11716,N_11564,N_11639);
and U11717 (N_11717,N_11614,N_11698);
xnor U11718 (N_11718,N_11560,N_11626);
nand U11719 (N_11719,N_11674,N_11647);
xor U11720 (N_11720,N_11687,N_11623);
and U11721 (N_11721,N_11678,N_11603);
nor U11722 (N_11722,N_11627,N_11609);
xnor U11723 (N_11723,N_11591,N_11569);
or U11724 (N_11724,N_11575,N_11620);
nand U11725 (N_11725,N_11659,N_11651);
or U11726 (N_11726,N_11593,N_11646);
and U11727 (N_11727,N_11633,N_11557);
or U11728 (N_11728,N_11568,N_11671);
nor U11729 (N_11729,N_11638,N_11582);
nand U11730 (N_11730,N_11691,N_11550);
nand U11731 (N_11731,N_11552,N_11694);
and U11732 (N_11732,N_11652,N_11600);
or U11733 (N_11733,N_11581,N_11655);
nand U11734 (N_11734,N_11562,N_11601);
or U11735 (N_11735,N_11645,N_11654);
xnor U11736 (N_11736,N_11697,N_11602);
and U11737 (N_11737,N_11672,N_11685);
xnor U11738 (N_11738,N_11634,N_11668);
nand U11739 (N_11739,N_11670,N_11606);
or U11740 (N_11740,N_11692,N_11649);
nand U11741 (N_11741,N_11598,N_11690);
or U11742 (N_11742,N_11644,N_11650);
nor U11743 (N_11743,N_11599,N_11635);
and U11744 (N_11744,N_11621,N_11555);
and U11745 (N_11745,N_11622,N_11636);
nor U11746 (N_11746,N_11612,N_11577);
nand U11747 (N_11747,N_11574,N_11629);
nand U11748 (N_11748,N_11616,N_11696);
xnor U11749 (N_11749,N_11567,N_11662);
xor U11750 (N_11750,N_11680,N_11641);
nand U11751 (N_11751,N_11558,N_11604);
nor U11752 (N_11752,N_11556,N_11563);
nand U11753 (N_11753,N_11667,N_11676);
or U11754 (N_11754,N_11615,N_11617);
nor U11755 (N_11755,N_11624,N_11684);
xor U11756 (N_11756,N_11628,N_11686);
nor U11757 (N_11757,N_11632,N_11561);
and U11758 (N_11758,N_11576,N_11571);
xnor U11759 (N_11759,N_11688,N_11653);
or U11760 (N_11760,N_11656,N_11607);
nor U11761 (N_11761,N_11637,N_11618);
xnor U11762 (N_11762,N_11608,N_11631);
nand U11763 (N_11763,N_11554,N_11584);
xor U11764 (N_11764,N_11592,N_11578);
or U11765 (N_11765,N_11553,N_11648);
or U11766 (N_11766,N_11605,N_11660);
nand U11767 (N_11767,N_11630,N_11677);
nor U11768 (N_11768,N_11586,N_11579);
and U11769 (N_11769,N_11594,N_11663);
or U11770 (N_11770,N_11675,N_11625);
and U11771 (N_11771,N_11669,N_11643);
xor U11772 (N_11772,N_11572,N_11559);
and U11773 (N_11773,N_11613,N_11597);
nor U11774 (N_11774,N_11695,N_11673);
or U11775 (N_11775,N_11639,N_11642);
and U11776 (N_11776,N_11678,N_11628);
nor U11777 (N_11777,N_11569,N_11578);
nor U11778 (N_11778,N_11630,N_11563);
nand U11779 (N_11779,N_11570,N_11673);
and U11780 (N_11780,N_11570,N_11582);
xor U11781 (N_11781,N_11695,N_11647);
nand U11782 (N_11782,N_11584,N_11616);
or U11783 (N_11783,N_11619,N_11553);
xor U11784 (N_11784,N_11631,N_11636);
xnor U11785 (N_11785,N_11604,N_11689);
nand U11786 (N_11786,N_11627,N_11690);
nor U11787 (N_11787,N_11642,N_11603);
nand U11788 (N_11788,N_11645,N_11627);
nor U11789 (N_11789,N_11571,N_11607);
nand U11790 (N_11790,N_11653,N_11697);
nand U11791 (N_11791,N_11658,N_11624);
and U11792 (N_11792,N_11679,N_11556);
nor U11793 (N_11793,N_11578,N_11590);
xnor U11794 (N_11794,N_11661,N_11646);
nand U11795 (N_11795,N_11599,N_11628);
nand U11796 (N_11796,N_11597,N_11636);
and U11797 (N_11797,N_11647,N_11639);
and U11798 (N_11798,N_11689,N_11652);
xnor U11799 (N_11799,N_11648,N_11685);
or U11800 (N_11800,N_11574,N_11572);
nor U11801 (N_11801,N_11642,N_11626);
or U11802 (N_11802,N_11593,N_11604);
nand U11803 (N_11803,N_11588,N_11650);
nor U11804 (N_11804,N_11552,N_11605);
xor U11805 (N_11805,N_11665,N_11603);
nand U11806 (N_11806,N_11693,N_11665);
xnor U11807 (N_11807,N_11570,N_11647);
and U11808 (N_11808,N_11693,N_11647);
or U11809 (N_11809,N_11592,N_11608);
and U11810 (N_11810,N_11639,N_11699);
and U11811 (N_11811,N_11580,N_11665);
nand U11812 (N_11812,N_11625,N_11591);
and U11813 (N_11813,N_11655,N_11651);
nor U11814 (N_11814,N_11553,N_11650);
nand U11815 (N_11815,N_11631,N_11607);
nor U11816 (N_11816,N_11681,N_11613);
or U11817 (N_11817,N_11628,N_11630);
or U11818 (N_11818,N_11664,N_11680);
nor U11819 (N_11819,N_11600,N_11683);
nor U11820 (N_11820,N_11554,N_11553);
xnor U11821 (N_11821,N_11697,N_11652);
nand U11822 (N_11822,N_11698,N_11653);
or U11823 (N_11823,N_11607,N_11646);
xnor U11824 (N_11824,N_11607,N_11694);
nand U11825 (N_11825,N_11550,N_11588);
and U11826 (N_11826,N_11587,N_11568);
nand U11827 (N_11827,N_11666,N_11557);
and U11828 (N_11828,N_11690,N_11619);
xnor U11829 (N_11829,N_11578,N_11691);
nor U11830 (N_11830,N_11650,N_11591);
and U11831 (N_11831,N_11577,N_11625);
nor U11832 (N_11832,N_11680,N_11578);
nand U11833 (N_11833,N_11611,N_11658);
xor U11834 (N_11834,N_11646,N_11589);
nand U11835 (N_11835,N_11589,N_11631);
nor U11836 (N_11836,N_11662,N_11592);
xnor U11837 (N_11837,N_11602,N_11630);
nor U11838 (N_11838,N_11646,N_11615);
and U11839 (N_11839,N_11578,N_11642);
xor U11840 (N_11840,N_11698,N_11599);
and U11841 (N_11841,N_11661,N_11636);
and U11842 (N_11842,N_11608,N_11629);
xnor U11843 (N_11843,N_11692,N_11628);
and U11844 (N_11844,N_11585,N_11611);
nand U11845 (N_11845,N_11615,N_11699);
and U11846 (N_11846,N_11645,N_11691);
and U11847 (N_11847,N_11693,N_11652);
nor U11848 (N_11848,N_11621,N_11617);
or U11849 (N_11849,N_11581,N_11592);
nor U11850 (N_11850,N_11804,N_11722);
and U11851 (N_11851,N_11737,N_11824);
and U11852 (N_11852,N_11814,N_11718);
or U11853 (N_11853,N_11759,N_11750);
and U11854 (N_11854,N_11786,N_11790);
nor U11855 (N_11855,N_11729,N_11841);
and U11856 (N_11856,N_11735,N_11740);
nand U11857 (N_11857,N_11796,N_11741);
or U11858 (N_11858,N_11721,N_11709);
xor U11859 (N_11859,N_11716,N_11736);
and U11860 (N_11860,N_11708,N_11762);
nor U11861 (N_11861,N_11701,N_11845);
and U11862 (N_11862,N_11755,N_11705);
xnor U11863 (N_11863,N_11800,N_11816);
and U11864 (N_11864,N_11840,N_11732);
or U11865 (N_11865,N_11767,N_11739);
nor U11866 (N_11866,N_11756,N_11712);
nor U11867 (N_11867,N_11760,N_11807);
xor U11868 (N_11868,N_11711,N_11748);
nor U11869 (N_11869,N_11823,N_11768);
nor U11870 (N_11870,N_11838,N_11725);
nand U11871 (N_11871,N_11733,N_11742);
nand U11872 (N_11872,N_11714,N_11749);
and U11873 (N_11873,N_11717,N_11842);
xor U11874 (N_11874,N_11761,N_11743);
nor U11875 (N_11875,N_11757,N_11764);
nand U11876 (N_11876,N_11753,N_11747);
nand U11877 (N_11877,N_11795,N_11789);
and U11878 (N_11878,N_11802,N_11798);
and U11879 (N_11879,N_11815,N_11769);
xnor U11880 (N_11880,N_11829,N_11746);
xor U11881 (N_11881,N_11730,N_11781);
nand U11882 (N_11882,N_11833,N_11754);
xor U11883 (N_11883,N_11763,N_11834);
and U11884 (N_11884,N_11821,N_11744);
nand U11885 (N_11885,N_11805,N_11723);
and U11886 (N_11886,N_11819,N_11825);
or U11887 (N_11887,N_11808,N_11782);
and U11888 (N_11888,N_11724,N_11783);
nand U11889 (N_11889,N_11775,N_11715);
nor U11890 (N_11890,N_11731,N_11710);
xnor U11891 (N_11891,N_11772,N_11704);
nor U11892 (N_11892,N_11799,N_11801);
or U11893 (N_11893,N_11832,N_11813);
nand U11894 (N_11894,N_11766,N_11818);
nand U11895 (N_11895,N_11848,N_11839);
nand U11896 (N_11896,N_11752,N_11774);
or U11897 (N_11897,N_11745,N_11791);
or U11898 (N_11898,N_11835,N_11751);
xnor U11899 (N_11899,N_11727,N_11831);
or U11900 (N_11900,N_11827,N_11828);
xnor U11901 (N_11901,N_11707,N_11738);
or U11902 (N_11902,N_11810,N_11779);
and U11903 (N_11903,N_11706,N_11806);
xor U11904 (N_11904,N_11849,N_11792);
nor U11905 (N_11905,N_11713,N_11771);
xnor U11906 (N_11906,N_11758,N_11720);
nand U11907 (N_11907,N_11700,N_11787);
or U11908 (N_11908,N_11780,N_11803);
and U11909 (N_11909,N_11770,N_11817);
xor U11910 (N_11910,N_11785,N_11784);
nand U11911 (N_11911,N_11794,N_11788);
nor U11912 (N_11912,N_11728,N_11719);
or U11913 (N_11913,N_11812,N_11793);
nand U11914 (N_11914,N_11778,N_11826);
nand U11915 (N_11915,N_11822,N_11777);
or U11916 (N_11916,N_11776,N_11734);
and U11917 (N_11917,N_11847,N_11726);
or U11918 (N_11918,N_11830,N_11844);
xor U11919 (N_11919,N_11703,N_11846);
or U11920 (N_11920,N_11702,N_11836);
xnor U11921 (N_11921,N_11811,N_11765);
xnor U11922 (N_11922,N_11797,N_11773);
nand U11923 (N_11923,N_11837,N_11809);
xnor U11924 (N_11924,N_11820,N_11843);
nor U11925 (N_11925,N_11838,N_11729);
and U11926 (N_11926,N_11718,N_11813);
xnor U11927 (N_11927,N_11785,N_11807);
nand U11928 (N_11928,N_11743,N_11832);
or U11929 (N_11929,N_11780,N_11758);
or U11930 (N_11930,N_11720,N_11743);
xor U11931 (N_11931,N_11721,N_11753);
or U11932 (N_11932,N_11757,N_11736);
or U11933 (N_11933,N_11736,N_11753);
xnor U11934 (N_11934,N_11793,N_11769);
nand U11935 (N_11935,N_11831,N_11782);
nor U11936 (N_11936,N_11773,N_11717);
nand U11937 (N_11937,N_11832,N_11836);
nor U11938 (N_11938,N_11835,N_11717);
nor U11939 (N_11939,N_11720,N_11813);
xor U11940 (N_11940,N_11771,N_11751);
or U11941 (N_11941,N_11769,N_11759);
nand U11942 (N_11942,N_11793,N_11724);
nor U11943 (N_11943,N_11792,N_11774);
nand U11944 (N_11944,N_11740,N_11805);
nand U11945 (N_11945,N_11733,N_11731);
xnor U11946 (N_11946,N_11743,N_11718);
or U11947 (N_11947,N_11766,N_11749);
and U11948 (N_11948,N_11732,N_11805);
xnor U11949 (N_11949,N_11740,N_11801);
or U11950 (N_11950,N_11789,N_11735);
or U11951 (N_11951,N_11776,N_11727);
xnor U11952 (N_11952,N_11803,N_11750);
and U11953 (N_11953,N_11845,N_11768);
and U11954 (N_11954,N_11739,N_11837);
nor U11955 (N_11955,N_11838,N_11710);
and U11956 (N_11956,N_11818,N_11847);
or U11957 (N_11957,N_11737,N_11825);
and U11958 (N_11958,N_11848,N_11849);
xnor U11959 (N_11959,N_11819,N_11722);
or U11960 (N_11960,N_11811,N_11837);
or U11961 (N_11961,N_11709,N_11846);
xor U11962 (N_11962,N_11771,N_11707);
nor U11963 (N_11963,N_11749,N_11779);
nor U11964 (N_11964,N_11725,N_11717);
xor U11965 (N_11965,N_11703,N_11761);
or U11966 (N_11966,N_11725,N_11815);
xor U11967 (N_11967,N_11817,N_11804);
and U11968 (N_11968,N_11722,N_11837);
or U11969 (N_11969,N_11782,N_11773);
nand U11970 (N_11970,N_11829,N_11787);
nand U11971 (N_11971,N_11815,N_11772);
nand U11972 (N_11972,N_11813,N_11830);
and U11973 (N_11973,N_11766,N_11831);
xnor U11974 (N_11974,N_11800,N_11821);
nand U11975 (N_11975,N_11792,N_11734);
xnor U11976 (N_11976,N_11772,N_11789);
nor U11977 (N_11977,N_11779,N_11764);
or U11978 (N_11978,N_11832,N_11716);
xor U11979 (N_11979,N_11710,N_11774);
nand U11980 (N_11980,N_11825,N_11713);
nor U11981 (N_11981,N_11840,N_11763);
xor U11982 (N_11982,N_11737,N_11768);
nor U11983 (N_11983,N_11738,N_11749);
or U11984 (N_11984,N_11754,N_11838);
and U11985 (N_11985,N_11793,N_11710);
or U11986 (N_11986,N_11741,N_11735);
or U11987 (N_11987,N_11709,N_11798);
and U11988 (N_11988,N_11768,N_11810);
nand U11989 (N_11989,N_11745,N_11712);
and U11990 (N_11990,N_11800,N_11846);
or U11991 (N_11991,N_11796,N_11743);
nand U11992 (N_11992,N_11733,N_11744);
and U11993 (N_11993,N_11803,N_11753);
or U11994 (N_11994,N_11809,N_11762);
xor U11995 (N_11995,N_11817,N_11701);
nor U11996 (N_11996,N_11823,N_11720);
nor U11997 (N_11997,N_11726,N_11817);
nor U11998 (N_11998,N_11758,N_11709);
xor U11999 (N_11999,N_11791,N_11752);
and U12000 (N_12000,N_11951,N_11943);
or U12001 (N_12001,N_11875,N_11898);
nand U12002 (N_12002,N_11979,N_11897);
or U12003 (N_12003,N_11861,N_11909);
nor U12004 (N_12004,N_11870,N_11894);
nor U12005 (N_12005,N_11891,N_11932);
and U12006 (N_12006,N_11964,N_11982);
and U12007 (N_12007,N_11944,N_11855);
nor U12008 (N_12008,N_11992,N_11987);
and U12009 (N_12009,N_11984,N_11873);
nor U12010 (N_12010,N_11955,N_11960);
or U12011 (N_12011,N_11997,N_11981);
and U12012 (N_12012,N_11863,N_11895);
nand U12013 (N_12013,N_11880,N_11953);
xnor U12014 (N_12014,N_11970,N_11949);
or U12015 (N_12015,N_11882,N_11945);
xnor U12016 (N_12016,N_11903,N_11852);
nor U12017 (N_12017,N_11874,N_11986);
xor U12018 (N_12018,N_11998,N_11884);
and U12019 (N_12019,N_11920,N_11927);
nor U12020 (N_12020,N_11919,N_11851);
xnor U12021 (N_12021,N_11869,N_11876);
or U12022 (N_12022,N_11978,N_11922);
nor U12023 (N_12023,N_11867,N_11893);
xnor U12024 (N_12024,N_11954,N_11988);
xnor U12025 (N_12025,N_11853,N_11887);
and U12026 (N_12026,N_11985,N_11877);
nor U12027 (N_12027,N_11974,N_11933);
xor U12028 (N_12028,N_11896,N_11879);
nand U12029 (N_12029,N_11957,N_11991);
xnor U12030 (N_12030,N_11888,N_11980);
nor U12031 (N_12031,N_11912,N_11993);
or U12032 (N_12032,N_11926,N_11856);
nor U12033 (N_12033,N_11976,N_11923);
xor U12034 (N_12034,N_11868,N_11913);
or U12035 (N_12035,N_11854,N_11892);
and U12036 (N_12036,N_11907,N_11999);
nand U12037 (N_12037,N_11935,N_11952);
nor U12038 (N_12038,N_11928,N_11939);
xnor U12039 (N_12039,N_11958,N_11946);
xor U12040 (N_12040,N_11940,N_11977);
and U12041 (N_12041,N_11934,N_11936);
nor U12042 (N_12042,N_11969,N_11965);
xnor U12043 (N_12043,N_11883,N_11941);
nor U12044 (N_12044,N_11990,N_11962);
nand U12045 (N_12045,N_11908,N_11862);
nand U12046 (N_12046,N_11917,N_11871);
nor U12047 (N_12047,N_11996,N_11931);
nor U12048 (N_12048,N_11857,N_11938);
and U12049 (N_12049,N_11950,N_11994);
or U12050 (N_12050,N_11967,N_11983);
nor U12051 (N_12051,N_11930,N_11995);
xor U12052 (N_12052,N_11989,N_11959);
or U12053 (N_12053,N_11878,N_11865);
and U12054 (N_12054,N_11968,N_11924);
or U12055 (N_12055,N_11905,N_11902);
or U12056 (N_12056,N_11889,N_11911);
nand U12057 (N_12057,N_11915,N_11942);
or U12058 (N_12058,N_11966,N_11948);
nand U12059 (N_12059,N_11937,N_11859);
and U12060 (N_12060,N_11872,N_11973);
or U12061 (N_12061,N_11929,N_11916);
nand U12062 (N_12062,N_11881,N_11961);
and U12063 (N_12063,N_11918,N_11906);
xnor U12064 (N_12064,N_11914,N_11925);
or U12065 (N_12065,N_11864,N_11947);
and U12066 (N_12066,N_11899,N_11885);
nor U12067 (N_12067,N_11910,N_11971);
and U12068 (N_12068,N_11956,N_11860);
xor U12069 (N_12069,N_11866,N_11886);
xnor U12070 (N_12070,N_11850,N_11900);
nand U12071 (N_12071,N_11972,N_11921);
xor U12072 (N_12072,N_11901,N_11975);
or U12073 (N_12073,N_11963,N_11858);
xnor U12074 (N_12074,N_11890,N_11904);
and U12075 (N_12075,N_11873,N_11868);
nand U12076 (N_12076,N_11952,N_11865);
xnor U12077 (N_12077,N_11877,N_11861);
xnor U12078 (N_12078,N_11893,N_11932);
nand U12079 (N_12079,N_11955,N_11918);
nor U12080 (N_12080,N_11964,N_11906);
nand U12081 (N_12081,N_11956,N_11929);
or U12082 (N_12082,N_11900,N_11966);
nor U12083 (N_12083,N_11873,N_11915);
and U12084 (N_12084,N_11976,N_11929);
nand U12085 (N_12085,N_11941,N_11956);
and U12086 (N_12086,N_11980,N_11868);
and U12087 (N_12087,N_11874,N_11870);
nor U12088 (N_12088,N_11900,N_11867);
xnor U12089 (N_12089,N_11958,N_11924);
or U12090 (N_12090,N_11898,N_11967);
nand U12091 (N_12091,N_11960,N_11944);
or U12092 (N_12092,N_11924,N_11953);
nor U12093 (N_12093,N_11894,N_11872);
nor U12094 (N_12094,N_11983,N_11945);
and U12095 (N_12095,N_11915,N_11916);
xor U12096 (N_12096,N_11953,N_11867);
or U12097 (N_12097,N_11949,N_11934);
and U12098 (N_12098,N_11877,N_11927);
xor U12099 (N_12099,N_11984,N_11943);
and U12100 (N_12100,N_11925,N_11997);
and U12101 (N_12101,N_11981,N_11929);
or U12102 (N_12102,N_11871,N_11866);
or U12103 (N_12103,N_11914,N_11893);
or U12104 (N_12104,N_11938,N_11983);
nor U12105 (N_12105,N_11921,N_11914);
nor U12106 (N_12106,N_11850,N_11879);
xnor U12107 (N_12107,N_11871,N_11853);
and U12108 (N_12108,N_11960,N_11898);
xor U12109 (N_12109,N_11923,N_11888);
or U12110 (N_12110,N_11868,N_11851);
xor U12111 (N_12111,N_11996,N_11927);
xor U12112 (N_12112,N_11877,N_11982);
xnor U12113 (N_12113,N_11858,N_11936);
or U12114 (N_12114,N_11927,N_11869);
nand U12115 (N_12115,N_11880,N_11917);
nand U12116 (N_12116,N_11949,N_11947);
or U12117 (N_12117,N_11950,N_11951);
nand U12118 (N_12118,N_11903,N_11885);
nor U12119 (N_12119,N_11942,N_11921);
or U12120 (N_12120,N_11913,N_11949);
nand U12121 (N_12121,N_11985,N_11919);
nor U12122 (N_12122,N_11920,N_11957);
xor U12123 (N_12123,N_11880,N_11865);
nor U12124 (N_12124,N_11915,N_11925);
nor U12125 (N_12125,N_11989,N_11987);
nor U12126 (N_12126,N_11938,N_11966);
nor U12127 (N_12127,N_11920,N_11970);
nand U12128 (N_12128,N_11932,N_11862);
and U12129 (N_12129,N_11942,N_11961);
and U12130 (N_12130,N_11981,N_11873);
nor U12131 (N_12131,N_11971,N_11900);
nand U12132 (N_12132,N_11996,N_11899);
or U12133 (N_12133,N_11949,N_11999);
nor U12134 (N_12134,N_11907,N_11870);
and U12135 (N_12135,N_11904,N_11993);
or U12136 (N_12136,N_11913,N_11959);
and U12137 (N_12137,N_11916,N_11994);
nor U12138 (N_12138,N_11903,N_11892);
nor U12139 (N_12139,N_11949,N_11861);
and U12140 (N_12140,N_11880,N_11983);
nor U12141 (N_12141,N_11964,N_11934);
and U12142 (N_12142,N_11930,N_11949);
nand U12143 (N_12143,N_11959,N_11886);
nand U12144 (N_12144,N_11974,N_11885);
nor U12145 (N_12145,N_11965,N_11957);
xnor U12146 (N_12146,N_11990,N_11878);
or U12147 (N_12147,N_11859,N_11921);
and U12148 (N_12148,N_11901,N_11928);
nand U12149 (N_12149,N_11956,N_11947);
xnor U12150 (N_12150,N_12092,N_12084);
nand U12151 (N_12151,N_12087,N_12041);
nand U12152 (N_12152,N_12046,N_12057);
xor U12153 (N_12153,N_12121,N_12111);
xnor U12154 (N_12154,N_12011,N_12102);
and U12155 (N_12155,N_12132,N_12123);
or U12156 (N_12156,N_12130,N_12058);
xor U12157 (N_12157,N_12086,N_12108);
nand U12158 (N_12158,N_12089,N_12112);
or U12159 (N_12159,N_12074,N_12016);
nor U12160 (N_12160,N_12068,N_12113);
or U12161 (N_12161,N_12035,N_12075);
and U12162 (N_12162,N_12119,N_12071);
xor U12163 (N_12163,N_12077,N_12053);
nor U12164 (N_12164,N_12097,N_12104);
xnor U12165 (N_12165,N_12145,N_12004);
or U12166 (N_12166,N_12007,N_12062);
or U12167 (N_12167,N_12002,N_12038);
and U12168 (N_12168,N_12096,N_12101);
xnor U12169 (N_12169,N_12014,N_12125);
nor U12170 (N_12170,N_12049,N_12144);
nor U12171 (N_12171,N_12103,N_12118);
nand U12172 (N_12172,N_12050,N_12063);
nor U12173 (N_12173,N_12072,N_12018);
xnor U12174 (N_12174,N_12031,N_12076);
xnor U12175 (N_12175,N_12142,N_12120);
xnor U12176 (N_12176,N_12134,N_12015);
nor U12177 (N_12177,N_12033,N_12009);
nand U12178 (N_12178,N_12017,N_12147);
nor U12179 (N_12179,N_12052,N_12146);
nor U12180 (N_12180,N_12055,N_12073);
or U12181 (N_12181,N_12005,N_12083);
nor U12182 (N_12182,N_12060,N_12107);
or U12183 (N_12183,N_12032,N_12021);
nand U12184 (N_12184,N_12027,N_12039);
nand U12185 (N_12185,N_12110,N_12012);
or U12186 (N_12186,N_12054,N_12067);
nand U12187 (N_12187,N_12090,N_12030);
or U12188 (N_12188,N_12034,N_12051);
and U12189 (N_12189,N_12098,N_12044);
nor U12190 (N_12190,N_12138,N_12122);
nand U12191 (N_12191,N_12003,N_12135);
nor U12192 (N_12192,N_12043,N_12069);
and U12193 (N_12193,N_12029,N_12023);
xnor U12194 (N_12194,N_12010,N_12028);
nand U12195 (N_12195,N_12127,N_12149);
nand U12196 (N_12196,N_12143,N_12114);
and U12197 (N_12197,N_12066,N_12136);
and U12198 (N_12198,N_12026,N_12020);
xor U12199 (N_12199,N_12006,N_12133);
and U12200 (N_12200,N_12064,N_12093);
nand U12201 (N_12201,N_12047,N_12079);
nand U12202 (N_12202,N_12115,N_12088);
nand U12203 (N_12203,N_12019,N_12045);
or U12204 (N_12204,N_12070,N_12116);
nor U12205 (N_12205,N_12124,N_12099);
nor U12206 (N_12206,N_12129,N_12008);
nand U12207 (N_12207,N_12025,N_12037);
nor U12208 (N_12208,N_12117,N_12085);
and U12209 (N_12209,N_12078,N_12065);
and U12210 (N_12210,N_12000,N_12105);
and U12211 (N_12211,N_12081,N_12059);
and U12212 (N_12212,N_12140,N_12106);
nor U12213 (N_12213,N_12040,N_12080);
and U12214 (N_12214,N_12128,N_12082);
or U12215 (N_12215,N_12056,N_12100);
and U12216 (N_12216,N_12036,N_12091);
or U12217 (N_12217,N_12137,N_12001);
and U12218 (N_12218,N_12131,N_12095);
and U12219 (N_12219,N_12013,N_12022);
nand U12220 (N_12220,N_12042,N_12024);
or U12221 (N_12221,N_12109,N_12139);
nor U12222 (N_12222,N_12048,N_12141);
xor U12223 (N_12223,N_12126,N_12061);
and U12224 (N_12224,N_12148,N_12094);
nand U12225 (N_12225,N_12111,N_12089);
nor U12226 (N_12226,N_12083,N_12029);
or U12227 (N_12227,N_12146,N_12114);
and U12228 (N_12228,N_12020,N_12034);
xnor U12229 (N_12229,N_12110,N_12142);
and U12230 (N_12230,N_12054,N_12040);
xor U12231 (N_12231,N_12146,N_12148);
and U12232 (N_12232,N_12002,N_12055);
nor U12233 (N_12233,N_12091,N_12035);
or U12234 (N_12234,N_12090,N_12019);
nor U12235 (N_12235,N_12007,N_12065);
and U12236 (N_12236,N_12049,N_12085);
and U12237 (N_12237,N_12089,N_12025);
or U12238 (N_12238,N_12143,N_12078);
or U12239 (N_12239,N_12133,N_12094);
nor U12240 (N_12240,N_12078,N_12088);
and U12241 (N_12241,N_12001,N_12010);
nand U12242 (N_12242,N_12091,N_12037);
nor U12243 (N_12243,N_12074,N_12129);
nand U12244 (N_12244,N_12078,N_12148);
nor U12245 (N_12245,N_12004,N_12075);
xor U12246 (N_12246,N_12142,N_12128);
nand U12247 (N_12247,N_12023,N_12021);
nor U12248 (N_12248,N_12064,N_12077);
nor U12249 (N_12249,N_12082,N_12040);
xnor U12250 (N_12250,N_12042,N_12048);
xor U12251 (N_12251,N_12102,N_12041);
xor U12252 (N_12252,N_12020,N_12115);
xnor U12253 (N_12253,N_12066,N_12004);
nor U12254 (N_12254,N_12053,N_12079);
and U12255 (N_12255,N_12103,N_12095);
and U12256 (N_12256,N_12097,N_12116);
nor U12257 (N_12257,N_12086,N_12020);
nand U12258 (N_12258,N_12077,N_12094);
nand U12259 (N_12259,N_12125,N_12076);
and U12260 (N_12260,N_12027,N_12128);
nand U12261 (N_12261,N_12013,N_12062);
and U12262 (N_12262,N_12112,N_12120);
nand U12263 (N_12263,N_12051,N_12084);
nand U12264 (N_12264,N_12104,N_12114);
nand U12265 (N_12265,N_12006,N_12033);
or U12266 (N_12266,N_12027,N_12064);
nor U12267 (N_12267,N_12145,N_12109);
nand U12268 (N_12268,N_12084,N_12038);
xor U12269 (N_12269,N_12062,N_12029);
xor U12270 (N_12270,N_12020,N_12146);
nand U12271 (N_12271,N_12025,N_12054);
or U12272 (N_12272,N_12018,N_12141);
xor U12273 (N_12273,N_12116,N_12092);
nor U12274 (N_12274,N_12025,N_12098);
and U12275 (N_12275,N_12047,N_12128);
nand U12276 (N_12276,N_12149,N_12042);
or U12277 (N_12277,N_12058,N_12012);
nor U12278 (N_12278,N_12064,N_12141);
xor U12279 (N_12279,N_12001,N_12110);
nand U12280 (N_12280,N_12006,N_12084);
nand U12281 (N_12281,N_12132,N_12087);
nand U12282 (N_12282,N_12032,N_12033);
nor U12283 (N_12283,N_12011,N_12068);
or U12284 (N_12284,N_12093,N_12025);
nor U12285 (N_12285,N_12091,N_12079);
and U12286 (N_12286,N_12000,N_12017);
nor U12287 (N_12287,N_12079,N_12111);
or U12288 (N_12288,N_12066,N_12140);
nor U12289 (N_12289,N_12058,N_12029);
xor U12290 (N_12290,N_12061,N_12082);
xor U12291 (N_12291,N_12133,N_12070);
xnor U12292 (N_12292,N_12077,N_12011);
or U12293 (N_12293,N_12130,N_12138);
nand U12294 (N_12294,N_12130,N_12129);
nand U12295 (N_12295,N_12068,N_12091);
nor U12296 (N_12296,N_12075,N_12107);
or U12297 (N_12297,N_12146,N_12016);
nor U12298 (N_12298,N_12041,N_12130);
or U12299 (N_12299,N_12053,N_12131);
xor U12300 (N_12300,N_12207,N_12267);
nor U12301 (N_12301,N_12156,N_12223);
nand U12302 (N_12302,N_12226,N_12153);
or U12303 (N_12303,N_12255,N_12164);
xor U12304 (N_12304,N_12299,N_12229);
or U12305 (N_12305,N_12192,N_12151);
nor U12306 (N_12306,N_12279,N_12215);
xnor U12307 (N_12307,N_12174,N_12196);
or U12308 (N_12308,N_12253,N_12231);
or U12309 (N_12309,N_12274,N_12193);
and U12310 (N_12310,N_12232,N_12205);
xor U12311 (N_12311,N_12158,N_12199);
nand U12312 (N_12312,N_12175,N_12282);
and U12313 (N_12313,N_12203,N_12177);
nand U12314 (N_12314,N_12296,N_12198);
xnor U12315 (N_12315,N_12217,N_12251);
nand U12316 (N_12316,N_12213,N_12165);
xnor U12317 (N_12317,N_12245,N_12297);
nor U12318 (N_12318,N_12210,N_12160);
xor U12319 (N_12319,N_12257,N_12161);
nor U12320 (N_12320,N_12277,N_12294);
nand U12321 (N_12321,N_12288,N_12167);
xor U12322 (N_12322,N_12269,N_12200);
xnor U12323 (N_12323,N_12230,N_12218);
nand U12324 (N_12324,N_12275,N_12208);
xnor U12325 (N_12325,N_12298,N_12271);
xor U12326 (N_12326,N_12202,N_12150);
nor U12327 (N_12327,N_12212,N_12220);
or U12328 (N_12328,N_12173,N_12219);
nand U12329 (N_12329,N_12256,N_12280);
xnor U12330 (N_12330,N_12190,N_12286);
xor U12331 (N_12331,N_12180,N_12284);
nand U12332 (N_12332,N_12206,N_12191);
nand U12333 (N_12333,N_12291,N_12163);
xnor U12334 (N_12334,N_12234,N_12189);
and U12335 (N_12335,N_12211,N_12246);
and U12336 (N_12336,N_12168,N_12157);
or U12337 (N_12337,N_12216,N_12242);
nand U12338 (N_12338,N_12228,N_12249);
nor U12339 (N_12339,N_12238,N_12262);
or U12340 (N_12340,N_12243,N_12260);
nand U12341 (N_12341,N_12268,N_12184);
or U12342 (N_12342,N_12195,N_12285);
and U12343 (N_12343,N_12250,N_12270);
and U12344 (N_12344,N_12278,N_12183);
or U12345 (N_12345,N_12264,N_12152);
and U12346 (N_12346,N_12172,N_12244);
nor U12347 (N_12347,N_12283,N_12287);
nor U12348 (N_12348,N_12254,N_12289);
xor U12349 (N_12349,N_12186,N_12235);
and U12350 (N_12350,N_12178,N_12224);
xor U12351 (N_12351,N_12273,N_12182);
and U12352 (N_12352,N_12179,N_12281);
nand U12353 (N_12353,N_12221,N_12162);
nor U12354 (N_12354,N_12227,N_12295);
and U12355 (N_12355,N_12170,N_12236);
nor U12356 (N_12356,N_12263,N_12181);
and U12357 (N_12357,N_12225,N_12261);
nor U12358 (N_12358,N_12214,N_12188);
nor U12359 (N_12359,N_12265,N_12154);
or U12360 (N_12360,N_12266,N_12290);
xnor U12361 (N_12361,N_12201,N_12209);
nand U12362 (N_12362,N_12187,N_12293);
nand U12363 (N_12363,N_12259,N_12292);
nor U12364 (N_12364,N_12171,N_12272);
or U12365 (N_12365,N_12159,N_12240);
nand U12366 (N_12366,N_12176,N_12166);
nand U12367 (N_12367,N_12233,N_12252);
and U12368 (N_12368,N_12237,N_12204);
nand U12369 (N_12369,N_12258,N_12241);
nor U12370 (N_12370,N_12239,N_12169);
xnor U12371 (N_12371,N_12248,N_12197);
nand U12372 (N_12372,N_12276,N_12185);
and U12373 (N_12373,N_12194,N_12247);
nand U12374 (N_12374,N_12155,N_12222);
nor U12375 (N_12375,N_12213,N_12280);
nor U12376 (N_12376,N_12197,N_12209);
xnor U12377 (N_12377,N_12181,N_12291);
nand U12378 (N_12378,N_12185,N_12232);
nor U12379 (N_12379,N_12187,N_12231);
nor U12380 (N_12380,N_12267,N_12169);
nor U12381 (N_12381,N_12277,N_12203);
xor U12382 (N_12382,N_12168,N_12170);
nand U12383 (N_12383,N_12175,N_12161);
nor U12384 (N_12384,N_12239,N_12278);
or U12385 (N_12385,N_12153,N_12255);
and U12386 (N_12386,N_12237,N_12219);
or U12387 (N_12387,N_12297,N_12183);
or U12388 (N_12388,N_12152,N_12206);
xnor U12389 (N_12389,N_12263,N_12250);
nor U12390 (N_12390,N_12201,N_12290);
nand U12391 (N_12391,N_12245,N_12257);
nor U12392 (N_12392,N_12152,N_12190);
and U12393 (N_12393,N_12281,N_12181);
nand U12394 (N_12394,N_12288,N_12285);
xnor U12395 (N_12395,N_12194,N_12186);
nand U12396 (N_12396,N_12150,N_12167);
nand U12397 (N_12397,N_12283,N_12211);
nand U12398 (N_12398,N_12274,N_12161);
xor U12399 (N_12399,N_12241,N_12205);
nand U12400 (N_12400,N_12172,N_12290);
xor U12401 (N_12401,N_12261,N_12153);
nand U12402 (N_12402,N_12217,N_12232);
or U12403 (N_12403,N_12200,N_12267);
nor U12404 (N_12404,N_12164,N_12253);
and U12405 (N_12405,N_12184,N_12252);
and U12406 (N_12406,N_12194,N_12156);
nand U12407 (N_12407,N_12175,N_12164);
or U12408 (N_12408,N_12264,N_12231);
nor U12409 (N_12409,N_12164,N_12170);
xnor U12410 (N_12410,N_12294,N_12271);
and U12411 (N_12411,N_12269,N_12221);
nor U12412 (N_12412,N_12244,N_12260);
nand U12413 (N_12413,N_12164,N_12264);
xnor U12414 (N_12414,N_12267,N_12240);
or U12415 (N_12415,N_12279,N_12226);
or U12416 (N_12416,N_12253,N_12285);
nand U12417 (N_12417,N_12151,N_12277);
and U12418 (N_12418,N_12246,N_12267);
nand U12419 (N_12419,N_12286,N_12275);
and U12420 (N_12420,N_12159,N_12211);
nand U12421 (N_12421,N_12156,N_12166);
and U12422 (N_12422,N_12276,N_12233);
or U12423 (N_12423,N_12281,N_12190);
nand U12424 (N_12424,N_12269,N_12207);
nor U12425 (N_12425,N_12221,N_12223);
and U12426 (N_12426,N_12160,N_12157);
xor U12427 (N_12427,N_12165,N_12238);
nand U12428 (N_12428,N_12271,N_12231);
xor U12429 (N_12429,N_12265,N_12251);
xnor U12430 (N_12430,N_12294,N_12183);
nand U12431 (N_12431,N_12284,N_12202);
or U12432 (N_12432,N_12269,N_12277);
nor U12433 (N_12433,N_12253,N_12158);
and U12434 (N_12434,N_12288,N_12210);
and U12435 (N_12435,N_12195,N_12294);
or U12436 (N_12436,N_12254,N_12279);
nor U12437 (N_12437,N_12217,N_12229);
xnor U12438 (N_12438,N_12166,N_12204);
or U12439 (N_12439,N_12206,N_12298);
and U12440 (N_12440,N_12289,N_12237);
nand U12441 (N_12441,N_12283,N_12180);
nor U12442 (N_12442,N_12293,N_12274);
nor U12443 (N_12443,N_12264,N_12274);
xnor U12444 (N_12444,N_12191,N_12265);
or U12445 (N_12445,N_12158,N_12286);
nand U12446 (N_12446,N_12202,N_12280);
and U12447 (N_12447,N_12260,N_12159);
xor U12448 (N_12448,N_12168,N_12280);
nand U12449 (N_12449,N_12238,N_12159);
nand U12450 (N_12450,N_12309,N_12432);
nor U12451 (N_12451,N_12346,N_12367);
and U12452 (N_12452,N_12359,N_12441);
and U12453 (N_12453,N_12429,N_12393);
xor U12454 (N_12454,N_12426,N_12320);
and U12455 (N_12455,N_12407,N_12412);
or U12456 (N_12456,N_12448,N_12446);
or U12457 (N_12457,N_12411,N_12406);
xor U12458 (N_12458,N_12365,N_12366);
or U12459 (N_12459,N_12338,N_12404);
or U12460 (N_12460,N_12356,N_12447);
or U12461 (N_12461,N_12347,N_12362);
and U12462 (N_12462,N_12357,N_12395);
or U12463 (N_12463,N_12301,N_12358);
xor U12464 (N_12464,N_12307,N_12415);
xor U12465 (N_12465,N_12302,N_12427);
nand U12466 (N_12466,N_12323,N_12431);
or U12467 (N_12467,N_12413,N_12384);
nor U12468 (N_12468,N_12425,N_12390);
and U12469 (N_12469,N_12391,N_12314);
nand U12470 (N_12470,N_12352,N_12315);
and U12471 (N_12471,N_12394,N_12434);
and U12472 (N_12472,N_12329,N_12363);
nand U12473 (N_12473,N_12423,N_12311);
nand U12474 (N_12474,N_12375,N_12354);
nor U12475 (N_12475,N_12360,N_12334);
nor U12476 (N_12476,N_12351,N_12319);
and U12477 (N_12477,N_12392,N_12408);
or U12478 (N_12478,N_12433,N_12353);
and U12479 (N_12479,N_12326,N_12439);
nand U12480 (N_12480,N_12306,N_12327);
xor U12481 (N_12481,N_12333,N_12436);
xnor U12482 (N_12482,N_12387,N_12325);
xor U12483 (N_12483,N_12377,N_12331);
nor U12484 (N_12484,N_12419,N_12373);
and U12485 (N_12485,N_12438,N_12364);
nand U12486 (N_12486,N_12378,N_12361);
xor U12487 (N_12487,N_12399,N_12402);
and U12488 (N_12488,N_12410,N_12383);
or U12489 (N_12489,N_12350,N_12380);
or U12490 (N_12490,N_12403,N_12321);
xor U12491 (N_12491,N_12414,N_12420);
nand U12492 (N_12492,N_12341,N_12444);
nor U12493 (N_12493,N_12322,N_12421);
xor U12494 (N_12494,N_12328,N_12335);
nand U12495 (N_12495,N_12417,N_12374);
nor U12496 (N_12496,N_12396,N_12304);
or U12497 (N_12497,N_12379,N_12371);
xor U12498 (N_12498,N_12418,N_12305);
xnor U12499 (N_12499,N_12386,N_12310);
xnor U12500 (N_12500,N_12316,N_12303);
xor U12501 (N_12501,N_12376,N_12437);
nor U12502 (N_12502,N_12389,N_12388);
nor U12503 (N_12503,N_12300,N_12332);
nand U12504 (N_12504,N_12435,N_12348);
and U12505 (N_12505,N_12401,N_12313);
nor U12506 (N_12506,N_12445,N_12355);
and U12507 (N_12507,N_12424,N_12318);
and U12508 (N_12508,N_12449,N_12324);
nand U12509 (N_12509,N_12372,N_12342);
xnor U12510 (N_12510,N_12442,N_12340);
nor U12511 (N_12511,N_12370,N_12368);
nor U12512 (N_12512,N_12312,N_12443);
xor U12513 (N_12513,N_12416,N_12330);
xnor U12514 (N_12514,N_12369,N_12430);
nand U12515 (N_12515,N_12422,N_12397);
nand U12516 (N_12516,N_12405,N_12440);
nor U12517 (N_12517,N_12349,N_12344);
or U12518 (N_12518,N_12381,N_12345);
or U12519 (N_12519,N_12385,N_12409);
nor U12520 (N_12520,N_12382,N_12339);
xor U12521 (N_12521,N_12428,N_12400);
or U12522 (N_12522,N_12343,N_12317);
nand U12523 (N_12523,N_12337,N_12398);
xnor U12524 (N_12524,N_12336,N_12308);
nor U12525 (N_12525,N_12356,N_12388);
and U12526 (N_12526,N_12365,N_12337);
and U12527 (N_12527,N_12381,N_12323);
nand U12528 (N_12528,N_12364,N_12320);
nand U12529 (N_12529,N_12378,N_12392);
nand U12530 (N_12530,N_12417,N_12405);
nor U12531 (N_12531,N_12367,N_12376);
and U12532 (N_12532,N_12383,N_12317);
xnor U12533 (N_12533,N_12351,N_12358);
nand U12534 (N_12534,N_12321,N_12327);
nand U12535 (N_12535,N_12439,N_12399);
or U12536 (N_12536,N_12307,N_12398);
and U12537 (N_12537,N_12343,N_12372);
nand U12538 (N_12538,N_12378,N_12389);
xnor U12539 (N_12539,N_12367,N_12395);
and U12540 (N_12540,N_12415,N_12340);
xnor U12541 (N_12541,N_12388,N_12301);
xnor U12542 (N_12542,N_12339,N_12391);
and U12543 (N_12543,N_12350,N_12437);
nand U12544 (N_12544,N_12438,N_12371);
nor U12545 (N_12545,N_12339,N_12319);
nand U12546 (N_12546,N_12418,N_12425);
nor U12547 (N_12547,N_12345,N_12365);
xnor U12548 (N_12548,N_12418,N_12337);
and U12549 (N_12549,N_12385,N_12372);
and U12550 (N_12550,N_12433,N_12313);
and U12551 (N_12551,N_12352,N_12328);
nor U12552 (N_12552,N_12404,N_12323);
and U12553 (N_12553,N_12337,N_12433);
xnor U12554 (N_12554,N_12338,N_12345);
nand U12555 (N_12555,N_12415,N_12440);
or U12556 (N_12556,N_12324,N_12357);
and U12557 (N_12557,N_12396,N_12402);
nand U12558 (N_12558,N_12352,N_12430);
nand U12559 (N_12559,N_12433,N_12414);
nor U12560 (N_12560,N_12383,N_12359);
or U12561 (N_12561,N_12345,N_12424);
xnor U12562 (N_12562,N_12311,N_12391);
nand U12563 (N_12563,N_12314,N_12323);
xnor U12564 (N_12564,N_12405,N_12381);
nand U12565 (N_12565,N_12406,N_12312);
nand U12566 (N_12566,N_12365,N_12411);
nand U12567 (N_12567,N_12414,N_12422);
or U12568 (N_12568,N_12444,N_12397);
nor U12569 (N_12569,N_12397,N_12419);
xnor U12570 (N_12570,N_12435,N_12408);
and U12571 (N_12571,N_12419,N_12439);
nand U12572 (N_12572,N_12390,N_12319);
and U12573 (N_12573,N_12339,N_12367);
xnor U12574 (N_12574,N_12325,N_12432);
or U12575 (N_12575,N_12332,N_12414);
or U12576 (N_12576,N_12302,N_12432);
xnor U12577 (N_12577,N_12430,N_12415);
and U12578 (N_12578,N_12409,N_12441);
xnor U12579 (N_12579,N_12317,N_12349);
or U12580 (N_12580,N_12386,N_12349);
nand U12581 (N_12581,N_12312,N_12431);
and U12582 (N_12582,N_12387,N_12396);
nor U12583 (N_12583,N_12417,N_12321);
or U12584 (N_12584,N_12348,N_12408);
xor U12585 (N_12585,N_12353,N_12371);
nand U12586 (N_12586,N_12391,N_12340);
nor U12587 (N_12587,N_12434,N_12413);
or U12588 (N_12588,N_12346,N_12357);
nor U12589 (N_12589,N_12366,N_12403);
or U12590 (N_12590,N_12370,N_12300);
or U12591 (N_12591,N_12387,N_12350);
nand U12592 (N_12592,N_12395,N_12317);
nand U12593 (N_12593,N_12448,N_12435);
nor U12594 (N_12594,N_12424,N_12444);
nand U12595 (N_12595,N_12372,N_12340);
and U12596 (N_12596,N_12406,N_12325);
and U12597 (N_12597,N_12345,N_12448);
nor U12598 (N_12598,N_12334,N_12389);
nor U12599 (N_12599,N_12447,N_12400);
and U12600 (N_12600,N_12562,N_12463);
and U12601 (N_12601,N_12501,N_12570);
nand U12602 (N_12602,N_12566,N_12568);
nand U12603 (N_12603,N_12481,N_12514);
xnor U12604 (N_12604,N_12498,N_12528);
and U12605 (N_12605,N_12457,N_12535);
nor U12606 (N_12606,N_12593,N_12475);
nor U12607 (N_12607,N_12541,N_12561);
xnor U12608 (N_12608,N_12526,N_12558);
xor U12609 (N_12609,N_12525,N_12546);
nor U12610 (N_12610,N_12458,N_12489);
and U12611 (N_12611,N_12557,N_12587);
nand U12612 (N_12612,N_12579,N_12565);
nor U12613 (N_12613,N_12563,N_12544);
and U12614 (N_12614,N_12581,N_12540);
or U12615 (N_12615,N_12508,N_12452);
xor U12616 (N_12616,N_12589,N_12536);
nor U12617 (N_12617,N_12496,N_12510);
xnor U12618 (N_12618,N_12504,N_12530);
nand U12619 (N_12619,N_12486,N_12450);
nand U12620 (N_12620,N_12513,N_12577);
xor U12621 (N_12621,N_12518,N_12473);
nor U12622 (N_12622,N_12506,N_12488);
nand U12623 (N_12623,N_12538,N_12572);
or U12624 (N_12624,N_12555,N_12453);
or U12625 (N_12625,N_12464,N_12479);
xor U12626 (N_12626,N_12578,N_12467);
nor U12627 (N_12627,N_12470,N_12474);
nand U12628 (N_12628,N_12454,N_12516);
nand U12629 (N_12629,N_12512,N_12519);
nand U12630 (N_12630,N_12485,N_12592);
xor U12631 (N_12631,N_12567,N_12527);
nand U12632 (N_12632,N_12576,N_12596);
xnor U12633 (N_12633,N_12552,N_12554);
nor U12634 (N_12634,N_12584,N_12517);
nor U12635 (N_12635,N_12594,N_12545);
and U12636 (N_12636,N_12560,N_12469);
nor U12637 (N_12637,N_12515,N_12553);
or U12638 (N_12638,N_12460,N_12548);
or U12639 (N_12639,N_12487,N_12597);
xor U12640 (N_12640,N_12591,N_12490);
xnor U12641 (N_12641,N_12582,N_12509);
xor U12642 (N_12642,N_12461,N_12556);
xnor U12643 (N_12643,N_12502,N_12550);
nand U12644 (N_12644,N_12505,N_12534);
xnor U12645 (N_12645,N_12573,N_12551);
or U12646 (N_12646,N_12559,N_12585);
xor U12647 (N_12647,N_12580,N_12520);
or U12648 (N_12648,N_12495,N_12493);
nand U12649 (N_12649,N_12466,N_12532);
nand U12650 (N_12650,N_12523,N_12468);
nand U12651 (N_12651,N_12459,N_12574);
xnor U12652 (N_12652,N_12455,N_12476);
nor U12653 (N_12653,N_12524,N_12471);
nand U12654 (N_12654,N_12521,N_12499);
or U12655 (N_12655,N_12569,N_12599);
nand U12656 (N_12656,N_12547,N_12533);
and U12657 (N_12657,N_12480,N_12507);
nand U12658 (N_12658,N_12529,N_12494);
xnor U12659 (N_12659,N_12477,N_12482);
xnor U12660 (N_12660,N_12484,N_12531);
and U12661 (N_12661,N_12491,N_12575);
xnor U12662 (N_12662,N_12539,N_12537);
or U12663 (N_12663,N_12588,N_12462);
xnor U12664 (N_12664,N_12497,N_12564);
nor U12665 (N_12665,N_12598,N_12543);
nand U12666 (N_12666,N_12542,N_12456);
or U12667 (N_12667,N_12595,N_12590);
and U12668 (N_12668,N_12586,N_12500);
and U12669 (N_12669,N_12465,N_12522);
nand U12670 (N_12670,N_12583,N_12472);
nor U12671 (N_12671,N_12511,N_12492);
and U12672 (N_12672,N_12451,N_12549);
or U12673 (N_12673,N_12483,N_12503);
or U12674 (N_12674,N_12571,N_12478);
nand U12675 (N_12675,N_12485,N_12542);
and U12676 (N_12676,N_12510,N_12543);
nand U12677 (N_12677,N_12500,N_12576);
xnor U12678 (N_12678,N_12589,N_12551);
xor U12679 (N_12679,N_12475,N_12462);
xor U12680 (N_12680,N_12596,N_12566);
nor U12681 (N_12681,N_12456,N_12518);
and U12682 (N_12682,N_12460,N_12510);
xor U12683 (N_12683,N_12576,N_12545);
and U12684 (N_12684,N_12526,N_12509);
xnor U12685 (N_12685,N_12567,N_12474);
nor U12686 (N_12686,N_12450,N_12512);
and U12687 (N_12687,N_12467,N_12519);
and U12688 (N_12688,N_12591,N_12571);
xnor U12689 (N_12689,N_12581,N_12506);
and U12690 (N_12690,N_12559,N_12545);
nand U12691 (N_12691,N_12478,N_12513);
nand U12692 (N_12692,N_12492,N_12499);
nor U12693 (N_12693,N_12457,N_12591);
nor U12694 (N_12694,N_12525,N_12552);
nand U12695 (N_12695,N_12489,N_12511);
and U12696 (N_12696,N_12538,N_12547);
and U12697 (N_12697,N_12523,N_12549);
and U12698 (N_12698,N_12554,N_12564);
nor U12699 (N_12699,N_12472,N_12532);
or U12700 (N_12700,N_12513,N_12538);
nor U12701 (N_12701,N_12542,N_12543);
and U12702 (N_12702,N_12465,N_12467);
or U12703 (N_12703,N_12572,N_12570);
xnor U12704 (N_12704,N_12513,N_12537);
nor U12705 (N_12705,N_12597,N_12541);
and U12706 (N_12706,N_12529,N_12484);
or U12707 (N_12707,N_12518,N_12596);
nor U12708 (N_12708,N_12493,N_12452);
xor U12709 (N_12709,N_12455,N_12587);
nor U12710 (N_12710,N_12586,N_12555);
nor U12711 (N_12711,N_12487,N_12569);
or U12712 (N_12712,N_12505,N_12568);
and U12713 (N_12713,N_12487,N_12588);
nand U12714 (N_12714,N_12560,N_12589);
nor U12715 (N_12715,N_12593,N_12582);
nand U12716 (N_12716,N_12509,N_12590);
xor U12717 (N_12717,N_12474,N_12555);
nand U12718 (N_12718,N_12563,N_12570);
nor U12719 (N_12719,N_12528,N_12497);
or U12720 (N_12720,N_12596,N_12475);
and U12721 (N_12721,N_12598,N_12529);
or U12722 (N_12722,N_12580,N_12515);
or U12723 (N_12723,N_12545,N_12454);
nor U12724 (N_12724,N_12594,N_12463);
nand U12725 (N_12725,N_12515,N_12535);
nand U12726 (N_12726,N_12472,N_12577);
nor U12727 (N_12727,N_12488,N_12584);
nand U12728 (N_12728,N_12456,N_12533);
nor U12729 (N_12729,N_12537,N_12559);
xnor U12730 (N_12730,N_12586,N_12513);
or U12731 (N_12731,N_12482,N_12572);
nor U12732 (N_12732,N_12522,N_12533);
and U12733 (N_12733,N_12538,N_12524);
nand U12734 (N_12734,N_12576,N_12468);
nor U12735 (N_12735,N_12474,N_12578);
or U12736 (N_12736,N_12568,N_12562);
or U12737 (N_12737,N_12575,N_12463);
nand U12738 (N_12738,N_12563,N_12481);
nor U12739 (N_12739,N_12482,N_12471);
or U12740 (N_12740,N_12579,N_12529);
or U12741 (N_12741,N_12489,N_12472);
nand U12742 (N_12742,N_12591,N_12471);
nor U12743 (N_12743,N_12581,N_12576);
nand U12744 (N_12744,N_12542,N_12565);
nor U12745 (N_12745,N_12583,N_12521);
nand U12746 (N_12746,N_12578,N_12589);
and U12747 (N_12747,N_12565,N_12514);
and U12748 (N_12748,N_12556,N_12478);
and U12749 (N_12749,N_12527,N_12494);
or U12750 (N_12750,N_12628,N_12635);
nor U12751 (N_12751,N_12749,N_12676);
nand U12752 (N_12752,N_12740,N_12624);
or U12753 (N_12753,N_12683,N_12620);
nor U12754 (N_12754,N_12691,N_12636);
or U12755 (N_12755,N_12603,N_12695);
and U12756 (N_12756,N_12614,N_12615);
nand U12757 (N_12757,N_12668,N_12675);
nor U12758 (N_12758,N_12722,N_12671);
and U12759 (N_12759,N_12726,N_12613);
or U12760 (N_12760,N_12602,N_12730);
nor U12761 (N_12761,N_12670,N_12634);
xor U12762 (N_12762,N_12721,N_12687);
and U12763 (N_12763,N_12682,N_12681);
and U12764 (N_12764,N_12746,N_12651);
nor U12765 (N_12765,N_12619,N_12640);
or U12766 (N_12766,N_12712,N_12650);
nor U12767 (N_12767,N_12659,N_12747);
or U12768 (N_12768,N_12652,N_12696);
xor U12769 (N_12769,N_12600,N_12700);
nand U12770 (N_12770,N_12710,N_12688);
nor U12771 (N_12771,N_12680,N_12653);
xor U12772 (N_12772,N_12632,N_12626);
or U12773 (N_12773,N_12701,N_12698);
or U12774 (N_12774,N_12741,N_12705);
nor U12775 (N_12775,N_12724,N_12631);
xor U12776 (N_12776,N_12667,N_12723);
or U12777 (N_12777,N_12649,N_12677);
nand U12778 (N_12778,N_12639,N_12699);
and U12779 (N_12779,N_12633,N_12669);
nand U12780 (N_12780,N_12658,N_12715);
and U12781 (N_12781,N_12692,N_12672);
and U12782 (N_12782,N_12684,N_12648);
nor U12783 (N_12783,N_12738,N_12657);
xnor U12784 (N_12784,N_12664,N_12604);
or U12785 (N_12785,N_12654,N_12733);
xnor U12786 (N_12786,N_12732,N_12716);
nor U12787 (N_12787,N_12627,N_12630);
xnor U12788 (N_12788,N_12641,N_12673);
and U12789 (N_12789,N_12729,N_12610);
and U12790 (N_12790,N_12714,N_12607);
xor U12791 (N_12791,N_12731,N_12739);
and U12792 (N_12792,N_12617,N_12706);
nor U12793 (N_12793,N_12611,N_12644);
nor U12794 (N_12794,N_12642,N_12665);
and U12795 (N_12795,N_12720,N_12625);
xnor U12796 (N_12796,N_12702,N_12717);
nand U12797 (N_12797,N_12690,N_12719);
nor U12798 (N_12798,N_12693,N_12679);
nand U12799 (N_12799,N_12703,N_12728);
nor U12800 (N_12800,N_12663,N_12735);
and U12801 (N_12801,N_12725,N_12656);
nand U12802 (N_12802,N_12645,N_12601);
nand U12803 (N_12803,N_12686,N_12736);
nor U12804 (N_12804,N_12608,N_12655);
nor U12805 (N_12805,N_12707,N_12737);
xor U12806 (N_12806,N_12629,N_12647);
and U12807 (N_12807,N_12713,N_12660);
nor U12808 (N_12808,N_12678,N_12697);
nand U12809 (N_12809,N_12743,N_12606);
xor U12810 (N_12810,N_12727,N_12718);
nor U12811 (N_12811,N_12734,N_12748);
nor U12812 (N_12812,N_12616,N_12621);
nor U12813 (N_12813,N_12638,N_12704);
nand U12814 (N_12814,N_12643,N_12605);
and U12815 (N_12815,N_12609,N_12637);
xor U12816 (N_12816,N_12694,N_12622);
xor U12817 (N_12817,N_12711,N_12744);
nand U12818 (N_12818,N_12661,N_12689);
and U12819 (N_12819,N_12708,N_12674);
nor U12820 (N_12820,N_12742,N_12745);
xor U12821 (N_12821,N_12612,N_12623);
and U12822 (N_12822,N_12662,N_12618);
and U12823 (N_12823,N_12709,N_12666);
xnor U12824 (N_12824,N_12685,N_12646);
or U12825 (N_12825,N_12631,N_12698);
and U12826 (N_12826,N_12664,N_12652);
nor U12827 (N_12827,N_12748,N_12613);
or U12828 (N_12828,N_12660,N_12710);
xor U12829 (N_12829,N_12711,N_12673);
and U12830 (N_12830,N_12662,N_12706);
xnor U12831 (N_12831,N_12729,N_12622);
nor U12832 (N_12832,N_12682,N_12673);
nand U12833 (N_12833,N_12631,N_12626);
nand U12834 (N_12834,N_12614,N_12634);
or U12835 (N_12835,N_12650,N_12634);
nand U12836 (N_12836,N_12612,N_12606);
nand U12837 (N_12837,N_12723,N_12698);
nand U12838 (N_12838,N_12736,N_12727);
xor U12839 (N_12839,N_12716,N_12664);
nand U12840 (N_12840,N_12649,N_12688);
or U12841 (N_12841,N_12605,N_12646);
and U12842 (N_12842,N_12601,N_12628);
xnor U12843 (N_12843,N_12639,N_12665);
xnor U12844 (N_12844,N_12694,N_12673);
nand U12845 (N_12845,N_12718,N_12735);
nand U12846 (N_12846,N_12641,N_12674);
nor U12847 (N_12847,N_12686,N_12727);
or U12848 (N_12848,N_12708,N_12679);
and U12849 (N_12849,N_12617,N_12625);
nand U12850 (N_12850,N_12709,N_12726);
and U12851 (N_12851,N_12643,N_12641);
nor U12852 (N_12852,N_12672,N_12746);
nand U12853 (N_12853,N_12680,N_12713);
nor U12854 (N_12854,N_12628,N_12706);
xor U12855 (N_12855,N_12673,N_12638);
xor U12856 (N_12856,N_12655,N_12674);
nor U12857 (N_12857,N_12702,N_12673);
and U12858 (N_12858,N_12715,N_12648);
or U12859 (N_12859,N_12636,N_12676);
xor U12860 (N_12860,N_12742,N_12740);
and U12861 (N_12861,N_12602,N_12616);
or U12862 (N_12862,N_12678,N_12652);
and U12863 (N_12863,N_12649,N_12700);
nor U12864 (N_12864,N_12639,N_12694);
and U12865 (N_12865,N_12639,N_12667);
and U12866 (N_12866,N_12685,N_12608);
and U12867 (N_12867,N_12690,N_12667);
nand U12868 (N_12868,N_12606,N_12641);
nand U12869 (N_12869,N_12644,N_12737);
or U12870 (N_12870,N_12609,N_12640);
or U12871 (N_12871,N_12632,N_12617);
or U12872 (N_12872,N_12684,N_12732);
xnor U12873 (N_12873,N_12647,N_12721);
xor U12874 (N_12874,N_12650,N_12680);
nor U12875 (N_12875,N_12742,N_12626);
xor U12876 (N_12876,N_12743,N_12699);
xor U12877 (N_12877,N_12682,N_12646);
nor U12878 (N_12878,N_12618,N_12600);
nand U12879 (N_12879,N_12643,N_12656);
xnor U12880 (N_12880,N_12648,N_12732);
and U12881 (N_12881,N_12610,N_12703);
nor U12882 (N_12882,N_12649,N_12713);
or U12883 (N_12883,N_12686,N_12644);
nand U12884 (N_12884,N_12747,N_12653);
nand U12885 (N_12885,N_12641,N_12621);
nand U12886 (N_12886,N_12743,N_12640);
xor U12887 (N_12887,N_12621,N_12619);
xnor U12888 (N_12888,N_12617,N_12655);
nor U12889 (N_12889,N_12622,N_12601);
xnor U12890 (N_12890,N_12670,N_12651);
and U12891 (N_12891,N_12610,N_12710);
or U12892 (N_12892,N_12744,N_12613);
nand U12893 (N_12893,N_12639,N_12602);
nor U12894 (N_12894,N_12749,N_12659);
and U12895 (N_12895,N_12740,N_12634);
nand U12896 (N_12896,N_12695,N_12616);
nand U12897 (N_12897,N_12668,N_12740);
and U12898 (N_12898,N_12748,N_12642);
nor U12899 (N_12899,N_12633,N_12671);
nand U12900 (N_12900,N_12855,N_12852);
or U12901 (N_12901,N_12781,N_12777);
or U12902 (N_12902,N_12804,N_12757);
nor U12903 (N_12903,N_12887,N_12778);
and U12904 (N_12904,N_12842,N_12839);
nor U12905 (N_12905,N_12774,N_12761);
or U12906 (N_12906,N_12846,N_12847);
and U12907 (N_12907,N_12869,N_12875);
nand U12908 (N_12908,N_12776,N_12764);
xor U12909 (N_12909,N_12835,N_12880);
nor U12910 (N_12910,N_12797,N_12895);
or U12911 (N_12911,N_12818,N_12888);
xnor U12912 (N_12912,N_12815,N_12786);
nand U12913 (N_12913,N_12832,N_12762);
xor U12914 (N_12914,N_12873,N_12760);
nand U12915 (N_12915,N_12876,N_12898);
or U12916 (N_12916,N_12826,N_12795);
nand U12917 (N_12917,N_12751,N_12822);
nor U12918 (N_12918,N_12783,N_12883);
nor U12919 (N_12919,N_12845,N_12856);
nor U12920 (N_12920,N_12836,N_12857);
and U12921 (N_12921,N_12755,N_12861);
nand U12922 (N_12922,N_12811,N_12814);
and U12923 (N_12923,N_12833,N_12882);
nor U12924 (N_12924,N_12807,N_12790);
and U12925 (N_12925,N_12854,N_12802);
xor U12926 (N_12926,N_12831,N_12868);
nor U12927 (N_12927,N_12763,N_12791);
nor U12928 (N_12928,N_12899,N_12771);
xor U12929 (N_12929,N_12858,N_12819);
and U12930 (N_12930,N_12794,N_12821);
xor U12931 (N_12931,N_12825,N_12896);
or U12932 (N_12932,N_12892,N_12840);
xnor U12933 (N_12933,N_12756,N_12810);
nor U12934 (N_12934,N_12801,N_12881);
nand U12935 (N_12935,N_12862,N_12784);
nor U12936 (N_12936,N_12788,N_12830);
and U12937 (N_12937,N_12808,N_12841);
or U12938 (N_12938,N_12780,N_12885);
nor U12939 (N_12939,N_12863,N_12800);
nand U12940 (N_12940,N_12829,N_12867);
xor U12941 (N_12941,N_12872,N_12828);
nor U12942 (N_12942,N_12812,N_12886);
nor U12943 (N_12943,N_12772,N_12893);
nor U12944 (N_12944,N_12793,N_12798);
nand U12945 (N_12945,N_12853,N_12827);
xnor U12946 (N_12946,N_12834,N_12809);
nor U12947 (N_12947,N_12843,N_12775);
or U12948 (N_12948,N_12759,N_12806);
nor U12949 (N_12949,N_12837,N_12750);
xnor U12950 (N_12950,N_12889,N_12792);
nor U12951 (N_12951,N_12782,N_12752);
nand U12952 (N_12952,N_12851,N_12758);
and U12953 (N_12953,N_12816,N_12817);
nor U12954 (N_12954,N_12890,N_12874);
and U12955 (N_12955,N_12770,N_12877);
nor U12956 (N_12956,N_12823,N_12767);
or U12957 (N_12957,N_12865,N_12773);
xnor U12958 (N_12958,N_12789,N_12866);
or U12959 (N_12959,N_12897,N_12768);
nor U12960 (N_12960,N_12820,N_12796);
nor U12961 (N_12961,N_12871,N_12878);
nor U12962 (N_12962,N_12864,N_12754);
nand U12963 (N_12963,N_12838,N_12870);
nor U12964 (N_12964,N_12813,N_12803);
nor U12965 (N_12965,N_12879,N_12850);
or U12966 (N_12966,N_12824,N_12844);
and U12967 (N_12967,N_12860,N_12765);
nand U12968 (N_12968,N_12894,N_12785);
nand U12969 (N_12969,N_12884,N_12805);
nor U12970 (N_12970,N_12849,N_12753);
xor U12971 (N_12971,N_12787,N_12891);
or U12972 (N_12972,N_12769,N_12779);
and U12973 (N_12973,N_12859,N_12799);
xnor U12974 (N_12974,N_12848,N_12766);
and U12975 (N_12975,N_12795,N_12868);
xnor U12976 (N_12976,N_12778,N_12786);
nand U12977 (N_12977,N_12872,N_12760);
xnor U12978 (N_12978,N_12799,N_12873);
nand U12979 (N_12979,N_12818,N_12885);
or U12980 (N_12980,N_12756,N_12836);
xnor U12981 (N_12981,N_12791,N_12800);
nand U12982 (N_12982,N_12810,N_12856);
nand U12983 (N_12983,N_12865,N_12898);
or U12984 (N_12984,N_12832,N_12860);
xor U12985 (N_12985,N_12874,N_12842);
nand U12986 (N_12986,N_12789,N_12880);
or U12987 (N_12987,N_12886,N_12834);
and U12988 (N_12988,N_12874,N_12778);
nor U12989 (N_12989,N_12777,N_12837);
nand U12990 (N_12990,N_12812,N_12821);
xnor U12991 (N_12991,N_12816,N_12806);
nor U12992 (N_12992,N_12779,N_12797);
xnor U12993 (N_12993,N_12832,N_12818);
and U12994 (N_12994,N_12884,N_12759);
nand U12995 (N_12995,N_12768,N_12844);
and U12996 (N_12996,N_12895,N_12795);
nand U12997 (N_12997,N_12807,N_12895);
or U12998 (N_12998,N_12799,N_12849);
xor U12999 (N_12999,N_12753,N_12870);
nand U13000 (N_13000,N_12857,N_12858);
and U13001 (N_13001,N_12892,N_12822);
nor U13002 (N_13002,N_12792,N_12815);
nand U13003 (N_13003,N_12770,N_12896);
nor U13004 (N_13004,N_12838,N_12840);
xnor U13005 (N_13005,N_12791,N_12860);
or U13006 (N_13006,N_12842,N_12885);
or U13007 (N_13007,N_12772,N_12888);
and U13008 (N_13008,N_12799,N_12856);
and U13009 (N_13009,N_12844,N_12804);
nor U13010 (N_13010,N_12791,N_12838);
xor U13011 (N_13011,N_12799,N_12827);
and U13012 (N_13012,N_12841,N_12881);
nor U13013 (N_13013,N_12816,N_12802);
and U13014 (N_13014,N_12860,N_12777);
xnor U13015 (N_13015,N_12841,N_12893);
or U13016 (N_13016,N_12795,N_12858);
or U13017 (N_13017,N_12824,N_12888);
nor U13018 (N_13018,N_12795,N_12799);
and U13019 (N_13019,N_12804,N_12792);
nand U13020 (N_13020,N_12787,N_12774);
nand U13021 (N_13021,N_12890,N_12877);
or U13022 (N_13022,N_12772,N_12805);
or U13023 (N_13023,N_12856,N_12850);
nor U13024 (N_13024,N_12864,N_12866);
xnor U13025 (N_13025,N_12823,N_12869);
and U13026 (N_13026,N_12838,N_12880);
xor U13027 (N_13027,N_12807,N_12810);
or U13028 (N_13028,N_12755,N_12832);
nand U13029 (N_13029,N_12868,N_12780);
nor U13030 (N_13030,N_12757,N_12855);
nand U13031 (N_13031,N_12771,N_12780);
xor U13032 (N_13032,N_12778,N_12812);
and U13033 (N_13033,N_12888,N_12803);
nor U13034 (N_13034,N_12807,N_12813);
nor U13035 (N_13035,N_12785,N_12881);
xor U13036 (N_13036,N_12789,N_12807);
or U13037 (N_13037,N_12853,N_12783);
and U13038 (N_13038,N_12801,N_12846);
and U13039 (N_13039,N_12811,N_12792);
nand U13040 (N_13040,N_12869,N_12782);
and U13041 (N_13041,N_12887,N_12761);
or U13042 (N_13042,N_12846,N_12861);
nand U13043 (N_13043,N_12850,N_12863);
nor U13044 (N_13044,N_12790,N_12770);
or U13045 (N_13045,N_12877,N_12792);
nand U13046 (N_13046,N_12857,N_12830);
or U13047 (N_13047,N_12788,N_12772);
nor U13048 (N_13048,N_12806,N_12752);
nor U13049 (N_13049,N_12880,N_12872);
nand U13050 (N_13050,N_12983,N_12904);
xor U13051 (N_13051,N_12934,N_13035);
or U13052 (N_13052,N_12972,N_12954);
nor U13053 (N_13053,N_12911,N_13013);
nand U13054 (N_13054,N_13032,N_12940);
nand U13055 (N_13055,N_12995,N_12919);
xor U13056 (N_13056,N_12909,N_13005);
xnor U13057 (N_13057,N_13016,N_13011);
or U13058 (N_13058,N_13006,N_13017);
nand U13059 (N_13059,N_13012,N_13027);
or U13060 (N_13060,N_12989,N_13039);
and U13061 (N_13061,N_12936,N_13023);
or U13062 (N_13062,N_13008,N_12969);
xor U13063 (N_13063,N_12959,N_12964);
xor U13064 (N_13064,N_12937,N_12963);
or U13065 (N_13065,N_12916,N_12952);
xor U13066 (N_13066,N_13003,N_13028);
nand U13067 (N_13067,N_13014,N_12961);
nand U13068 (N_13068,N_12902,N_12912);
or U13069 (N_13069,N_12933,N_12920);
nand U13070 (N_13070,N_12926,N_12988);
xnor U13071 (N_13071,N_12927,N_12976);
nand U13072 (N_13072,N_13045,N_12953);
and U13073 (N_13073,N_12985,N_12924);
nor U13074 (N_13074,N_13000,N_12977);
nand U13075 (N_13075,N_12950,N_13024);
or U13076 (N_13076,N_13046,N_12944);
nand U13077 (N_13077,N_12907,N_12984);
nor U13078 (N_13078,N_13020,N_12903);
and U13079 (N_13079,N_12962,N_12923);
nand U13080 (N_13080,N_13049,N_13030);
nand U13081 (N_13081,N_13007,N_13010);
xnor U13082 (N_13082,N_12979,N_12935);
and U13083 (N_13083,N_13026,N_12941);
xor U13084 (N_13084,N_12922,N_13042);
nor U13085 (N_13085,N_12967,N_13037);
nor U13086 (N_13086,N_12978,N_13001);
or U13087 (N_13087,N_12982,N_12973);
and U13088 (N_13088,N_13040,N_12914);
xnor U13089 (N_13089,N_12946,N_13002);
and U13090 (N_13090,N_13025,N_12913);
and U13091 (N_13091,N_12996,N_12993);
xnor U13092 (N_13092,N_13048,N_12947);
and U13093 (N_13093,N_12921,N_12999);
nor U13094 (N_13094,N_12997,N_12929);
nand U13095 (N_13095,N_13015,N_12932);
nor U13096 (N_13096,N_12928,N_12992);
xor U13097 (N_13097,N_12948,N_12930);
nor U13098 (N_13098,N_12970,N_13019);
or U13099 (N_13099,N_12949,N_12971);
nor U13100 (N_13100,N_12975,N_13034);
or U13101 (N_13101,N_12968,N_13033);
xnor U13102 (N_13102,N_13044,N_13021);
nand U13103 (N_13103,N_12957,N_12945);
nand U13104 (N_13104,N_12900,N_12956);
or U13105 (N_13105,N_12980,N_13047);
nand U13106 (N_13106,N_12960,N_12931);
nand U13107 (N_13107,N_13018,N_13041);
and U13108 (N_13108,N_12942,N_13031);
xor U13109 (N_13109,N_13036,N_12986);
nand U13110 (N_13110,N_12906,N_12998);
nand U13111 (N_13111,N_12955,N_12905);
or U13112 (N_13112,N_13022,N_12958);
nand U13113 (N_13113,N_13038,N_12939);
nand U13114 (N_13114,N_12917,N_12910);
xor U13115 (N_13115,N_12938,N_12994);
nor U13116 (N_13116,N_13029,N_12974);
nor U13117 (N_13117,N_12966,N_12915);
nor U13118 (N_13118,N_12925,N_13004);
nor U13119 (N_13119,N_12987,N_12965);
nand U13120 (N_13120,N_13009,N_12990);
and U13121 (N_13121,N_12981,N_12908);
or U13122 (N_13122,N_12991,N_13043);
or U13123 (N_13123,N_12901,N_12918);
or U13124 (N_13124,N_12943,N_12951);
and U13125 (N_13125,N_12980,N_12967);
nor U13126 (N_13126,N_12997,N_13046);
or U13127 (N_13127,N_13035,N_12957);
nor U13128 (N_13128,N_12973,N_13011);
xor U13129 (N_13129,N_12986,N_13023);
nor U13130 (N_13130,N_12971,N_12952);
xnor U13131 (N_13131,N_13028,N_12981);
or U13132 (N_13132,N_13020,N_12991);
xor U13133 (N_13133,N_12923,N_12909);
or U13134 (N_13134,N_12902,N_12903);
nand U13135 (N_13135,N_13021,N_12926);
nor U13136 (N_13136,N_13040,N_13035);
or U13137 (N_13137,N_13015,N_13002);
or U13138 (N_13138,N_13026,N_12978);
nor U13139 (N_13139,N_13037,N_12902);
nand U13140 (N_13140,N_12971,N_12975);
nand U13141 (N_13141,N_12946,N_12950);
and U13142 (N_13142,N_12913,N_13035);
xor U13143 (N_13143,N_12928,N_12920);
and U13144 (N_13144,N_13011,N_12917);
or U13145 (N_13145,N_12944,N_12980);
or U13146 (N_13146,N_12905,N_12965);
nor U13147 (N_13147,N_12949,N_12969);
xor U13148 (N_13148,N_12929,N_13047);
and U13149 (N_13149,N_13008,N_13003);
nand U13150 (N_13150,N_12950,N_13012);
nand U13151 (N_13151,N_12955,N_13040);
nand U13152 (N_13152,N_12953,N_13015);
and U13153 (N_13153,N_12942,N_12967);
xor U13154 (N_13154,N_12996,N_12908);
and U13155 (N_13155,N_12969,N_12987);
or U13156 (N_13156,N_13011,N_12908);
xnor U13157 (N_13157,N_12981,N_13035);
and U13158 (N_13158,N_13021,N_12989);
nor U13159 (N_13159,N_12986,N_13021);
xor U13160 (N_13160,N_13036,N_12946);
and U13161 (N_13161,N_13013,N_13018);
and U13162 (N_13162,N_12986,N_12910);
nor U13163 (N_13163,N_12923,N_13033);
or U13164 (N_13164,N_12980,N_12954);
and U13165 (N_13165,N_13001,N_12947);
and U13166 (N_13166,N_12931,N_13016);
nor U13167 (N_13167,N_13003,N_12979);
nor U13168 (N_13168,N_12904,N_13005);
and U13169 (N_13169,N_12987,N_12922);
nand U13170 (N_13170,N_12992,N_13020);
nor U13171 (N_13171,N_13011,N_12901);
and U13172 (N_13172,N_13026,N_13015);
or U13173 (N_13173,N_12953,N_12914);
nor U13174 (N_13174,N_12998,N_13011);
nand U13175 (N_13175,N_12962,N_12972);
and U13176 (N_13176,N_12918,N_13013);
xor U13177 (N_13177,N_13011,N_13044);
and U13178 (N_13178,N_12954,N_12940);
nor U13179 (N_13179,N_12945,N_12983);
nor U13180 (N_13180,N_12963,N_13001);
nor U13181 (N_13181,N_12989,N_12904);
nor U13182 (N_13182,N_12929,N_12975);
or U13183 (N_13183,N_13019,N_13021);
and U13184 (N_13184,N_12969,N_13041);
xnor U13185 (N_13185,N_12950,N_12967);
nor U13186 (N_13186,N_13002,N_13004);
nor U13187 (N_13187,N_12965,N_12903);
or U13188 (N_13188,N_12981,N_12960);
xor U13189 (N_13189,N_12987,N_12997);
nor U13190 (N_13190,N_12998,N_12949);
or U13191 (N_13191,N_12961,N_13020);
nand U13192 (N_13192,N_13012,N_12993);
or U13193 (N_13193,N_12923,N_13034);
and U13194 (N_13194,N_12983,N_12932);
xnor U13195 (N_13195,N_12957,N_12962);
xor U13196 (N_13196,N_12968,N_12938);
nand U13197 (N_13197,N_13000,N_12973);
nor U13198 (N_13198,N_12960,N_13025);
nor U13199 (N_13199,N_12979,N_12956);
or U13200 (N_13200,N_13145,N_13188);
nor U13201 (N_13201,N_13055,N_13162);
and U13202 (N_13202,N_13153,N_13062);
nand U13203 (N_13203,N_13111,N_13135);
and U13204 (N_13204,N_13097,N_13142);
xor U13205 (N_13205,N_13167,N_13138);
nand U13206 (N_13206,N_13171,N_13098);
nand U13207 (N_13207,N_13181,N_13106);
xor U13208 (N_13208,N_13050,N_13095);
nor U13209 (N_13209,N_13114,N_13078);
or U13210 (N_13210,N_13184,N_13169);
or U13211 (N_13211,N_13179,N_13122);
or U13212 (N_13212,N_13096,N_13063);
xor U13213 (N_13213,N_13189,N_13126);
xor U13214 (N_13214,N_13185,N_13118);
nand U13215 (N_13215,N_13128,N_13132);
nand U13216 (N_13216,N_13084,N_13140);
and U13217 (N_13217,N_13087,N_13182);
and U13218 (N_13218,N_13100,N_13147);
and U13219 (N_13219,N_13198,N_13081);
xnor U13220 (N_13220,N_13108,N_13115);
and U13221 (N_13221,N_13121,N_13168);
or U13222 (N_13222,N_13061,N_13148);
nor U13223 (N_13223,N_13089,N_13119);
xnor U13224 (N_13224,N_13131,N_13161);
nor U13225 (N_13225,N_13064,N_13065);
xnor U13226 (N_13226,N_13123,N_13165);
nor U13227 (N_13227,N_13112,N_13074);
and U13228 (N_13228,N_13116,N_13125);
nor U13229 (N_13229,N_13066,N_13175);
nand U13230 (N_13230,N_13129,N_13173);
nor U13231 (N_13231,N_13052,N_13152);
nand U13232 (N_13232,N_13192,N_13177);
xor U13233 (N_13233,N_13083,N_13154);
nor U13234 (N_13234,N_13183,N_13059);
nand U13235 (N_13235,N_13102,N_13105);
and U13236 (N_13236,N_13190,N_13104);
nor U13237 (N_13237,N_13159,N_13054);
xnor U13238 (N_13238,N_13107,N_13178);
nand U13239 (N_13239,N_13070,N_13130);
or U13240 (N_13240,N_13150,N_13156);
xnor U13241 (N_13241,N_13149,N_13146);
nand U13242 (N_13242,N_13163,N_13199);
or U13243 (N_13243,N_13186,N_13093);
xnor U13244 (N_13244,N_13197,N_13174);
nor U13245 (N_13245,N_13109,N_13164);
nand U13246 (N_13246,N_13071,N_13155);
nand U13247 (N_13247,N_13110,N_13172);
or U13248 (N_13248,N_13144,N_13139);
nor U13249 (N_13249,N_13193,N_13073);
nand U13250 (N_13250,N_13053,N_13127);
nand U13251 (N_13251,N_13091,N_13137);
or U13252 (N_13252,N_13079,N_13117);
nor U13253 (N_13253,N_13090,N_13151);
and U13254 (N_13254,N_13088,N_13158);
xnor U13255 (N_13255,N_13166,N_13191);
xor U13256 (N_13256,N_13060,N_13051);
or U13257 (N_13257,N_13056,N_13094);
nand U13258 (N_13258,N_13170,N_13076);
xor U13259 (N_13259,N_13176,N_13082);
xor U13260 (N_13260,N_13136,N_13103);
nand U13261 (N_13261,N_13134,N_13120);
or U13262 (N_13262,N_13157,N_13057);
xor U13263 (N_13263,N_13077,N_13067);
xnor U13264 (N_13264,N_13086,N_13187);
nor U13265 (N_13265,N_13069,N_13143);
nor U13266 (N_13266,N_13141,N_13160);
nor U13267 (N_13267,N_13195,N_13196);
and U13268 (N_13268,N_13101,N_13113);
nor U13269 (N_13269,N_13133,N_13194);
and U13270 (N_13270,N_13080,N_13124);
and U13271 (N_13271,N_13092,N_13180);
and U13272 (N_13272,N_13058,N_13099);
nand U13273 (N_13273,N_13085,N_13072);
xnor U13274 (N_13274,N_13075,N_13068);
xor U13275 (N_13275,N_13076,N_13140);
nand U13276 (N_13276,N_13051,N_13168);
or U13277 (N_13277,N_13179,N_13173);
xor U13278 (N_13278,N_13169,N_13116);
xor U13279 (N_13279,N_13157,N_13180);
nor U13280 (N_13280,N_13101,N_13162);
and U13281 (N_13281,N_13189,N_13148);
or U13282 (N_13282,N_13134,N_13140);
or U13283 (N_13283,N_13058,N_13145);
or U13284 (N_13284,N_13054,N_13051);
and U13285 (N_13285,N_13150,N_13078);
nand U13286 (N_13286,N_13144,N_13113);
nand U13287 (N_13287,N_13115,N_13179);
nor U13288 (N_13288,N_13111,N_13140);
nand U13289 (N_13289,N_13081,N_13101);
and U13290 (N_13290,N_13063,N_13146);
or U13291 (N_13291,N_13161,N_13184);
nor U13292 (N_13292,N_13162,N_13082);
xor U13293 (N_13293,N_13119,N_13077);
xnor U13294 (N_13294,N_13093,N_13122);
or U13295 (N_13295,N_13115,N_13164);
nand U13296 (N_13296,N_13057,N_13145);
xnor U13297 (N_13297,N_13092,N_13183);
nand U13298 (N_13298,N_13155,N_13157);
or U13299 (N_13299,N_13152,N_13169);
nand U13300 (N_13300,N_13081,N_13177);
xnor U13301 (N_13301,N_13093,N_13070);
nor U13302 (N_13302,N_13102,N_13130);
or U13303 (N_13303,N_13083,N_13147);
nand U13304 (N_13304,N_13185,N_13120);
nor U13305 (N_13305,N_13148,N_13164);
or U13306 (N_13306,N_13177,N_13096);
nand U13307 (N_13307,N_13104,N_13194);
nand U13308 (N_13308,N_13084,N_13149);
nand U13309 (N_13309,N_13082,N_13065);
nor U13310 (N_13310,N_13071,N_13125);
nor U13311 (N_13311,N_13077,N_13063);
and U13312 (N_13312,N_13161,N_13098);
and U13313 (N_13313,N_13152,N_13164);
or U13314 (N_13314,N_13051,N_13192);
or U13315 (N_13315,N_13189,N_13156);
xnor U13316 (N_13316,N_13053,N_13118);
and U13317 (N_13317,N_13162,N_13099);
and U13318 (N_13318,N_13090,N_13168);
nor U13319 (N_13319,N_13153,N_13133);
nand U13320 (N_13320,N_13193,N_13134);
and U13321 (N_13321,N_13077,N_13157);
nand U13322 (N_13322,N_13195,N_13148);
nand U13323 (N_13323,N_13164,N_13198);
xnor U13324 (N_13324,N_13099,N_13123);
and U13325 (N_13325,N_13159,N_13168);
nor U13326 (N_13326,N_13163,N_13194);
nor U13327 (N_13327,N_13176,N_13162);
nor U13328 (N_13328,N_13193,N_13150);
nor U13329 (N_13329,N_13090,N_13098);
or U13330 (N_13330,N_13125,N_13120);
nor U13331 (N_13331,N_13110,N_13134);
nor U13332 (N_13332,N_13186,N_13106);
and U13333 (N_13333,N_13070,N_13143);
nor U13334 (N_13334,N_13108,N_13107);
nor U13335 (N_13335,N_13117,N_13056);
xnor U13336 (N_13336,N_13175,N_13128);
xnor U13337 (N_13337,N_13063,N_13167);
or U13338 (N_13338,N_13145,N_13182);
or U13339 (N_13339,N_13143,N_13125);
and U13340 (N_13340,N_13199,N_13194);
nor U13341 (N_13341,N_13142,N_13060);
or U13342 (N_13342,N_13180,N_13145);
nor U13343 (N_13343,N_13104,N_13170);
nand U13344 (N_13344,N_13070,N_13056);
or U13345 (N_13345,N_13150,N_13057);
or U13346 (N_13346,N_13169,N_13067);
nand U13347 (N_13347,N_13084,N_13137);
or U13348 (N_13348,N_13175,N_13095);
nand U13349 (N_13349,N_13144,N_13189);
nor U13350 (N_13350,N_13258,N_13239);
and U13351 (N_13351,N_13333,N_13341);
xor U13352 (N_13352,N_13306,N_13284);
nor U13353 (N_13353,N_13238,N_13346);
or U13354 (N_13354,N_13293,N_13233);
nand U13355 (N_13355,N_13254,N_13231);
nor U13356 (N_13356,N_13323,N_13281);
and U13357 (N_13357,N_13348,N_13286);
xnor U13358 (N_13358,N_13222,N_13225);
nor U13359 (N_13359,N_13344,N_13328);
and U13360 (N_13360,N_13315,N_13202);
or U13361 (N_13361,N_13305,N_13287);
and U13362 (N_13362,N_13329,N_13327);
and U13363 (N_13363,N_13252,N_13249);
nand U13364 (N_13364,N_13331,N_13257);
xnor U13365 (N_13365,N_13265,N_13312);
and U13366 (N_13366,N_13277,N_13299);
or U13367 (N_13367,N_13313,N_13227);
nor U13368 (N_13368,N_13342,N_13269);
xor U13369 (N_13369,N_13274,N_13235);
or U13370 (N_13370,N_13263,N_13345);
nand U13371 (N_13371,N_13326,N_13273);
nor U13372 (N_13372,N_13336,N_13237);
nor U13373 (N_13373,N_13212,N_13217);
or U13374 (N_13374,N_13279,N_13247);
nand U13375 (N_13375,N_13285,N_13295);
nor U13376 (N_13376,N_13275,N_13278);
and U13377 (N_13377,N_13349,N_13325);
nor U13378 (N_13378,N_13241,N_13259);
nand U13379 (N_13379,N_13322,N_13206);
nand U13380 (N_13380,N_13207,N_13297);
and U13381 (N_13381,N_13256,N_13210);
and U13382 (N_13382,N_13260,N_13298);
nor U13383 (N_13383,N_13203,N_13221);
nand U13384 (N_13384,N_13282,N_13264);
nor U13385 (N_13385,N_13316,N_13208);
and U13386 (N_13386,N_13245,N_13223);
xnor U13387 (N_13387,N_13334,N_13300);
nand U13388 (N_13388,N_13229,N_13304);
nor U13389 (N_13389,N_13292,N_13253);
xnor U13390 (N_13390,N_13337,N_13209);
or U13391 (N_13391,N_13251,N_13340);
nor U13392 (N_13392,N_13219,N_13332);
xor U13393 (N_13393,N_13215,N_13204);
nor U13394 (N_13394,N_13224,N_13214);
nand U13395 (N_13395,N_13220,N_13216);
xnor U13396 (N_13396,N_13213,N_13244);
and U13397 (N_13397,N_13320,N_13271);
or U13398 (N_13398,N_13319,N_13347);
nor U13399 (N_13399,N_13294,N_13262);
and U13400 (N_13400,N_13226,N_13283);
nand U13401 (N_13401,N_13311,N_13267);
and U13402 (N_13402,N_13291,N_13230);
nand U13403 (N_13403,N_13242,N_13270);
nor U13404 (N_13404,N_13310,N_13308);
or U13405 (N_13405,N_13218,N_13288);
and U13406 (N_13406,N_13324,N_13314);
or U13407 (N_13407,N_13211,N_13205);
and U13408 (N_13408,N_13303,N_13268);
nor U13409 (N_13409,N_13201,N_13330);
nor U13410 (N_13410,N_13289,N_13296);
and U13411 (N_13411,N_13276,N_13234);
and U13412 (N_13412,N_13321,N_13339);
or U13413 (N_13413,N_13240,N_13301);
nand U13414 (N_13414,N_13343,N_13309);
nor U13415 (N_13415,N_13280,N_13335);
and U13416 (N_13416,N_13236,N_13290);
or U13417 (N_13417,N_13317,N_13266);
xnor U13418 (N_13418,N_13243,N_13248);
xor U13419 (N_13419,N_13272,N_13261);
nand U13420 (N_13420,N_13302,N_13246);
xor U13421 (N_13421,N_13255,N_13228);
nor U13422 (N_13422,N_13307,N_13338);
or U13423 (N_13423,N_13232,N_13318);
nor U13424 (N_13424,N_13250,N_13200);
and U13425 (N_13425,N_13290,N_13287);
or U13426 (N_13426,N_13291,N_13347);
xnor U13427 (N_13427,N_13207,N_13220);
nand U13428 (N_13428,N_13313,N_13231);
nand U13429 (N_13429,N_13257,N_13282);
nor U13430 (N_13430,N_13312,N_13325);
xnor U13431 (N_13431,N_13215,N_13208);
and U13432 (N_13432,N_13271,N_13222);
nor U13433 (N_13433,N_13336,N_13327);
nand U13434 (N_13434,N_13333,N_13320);
xnor U13435 (N_13435,N_13275,N_13336);
nand U13436 (N_13436,N_13257,N_13336);
and U13437 (N_13437,N_13314,N_13302);
nand U13438 (N_13438,N_13284,N_13258);
or U13439 (N_13439,N_13293,N_13227);
xor U13440 (N_13440,N_13329,N_13283);
or U13441 (N_13441,N_13331,N_13297);
xnor U13442 (N_13442,N_13204,N_13292);
xnor U13443 (N_13443,N_13239,N_13266);
nor U13444 (N_13444,N_13346,N_13275);
nor U13445 (N_13445,N_13221,N_13334);
nand U13446 (N_13446,N_13219,N_13215);
nor U13447 (N_13447,N_13300,N_13263);
xor U13448 (N_13448,N_13233,N_13248);
nor U13449 (N_13449,N_13328,N_13217);
xor U13450 (N_13450,N_13297,N_13312);
or U13451 (N_13451,N_13235,N_13256);
and U13452 (N_13452,N_13287,N_13223);
nand U13453 (N_13453,N_13304,N_13291);
xnor U13454 (N_13454,N_13321,N_13332);
and U13455 (N_13455,N_13261,N_13226);
nor U13456 (N_13456,N_13341,N_13303);
xnor U13457 (N_13457,N_13347,N_13216);
and U13458 (N_13458,N_13275,N_13296);
and U13459 (N_13459,N_13344,N_13306);
nor U13460 (N_13460,N_13310,N_13314);
nand U13461 (N_13461,N_13312,N_13264);
xnor U13462 (N_13462,N_13204,N_13276);
or U13463 (N_13463,N_13317,N_13315);
nand U13464 (N_13464,N_13234,N_13335);
nand U13465 (N_13465,N_13244,N_13328);
nor U13466 (N_13466,N_13298,N_13310);
nand U13467 (N_13467,N_13278,N_13291);
xnor U13468 (N_13468,N_13201,N_13240);
xnor U13469 (N_13469,N_13302,N_13248);
nand U13470 (N_13470,N_13221,N_13315);
nor U13471 (N_13471,N_13273,N_13249);
nor U13472 (N_13472,N_13348,N_13287);
xor U13473 (N_13473,N_13318,N_13308);
xnor U13474 (N_13474,N_13250,N_13304);
and U13475 (N_13475,N_13299,N_13260);
or U13476 (N_13476,N_13290,N_13241);
nor U13477 (N_13477,N_13311,N_13209);
xor U13478 (N_13478,N_13267,N_13225);
and U13479 (N_13479,N_13337,N_13330);
xor U13480 (N_13480,N_13272,N_13326);
or U13481 (N_13481,N_13300,N_13268);
or U13482 (N_13482,N_13312,N_13273);
and U13483 (N_13483,N_13268,N_13312);
and U13484 (N_13484,N_13250,N_13223);
nor U13485 (N_13485,N_13292,N_13305);
nor U13486 (N_13486,N_13215,N_13302);
xor U13487 (N_13487,N_13229,N_13255);
nor U13488 (N_13488,N_13295,N_13243);
nand U13489 (N_13489,N_13242,N_13334);
and U13490 (N_13490,N_13328,N_13234);
nor U13491 (N_13491,N_13234,N_13232);
nor U13492 (N_13492,N_13215,N_13209);
or U13493 (N_13493,N_13292,N_13299);
and U13494 (N_13494,N_13236,N_13221);
nand U13495 (N_13495,N_13235,N_13262);
and U13496 (N_13496,N_13220,N_13310);
xnor U13497 (N_13497,N_13289,N_13298);
nor U13498 (N_13498,N_13203,N_13342);
and U13499 (N_13499,N_13257,N_13292);
xor U13500 (N_13500,N_13388,N_13461);
nor U13501 (N_13501,N_13493,N_13387);
or U13502 (N_13502,N_13409,N_13450);
and U13503 (N_13503,N_13437,N_13359);
nand U13504 (N_13504,N_13438,N_13463);
nor U13505 (N_13505,N_13404,N_13423);
nand U13506 (N_13506,N_13458,N_13466);
and U13507 (N_13507,N_13371,N_13453);
or U13508 (N_13508,N_13370,N_13369);
xnor U13509 (N_13509,N_13407,N_13383);
and U13510 (N_13510,N_13478,N_13403);
xor U13511 (N_13511,N_13491,N_13352);
or U13512 (N_13512,N_13376,N_13467);
or U13513 (N_13513,N_13373,N_13397);
or U13514 (N_13514,N_13468,N_13406);
and U13515 (N_13515,N_13424,N_13457);
nand U13516 (N_13516,N_13364,N_13497);
nand U13517 (N_13517,N_13474,N_13431);
nor U13518 (N_13518,N_13413,N_13402);
xor U13519 (N_13519,N_13480,N_13494);
nand U13520 (N_13520,N_13429,N_13469);
and U13521 (N_13521,N_13483,N_13390);
xnor U13522 (N_13522,N_13433,N_13385);
nor U13523 (N_13523,N_13356,N_13486);
nand U13524 (N_13524,N_13355,N_13477);
xnor U13525 (N_13525,N_13354,N_13363);
nand U13526 (N_13526,N_13412,N_13394);
xnor U13527 (N_13527,N_13482,N_13396);
nor U13528 (N_13528,N_13445,N_13451);
xor U13529 (N_13529,N_13464,N_13426);
xor U13530 (N_13530,N_13441,N_13484);
nand U13531 (N_13531,N_13471,N_13470);
xnor U13532 (N_13532,N_13473,N_13417);
nor U13533 (N_13533,N_13416,N_13420);
nor U13534 (N_13534,N_13411,N_13414);
nand U13535 (N_13535,N_13479,N_13380);
xnor U13536 (N_13536,N_13487,N_13395);
nor U13537 (N_13537,N_13350,N_13361);
or U13538 (N_13538,N_13456,N_13442);
nor U13539 (N_13539,N_13428,N_13408);
or U13540 (N_13540,N_13365,N_13489);
nor U13541 (N_13541,N_13384,N_13372);
nor U13542 (N_13542,N_13422,N_13435);
nand U13543 (N_13543,N_13386,N_13398);
xnor U13544 (N_13544,N_13440,N_13400);
nand U13545 (N_13545,N_13377,N_13462);
or U13546 (N_13546,N_13434,N_13382);
and U13547 (N_13547,N_13454,N_13446);
or U13548 (N_13548,N_13360,N_13391);
nand U13549 (N_13549,N_13472,N_13410);
nand U13550 (N_13550,N_13436,N_13379);
xnor U13551 (N_13551,N_13476,N_13358);
nor U13552 (N_13552,N_13465,N_13375);
nor U13553 (N_13553,N_13392,N_13378);
nand U13554 (N_13554,N_13374,N_13492);
nand U13555 (N_13555,N_13460,N_13439);
or U13556 (N_13556,N_13389,N_13393);
nand U13557 (N_13557,N_13490,N_13401);
or U13558 (N_13558,N_13447,N_13427);
xnor U13559 (N_13559,N_13481,N_13368);
or U13560 (N_13560,N_13475,N_13351);
nor U13561 (N_13561,N_13357,N_13448);
or U13562 (N_13562,N_13499,N_13399);
or U13563 (N_13563,N_13459,N_13498);
and U13564 (N_13564,N_13425,N_13353);
and U13565 (N_13565,N_13381,N_13367);
nand U13566 (N_13566,N_13418,N_13449);
xor U13567 (N_13567,N_13366,N_13455);
nand U13568 (N_13568,N_13362,N_13405);
xnor U13569 (N_13569,N_13443,N_13419);
xnor U13570 (N_13570,N_13430,N_13488);
nand U13571 (N_13571,N_13452,N_13415);
and U13572 (N_13572,N_13432,N_13495);
nor U13573 (N_13573,N_13421,N_13485);
nand U13574 (N_13574,N_13444,N_13496);
xor U13575 (N_13575,N_13409,N_13404);
nand U13576 (N_13576,N_13499,N_13364);
xor U13577 (N_13577,N_13472,N_13355);
or U13578 (N_13578,N_13359,N_13460);
and U13579 (N_13579,N_13368,N_13447);
or U13580 (N_13580,N_13361,N_13381);
and U13581 (N_13581,N_13376,N_13473);
xor U13582 (N_13582,N_13432,N_13350);
or U13583 (N_13583,N_13480,N_13459);
and U13584 (N_13584,N_13391,N_13378);
or U13585 (N_13585,N_13355,N_13461);
xnor U13586 (N_13586,N_13375,N_13448);
xnor U13587 (N_13587,N_13480,N_13491);
or U13588 (N_13588,N_13408,N_13363);
nand U13589 (N_13589,N_13479,N_13456);
nand U13590 (N_13590,N_13368,N_13397);
and U13591 (N_13591,N_13377,N_13469);
nand U13592 (N_13592,N_13433,N_13382);
nand U13593 (N_13593,N_13395,N_13368);
xnor U13594 (N_13594,N_13371,N_13499);
xor U13595 (N_13595,N_13387,N_13421);
and U13596 (N_13596,N_13402,N_13423);
and U13597 (N_13597,N_13437,N_13442);
or U13598 (N_13598,N_13439,N_13382);
nand U13599 (N_13599,N_13411,N_13364);
and U13600 (N_13600,N_13372,N_13409);
or U13601 (N_13601,N_13477,N_13424);
or U13602 (N_13602,N_13472,N_13401);
nor U13603 (N_13603,N_13351,N_13476);
nand U13604 (N_13604,N_13497,N_13477);
xor U13605 (N_13605,N_13371,N_13420);
nand U13606 (N_13606,N_13353,N_13393);
nand U13607 (N_13607,N_13439,N_13437);
nand U13608 (N_13608,N_13487,N_13389);
nor U13609 (N_13609,N_13362,N_13402);
xor U13610 (N_13610,N_13366,N_13489);
xor U13611 (N_13611,N_13423,N_13377);
and U13612 (N_13612,N_13442,N_13475);
nor U13613 (N_13613,N_13476,N_13440);
xnor U13614 (N_13614,N_13467,N_13454);
or U13615 (N_13615,N_13408,N_13497);
nor U13616 (N_13616,N_13480,N_13359);
nand U13617 (N_13617,N_13355,N_13439);
nor U13618 (N_13618,N_13350,N_13447);
nand U13619 (N_13619,N_13474,N_13396);
xnor U13620 (N_13620,N_13499,N_13362);
nor U13621 (N_13621,N_13378,N_13421);
and U13622 (N_13622,N_13497,N_13480);
nor U13623 (N_13623,N_13371,N_13387);
nor U13624 (N_13624,N_13376,N_13474);
and U13625 (N_13625,N_13369,N_13465);
xor U13626 (N_13626,N_13472,N_13354);
and U13627 (N_13627,N_13476,N_13382);
and U13628 (N_13628,N_13491,N_13397);
and U13629 (N_13629,N_13407,N_13473);
nand U13630 (N_13630,N_13491,N_13355);
and U13631 (N_13631,N_13428,N_13374);
nand U13632 (N_13632,N_13354,N_13375);
xor U13633 (N_13633,N_13416,N_13378);
nor U13634 (N_13634,N_13401,N_13363);
xor U13635 (N_13635,N_13355,N_13372);
nand U13636 (N_13636,N_13420,N_13358);
nor U13637 (N_13637,N_13398,N_13385);
nor U13638 (N_13638,N_13378,N_13351);
xnor U13639 (N_13639,N_13397,N_13367);
nand U13640 (N_13640,N_13355,N_13357);
nor U13641 (N_13641,N_13454,N_13438);
or U13642 (N_13642,N_13385,N_13389);
nor U13643 (N_13643,N_13429,N_13383);
xnor U13644 (N_13644,N_13391,N_13413);
and U13645 (N_13645,N_13370,N_13404);
nor U13646 (N_13646,N_13420,N_13359);
or U13647 (N_13647,N_13487,N_13430);
nor U13648 (N_13648,N_13479,N_13426);
nand U13649 (N_13649,N_13415,N_13449);
nor U13650 (N_13650,N_13589,N_13509);
xor U13651 (N_13651,N_13588,N_13501);
xnor U13652 (N_13652,N_13599,N_13641);
nor U13653 (N_13653,N_13594,N_13633);
nand U13654 (N_13654,N_13643,N_13518);
or U13655 (N_13655,N_13598,N_13563);
nor U13656 (N_13656,N_13549,N_13559);
xnor U13657 (N_13657,N_13502,N_13521);
or U13658 (N_13658,N_13620,N_13625);
or U13659 (N_13659,N_13531,N_13503);
xor U13660 (N_13660,N_13606,N_13603);
xnor U13661 (N_13661,N_13539,N_13601);
nor U13662 (N_13662,N_13542,N_13635);
and U13663 (N_13663,N_13565,N_13578);
xor U13664 (N_13664,N_13617,N_13622);
xor U13665 (N_13665,N_13611,N_13607);
nand U13666 (N_13666,N_13519,N_13616);
xor U13667 (N_13667,N_13591,N_13645);
xor U13668 (N_13668,N_13555,N_13592);
nand U13669 (N_13669,N_13574,N_13582);
xnor U13670 (N_13670,N_13567,N_13514);
nand U13671 (N_13671,N_13564,N_13560);
nor U13672 (N_13672,N_13571,N_13543);
nor U13673 (N_13673,N_13642,N_13553);
nor U13674 (N_13674,N_13538,N_13596);
nor U13675 (N_13675,N_13528,N_13638);
nor U13676 (N_13676,N_13546,N_13587);
and U13677 (N_13677,N_13536,N_13644);
nand U13678 (N_13678,N_13551,N_13597);
nand U13679 (N_13679,N_13628,N_13586);
nor U13680 (N_13680,N_13580,N_13516);
xor U13681 (N_13681,N_13605,N_13585);
nor U13682 (N_13682,N_13508,N_13634);
and U13683 (N_13683,N_13557,N_13590);
or U13684 (N_13684,N_13513,N_13612);
or U13685 (N_13685,N_13547,N_13602);
or U13686 (N_13686,N_13604,N_13523);
or U13687 (N_13687,N_13629,N_13554);
and U13688 (N_13688,N_13600,N_13627);
xor U13689 (N_13689,N_13529,N_13530);
xnor U13690 (N_13690,N_13608,N_13515);
or U13691 (N_13691,N_13630,N_13526);
nand U13692 (N_13692,N_13632,N_13570);
nand U13693 (N_13693,N_13584,N_13639);
and U13694 (N_13694,N_13637,N_13505);
nand U13695 (N_13695,N_13581,N_13506);
nand U13696 (N_13696,N_13613,N_13533);
xor U13697 (N_13697,N_13540,N_13534);
nand U13698 (N_13698,N_13647,N_13576);
nand U13699 (N_13699,N_13512,N_13572);
or U13700 (N_13700,N_13541,N_13626);
nand U13701 (N_13701,N_13621,N_13568);
xnor U13702 (N_13702,N_13558,N_13579);
or U13703 (N_13703,N_13552,N_13562);
and U13704 (N_13704,N_13544,N_13636);
nand U13705 (N_13705,N_13561,N_13583);
xor U13706 (N_13706,N_13537,N_13510);
and U13707 (N_13707,N_13648,N_13504);
nand U13708 (N_13708,N_13615,N_13610);
and U13709 (N_13709,N_13573,N_13619);
nor U13710 (N_13710,N_13525,N_13566);
and U13711 (N_13711,N_13624,N_13507);
or U13712 (N_13712,N_13623,N_13646);
nor U13713 (N_13713,N_13614,N_13556);
nand U13714 (N_13714,N_13640,N_13527);
nor U13715 (N_13715,N_13569,N_13593);
and U13716 (N_13716,N_13524,N_13649);
or U13717 (N_13717,N_13609,N_13511);
nor U13718 (N_13718,N_13618,N_13631);
nand U13719 (N_13719,N_13595,N_13535);
and U13720 (N_13720,N_13575,N_13500);
nand U13721 (N_13721,N_13545,N_13550);
and U13722 (N_13722,N_13548,N_13532);
nor U13723 (N_13723,N_13522,N_13517);
nor U13724 (N_13724,N_13577,N_13520);
nand U13725 (N_13725,N_13607,N_13536);
and U13726 (N_13726,N_13511,N_13578);
and U13727 (N_13727,N_13624,N_13616);
nor U13728 (N_13728,N_13521,N_13576);
nor U13729 (N_13729,N_13517,N_13614);
or U13730 (N_13730,N_13603,N_13500);
and U13731 (N_13731,N_13637,N_13600);
or U13732 (N_13732,N_13627,N_13609);
or U13733 (N_13733,N_13587,N_13645);
nand U13734 (N_13734,N_13522,N_13587);
nand U13735 (N_13735,N_13633,N_13606);
nor U13736 (N_13736,N_13516,N_13605);
or U13737 (N_13737,N_13597,N_13585);
and U13738 (N_13738,N_13585,N_13548);
xor U13739 (N_13739,N_13594,N_13549);
xnor U13740 (N_13740,N_13606,N_13621);
nand U13741 (N_13741,N_13640,N_13553);
nor U13742 (N_13742,N_13528,N_13570);
xor U13743 (N_13743,N_13528,N_13531);
xnor U13744 (N_13744,N_13586,N_13541);
and U13745 (N_13745,N_13555,N_13547);
and U13746 (N_13746,N_13572,N_13513);
and U13747 (N_13747,N_13559,N_13622);
nor U13748 (N_13748,N_13557,N_13580);
nor U13749 (N_13749,N_13551,N_13598);
nor U13750 (N_13750,N_13564,N_13573);
or U13751 (N_13751,N_13625,N_13525);
or U13752 (N_13752,N_13546,N_13509);
nand U13753 (N_13753,N_13644,N_13531);
nor U13754 (N_13754,N_13615,N_13504);
and U13755 (N_13755,N_13580,N_13508);
nand U13756 (N_13756,N_13631,N_13531);
nand U13757 (N_13757,N_13592,N_13596);
xnor U13758 (N_13758,N_13585,N_13554);
nor U13759 (N_13759,N_13622,N_13618);
nand U13760 (N_13760,N_13537,N_13543);
or U13761 (N_13761,N_13592,N_13606);
or U13762 (N_13762,N_13534,N_13616);
nand U13763 (N_13763,N_13555,N_13537);
and U13764 (N_13764,N_13508,N_13581);
nor U13765 (N_13765,N_13517,N_13572);
and U13766 (N_13766,N_13587,N_13603);
nor U13767 (N_13767,N_13605,N_13572);
nand U13768 (N_13768,N_13568,N_13615);
nor U13769 (N_13769,N_13605,N_13511);
xor U13770 (N_13770,N_13509,N_13648);
or U13771 (N_13771,N_13545,N_13580);
or U13772 (N_13772,N_13620,N_13515);
nand U13773 (N_13773,N_13523,N_13553);
and U13774 (N_13774,N_13543,N_13519);
nand U13775 (N_13775,N_13606,N_13530);
or U13776 (N_13776,N_13592,N_13593);
nand U13777 (N_13777,N_13573,N_13516);
nor U13778 (N_13778,N_13569,N_13622);
and U13779 (N_13779,N_13547,N_13549);
nor U13780 (N_13780,N_13619,N_13644);
nand U13781 (N_13781,N_13507,N_13563);
nand U13782 (N_13782,N_13538,N_13591);
nor U13783 (N_13783,N_13546,N_13545);
xnor U13784 (N_13784,N_13522,N_13516);
nand U13785 (N_13785,N_13600,N_13632);
and U13786 (N_13786,N_13614,N_13617);
nand U13787 (N_13787,N_13571,N_13514);
and U13788 (N_13788,N_13508,N_13509);
and U13789 (N_13789,N_13585,N_13517);
nand U13790 (N_13790,N_13634,N_13633);
nor U13791 (N_13791,N_13618,N_13642);
and U13792 (N_13792,N_13570,N_13641);
and U13793 (N_13793,N_13558,N_13525);
and U13794 (N_13794,N_13554,N_13608);
and U13795 (N_13795,N_13514,N_13570);
nor U13796 (N_13796,N_13644,N_13618);
or U13797 (N_13797,N_13630,N_13538);
or U13798 (N_13798,N_13611,N_13531);
nand U13799 (N_13799,N_13635,N_13596);
or U13800 (N_13800,N_13690,N_13651);
xnor U13801 (N_13801,N_13662,N_13657);
xor U13802 (N_13802,N_13789,N_13756);
or U13803 (N_13803,N_13736,N_13747);
nor U13804 (N_13804,N_13696,N_13770);
nor U13805 (N_13805,N_13672,N_13675);
nand U13806 (N_13806,N_13735,N_13779);
and U13807 (N_13807,N_13658,N_13741);
and U13808 (N_13808,N_13763,N_13692);
or U13809 (N_13809,N_13667,N_13781);
and U13810 (N_13810,N_13653,N_13728);
or U13811 (N_13811,N_13794,N_13785);
nor U13812 (N_13812,N_13768,N_13689);
xor U13813 (N_13813,N_13740,N_13684);
or U13814 (N_13814,N_13720,N_13787);
xnor U13815 (N_13815,N_13784,N_13687);
and U13816 (N_13816,N_13704,N_13655);
or U13817 (N_13817,N_13703,N_13745);
and U13818 (N_13818,N_13721,N_13691);
or U13819 (N_13819,N_13668,N_13674);
nand U13820 (N_13820,N_13712,N_13737);
or U13821 (N_13821,N_13759,N_13798);
and U13822 (N_13822,N_13778,N_13783);
xnor U13823 (N_13823,N_13769,N_13782);
or U13824 (N_13824,N_13697,N_13700);
and U13825 (N_13825,N_13670,N_13760);
xnor U13826 (N_13826,N_13757,N_13765);
or U13827 (N_13827,N_13719,N_13652);
nor U13828 (N_13828,N_13699,N_13780);
nor U13829 (N_13829,N_13766,N_13773);
nand U13830 (N_13830,N_13748,N_13762);
or U13831 (N_13831,N_13799,N_13677);
or U13832 (N_13832,N_13775,N_13659);
or U13833 (N_13833,N_13707,N_13742);
and U13834 (N_13834,N_13732,N_13679);
or U13835 (N_13835,N_13733,N_13795);
xor U13836 (N_13836,N_13758,N_13722);
nor U13837 (N_13837,N_13686,N_13676);
or U13838 (N_13838,N_13680,N_13706);
nand U13839 (N_13839,N_13705,N_13788);
or U13840 (N_13840,N_13750,N_13723);
nand U13841 (N_13841,N_13663,N_13793);
or U13842 (N_13842,N_13739,N_13749);
or U13843 (N_13843,N_13682,N_13688);
or U13844 (N_13844,N_13725,N_13701);
or U13845 (N_13845,N_13738,N_13755);
nand U13846 (N_13846,N_13771,N_13729);
nand U13847 (N_13847,N_13665,N_13772);
xor U13848 (N_13848,N_13767,N_13792);
or U13849 (N_13849,N_13650,N_13761);
nand U13850 (N_13850,N_13713,N_13754);
or U13851 (N_13851,N_13695,N_13751);
and U13852 (N_13852,N_13726,N_13678);
xnor U13853 (N_13853,N_13654,N_13710);
or U13854 (N_13854,N_13685,N_13671);
xnor U13855 (N_13855,N_13790,N_13718);
or U13856 (N_13856,N_13731,N_13743);
and U13857 (N_13857,N_13774,N_13727);
nor U13858 (N_13858,N_13664,N_13752);
or U13859 (N_13859,N_13730,N_13698);
and U13860 (N_13860,N_13660,N_13708);
nand U13861 (N_13861,N_13702,N_13716);
nand U13862 (N_13862,N_13746,N_13796);
nor U13863 (N_13863,N_13693,N_13715);
and U13864 (N_13864,N_13734,N_13714);
nor U13865 (N_13865,N_13656,N_13724);
or U13866 (N_13866,N_13753,N_13764);
nor U13867 (N_13867,N_13694,N_13744);
nor U13868 (N_13868,N_13661,N_13797);
nor U13869 (N_13869,N_13681,N_13666);
or U13870 (N_13870,N_13791,N_13683);
and U13871 (N_13871,N_13669,N_13717);
xor U13872 (N_13872,N_13709,N_13711);
or U13873 (N_13873,N_13777,N_13786);
nand U13874 (N_13874,N_13673,N_13776);
and U13875 (N_13875,N_13740,N_13659);
xnor U13876 (N_13876,N_13795,N_13758);
or U13877 (N_13877,N_13753,N_13793);
nor U13878 (N_13878,N_13741,N_13770);
nand U13879 (N_13879,N_13773,N_13669);
or U13880 (N_13880,N_13691,N_13670);
and U13881 (N_13881,N_13769,N_13714);
nand U13882 (N_13882,N_13792,N_13701);
xnor U13883 (N_13883,N_13787,N_13766);
or U13884 (N_13884,N_13688,N_13659);
xor U13885 (N_13885,N_13777,N_13729);
and U13886 (N_13886,N_13783,N_13650);
or U13887 (N_13887,N_13793,N_13681);
xnor U13888 (N_13888,N_13768,N_13684);
or U13889 (N_13889,N_13775,N_13681);
and U13890 (N_13890,N_13797,N_13728);
xnor U13891 (N_13891,N_13668,N_13695);
xnor U13892 (N_13892,N_13703,N_13677);
nor U13893 (N_13893,N_13742,N_13774);
nand U13894 (N_13894,N_13679,N_13778);
nor U13895 (N_13895,N_13671,N_13704);
or U13896 (N_13896,N_13757,N_13685);
nor U13897 (N_13897,N_13717,N_13670);
nand U13898 (N_13898,N_13746,N_13759);
nand U13899 (N_13899,N_13753,N_13763);
and U13900 (N_13900,N_13741,N_13662);
and U13901 (N_13901,N_13741,N_13714);
nor U13902 (N_13902,N_13691,N_13720);
and U13903 (N_13903,N_13745,N_13717);
nand U13904 (N_13904,N_13664,N_13791);
xnor U13905 (N_13905,N_13744,N_13690);
xor U13906 (N_13906,N_13760,N_13779);
nor U13907 (N_13907,N_13739,N_13761);
nand U13908 (N_13908,N_13698,N_13775);
nand U13909 (N_13909,N_13736,N_13716);
or U13910 (N_13910,N_13660,N_13666);
or U13911 (N_13911,N_13774,N_13741);
nor U13912 (N_13912,N_13771,N_13747);
and U13913 (N_13913,N_13699,N_13797);
nor U13914 (N_13914,N_13777,N_13732);
or U13915 (N_13915,N_13783,N_13699);
and U13916 (N_13916,N_13758,N_13696);
and U13917 (N_13917,N_13734,N_13666);
or U13918 (N_13918,N_13660,N_13671);
nand U13919 (N_13919,N_13796,N_13794);
nand U13920 (N_13920,N_13706,N_13653);
or U13921 (N_13921,N_13762,N_13785);
and U13922 (N_13922,N_13751,N_13793);
and U13923 (N_13923,N_13731,N_13741);
nand U13924 (N_13924,N_13676,N_13712);
nand U13925 (N_13925,N_13788,N_13791);
xor U13926 (N_13926,N_13799,N_13657);
and U13927 (N_13927,N_13714,N_13735);
or U13928 (N_13928,N_13751,N_13670);
xnor U13929 (N_13929,N_13678,N_13684);
nor U13930 (N_13930,N_13743,N_13700);
and U13931 (N_13931,N_13711,N_13763);
or U13932 (N_13932,N_13780,N_13707);
and U13933 (N_13933,N_13797,N_13678);
and U13934 (N_13934,N_13797,N_13768);
nor U13935 (N_13935,N_13718,N_13710);
nand U13936 (N_13936,N_13661,N_13714);
xnor U13937 (N_13937,N_13725,N_13750);
nand U13938 (N_13938,N_13789,N_13778);
nand U13939 (N_13939,N_13782,N_13717);
or U13940 (N_13940,N_13705,N_13795);
and U13941 (N_13941,N_13685,N_13691);
nand U13942 (N_13942,N_13777,N_13721);
nor U13943 (N_13943,N_13768,N_13673);
or U13944 (N_13944,N_13766,N_13695);
nor U13945 (N_13945,N_13773,N_13745);
nand U13946 (N_13946,N_13773,N_13667);
nor U13947 (N_13947,N_13749,N_13793);
and U13948 (N_13948,N_13704,N_13697);
nor U13949 (N_13949,N_13731,N_13722);
nand U13950 (N_13950,N_13867,N_13825);
nor U13951 (N_13951,N_13841,N_13908);
and U13952 (N_13952,N_13856,N_13886);
and U13953 (N_13953,N_13895,N_13885);
nand U13954 (N_13954,N_13833,N_13899);
nor U13955 (N_13955,N_13923,N_13882);
and U13956 (N_13956,N_13861,N_13806);
xnor U13957 (N_13957,N_13918,N_13928);
nand U13958 (N_13958,N_13868,N_13824);
or U13959 (N_13959,N_13843,N_13801);
nand U13960 (N_13960,N_13881,N_13898);
nand U13961 (N_13961,N_13831,N_13900);
and U13962 (N_13962,N_13820,N_13857);
or U13963 (N_13963,N_13887,N_13871);
or U13964 (N_13964,N_13909,N_13817);
and U13965 (N_13965,N_13830,N_13925);
nor U13966 (N_13966,N_13838,N_13828);
and U13967 (N_13967,N_13926,N_13829);
and U13968 (N_13968,N_13863,N_13920);
or U13969 (N_13969,N_13805,N_13903);
or U13970 (N_13970,N_13823,N_13924);
nand U13971 (N_13971,N_13858,N_13800);
or U13972 (N_13972,N_13854,N_13864);
nor U13973 (N_13973,N_13891,N_13810);
nand U13974 (N_13974,N_13901,N_13803);
xnor U13975 (N_13975,N_13818,N_13815);
or U13976 (N_13976,N_13847,N_13807);
nand U13977 (N_13977,N_13877,N_13879);
xnor U13978 (N_13978,N_13938,N_13939);
nand U13979 (N_13979,N_13893,N_13822);
xor U13980 (N_13980,N_13894,N_13880);
nand U13981 (N_13981,N_13816,N_13905);
xnor U13982 (N_13982,N_13846,N_13859);
nor U13983 (N_13983,N_13804,N_13851);
nor U13984 (N_13984,N_13919,N_13947);
and U13985 (N_13985,N_13929,N_13840);
xnor U13986 (N_13986,N_13916,N_13819);
nor U13987 (N_13987,N_13875,N_13883);
nand U13988 (N_13988,N_13835,N_13933);
and U13989 (N_13989,N_13848,N_13874);
and U13990 (N_13990,N_13913,N_13915);
or U13991 (N_13991,N_13937,N_13809);
nand U13992 (N_13992,N_13945,N_13904);
nand U13993 (N_13993,N_13942,N_13906);
xor U13994 (N_13994,N_13892,N_13860);
nand U13995 (N_13995,N_13907,N_13808);
and U13996 (N_13996,N_13902,N_13935);
and U13997 (N_13997,N_13914,N_13888);
and U13998 (N_13998,N_13890,N_13897);
and U13999 (N_13999,N_13827,N_13845);
nor U14000 (N_14000,N_13910,N_13917);
or U14001 (N_14001,N_13872,N_13865);
nand U14002 (N_14002,N_13814,N_13844);
xor U14003 (N_14003,N_13853,N_13869);
nor U14004 (N_14004,N_13876,N_13855);
or U14005 (N_14005,N_13921,N_13832);
and U14006 (N_14006,N_13940,N_13946);
nand U14007 (N_14007,N_13813,N_13836);
nor U14008 (N_14008,N_13837,N_13927);
and U14009 (N_14009,N_13842,N_13839);
nand U14010 (N_14010,N_13802,N_13941);
nand U14011 (N_14011,N_13884,N_13812);
nand U14012 (N_14012,N_13930,N_13873);
and U14013 (N_14013,N_13852,N_13850);
and U14014 (N_14014,N_13943,N_13866);
xnor U14015 (N_14015,N_13870,N_13934);
and U14016 (N_14016,N_13811,N_13878);
nor U14017 (N_14017,N_13896,N_13931);
and U14018 (N_14018,N_13821,N_13889);
xor U14019 (N_14019,N_13944,N_13834);
nor U14020 (N_14020,N_13948,N_13826);
xor U14021 (N_14021,N_13912,N_13932);
nor U14022 (N_14022,N_13922,N_13849);
or U14023 (N_14023,N_13949,N_13862);
or U14024 (N_14024,N_13911,N_13936);
xor U14025 (N_14025,N_13829,N_13800);
or U14026 (N_14026,N_13900,N_13931);
nand U14027 (N_14027,N_13909,N_13811);
and U14028 (N_14028,N_13907,N_13842);
xnor U14029 (N_14029,N_13850,N_13807);
or U14030 (N_14030,N_13893,N_13889);
and U14031 (N_14031,N_13921,N_13811);
and U14032 (N_14032,N_13841,N_13894);
nor U14033 (N_14033,N_13878,N_13940);
nand U14034 (N_14034,N_13812,N_13921);
and U14035 (N_14035,N_13822,N_13821);
or U14036 (N_14036,N_13852,N_13929);
or U14037 (N_14037,N_13858,N_13920);
xnor U14038 (N_14038,N_13920,N_13900);
nand U14039 (N_14039,N_13864,N_13815);
nand U14040 (N_14040,N_13943,N_13829);
and U14041 (N_14041,N_13845,N_13841);
nor U14042 (N_14042,N_13839,N_13945);
and U14043 (N_14043,N_13897,N_13822);
and U14044 (N_14044,N_13804,N_13867);
or U14045 (N_14045,N_13940,N_13933);
or U14046 (N_14046,N_13909,N_13810);
and U14047 (N_14047,N_13829,N_13806);
nand U14048 (N_14048,N_13946,N_13921);
or U14049 (N_14049,N_13894,N_13832);
nand U14050 (N_14050,N_13878,N_13860);
and U14051 (N_14051,N_13904,N_13859);
or U14052 (N_14052,N_13815,N_13921);
and U14053 (N_14053,N_13828,N_13863);
xor U14054 (N_14054,N_13934,N_13825);
nor U14055 (N_14055,N_13875,N_13831);
nor U14056 (N_14056,N_13866,N_13915);
nand U14057 (N_14057,N_13859,N_13844);
xor U14058 (N_14058,N_13800,N_13918);
xor U14059 (N_14059,N_13911,N_13810);
xor U14060 (N_14060,N_13824,N_13947);
and U14061 (N_14061,N_13924,N_13821);
xnor U14062 (N_14062,N_13857,N_13834);
nand U14063 (N_14063,N_13848,N_13867);
xor U14064 (N_14064,N_13821,N_13878);
or U14065 (N_14065,N_13821,N_13909);
or U14066 (N_14066,N_13843,N_13819);
xnor U14067 (N_14067,N_13905,N_13825);
and U14068 (N_14068,N_13863,N_13850);
or U14069 (N_14069,N_13920,N_13816);
nor U14070 (N_14070,N_13901,N_13884);
and U14071 (N_14071,N_13894,N_13940);
nor U14072 (N_14072,N_13911,N_13913);
nand U14073 (N_14073,N_13822,N_13889);
or U14074 (N_14074,N_13816,N_13924);
nand U14075 (N_14075,N_13928,N_13897);
or U14076 (N_14076,N_13925,N_13945);
and U14077 (N_14077,N_13929,N_13916);
nor U14078 (N_14078,N_13875,N_13902);
nand U14079 (N_14079,N_13855,N_13837);
or U14080 (N_14080,N_13943,N_13934);
xor U14081 (N_14081,N_13894,N_13882);
xnor U14082 (N_14082,N_13942,N_13846);
nand U14083 (N_14083,N_13868,N_13853);
and U14084 (N_14084,N_13907,N_13811);
nand U14085 (N_14085,N_13921,N_13893);
or U14086 (N_14086,N_13857,N_13840);
xor U14087 (N_14087,N_13872,N_13904);
or U14088 (N_14088,N_13924,N_13869);
nor U14089 (N_14089,N_13908,N_13820);
nand U14090 (N_14090,N_13933,N_13864);
nand U14091 (N_14091,N_13826,N_13925);
nand U14092 (N_14092,N_13856,N_13899);
or U14093 (N_14093,N_13865,N_13818);
or U14094 (N_14094,N_13940,N_13802);
and U14095 (N_14095,N_13865,N_13884);
nor U14096 (N_14096,N_13892,N_13854);
nand U14097 (N_14097,N_13828,N_13878);
xor U14098 (N_14098,N_13925,N_13831);
xor U14099 (N_14099,N_13897,N_13923);
nand U14100 (N_14100,N_14058,N_13959);
nor U14101 (N_14101,N_13979,N_14016);
and U14102 (N_14102,N_14087,N_14015);
and U14103 (N_14103,N_14051,N_13978);
xnor U14104 (N_14104,N_14006,N_13976);
nor U14105 (N_14105,N_14069,N_14012);
and U14106 (N_14106,N_14072,N_14019);
or U14107 (N_14107,N_13965,N_13964);
xor U14108 (N_14108,N_14007,N_13961);
or U14109 (N_14109,N_14041,N_14044);
nor U14110 (N_14110,N_13974,N_14032);
and U14111 (N_14111,N_14045,N_13956);
nor U14112 (N_14112,N_13986,N_14024);
and U14113 (N_14113,N_13997,N_14085);
nand U14114 (N_14114,N_14017,N_14040);
xnor U14115 (N_14115,N_14054,N_14097);
nor U14116 (N_14116,N_13951,N_13981);
and U14117 (N_14117,N_13955,N_14008);
or U14118 (N_14118,N_13973,N_14098);
nor U14119 (N_14119,N_14060,N_13983);
xnor U14120 (N_14120,N_13998,N_14023);
and U14121 (N_14121,N_13975,N_14005);
and U14122 (N_14122,N_14037,N_13968);
xnor U14123 (N_14123,N_14003,N_14056);
nand U14124 (N_14124,N_14073,N_14013);
nand U14125 (N_14125,N_13994,N_14094);
and U14126 (N_14126,N_14062,N_14088);
nor U14127 (N_14127,N_14010,N_14084);
xnor U14128 (N_14128,N_14009,N_14028);
or U14129 (N_14129,N_13988,N_14053);
xnor U14130 (N_14130,N_14092,N_14035);
nor U14131 (N_14131,N_14048,N_13980);
xor U14132 (N_14132,N_14090,N_14011);
or U14133 (N_14133,N_14068,N_13977);
or U14134 (N_14134,N_13989,N_13952);
nor U14135 (N_14135,N_13963,N_13969);
nor U14136 (N_14136,N_14050,N_14020);
nand U14137 (N_14137,N_14077,N_14079);
xnor U14138 (N_14138,N_14029,N_14047);
nor U14139 (N_14139,N_13971,N_14057);
nand U14140 (N_14140,N_13992,N_13966);
or U14141 (N_14141,N_14089,N_14066);
or U14142 (N_14142,N_13996,N_14001);
xnor U14143 (N_14143,N_14018,N_14049);
xnor U14144 (N_14144,N_13950,N_14076);
xor U14145 (N_14145,N_14000,N_13995);
and U14146 (N_14146,N_13967,N_14052);
and U14147 (N_14147,N_14042,N_14080);
nor U14148 (N_14148,N_14033,N_14014);
xor U14149 (N_14149,N_14039,N_14055);
or U14150 (N_14150,N_14065,N_14074);
or U14151 (N_14151,N_14038,N_14063);
nand U14152 (N_14152,N_14059,N_13960);
and U14153 (N_14153,N_13993,N_13962);
or U14154 (N_14154,N_14021,N_14086);
nand U14155 (N_14155,N_14061,N_13984);
nand U14156 (N_14156,N_13985,N_14096);
nand U14157 (N_14157,N_13982,N_14022);
nor U14158 (N_14158,N_13957,N_13990);
and U14159 (N_14159,N_14034,N_13958);
nand U14160 (N_14160,N_14046,N_14075);
and U14161 (N_14161,N_14030,N_14036);
nor U14162 (N_14162,N_13970,N_14064);
nor U14163 (N_14163,N_14070,N_14078);
nand U14164 (N_14164,N_14027,N_14091);
nor U14165 (N_14165,N_14043,N_13954);
and U14166 (N_14166,N_14067,N_14004);
nand U14167 (N_14167,N_14025,N_14082);
nor U14168 (N_14168,N_14093,N_13991);
nand U14169 (N_14169,N_14081,N_13987);
and U14170 (N_14170,N_14095,N_13999);
nand U14171 (N_14171,N_14071,N_14002);
or U14172 (N_14172,N_14099,N_14083);
nand U14173 (N_14173,N_14026,N_14031);
nand U14174 (N_14174,N_13953,N_13972);
or U14175 (N_14175,N_14059,N_14037);
and U14176 (N_14176,N_13999,N_14039);
and U14177 (N_14177,N_14013,N_14074);
and U14178 (N_14178,N_13979,N_14076);
xnor U14179 (N_14179,N_13986,N_14042);
nand U14180 (N_14180,N_14054,N_14029);
nand U14181 (N_14181,N_14011,N_13977);
and U14182 (N_14182,N_13998,N_14060);
xor U14183 (N_14183,N_14088,N_14000);
nor U14184 (N_14184,N_13985,N_14024);
xor U14185 (N_14185,N_14055,N_13960);
xor U14186 (N_14186,N_14043,N_14091);
and U14187 (N_14187,N_14061,N_14058);
and U14188 (N_14188,N_14045,N_13960);
nand U14189 (N_14189,N_14015,N_14079);
and U14190 (N_14190,N_14018,N_13953);
and U14191 (N_14191,N_13998,N_14022);
xnor U14192 (N_14192,N_13986,N_14018);
nand U14193 (N_14193,N_13993,N_13976);
and U14194 (N_14194,N_13998,N_13984);
nand U14195 (N_14195,N_14084,N_14040);
xor U14196 (N_14196,N_13976,N_14002);
xor U14197 (N_14197,N_14012,N_13962);
or U14198 (N_14198,N_13955,N_13994);
nand U14199 (N_14199,N_14087,N_13966);
and U14200 (N_14200,N_14052,N_14040);
and U14201 (N_14201,N_14024,N_14082);
xor U14202 (N_14202,N_14090,N_14015);
nand U14203 (N_14203,N_14082,N_14092);
xor U14204 (N_14204,N_14000,N_14030);
or U14205 (N_14205,N_13976,N_14083);
nor U14206 (N_14206,N_13996,N_14039);
nand U14207 (N_14207,N_14069,N_14018);
nand U14208 (N_14208,N_14072,N_14045);
nor U14209 (N_14209,N_14061,N_13970);
xnor U14210 (N_14210,N_13977,N_14084);
nand U14211 (N_14211,N_13987,N_13950);
and U14212 (N_14212,N_14014,N_13969);
xnor U14213 (N_14213,N_14023,N_13997);
and U14214 (N_14214,N_13983,N_14085);
nand U14215 (N_14215,N_14045,N_13994);
xnor U14216 (N_14216,N_13956,N_13990);
and U14217 (N_14217,N_14029,N_14031);
and U14218 (N_14218,N_14069,N_13953);
xnor U14219 (N_14219,N_14000,N_14061);
nor U14220 (N_14220,N_13996,N_14090);
xnor U14221 (N_14221,N_13965,N_14001);
nor U14222 (N_14222,N_14098,N_14017);
and U14223 (N_14223,N_13993,N_14082);
nor U14224 (N_14224,N_14091,N_14066);
nor U14225 (N_14225,N_14005,N_14070);
xor U14226 (N_14226,N_13978,N_13962);
nor U14227 (N_14227,N_14083,N_14050);
nand U14228 (N_14228,N_14018,N_14086);
or U14229 (N_14229,N_14076,N_13969);
and U14230 (N_14230,N_14002,N_13977);
xor U14231 (N_14231,N_13986,N_13976);
and U14232 (N_14232,N_13980,N_13985);
and U14233 (N_14233,N_14032,N_14015);
or U14234 (N_14234,N_14047,N_14001);
nand U14235 (N_14235,N_14049,N_14047);
or U14236 (N_14236,N_14073,N_14014);
and U14237 (N_14237,N_13964,N_14041);
nor U14238 (N_14238,N_14025,N_14004);
and U14239 (N_14239,N_14048,N_14047);
xnor U14240 (N_14240,N_14070,N_14097);
and U14241 (N_14241,N_14046,N_13969);
and U14242 (N_14242,N_13995,N_13977);
xnor U14243 (N_14243,N_13953,N_14074);
nor U14244 (N_14244,N_14037,N_13963);
xnor U14245 (N_14245,N_14076,N_14038);
xnor U14246 (N_14246,N_13996,N_13963);
nor U14247 (N_14247,N_14019,N_14010);
nand U14248 (N_14248,N_14046,N_13977);
xnor U14249 (N_14249,N_14092,N_13966);
or U14250 (N_14250,N_14227,N_14127);
nor U14251 (N_14251,N_14186,N_14125);
or U14252 (N_14252,N_14135,N_14102);
xor U14253 (N_14253,N_14239,N_14152);
xnor U14254 (N_14254,N_14244,N_14177);
xor U14255 (N_14255,N_14183,N_14214);
and U14256 (N_14256,N_14113,N_14243);
and U14257 (N_14257,N_14213,N_14195);
and U14258 (N_14258,N_14208,N_14164);
nand U14259 (N_14259,N_14248,N_14151);
xor U14260 (N_14260,N_14169,N_14228);
nor U14261 (N_14261,N_14111,N_14144);
xnor U14262 (N_14262,N_14124,N_14118);
and U14263 (N_14263,N_14187,N_14150);
nand U14264 (N_14264,N_14104,N_14171);
nand U14265 (N_14265,N_14112,N_14200);
nand U14266 (N_14266,N_14160,N_14201);
or U14267 (N_14267,N_14184,N_14210);
xnor U14268 (N_14268,N_14233,N_14222);
xnor U14269 (N_14269,N_14162,N_14116);
nor U14270 (N_14270,N_14123,N_14237);
and U14271 (N_14271,N_14121,N_14140);
nor U14272 (N_14272,N_14193,N_14138);
nand U14273 (N_14273,N_14126,N_14232);
xnor U14274 (N_14274,N_14190,N_14246);
xor U14275 (N_14275,N_14207,N_14223);
nor U14276 (N_14276,N_14147,N_14212);
nand U14277 (N_14277,N_14109,N_14166);
or U14278 (N_14278,N_14130,N_14149);
and U14279 (N_14279,N_14173,N_14179);
or U14280 (N_14280,N_14159,N_14220);
nor U14281 (N_14281,N_14119,N_14181);
xnor U14282 (N_14282,N_14229,N_14202);
nand U14283 (N_14283,N_14129,N_14234);
nor U14284 (N_14284,N_14114,N_14178);
nor U14285 (N_14285,N_14247,N_14203);
or U14286 (N_14286,N_14146,N_14194);
nor U14287 (N_14287,N_14153,N_14180);
or U14288 (N_14288,N_14136,N_14215);
nor U14289 (N_14289,N_14192,N_14131);
nand U14290 (N_14290,N_14226,N_14141);
nand U14291 (N_14291,N_14156,N_14219);
xor U14292 (N_14292,N_14199,N_14134);
nor U14293 (N_14293,N_14108,N_14217);
and U14294 (N_14294,N_14174,N_14185);
or U14295 (N_14295,N_14122,N_14107);
and U14296 (N_14296,N_14106,N_14161);
or U14297 (N_14297,N_14196,N_14249);
or U14298 (N_14298,N_14206,N_14189);
xnor U14299 (N_14299,N_14168,N_14188);
nand U14300 (N_14300,N_14197,N_14216);
or U14301 (N_14301,N_14245,N_14165);
or U14302 (N_14302,N_14103,N_14142);
nor U14303 (N_14303,N_14221,N_14218);
and U14304 (N_14304,N_14198,N_14175);
and U14305 (N_14305,N_14241,N_14238);
xor U14306 (N_14306,N_14167,N_14176);
or U14307 (N_14307,N_14100,N_14182);
and U14308 (N_14308,N_14235,N_14231);
nor U14309 (N_14309,N_14191,N_14132);
or U14310 (N_14310,N_14133,N_14154);
and U14311 (N_14311,N_14211,N_14120);
and U14312 (N_14312,N_14148,N_14225);
xor U14313 (N_14313,N_14163,N_14117);
nand U14314 (N_14314,N_14145,N_14242);
and U14315 (N_14315,N_14230,N_14143);
nor U14316 (N_14316,N_14115,N_14110);
or U14317 (N_14317,N_14101,N_14205);
nor U14318 (N_14318,N_14157,N_14139);
nor U14319 (N_14319,N_14158,N_14209);
xnor U14320 (N_14320,N_14204,N_14236);
and U14321 (N_14321,N_14170,N_14128);
nor U14322 (N_14322,N_14105,N_14240);
nand U14323 (N_14323,N_14155,N_14224);
or U14324 (N_14324,N_14137,N_14172);
xor U14325 (N_14325,N_14165,N_14156);
nand U14326 (N_14326,N_14155,N_14191);
nor U14327 (N_14327,N_14158,N_14105);
xnor U14328 (N_14328,N_14221,N_14171);
nor U14329 (N_14329,N_14202,N_14215);
or U14330 (N_14330,N_14156,N_14213);
and U14331 (N_14331,N_14217,N_14146);
nand U14332 (N_14332,N_14116,N_14200);
and U14333 (N_14333,N_14213,N_14115);
nor U14334 (N_14334,N_14108,N_14138);
nor U14335 (N_14335,N_14121,N_14228);
nand U14336 (N_14336,N_14242,N_14191);
and U14337 (N_14337,N_14140,N_14245);
and U14338 (N_14338,N_14186,N_14166);
and U14339 (N_14339,N_14217,N_14201);
nor U14340 (N_14340,N_14134,N_14137);
nand U14341 (N_14341,N_14234,N_14232);
and U14342 (N_14342,N_14129,N_14205);
xor U14343 (N_14343,N_14197,N_14223);
and U14344 (N_14344,N_14126,N_14184);
xnor U14345 (N_14345,N_14184,N_14114);
or U14346 (N_14346,N_14216,N_14201);
xnor U14347 (N_14347,N_14108,N_14226);
nor U14348 (N_14348,N_14220,N_14202);
xnor U14349 (N_14349,N_14109,N_14244);
nor U14350 (N_14350,N_14171,N_14247);
xnor U14351 (N_14351,N_14171,N_14164);
or U14352 (N_14352,N_14122,N_14159);
nand U14353 (N_14353,N_14133,N_14145);
nand U14354 (N_14354,N_14119,N_14152);
xor U14355 (N_14355,N_14145,N_14223);
nand U14356 (N_14356,N_14219,N_14208);
nor U14357 (N_14357,N_14245,N_14232);
or U14358 (N_14358,N_14141,N_14160);
or U14359 (N_14359,N_14215,N_14245);
xnor U14360 (N_14360,N_14239,N_14117);
nand U14361 (N_14361,N_14200,N_14145);
xor U14362 (N_14362,N_14182,N_14214);
nor U14363 (N_14363,N_14232,N_14190);
or U14364 (N_14364,N_14236,N_14191);
or U14365 (N_14365,N_14198,N_14127);
nand U14366 (N_14366,N_14124,N_14112);
and U14367 (N_14367,N_14246,N_14132);
nor U14368 (N_14368,N_14204,N_14116);
nand U14369 (N_14369,N_14174,N_14223);
or U14370 (N_14370,N_14160,N_14176);
xnor U14371 (N_14371,N_14100,N_14151);
or U14372 (N_14372,N_14245,N_14243);
nand U14373 (N_14373,N_14246,N_14180);
or U14374 (N_14374,N_14165,N_14223);
or U14375 (N_14375,N_14123,N_14224);
nand U14376 (N_14376,N_14246,N_14247);
nor U14377 (N_14377,N_14159,N_14185);
nor U14378 (N_14378,N_14234,N_14199);
and U14379 (N_14379,N_14208,N_14239);
nor U14380 (N_14380,N_14104,N_14143);
and U14381 (N_14381,N_14184,N_14112);
xor U14382 (N_14382,N_14223,N_14220);
and U14383 (N_14383,N_14246,N_14232);
nand U14384 (N_14384,N_14195,N_14153);
nand U14385 (N_14385,N_14170,N_14195);
nand U14386 (N_14386,N_14128,N_14235);
nor U14387 (N_14387,N_14196,N_14139);
xor U14388 (N_14388,N_14219,N_14225);
or U14389 (N_14389,N_14230,N_14136);
nor U14390 (N_14390,N_14136,N_14205);
nand U14391 (N_14391,N_14242,N_14101);
nand U14392 (N_14392,N_14197,N_14119);
nand U14393 (N_14393,N_14207,N_14175);
or U14394 (N_14394,N_14105,N_14190);
or U14395 (N_14395,N_14203,N_14226);
nand U14396 (N_14396,N_14224,N_14172);
nor U14397 (N_14397,N_14106,N_14196);
nand U14398 (N_14398,N_14215,N_14168);
nor U14399 (N_14399,N_14186,N_14182);
nor U14400 (N_14400,N_14339,N_14361);
or U14401 (N_14401,N_14366,N_14399);
xnor U14402 (N_14402,N_14253,N_14360);
xor U14403 (N_14403,N_14315,N_14342);
xnor U14404 (N_14404,N_14334,N_14381);
xnor U14405 (N_14405,N_14295,N_14269);
or U14406 (N_14406,N_14362,N_14260);
xnor U14407 (N_14407,N_14394,N_14265);
or U14408 (N_14408,N_14278,N_14291);
nor U14409 (N_14409,N_14390,N_14392);
xor U14410 (N_14410,N_14396,N_14282);
nor U14411 (N_14411,N_14388,N_14325);
nand U14412 (N_14412,N_14302,N_14344);
xnor U14413 (N_14413,N_14254,N_14250);
and U14414 (N_14414,N_14335,N_14397);
xor U14415 (N_14415,N_14270,N_14353);
nor U14416 (N_14416,N_14287,N_14273);
xnor U14417 (N_14417,N_14276,N_14307);
and U14418 (N_14418,N_14283,N_14332);
or U14419 (N_14419,N_14303,N_14393);
nand U14420 (N_14420,N_14293,N_14330);
and U14421 (N_14421,N_14320,N_14380);
xor U14422 (N_14422,N_14395,N_14311);
or U14423 (N_14423,N_14300,N_14301);
and U14424 (N_14424,N_14314,N_14357);
nand U14425 (N_14425,N_14343,N_14376);
or U14426 (N_14426,N_14351,N_14251);
nand U14427 (N_14427,N_14354,N_14365);
or U14428 (N_14428,N_14288,N_14255);
nor U14429 (N_14429,N_14391,N_14304);
and U14430 (N_14430,N_14324,N_14305);
nand U14431 (N_14431,N_14386,N_14297);
or U14432 (N_14432,N_14369,N_14309);
and U14433 (N_14433,N_14389,N_14290);
nand U14434 (N_14434,N_14279,N_14346);
or U14435 (N_14435,N_14371,N_14358);
nand U14436 (N_14436,N_14271,N_14356);
xor U14437 (N_14437,N_14319,N_14292);
or U14438 (N_14438,N_14373,N_14316);
xnor U14439 (N_14439,N_14328,N_14398);
nand U14440 (N_14440,N_14299,N_14322);
and U14441 (N_14441,N_14331,N_14341);
nor U14442 (N_14442,N_14313,N_14284);
and U14443 (N_14443,N_14382,N_14310);
and U14444 (N_14444,N_14350,N_14379);
or U14445 (N_14445,N_14364,N_14275);
nor U14446 (N_14446,N_14252,N_14298);
nor U14447 (N_14447,N_14370,N_14267);
xnor U14448 (N_14448,N_14262,N_14387);
or U14449 (N_14449,N_14277,N_14352);
nor U14450 (N_14450,N_14385,N_14258);
or U14451 (N_14451,N_14321,N_14306);
nand U14452 (N_14452,N_14383,N_14337);
nor U14453 (N_14453,N_14349,N_14340);
or U14454 (N_14454,N_14317,N_14363);
and U14455 (N_14455,N_14266,N_14347);
nor U14456 (N_14456,N_14367,N_14336);
and U14457 (N_14457,N_14274,N_14355);
and U14458 (N_14458,N_14377,N_14338);
and U14459 (N_14459,N_14264,N_14281);
nor U14460 (N_14460,N_14261,N_14375);
or U14461 (N_14461,N_14268,N_14259);
nand U14462 (N_14462,N_14286,N_14294);
xor U14463 (N_14463,N_14308,N_14323);
or U14464 (N_14464,N_14257,N_14263);
nand U14465 (N_14465,N_14329,N_14368);
xor U14466 (N_14466,N_14374,N_14372);
and U14467 (N_14467,N_14280,N_14312);
nor U14468 (N_14468,N_14326,N_14285);
or U14469 (N_14469,N_14333,N_14318);
nand U14470 (N_14470,N_14289,N_14348);
xor U14471 (N_14471,N_14327,N_14345);
or U14472 (N_14472,N_14272,N_14384);
xor U14473 (N_14473,N_14296,N_14378);
nand U14474 (N_14474,N_14359,N_14256);
and U14475 (N_14475,N_14259,N_14381);
nor U14476 (N_14476,N_14267,N_14372);
or U14477 (N_14477,N_14359,N_14294);
nor U14478 (N_14478,N_14397,N_14307);
or U14479 (N_14479,N_14392,N_14269);
xor U14480 (N_14480,N_14328,N_14291);
and U14481 (N_14481,N_14336,N_14362);
nand U14482 (N_14482,N_14366,N_14378);
nand U14483 (N_14483,N_14329,N_14352);
nand U14484 (N_14484,N_14259,N_14374);
nor U14485 (N_14485,N_14299,N_14332);
nor U14486 (N_14486,N_14268,N_14340);
xnor U14487 (N_14487,N_14286,N_14380);
xnor U14488 (N_14488,N_14297,N_14343);
nor U14489 (N_14489,N_14342,N_14265);
nand U14490 (N_14490,N_14315,N_14301);
nand U14491 (N_14491,N_14365,N_14276);
or U14492 (N_14492,N_14275,N_14393);
nand U14493 (N_14493,N_14386,N_14261);
and U14494 (N_14494,N_14399,N_14347);
and U14495 (N_14495,N_14298,N_14377);
and U14496 (N_14496,N_14385,N_14250);
nand U14497 (N_14497,N_14344,N_14301);
or U14498 (N_14498,N_14333,N_14393);
nand U14499 (N_14499,N_14395,N_14290);
nand U14500 (N_14500,N_14262,N_14359);
and U14501 (N_14501,N_14286,N_14328);
xnor U14502 (N_14502,N_14282,N_14360);
xnor U14503 (N_14503,N_14389,N_14337);
or U14504 (N_14504,N_14352,N_14258);
nor U14505 (N_14505,N_14397,N_14264);
nor U14506 (N_14506,N_14280,N_14325);
nand U14507 (N_14507,N_14345,N_14362);
or U14508 (N_14508,N_14251,N_14396);
or U14509 (N_14509,N_14345,N_14357);
nand U14510 (N_14510,N_14361,N_14360);
and U14511 (N_14511,N_14347,N_14328);
xor U14512 (N_14512,N_14323,N_14261);
and U14513 (N_14513,N_14288,N_14274);
nor U14514 (N_14514,N_14351,N_14273);
nand U14515 (N_14515,N_14372,N_14268);
or U14516 (N_14516,N_14287,N_14257);
nor U14517 (N_14517,N_14273,N_14303);
and U14518 (N_14518,N_14292,N_14329);
nand U14519 (N_14519,N_14264,N_14344);
nor U14520 (N_14520,N_14383,N_14353);
nor U14521 (N_14521,N_14340,N_14273);
xnor U14522 (N_14522,N_14391,N_14363);
xnor U14523 (N_14523,N_14300,N_14381);
nor U14524 (N_14524,N_14398,N_14333);
nor U14525 (N_14525,N_14302,N_14307);
and U14526 (N_14526,N_14351,N_14291);
or U14527 (N_14527,N_14310,N_14365);
nand U14528 (N_14528,N_14330,N_14397);
nor U14529 (N_14529,N_14374,N_14324);
xnor U14530 (N_14530,N_14251,N_14360);
xor U14531 (N_14531,N_14264,N_14291);
xnor U14532 (N_14532,N_14252,N_14284);
or U14533 (N_14533,N_14319,N_14394);
xor U14534 (N_14534,N_14293,N_14301);
or U14535 (N_14535,N_14335,N_14344);
or U14536 (N_14536,N_14326,N_14397);
nand U14537 (N_14537,N_14389,N_14398);
nand U14538 (N_14538,N_14376,N_14334);
nand U14539 (N_14539,N_14286,N_14256);
nand U14540 (N_14540,N_14372,N_14350);
xor U14541 (N_14541,N_14282,N_14317);
or U14542 (N_14542,N_14399,N_14336);
xnor U14543 (N_14543,N_14274,N_14299);
and U14544 (N_14544,N_14252,N_14304);
xor U14545 (N_14545,N_14295,N_14399);
and U14546 (N_14546,N_14292,N_14310);
and U14547 (N_14547,N_14287,N_14309);
and U14548 (N_14548,N_14285,N_14308);
nor U14549 (N_14549,N_14304,N_14329);
nor U14550 (N_14550,N_14401,N_14430);
and U14551 (N_14551,N_14538,N_14527);
xnor U14552 (N_14552,N_14416,N_14543);
nor U14553 (N_14553,N_14474,N_14536);
nor U14554 (N_14554,N_14422,N_14466);
nor U14555 (N_14555,N_14460,N_14509);
and U14556 (N_14556,N_14435,N_14410);
nand U14557 (N_14557,N_14456,N_14468);
or U14558 (N_14558,N_14443,N_14486);
xor U14559 (N_14559,N_14471,N_14447);
xnor U14560 (N_14560,N_14437,N_14433);
or U14561 (N_14561,N_14530,N_14514);
nand U14562 (N_14562,N_14504,N_14525);
nand U14563 (N_14563,N_14485,N_14439);
and U14564 (N_14564,N_14415,N_14444);
and U14565 (N_14565,N_14408,N_14421);
or U14566 (N_14566,N_14516,N_14499);
nand U14567 (N_14567,N_14533,N_14450);
xnor U14568 (N_14568,N_14495,N_14477);
nor U14569 (N_14569,N_14406,N_14463);
xnor U14570 (N_14570,N_14492,N_14500);
nand U14571 (N_14571,N_14417,N_14512);
xor U14572 (N_14572,N_14541,N_14489);
nor U14573 (N_14573,N_14482,N_14521);
xor U14574 (N_14574,N_14501,N_14458);
and U14575 (N_14575,N_14442,N_14479);
and U14576 (N_14576,N_14470,N_14452);
nand U14577 (N_14577,N_14457,N_14453);
nor U14578 (N_14578,N_14413,N_14490);
nor U14579 (N_14579,N_14424,N_14547);
xnor U14580 (N_14580,N_14407,N_14469);
and U14581 (N_14581,N_14425,N_14531);
or U14582 (N_14582,N_14446,N_14455);
or U14583 (N_14583,N_14451,N_14502);
or U14584 (N_14584,N_14481,N_14403);
and U14585 (N_14585,N_14423,N_14449);
nand U14586 (N_14586,N_14432,N_14478);
xor U14587 (N_14587,N_14526,N_14519);
nor U14588 (N_14588,N_14454,N_14532);
nor U14589 (N_14589,N_14402,N_14517);
or U14590 (N_14590,N_14418,N_14497);
and U14591 (N_14591,N_14475,N_14441);
nand U14592 (N_14592,N_14462,N_14496);
or U14593 (N_14593,N_14465,N_14483);
or U14594 (N_14594,N_14549,N_14411);
nor U14595 (N_14595,N_14461,N_14428);
xnor U14596 (N_14596,N_14498,N_14473);
and U14597 (N_14597,N_14440,N_14438);
or U14598 (N_14598,N_14434,N_14520);
nor U14599 (N_14599,N_14476,N_14472);
or U14600 (N_14600,N_14518,N_14545);
and U14601 (N_14601,N_14534,N_14414);
and U14602 (N_14602,N_14431,N_14539);
xor U14603 (N_14603,N_14537,N_14420);
nor U14604 (N_14604,N_14467,N_14510);
xnor U14605 (N_14605,N_14436,N_14445);
xor U14606 (N_14606,N_14412,N_14409);
nor U14607 (N_14607,N_14515,N_14426);
and U14608 (N_14608,N_14535,N_14427);
nor U14609 (N_14609,N_14507,N_14491);
and U14610 (N_14610,N_14487,N_14506);
or U14611 (N_14611,N_14404,N_14529);
xnor U14612 (N_14612,N_14523,N_14528);
and U14613 (N_14613,N_14508,N_14480);
and U14614 (N_14614,N_14548,N_14546);
nor U14615 (N_14615,N_14542,N_14544);
or U14616 (N_14616,N_14505,N_14494);
nand U14617 (N_14617,N_14522,N_14405);
nor U14618 (N_14618,N_14459,N_14513);
nand U14619 (N_14619,N_14448,N_14400);
nor U14620 (N_14620,N_14464,N_14493);
nor U14621 (N_14621,N_14524,N_14484);
nor U14622 (N_14622,N_14419,N_14540);
nor U14623 (N_14623,N_14429,N_14511);
nor U14624 (N_14624,N_14503,N_14488);
nor U14625 (N_14625,N_14515,N_14510);
nand U14626 (N_14626,N_14438,N_14476);
or U14627 (N_14627,N_14504,N_14515);
or U14628 (N_14628,N_14506,N_14498);
xor U14629 (N_14629,N_14532,N_14512);
nand U14630 (N_14630,N_14448,N_14529);
nor U14631 (N_14631,N_14541,N_14539);
or U14632 (N_14632,N_14460,N_14536);
nand U14633 (N_14633,N_14482,N_14469);
and U14634 (N_14634,N_14506,N_14465);
and U14635 (N_14635,N_14425,N_14546);
and U14636 (N_14636,N_14488,N_14456);
or U14637 (N_14637,N_14402,N_14467);
and U14638 (N_14638,N_14405,N_14444);
or U14639 (N_14639,N_14533,N_14522);
nor U14640 (N_14640,N_14526,N_14416);
and U14641 (N_14641,N_14403,N_14502);
nor U14642 (N_14642,N_14490,N_14535);
and U14643 (N_14643,N_14422,N_14471);
nand U14644 (N_14644,N_14407,N_14432);
and U14645 (N_14645,N_14449,N_14460);
and U14646 (N_14646,N_14491,N_14534);
and U14647 (N_14647,N_14429,N_14435);
and U14648 (N_14648,N_14477,N_14544);
or U14649 (N_14649,N_14442,N_14416);
nand U14650 (N_14650,N_14471,N_14434);
and U14651 (N_14651,N_14414,N_14533);
and U14652 (N_14652,N_14521,N_14457);
and U14653 (N_14653,N_14451,N_14469);
nand U14654 (N_14654,N_14403,N_14463);
and U14655 (N_14655,N_14534,N_14522);
or U14656 (N_14656,N_14487,N_14500);
nor U14657 (N_14657,N_14427,N_14448);
xor U14658 (N_14658,N_14428,N_14412);
xnor U14659 (N_14659,N_14474,N_14493);
or U14660 (N_14660,N_14528,N_14466);
xnor U14661 (N_14661,N_14420,N_14444);
or U14662 (N_14662,N_14549,N_14437);
xor U14663 (N_14663,N_14460,N_14518);
xnor U14664 (N_14664,N_14507,N_14522);
xor U14665 (N_14665,N_14437,N_14519);
nand U14666 (N_14666,N_14510,N_14516);
and U14667 (N_14667,N_14473,N_14525);
xnor U14668 (N_14668,N_14486,N_14484);
nand U14669 (N_14669,N_14491,N_14453);
and U14670 (N_14670,N_14443,N_14405);
nor U14671 (N_14671,N_14531,N_14451);
nand U14672 (N_14672,N_14476,N_14516);
nand U14673 (N_14673,N_14421,N_14414);
nand U14674 (N_14674,N_14530,N_14500);
or U14675 (N_14675,N_14418,N_14511);
or U14676 (N_14676,N_14549,N_14430);
xor U14677 (N_14677,N_14488,N_14467);
and U14678 (N_14678,N_14439,N_14505);
xor U14679 (N_14679,N_14537,N_14465);
and U14680 (N_14680,N_14488,N_14549);
xnor U14681 (N_14681,N_14504,N_14473);
or U14682 (N_14682,N_14464,N_14524);
nand U14683 (N_14683,N_14543,N_14430);
xor U14684 (N_14684,N_14546,N_14501);
or U14685 (N_14685,N_14514,N_14498);
and U14686 (N_14686,N_14407,N_14479);
xor U14687 (N_14687,N_14521,N_14450);
nand U14688 (N_14688,N_14465,N_14445);
or U14689 (N_14689,N_14419,N_14417);
nor U14690 (N_14690,N_14448,N_14443);
nor U14691 (N_14691,N_14480,N_14427);
or U14692 (N_14692,N_14422,N_14487);
xor U14693 (N_14693,N_14456,N_14430);
or U14694 (N_14694,N_14443,N_14512);
xnor U14695 (N_14695,N_14501,N_14494);
nand U14696 (N_14696,N_14450,N_14512);
nand U14697 (N_14697,N_14535,N_14538);
or U14698 (N_14698,N_14410,N_14400);
nand U14699 (N_14699,N_14534,N_14456);
and U14700 (N_14700,N_14594,N_14681);
or U14701 (N_14701,N_14620,N_14633);
nor U14702 (N_14702,N_14656,N_14698);
nand U14703 (N_14703,N_14602,N_14603);
nor U14704 (N_14704,N_14664,N_14563);
xor U14705 (N_14705,N_14635,N_14608);
and U14706 (N_14706,N_14622,N_14584);
and U14707 (N_14707,N_14640,N_14554);
and U14708 (N_14708,N_14616,N_14659);
and U14709 (N_14709,N_14565,N_14689);
and U14710 (N_14710,N_14680,N_14574);
and U14711 (N_14711,N_14596,N_14694);
nor U14712 (N_14712,N_14618,N_14683);
and U14713 (N_14713,N_14636,N_14674);
or U14714 (N_14714,N_14637,N_14578);
nand U14715 (N_14715,N_14638,N_14685);
xnor U14716 (N_14716,N_14573,N_14609);
xnor U14717 (N_14717,N_14621,N_14677);
and U14718 (N_14718,N_14592,N_14655);
nand U14719 (N_14719,N_14629,N_14590);
and U14720 (N_14720,N_14614,N_14652);
xor U14721 (N_14721,N_14582,N_14593);
or U14722 (N_14722,N_14668,N_14551);
nor U14723 (N_14723,N_14556,N_14583);
xor U14724 (N_14724,N_14690,N_14628);
and U14725 (N_14725,N_14661,N_14581);
xor U14726 (N_14726,N_14691,N_14610);
xor U14727 (N_14727,N_14571,N_14606);
nand U14728 (N_14728,N_14634,N_14639);
xnor U14729 (N_14729,N_14564,N_14693);
or U14730 (N_14730,N_14644,N_14686);
nor U14731 (N_14731,N_14576,N_14619);
nor U14732 (N_14732,N_14632,N_14678);
nor U14733 (N_14733,N_14552,N_14630);
nand U14734 (N_14734,N_14588,N_14612);
nor U14735 (N_14735,N_14660,N_14676);
nor U14736 (N_14736,N_14558,N_14649);
or U14737 (N_14737,N_14617,N_14658);
nand U14738 (N_14738,N_14607,N_14647);
and U14739 (N_14739,N_14692,N_14697);
and U14740 (N_14740,N_14587,N_14580);
xor U14741 (N_14741,N_14695,N_14654);
or U14742 (N_14742,N_14631,N_14666);
and U14743 (N_14743,N_14560,N_14568);
nor U14744 (N_14744,N_14646,N_14579);
nor U14745 (N_14745,N_14553,N_14600);
nor U14746 (N_14746,N_14669,N_14645);
nor U14747 (N_14747,N_14572,N_14662);
nand U14748 (N_14748,N_14696,N_14642);
and U14749 (N_14749,N_14665,N_14570);
or U14750 (N_14750,N_14648,N_14557);
nand U14751 (N_14751,N_14559,N_14699);
and U14752 (N_14752,N_14653,N_14561);
or U14753 (N_14753,N_14641,N_14627);
nand U14754 (N_14754,N_14604,N_14643);
or U14755 (N_14755,N_14670,N_14605);
and U14756 (N_14756,N_14589,N_14597);
nor U14757 (N_14757,N_14625,N_14675);
nand U14758 (N_14758,N_14575,N_14550);
nand U14759 (N_14759,N_14577,N_14623);
nor U14760 (N_14760,N_14586,N_14657);
nor U14761 (N_14761,N_14650,N_14555);
nand U14762 (N_14762,N_14671,N_14601);
or U14763 (N_14763,N_14679,N_14599);
nor U14764 (N_14764,N_14673,N_14569);
and U14765 (N_14765,N_14688,N_14682);
nor U14766 (N_14766,N_14567,N_14626);
nand U14767 (N_14767,N_14598,N_14613);
nand U14768 (N_14768,N_14667,N_14595);
nor U14769 (N_14769,N_14591,N_14687);
nand U14770 (N_14770,N_14684,N_14615);
xnor U14771 (N_14771,N_14624,N_14611);
nand U14772 (N_14772,N_14651,N_14562);
xor U14773 (N_14773,N_14672,N_14663);
or U14774 (N_14774,N_14566,N_14585);
or U14775 (N_14775,N_14606,N_14673);
nor U14776 (N_14776,N_14635,N_14662);
or U14777 (N_14777,N_14649,N_14600);
nor U14778 (N_14778,N_14615,N_14643);
nand U14779 (N_14779,N_14669,N_14671);
nand U14780 (N_14780,N_14624,N_14618);
or U14781 (N_14781,N_14687,N_14618);
or U14782 (N_14782,N_14619,N_14660);
nor U14783 (N_14783,N_14575,N_14584);
nand U14784 (N_14784,N_14661,N_14563);
xnor U14785 (N_14785,N_14595,N_14552);
or U14786 (N_14786,N_14604,N_14636);
or U14787 (N_14787,N_14659,N_14665);
xor U14788 (N_14788,N_14599,N_14595);
xnor U14789 (N_14789,N_14593,N_14625);
or U14790 (N_14790,N_14696,N_14693);
or U14791 (N_14791,N_14672,N_14569);
nand U14792 (N_14792,N_14655,N_14699);
and U14793 (N_14793,N_14615,N_14667);
and U14794 (N_14794,N_14675,N_14588);
nor U14795 (N_14795,N_14600,N_14669);
nor U14796 (N_14796,N_14673,N_14566);
and U14797 (N_14797,N_14553,N_14655);
and U14798 (N_14798,N_14552,N_14698);
or U14799 (N_14799,N_14651,N_14576);
and U14800 (N_14800,N_14687,N_14609);
nor U14801 (N_14801,N_14554,N_14558);
or U14802 (N_14802,N_14621,N_14577);
nor U14803 (N_14803,N_14568,N_14691);
xnor U14804 (N_14804,N_14570,N_14628);
or U14805 (N_14805,N_14678,N_14593);
and U14806 (N_14806,N_14679,N_14568);
nor U14807 (N_14807,N_14680,N_14629);
xnor U14808 (N_14808,N_14607,N_14634);
xnor U14809 (N_14809,N_14618,N_14638);
and U14810 (N_14810,N_14646,N_14575);
nor U14811 (N_14811,N_14592,N_14591);
nand U14812 (N_14812,N_14602,N_14568);
and U14813 (N_14813,N_14624,N_14567);
xor U14814 (N_14814,N_14673,N_14614);
xnor U14815 (N_14815,N_14659,N_14585);
or U14816 (N_14816,N_14600,N_14640);
xnor U14817 (N_14817,N_14639,N_14561);
nand U14818 (N_14818,N_14695,N_14635);
nand U14819 (N_14819,N_14678,N_14667);
nand U14820 (N_14820,N_14633,N_14597);
nor U14821 (N_14821,N_14660,N_14558);
nand U14822 (N_14822,N_14650,N_14634);
or U14823 (N_14823,N_14582,N_14561);
and U14824 (N_14824,N_14655,N_14669);
nor U14825 (N_14825,N_14696,N_14667);
nor U14826 (N_14826,N_14574,N_14570);
nor U14827 (N_14827,N_14651,N_14597);
nor U14828 (N_14828,N_14699,N_14597);
or U14829 (N_14829,N_14669,N_14594);
xnor U14830 (N_14830,N_14608,N_14598);
nor U14831 (N_14831,N_14555,N_14693);
and U14832 (N_14832,N_14600,N_14555);
or U14833 (N_14833,N_14603,N_14574);
xnor U14834 (N_14834,N_14595,N_14551);
nand U14835 (N_14835,N_14644,N_14668);
xor U14836 (N_14836,N_14610,N_14696);
or U14837 (N_14837,N_14652,N_14661);
nand U14838 (N_14838,N_14551,N_14557);
nand U14839 (N_14839,N_14625,N_14630);
and U14840 (N_14840,N_14630,N_14577);
nand U14841 (N_14841,N_14603,N_14667);
nor U14842 (N_14842,N_14589,N_14666);
or U14843 (N_14843,N_14690,N_14613);
nand U14844 (N_14844,N_14673,N_14556);
or U14845 (N_14845,N_14698,N_14655);
xor U14846 (N_14846,N_14589,N_14613);
xnor U14847 (N_14847,N_14644,N_14591);
or U14848 (N_14848,N_14610,N_14663);
nand U14849 (N_14849,N_14568,N_14636);
xor U14850 (N_14850,N_14789,N_14767);
nor U14851 (N_14851,N_14746,N_14747);
nor U14852 (N_14852,N_14814,N_14772);
and U14853 (N_14853,N_14798,N_14731);
nor U14854 (N_14854,N_14782,N_14724);
nor U14855 (N_14855,N_14769,N_14784);
nor U14856 (N_14856,N_14761,N_14739);
xor U14857 (N_14857,N_14708,N_14804);
or U14858 (N_14858,N_14743,N_14725);
or U14859 (N_14859,N_14827,N_14790);
nor U14860 (N_14860,N_14733,N_14757);
and U14861 (N_14861,N_14750,N_14794);
and U14862 (N_14862,N_14833,N_14728);
or U14863 (N_14863,N_14763,N_14726);
nor U14864 (N_14864,N_14707,N_14751);
or U14865 (N_14865,N_14842,N_14783);
nor U14866 (N_14866,N_14738,N_14745);
and U14867 (N_14867,N_14844,N_14777);
or U14868 (N_14868,N_14836,N_14826);
nand U14869 (N_14869,N_14825,N_14758);
and U14870 (N_14870,N_14792,N_14702);
and U14871 (N_14871,N_14796,N_14727);
and U14872 (N_14872,N_14785,N_14841);
nor U14873 (N_14873,N_14832,N_14760);
xor U14874 (N_14874,N_14752,N_14712);
nand U14875 (N_14875,N_14834,N_14754);
and U14876 (N_14876,N_14820,N_14720);
nor U14877 (N_14877,N_14781,N_14764);
and U14878 (N_14878,N_14709,N_14723);
xnor U14879 (N_14879,N_14714,N_14806);
or U14880 (N_14880,N_14801,N_14721);
or U14881 (N_14881,N_14729,N_14831);
and U14882 (N_14882,N_14737,N_14701);
nand U14883 (N_14883,N_14773,N_14713);
or U14884 (N_14884,N_14776,N_14815);
or U14885 (N_14885,N_14821,N_14716);
nor U14886 (N_14886,N_14847,N_14744);
and U14887 (N_14887,N_14816,N_14732);
or U14888 (N_14888,N_14791,N_14765);
nor U14889 (N_14889,N_14749,N_14819);
xnor U14890 (N_14890,N_14722,N_14775);
and U14891 (N_14891,N_14812,N_14805);
and U14892 (N_14892,N_14771,N_14809);
xor U14893 (N_14893,N_14710,N_14755);
and U14894 (N_14894,N_14787,N_14706);
and U14895 (N_14895,N_14803,N_14700);
nand U14896 (N_14896,N_14719,N_14788);
xnor U14897 (N_14897,N_14797,N_14849);
nor U14898 (N_14898,N_14811,N_14807);
nor U14899 (N_14899,N_14734,N_14759);
and U14900 (N_14900,N_14843,N_14824);
nor U14901 (N_14901,N_14813,N_14810);
nor U14902 (N_14902,N_14780,N_14778);
nand U14903 (N_14903,N_14770,N_14735);
xor U14904 (N_14904,N_14740,N_14848);
nor U14905 (N_14905,N_14829,N_14817);
and U14906 (N_14906,N_14846,N_14799);
or U14907 (N_14907,N_14835,N_14774);
xnor U14908 (N_14908,N_14838,N_14818);
xnor U14909 (N_14909,N_14800,N_14718);
xor U14910 (N_14910,N_14736,N_14705);
or U14911 (N_14911,N_14779,N_14837);
nand U14912 (N_14912,N_14715,N_14753);
and U14913 (N_14913,N_14822,N_14845);
nand U14914 (N_14914,N_14748,N_14742);
and U14915 (N_14915,N_14768,N_14703);
and U14916 (N_14916,N_14823,N_14839);
xnor U14917 (N_14917,N_14762,N_14717);
and U14918 (N_14918,N_14711,N_14756);
and U14919 (N_14919,N_14704,N_14766);
and U14920 (N_14920,N_14828,N_14840);
nor U14921 (N_14921,N_14808,N_14795);
nand U14922 (N_14922,N_14741,N_14830);
and U14923 (N_14923,N_14730,N_14786);
xnor U14924 (N_14924,N_14802,N_14793);
nand U14925 (N_14925,N_14839,N_14810);
nand U14926 (N_14926,N_14826,N_14782);
nor U14927 (N_14927,N_14789,N_14849);
and U14928 (N_14928,N_14842,N_14708);
xor U14929 (N_14929,N_14764,N_14704);
xnor U14930 (N_14930,N_14792,N_14737);
xor U14931 (N_14931,N_14821,N_14705);
and U14932 (N_14932,N_14825,N_14761);
xnor U14933 (N_14933,N_14820,N_14723);
nor U14934 (N_14934,N_14774,N_14831);
nand U14935 (N_14935,N_14791,N_14842);
or U14936 (N_14936,N_14766,N_14779);
xor U14937 (N_14937,N_14732,N_14758);
nand U14938 (N_14938,N_14804,N_14833);
or U14939 (N_14939,N_14740,N_14809);
nand U14940 (N_14940,N_14726,N_14820);
or U14941 (N_14941,N_14838,N_14781);
and U14942 (N_14942,N_14825,N_14752);
and U14943 (N_14943,N_14756,N_14765);
and U14944 (N_14944,N_14793,N_14817);
or U14945 (N_14945,N_14766,N_14714);
xnor U14946 (N_14946,N_14807,N_14834);
nor U14947 (N_14947,N_14749,N_14802);
and U14948 (N_14948,N_14727,N_14701);
nor U14949 (N_14949,N_14757,N_14721);
xnor U14950 (N_14950,N_14769,N_14849);
xnor U14951 (N_14951,N_14743,N_14800);
nor U14952 (N_14952,N_14782,N_14834);
and U14953 (N_14953,N_14715,N_14725);
and U14954 (N_14954,N_14756,N_14705);
or U14955 (N_14955,N_14774,N_14776);
or U14956 (N_14956,N_14845,N_14843);
nor U14957 (N_14957,N_14801,N_14760);
xnor U14958 (N_14958,N_14832,N_14743);
or U14959 (N_14959,N_14722,N_14740);
nand U14960 (N_14960,N_14818,N_14739);
nand U14961 (N_14961,N_14741,N_14727);
and U14962 (N_14962,N_14786,N_14804);
and U14963 (N_14963,N_14795,N_14720);
nor U14964 (N_14964,N_14794,N_14838);
or U14965 (N_14965,N_14763,N_14786);
or U14966 (N_14966,N_14739,N_14737);
nor U14967 (N_14967,N_14776,N_14771);
nand U14968 (N_14968,N_14735,N_14728);
or U14969 (N_14969,N_14712,N_14793);
nor U14970 (N_14970,N_14795,N_14750);
and U14971 (N_14971,N_14810,N_14803);
nor U14972 (N_14972,N_14810,N_14769);
or U14973 (N_14973,N_14814,N_14763);
nand U14974 (N_14974,N_14840,N_14775);
or U14975 (N_14975,N_14727,N_14762);
and U14976 (N_14976,N_14793,N_14726);
xor U14977 (N_14977,N_14792,N_14809);
nand U14978 (N_14978,N_14752,N_14838);
xor U14979 (N_14979,N_14791,N_14749);
nor U14980 (N_14980,N_14718,N_14829);
and U14981 (N_14981,N_14810,N_14791);
nand U14982 (N_14982,N_14792,N_14786);
or U14983 (N_14983,N_14803,N_14824);
nor U14984 (N_14984,N_14842,N_14817);
xnor U14985 (N_14985,N_14773,N_14848);
nand U14986 (N_14986,N_14720,N_14729);
nand U14987 (N_14987,N_14820,N_14781);
or U14988 (N_14988,N_14840,N_14729);
nor U14989 (N_14989,N_14767,N_14722);
nor U14990 (N_14990,N_14718,N_14788);
or U14991 (N_14991,N_14735,N_14749);
and U14992 (N_14992,N_14755,N_14736);
and U14993 (N_14993,N_14767,N_14727);
xnor U14994 (N_14994,N_14749,N_14705);
xnor U14995 (N_14995,N_14727,N_14735);
nand U14996 (N_14996,N_14761,N_14748);
and U14997 (N_14997,N_14769,N_14830);
and U14998 (N_14998,N_14756,N_14703);
and U14999 (N_14999,N_14788,N_14843);
nand UO_0 (O_0,N_14859,N_14971);
nor UO_1 (O_1,N_14852,N_14895);
or UO_2 (O_2,N_14894,N_14939);
or UO_3 (O_3,N_14862,N_14860);
nand UO_4 (O_4,N_14997,N_14910);
and UO_5 (O_5,N_14865,N_14934);
or UO_6 (O_6,N_14941,N_14913);
and UO_7 (O_7,N_14986,N_14912);
or UO_8 (O_8,N_14962,N_14976);
or UO_9 (O_9,N_14903,N_14870);
or UO_10 (O_10,N_14888,N_14901);
or UO_11 (O_11,N_14940,N_14923);
and UO_12 (O_12,N_14980,N_14871);
xor UO_13 (O_13,N_14964,N_14953);
nor UO_14 (O_14,N_14983,N_14907);
nor UO_15 (O_15,N_14970,N_14911);
nand UO_16 (O_16,N_14909,N_14973);
and UO_17 (O_17,N_14946,N_14998);
or UO_18 (O_18,N_14853,N_14904);
xor UO_19 (O_19,N_14930,N_14929);
nor UO_20 (O_20,N_14950,N_14921);
nand UO_21 (O_21,N_14958,N_14883);
xnor UO_22 (O_22,N_14948,N_14977);
nor UO_23 (O_23,N_14960,N_14879);
and UO_24 (O_24,N_14979,N_14896);
or UO_25 (O_25,N_14906,N_14861);
xor UO_26 (O_26,N_14874,N_14996);
and UO_27 (O_27,N_14917,N_14931);
or UO_28 (O_28,N_14981,N_14876);
or UO_29 (O_29,N_14855,N_14937);
nor UO_30 (O_30,N_14886,N_14952);
or UO_31 (O_31,N_14945,N_14850);
nand UO_32 (O_32,N_14943,N_14916);
and UO_33 (O_33,N_14873,N_14932);
nand UO_34 (O_34,N_14972,N_14900);
nor UO_35 (O_35,N_14957,N_14951);
xnor UO_36 (O_36,N_14928,N_14897);
and UO_37 (O_37,N_14914,N_14864);
nor UO_38 (O_38,N_14905,N_14967);
and UO_39 (O_39,N_14956,N_14968);
nand UO_40 (O_40,N_14990,N_14959);
nand UO_41 (O_41,N_14891,N_14994);
nand UO_42 (O_42,N_14887,N_14995);
and UO_43 (O_43,N_14892,N_14863);
or UO_44 (O_44,N_14947,N_14987);
or UO_45 (O_45,N_14868,N_14908);
nor UO_46 (O_46,N_14854,N_14875);
nor UO_47 (O_47,N_14978,N_14869);
or UO_48 (O_48,N_14867,N_14857);
nor UO_49 (O_49,N_14924,N_14898);
or UO_50 (O_50,N_14984,N_14889);
and UO_51 (O_51,N_14974,N_14993);
nor UO_52 (O_52,N_14915,N_14936);
nand UO_53 (O_53,N_14988,N_14919);
xnor UO_54 (O_54,N_14938,N_14949);
or UO_55 (O_55,N_14872,N_14985);
nand UO_56 (O_56,N_14878,N_14942);
and UO_57 (O_57,N_14920,N_14961);
and UO_58 (O_58,N_14963,N_14989);
or UO_59 (O_59,N_14882,N_14935);
and UO_60 (O_60,N_14982,N_14933);
and UO_61 (O_61,N_14877,N_14927);
nand UO_62 (O_62,N_14992,N_14965);
nand UO_63 (O_63,N_14851,N_14893);
nand UO_64 (O_64,N_14944,N_14925);
nor UO_65 (O_65,N_14856,N_14866);
xnor UO_66 (O_66,N_14881,N_14955);
nand UO_67 (O_67,N_14918,N_14999);
nor UO_68 (O_68,N_14885,N_14954);
xnor UO_69 (O_69,N_14890,N_14884);
nor UO_70 (O_70,N_14966,N_14858);
nand UO_71 (O_71,N_14991,N_14969);
nand UO_72 (O_72,N_14880,N_14899);
nor UO_73 (O_73,N_14926,N_14922);
nand UO_74 (O_74,N_14902,N_14975);
or UO_75 (O_75,N_14878,N_14853);
nand UO_76 (O_76,N_14955,N_14921);
xnor UO_77 (O_77,N_14893,N_14876);
nand UO_78 (O_78,N_14880,N_14884);
xor UO_79 (O_79,N_14908,N_14902);
or UO_80 (O_80,N_14968,N_14966);
or UO_81 (O_81,N_14957,N_14950);
nand UO_82 (O_82,N_14903,N_14941);
and UO_83 (O_83,N_14965,N_14852);
xor UO_84 (O_84,N_14976,N_14998);
nand UO_85 (O_85,N_14921,N_14905);
or UO_86 (O_86,N_14871,N_14934);
and UO_87 (O_87,N_14857,N_14972);
and UO_88 (O_88,N_14876,N_14932);
and UO_89 (O_89,N_14991,N_14899);
nand UO_90 (O_90,N_14940,N_14941);
nand UO_91 (O_91,N_14923,N_14971);
nor UO_92 (O_92,N_14946,N_14854);
xor UO_93 (O_93,N_14976,N_14856);
nand UO_94 (O_94,N_14972,N_14874);
xor UO_95 (O_95,N_14959,N_14930);
and UO_96 (O_96,N_14910,N_14861);
or UO_97 (O_97,N_14889,N_14949);
and UO_98 (O_98,N_14853,N_14975);
xnor UO_99 (O_99,N_14933,N_14850);
or UO_100 (O_100,N_14941,N_14871);
nand UO_101 (O_101,N_14876,N_14997);
xor UO_102 (O_102,N_14917,N_14972);
nand UO_103 (O_103,N_14903,N_14959);
nor UO_104 (O_104,N_14939,N_14918);
or UO_105 (O_105,N_14986,N_14853);
and UO_106 (O_106,N_14912,N_14922);
xor UO_107 (O_107,N_14953,N_14859);
or UO_108 (O_108,N_14927,N_14856);
nor UO_109 (O_109,N_14913,N_14903);
xnor UO_110 (O_110,N_14923,N_14968);
and UO_111 (O_111,N_14947,N_14970);
nand UO_112 (O_112,N_14967,N_14973);
or UO_113 (O_113,N_14863,N_14929);
xnor UO_114 (O_114,N_14934,N_14997);
or UO_115 (O_115,N_14877,N_14987);
nor UO_116 (O_116,N_14859,N_14912);
nor UO_117 (O_117,N_14986,N_14974);
xor UO_118 (O_118,N_14943,N_14989);
nor UO_119 (O_119,N_14907,N_14954);
nor UO_120 (O_120,N_14867,N_14961);
and UO_121 (O_121,N_14879,N_14863);
nor UO_122 (O_122,N_14862,N_14928);
xnor UO_123 (O_123,N_14860,N_14868);
nor UO_124 (O_124,N_14905,N_14869);
xor UO_125 (O_125,N_14933,N_14901);
or UO_126 (O_126,N_14897,N_14951);
or UO_127 (O_127,N_14878,N_14867);
nor UO_128 (O_128,N_14851,N_14939);
or UO_129 (O_129,N_14900,N_14881);
xnor UO_130 (O_130,N_14882,N_14904);
xnor UO_131 (O_131,N_14967,N_14853);
or UO_132 (O_132,N_14894,N_14984);
nand UO_133 (O_133,N_14939,N_14873);
and UO_134 (O_134,N_14956,N_14979);
nand UO_135 (O_135,N_14961,N_14995);
or UO_136 (O_136,N_14932,N_14858);
xor UO_137 (O_137,N_14989,N_14896);
and UO_138 (O_138,N_14993,N_14977);
nor UO_139 (O_139,N_14870,N_14921);
xor UO_140 (O_140,N_14864,N_14869);
and UO_141 (O_141,N_14869,N_14886);
nor UO_142 (O_142,N_14965,N_14927);
xnor UO_143 (O_143,N_14914,N_14934);
nor UO_144 (O_144,N_14942,N_14867);
nor UO_145 (O_145,N_14927,N_14885);
or UO_146 (O_146,N_14852,N_14883);
nand UO_147 (O_147,N_14876,N_14957);
xnor UO_148 (O_148,N_14972,N_14867);
and UO_149 (O_149,N_14881,N_14858);
nand UO_150 (O_150,N_14884,N_14935);
nand UO_151 (O_151,N_14904,N_14984);
nor UO_152 (O_152,N_14895,N_14860);
nand UO_153 (O_153,N_14854,N_14868);
nor UO_154 (O_154,N_14865,N_14998);
xor UO_155 (O_155,N_14957,N_14858);
xnor UO_156 (O_156,N_14996,N_14975);
nor UO_157 (O_157,N_14903,N_14926);
xnor UO_158 (O_158,N_14863,N_14984);
nand UO_159 (O_159,N_14850,N_14855);
nor UO_160 (O_160,N_14899,N_14869);
and UO_161 (O_161,N_14898,N_14919);
and UO_162 (O_162,N_14982,N_14935);
nand UO_163 (O_163,N_14940,N_14970);
nor UO_164 (O_164,N_14973,N_14959);
and UO_165 (O_165,N_14885,N_14999);
or UO_166 (O_166,N_14978,N_14924);
xor UO_167 (O_167,N_14884,N_14934);
and UO_168 (O_168,N_14908,N_14992);
or UO_169 (O_169,N_14884,N_14873);
nand UO_170 (O_170,N_14948,N_14860);
and UO_171 (O_171,N_14860,N_14987);
nor UO_172 (O_172,N_14949,N_14854);
xor UO_173 (O_173,N_14947,N_14922);
nor UO_174 (O_174,N_14957,N_14952);
and UO_175 (O_175,N_14882,N_14850);
or UO_176 (O_176,N_14994,N_14946);
and UO_177 (O_177,N_14927,N_14875);
and UO_178 (O_178,N_14892,N_14893);
nand UO_179 (O_179,N_14867,N_14854);
or UO_180 (O_180,N_14993,N_14960);
xor UO_181 (O_181,N_14884,N_14938);
nor UO_182 (O_182,N_14903,N_14857);
and UO_183 (O_183,N_14902,N_14873);
nand UO_184 (O_184,N_14968,N_14917);
nor UO_185 (O_185,N_14885,N_14907);
nand UO_186 (O_186,N_14862,N_14917);
nor UO_187 (O_187,N_14927,N_14978);
and UO_188 (O_188,N_14933,N_14904);
xnor UO_189 (O_189,N_14950,N_14933);
xor UO_190 (O_190,N_14990,N_14976);
nand UO_191 (O_191,N_14952,N_14914);
xor UO_192 (O_192,N_14901,N_14988);
nor UO_193 (O_193,N_14851,N_14935);
and UO_194 (O_194,N_14901,N_14870);
or UO_195 (O_195,N_14975,N_14966);
nand UO_196 (O_196,N_14916,N_14893);
or UO_197 (O_197,N_14932,N_14957);
nand UO_198 (O_198,N_14892,N_14944);
nand UO_199 (O_199,N_14997,N_14900);
xor UO_200 (O_200,N_14928,N_14914);
or UO_201 (O_201,N_14957,N_14904);
nand UO_202 (O_202,N_14851,N_14889);
and UO_203 (O_203,N_14860,N_14890);
xor UO_204 (O_204,N_14963,N_14927);
or UO_205 (O_205,N_14958,N_14850);
nor UO_206 (O_206,N_14857,N_14963);
nand UO_207 (O_207,N_14956,N_14953);
or UO_208 (O_208,N_14892,N_14864);
or UO_209 (O_209,N_14984,N_14907);
xor UO_210 (O_210,N_14852,N_14904);
or UO_211 (O_211,N_14862,N_14881);
and UO_212 (O_212,N_14878,N_14950);
nor UO_213 (O_213,N_14990,N_14923);
nor UO_214 (O_214,N_14897,N_14860);
and UO_215 (O_215,N_14859,N_14878);
xor UO_216 (O_216,N_14931,N_14969);
xor UO_217 (O_217,N_14991,N_14973);
xnor UO_218 (O_218,N_14935,N_14916);
and UO_219 (O_219,N_14881,N_14935);
nand UO_220 (O_220,N_14893,N_14993);
nand UO_221 (O_221,N_14984,N_14921);
xnor UO_222 (O_222,N_14911,N_14942);
nor UO_223 (O_223,N_14919,N_14939);
nor UO_224 (O_224,N_14905,N_14911);
xnor UO_225 (O_225,N_14922,N_14890);
nand UO_226 (O_226,N_14887,N_14945);
xor UO_227 (O_227,N_14969,N_14890);
nor UO_228 (O_228,N_14945,N_14928);
nand UO_229 (O_229,N_14915,N_14928);
nor UO_230 (O_230,N_14852,N_14987);
and UO_231 (O_231,N_14983,N_14943);
and UO_232 (O_232,N_14920,N_14879);
and UO_233 (O_233,N_14985,N_14939);
nor UO_234 (O_234,N_14985,N_14891);
nor UO_235 (O_235,N_14939,N_14883);
nor UO_236 (O_236,N_14915,N_14866);
nor UO_237 (O_237,N_14900,N_14923);
nand UO_238 (O_238,N_14923,N_14975);
xor UO_239 (O_239,N_14856,N_14876);
xnor UO_240 (O_240,N_14965,N_14997);
and UO_241 (O_241,N_14931,N_14916);
or UO_242 (O_242,N_14933,N_14956);
and UO_243 (O_243,N_14968,N_14971);
nor UO_244 (O_244,N_14877,N_14906);
or UO_245 (O_245,N_14859,N_14945);
and UO_246 (O_246,N_14876,N_14909);
nand UO_247 (O_247,N_14925,N_14873);
or UO_248 (O_248,N_14936,N_14986);
xnor UO_249 (O_249,N_14981,N_14896);
xor UO_250 (O_250,N_14987,N_14970);
xnor UO_251 (O_251,N_14933,N_14945);
or UO_252 (O_252,N_14994,N_14894);
and UO_253 (O_253,N_14929,N_14994);
nand UO_254 (O_254,N_14920,N_14870);
and UO_255 (O_255,N_14998,N_14897);
or UO_256 (O_256,N_14912,N_14876);
xor UO_257 (O_257,N_14851,N_14937);
and UO_258 (O_258,N_14997,N_14893);
or UO_259 (O_259,N_14924,N_14891);
nand UO_260 (O_260,N_14973,N_14865);
nor UO_261 (O_261,N_14857,N_14886);
nand UO_262 (O_262,N_14981,N_14958);
or UO_263 (O_263,N_14996,N_14892);
xor UO_264 (O_264,N_14990,N_14962);
xnor UO_265 (O_265,N_14958,N_14966);
and UO_266 (O_266,N_14997,N_14950);
nor UO_267 (O_267,N_14968,N_14964);
or UO_268 (O_268,N_14920,N_14880);
nand UO_269 (O_269,N_14983,N_14997);
and UO_270 (O_270,N_14854,N_14984);
nor UO_271 (O_271,N_14877,N_14991);
or UO_272 (O_272,N_14956,N_14971);
nor UO_273 (O_273,N_14859,N_14935);
nand UO_274 (O_274,N_14954,N_14883);
and UO_275 (O_275,N_14922,N_14880);
and UO_276 (O_276,N_14937,N_14905);
nand UO_277 (O_277,N_14978,N_14971);
or UO_278 (O_278,N_14972,N_14889);
xor UO_279 (O_279,N_14933,N_14972);
nand UO_280 (O_280,N_14908,N_14987);
nor UO_281 (O_281,N_14902,N_14889);
xor UO_282 (O_282,N_14915,N_14850);
or UO_283 (O_283,N_14942,N_14892);
xnor UO_284 (O_284,N_14850,N_14954);
nor UO_285 (O_285,N_14918,N_14867);
or UO_286 (O_286,N_14971,N_14977);
nor UO_287 (O_287,N_14922,N_14862);
and UO_288 (O_288,N_14891,N_14988);
and UO_289 (O_289,N_14939,N_14933);
xor UO_290 (O_290,N_14994,N_14855);
or UO_291 (O_291,N_14928,N_14886);
nor UO_292 (O_292,N_14945,N_14878);
or UO_293 (O_293,N_14978,N_14887);
nor UO_294 (O_294,N_14934,N_14956);
nor UO_295 (O_295,N_14870,N_14862);
nor UO_296 (O_296,N_14901,N_14872);
or UO_297 (O_297,N_14927,N_14910);
xor UO_298 (O_298,N_14952,N_14889);
xor UO_299 (O_299,N_14913,N_14915);
nand UO_300 (O_300,N_14971,N_14989);
nor UO_301 (O_301,N_14984,N_14870);
or UO_302 (O_302,N_14898,N_14972);
xor UO_303 (O_303,N_14986,N_14962);
and UO_304 (O_304,N_14973,N_14972);
or UO_305 (O_305,N_14923,N_14942);
xor UO_306 (O_306,N_14979,N_14968);
nand UO_307 (O_307,N_14985,N_14968);
nor UO_308 (O_308,N_14979,N_14859);
nand UO_309 (O_309,N_14912,N_14999);
nand UO_310 (O_310,N_14916,N_14853);
nor UO_311 (O_311,N_14866,N_14985);
and UO_312 (O_312,N_14908,N_14998);
nor UO_313 (O_313,N_14873,N_14898);
nand UO_314 (O_314,N_14986,N_14881);
xor UO_315 (O_315,N_14877,N_14992);
or UO_316 (O_316,N_14927,N_14950);
nor UO_317 (O_317,N_14990,N_14983);
nor UO_318 (O_318,N_14903,N_14995);
xnor UO_319 (O_319,N_14890,N_14992);
nand UO_320 (O_320,N_14945,N_14899);
nand UO_321 (O_321,N_14881,N_14861);
nor UO_322 (O_322,N_14913,N_14923);
xor UO_323 (O_323,N_14922,N_14936);
and UO_324 (O_324,N_14894,N_14916);
or UO_325 (O_325,N_14936,N_14983);
and UO_326 (O_326,N_14857,N_14985);
nand UO_327 (O_327,N_14939,N_14871);
nor UO_328 (O_328,N_14889,N_14895);
and UO_329 (O_329,N_14996,N_14999);
nand UO_330 (O_330,N_14926,N_14998);
xor UO_331 (O_331,N_14974,N_14851);
or UO_332 (O_332,N_14969,N_14971);
nand UO_333 (O_333,N_14941,N_14912);
or UO_334 (O_334,N_14958,N_14913);
nand UO_335 (O_335,N_14924,N_14853);
or UO_336 (O_336,N_14891,N_14887);
and UO_337 (O_337,N_14895,N_14868);
or UO_338 (O_338,N_14905,N_14956);
nand UO_339 (O_339,N_14972,N_14877);
xnor UO_340 (O_340,N_14886,N_14974);
nand UO_341 (O_341,N_14906,N_14954);
and UO_342 (O_342,N_14868,N_14858);
nand UO_343 (O_343,N_14959,N_14894);
nand UO_344 (O_344,N_14976,N_14963);
nor UO_345 (O_345,N_14914,N_14879);
nand UO_346 (O_346,N_14898,N_14903);
nand UO_347 (O_347,N_14879,N_14874);
nor UO_348 (O_348,N_14979,N_14862);
xnor UO_349 (O_349,N_14951,N_14991);
and UO_350 (O_350,N_14858,N_14903);
xnor UO_351 (O_351,N_14896,N_14904);
nor UO_352 (O_352,N_14944,N_14949);
xor UO_353 (O_353,N_14881,N_14913);
or UO_354 (O_354,N_14922,N_14986);
xnor UO_355 (O_355,N_14853,N_14910);
nand UO_356 (O_356,N_14958,N_14975);
xnor UO_357 (O_357,N_14992,N_14955);
nor UO_358 (O_358,N_14960,N_14908);
nand UO_359 (O_359,N_14954,N_14923);
and UO_360 (O_360,N_14929,N_14958);
xor UO_361 (O_361,N_14910,N_14955);
nor UO_362 (O_362,N_14999,N_14954);
xor UO_363 (O_363,N_14872,N_14939);
or UO_364 (O_364,N_14934,N_14907);
xnor UO_365 (O_365,N_14881,N_14872);
nand UO_366 (O_366,N_14988,N_14981);
nor UO_367 (O_367,N_14995,N_14970);
nand UO_368 (O_368,N_14936,N_14949);
or UO_369 (O_369,N_14975,N_14981);
nand UO_370 (O_370,N_14869,N_14967);
xnor UO_371 (O_371,N_14956,N_14947);
nand UO_372 (O_372,N_14880,N_14856);
xor UO_373 (O_373,N_14966,N_14900);
xor UO_374 (O_374,N_14948,N_14932);
nand UO_375 (O_375,N_14996,N_14940);
or UO_376 (O_376,N_14923,N_14928);
and UO_377 (O_377,N_14855,N_14987);
nand UO_378 (O_378,N_14977,N_14894);
nand UO_379 (O_379,N_14902,N_14958);
or UO_380 (O_380,N_14967,N_14965);
nand UO_381 (O_381,N_14970,N_14905);
nand UO_382 (O_382,N_14897,N_14859);
and UO_383 (O_383,N_14895,N_14997);
and UO_384 (O_384,N_14970,N_14953);
or UO_385 (O_385,N_14869,N_14904);
or UO_386 (O_386,N_14864,N_14990);
xor UO_387 (O_387,N_14978,N_14915);
nand UO_388 (O_388,N_14976,N_14863);
xnor UO_389 (O_389,N_14992,N_14893);
nand UO_390 (O_390,N_14883,N_14948);
nor UO_391 (O_391,N_14953,N_14921);
nand UO_392 (O_392,N_14886,N_14933);
nor UO_393 (O_393,N_14935,N_14862);
or UO_394 (O_394,N_14878,N_14926);
nor UO_395 (O_395,N_14954,N_14937);
and UO_396 (O_396,N_14907,N_14867);
nand UO_397 (O_397,N_14879,N_14873);
and UO_398 (O_398,N_14919,N_14976);
nand UO_399 (O_399,N_14999,N_14997);
nor UO_400 (O_400,N_14957,N_14974);
nand UO_401 (O_401,N_14876,N_14935);
nand UO_402 (O_402,N_14961,N_14875);
nor UO_403 (O_403,N_14916,N_14985);
and UO_404 (O_404,N_14919,N_14971);
xor UO_405 (O_405,N_14899,N_14967);
nor UO_406 (O_406,N_14910,N_14913);
nand UO_407 (O_407,N_14893,N_14903);
nor UO_408 (O_408,N_14906,N_14942);
or UO_409 (O_409,N_14965,N_14851);
and UO_410 (O_410,N_14851,N_14949);
and UO_411 (O_411,N_14902,N_14883);
and UO_412 (O_412,N_14992,N_14870);
xor UO_413 (O_413,N_14922,N_14952);
and UO_414 (O_414,N_14921,N_14954);
and UO_415 (O_415,N_14945,N_14897);
xor UO_416 (O_416,N_14937,N_14902);
or UO_417 (O_417,N_14857,N_14864);
and UO_418 (O_418,N_14906,N_14973);
nand UO_419 (O_419,N_14907,N_14855);
or UO_420 (O_420,N_14897,N_14932);
xnor UO_421 (O_421,N_14851,N_14966);
nor UO_422 (O_422,N_14923,N_14903);
xnor UO_423 (O_423,N_14875,N_14966);
xnor UO_424 (O_424,N_14866,N_14969);
or UO_425 (O_425,N_14982,N_14930);
and UO_426 (O_426,N_14927,N_14997);
or UO_427 (O_427,N_14903,N_14936);
and UO_428 (O_428,N_14942,N_14884);
nand UO_429 (O_429,N_14986,N_14965);
or UO_430 (O_430,N_14995,N_14852);
or UO_431 (O_431,N_14859,N_14910);
and UO_432 (O_432,N_14963,N_14871);
or UO_433 (O_433,N_14961,N_14930);
xor UO_434 (O_434,N_14994,N_14890);
nand UO_435 (O_435,N_14968,N_14990);
nor UO_436 (O_436,N_14915,N_14870);
or UO_437 (O_437,N_14983,N_14899);
or UO_438 (O_438,N_14971,N_14850);
xor UO_439 (O_439,N_14924,N_14851);
nand UO_440 (O_440,N_14987,N_14932);
or UO_441 (O_441,N_14971,N_14947);
and UO_442 (O_442,N_14979,N_14877);
nor UO_443 (O_443,N_14865,N_14886);
xnor UO_444 (O_444,N_14851,N_14912);
nand UO_445 (O_445,N_14861,N_14876);
or UO_446 (O_446,N_14992,N_14862);
or UO_447 (O_447,N_14991,N_14992);
xor UO_448 (O_448,N_14871,N_14970);
xnor UO_449 (O_449,N_14905,N_14857);
nor UO_450 (O_450,N_14859,N_14980);
and UO_451 (O_451,N_14860,N_14988);
or UO_452 (O_452,N_14985,N_14958);
nand UO_453 (O_453,N_14954,N_14979);
nor UO_454 (O_454,N_14856,N_14942);
nand UO_455 (O_455,N_14971,N_14893);
or UO_456 (O_456,N_14977,N_14877);
nand UO_457 (O_457,N_14949,N_14971);
xnor UO_458 (O_458,N_14944,N_14966);
xor UO_459 (O_459,N_14936,N_14908);
and UO_460 (O_460,N_14872,N_14934);
nor UO_461 (O_461,N_14973,N_14942);
xor UO_462 (O_462,N_14967,N_14871);
and UO_463 (O_463,N_14966,N_14887);
xor UO_464 (O_464,N_14958,N_14921);
xor UO_465 (O_465,N_14936,N_14977);
xor UO_466 (O_466,N_14984,N_14966);
xor UO_467 (O_467,N_14881,N_14984);
xor UO_468 (O_468,N_14994,N_14856);
or UO_469 (O_469,N_14991,N_14850);
xnor UO_470 (O_470,N_14854,N_14939);
xor UO_471 (O_471,N_14885,N_14869);
and UO_472 (O_472,N_14962,N_14881);
and UO_473 (O_473,N_14916,N_14954);
nand UO_474 (O_474,N_14901,N_14853);
and UO_475 (O_475,N_14965,N_14978);
nor UO_476 (O_476,N_14978,N_14990);
nand UO_477 (O_477,N_14964,N_14864);
nand UO_478 (O_478,N_14880,N_14964);
xnor UO_479 (O_479,N_14927,N_14933);
nor UO_480 (O_480,N_14984,N_14968);
xor UO_481 (O_481,N_14879,N_14966);
or UO_482 (O_482,N_14999,N_14893);
nor UO_483 (O_483,N_14870,N_14896);
and UO_484 (O_484,N_14887,N_14870);
xor UO_485 (O_485,N_14922,N_14971);
nor UO_486 (O_486,N_14986,N_14879);
and UO_487 (O_487,N_14982,N_14957);
nand UO_488 (O_488,N_14940,N_14928);
xor UO_489 (O_489,N_14854,N_14921);
xnor UO_490 (O_490,N_14889,N_14907);
and UO_491 (O_491,N_14916,N_14996);
nand UO_492 (O_492,N_14854,N_14998);
nor UO_493 (O_493,N_14859,N_14959);
xor UO_494 (O_494,N_14851,N_14999);
nand UO_495 (O_495,N_14976,N_14968);
or UO_496 (O_496,N_14877,N_14889);
nor UO_497 (O_497,N_14881,N_14998);
and UO_498 (O_498,N_14930,N_14927);
nor UO_499 (O_499,N_14955,N_14929);
xor UO_500 (O_500,N_14894,N_14868);
and UO_501 (O_501,N_14955,N_14989);
xor UO_502 (O_502,N_14941,N_14894);
xor UO_503 (O_503,N_14850,N_14953);
nand UO_504 (O_504,N_14980,N_14976);
nor UO_505 (O_505,N_14928,N_14958);
and UO_506 (O_506,N_14854,N_14850);
nor UO_507 (O_507,N_14920,N_14992);
nor UO_508 (O_508,N_14934,N_14988);
nor UO_509 (O_509,N_14889,N_14989);
and UO_510 (O_510,N_14960,N_14967);
nand UO_511 (O_511,N_14971,N_14887);
nor UO_512 (O_512,N_14949,N_14858);
or UO_513 (O_513,N_14889,N_14946);
or UO_514 (O_514,N_14930,N_14953);
and UO_515 (O_515,N_14998,N_14965);
nand UO_516 (O_516,N_14913,N_14886);
and UO_517 (O_517,N_14851,N_14907);
nand UO_518 (O_518,N_14876,N_14940);
nand UO_519 (O_519,N_14880,N_14985);
nor UO_520 (O_520,N_14898,N_14857);
xor UO_521 (O_521,N_14880,N_14911);
nand UO_522 (O_522,N_14889,N_14881);
or UO_523 (O_523,N_14883,N_14878);
nand UO_524 (O_524,N_14953,N_14933);
and UO_525 (O_525,N_14853,N_14890);
nand UO_526 (O_526,N_14920,N_14997);
or UO_527 (O_527,N_14974,N_14870);
xor UO_528 (O_528,N_14921,N_14861);
or UO_529 (O_529,N_14884,N_14850);
or UO_530 (O_530,N_14892,N_14957);
nand UO_531 (O_531,N_14990,N_14918);
xnor UO_532 (O_532,N_14958,N_14926);
nor UO_533 (O_533,N_14860,N_14982);
nand UO_534 (O_534,N_14897,N_14942);
and UO_535 (O_535,N_14902,N_14924);
nor UO_536 (O_536,N_14954,N_14969);
nand UO_537 (O_537,N_14988,N_14969);
xnor UO_538 (O_538,N_14937,N_14901);
or UO_539 (O_539,N_14874,N_14864);
or UO_540 (O_540,N_14873,N_14907);
nor UO_541 (O_541,N_14971,N_14876);
nand UO_542 (O_542,N_14860,N_14888);
nor UO_543 (O_543,N_14940,N_14917);
nor UO_544 (O_544,N_14991,N_14952);
xor UO_545 (O_545,N_14913,N_14865);
nor UO_546 (O_546,N_14932,N_14965);
nand UO_547 (O_547,N_14956,N_14996);
xor UO_548 (O_548,N_14866,N_14884);
nor UO_549 (O_549,N_14994,N_14997);
and UO_550 (O_550,N_14958,N_14909);
and UO_551 (O_551,N_14870,N_14932);
nand UO_552 (O_552,N_14948,N_14870);
and UO_553 (O_553,N_14870,N_14963);
nor UO_554 (O_554,N_14881,N_14867);
and UO_555 (O_555,N_14999,N_14894);
nand UO_556 (O_556,N_14951,N_14871);
nor UO_557 (O_557,N_14982,N_14955);
nand UO_558 (O_558,N_14945,N_14895);
nor UO_559 (O_559,N_14991,N_14883);
nor UO_560 (O_560,N_14916,N_14881);
and UO_561 (O_561,N_14865,N_14929);
nor UO_562 (O_562,N_14969,N_14993);
nor UO_563 (O_563,N_14981,N_14861);
or UO_564 (O_564,N_14871,N_14877);
nand UO_565 (O_565,N_14967,N_14948);
or UO_566 (O_566,N_14863,N_14904);
nand UO_567 (O_567,N_14959,N_14944);
nand UO_568 (O_568,N_14939,N_14914);
or UO_569 (O_569,N_14910,N_14851);
nor UO_570 (O_570,N_14894,N_14974);
xnor UO_571 (O_571,N_14941,N_14975);
and UO_572 (O_572,N_14850,N_14987);
nor UO_573 (O_573,N_14854,N_14896);
nor UO_574 (O_574,N_14863,N_14953);
or UO_575 (O_575,N_14916,N_14902);
nor UO_576 (O_576,N_14884,N_14995);
and UO_577 (O_577,N_14886,N_14890);
xor UO_578 (O_578,N_14975,N_14957);
xor UO_579 (O_579,N_14853,N_14895);
nand UO_580 (O_580,N_14884,N_14970);
xnor UO_581 (O_581,N_14958,N_14950);
nor UO_582 (O_582,N_14904,N_14964);
nand UO_583 (O_583,N_14914,N_14965);
nand UO_584 (O_584,N_14915,N_14882);
nor UO_585 (O_585,N_14894,N_14866);
or UO_586 (O_586,N_14984,N_14972);
and UO_587 (O_587,N_14965,N_14948);
xnor UO_588 (O_588,N_14986,N_14951);
and UO_589 (O_589,N_14855,N_14984);
and UO_590 (O_590,N_14902,N_14868);
nand UO_591 (O_591,N_14911,N_14903);
or UO_592 (O_592,N_14875,N_14867);
and UO_593 (O_593,N_14900,N_14994);
xor UO_594 (O_594,N_14876,N_14966);
or UO_595 (O_595,N_14921,N_14994);
and UO_596 (O_596,N_14921,N_14890);
and UO_597 (O_597,N_14854,N_14954);
nand UO_598 (O_598,N_14957,N_14960);
or UO_599 (O_599,N_14939,N_14905);
xnor UO_600 (O_600,N_14931,N_14980);
nand UO_601 (O_601,N_14873,N_14895);
or UO_602 (O_602,N_14892,N_14856);
nand UO_603 (O_603,N_14875,N_14899);
nor UO_604 (O_604,N_14913,N_14901);
and UO_605 (O_605,N_14889,N_14951);
xor UO_606 (O_606,N_14903,N_14889);
nor UO_607 (O_607,N_14918,N_14927);
and UO_608 (O_608,N_14885,N_14901);
xor UO_609 (O_609,N_14891,N_14861);
or UO_610 (O_610,N_14992,N_14939);
nand UO_611 (O_611,N_14867,N_14979);
and UO_612 (O_612,N_14913,N_14918);
nand UO_613 (O_613,N_14989,N_14972);
and UO_614 (O_614,N_14921,N_14996);
nor UO_615 (O_615,N_14975,N_14909);
xor UO_616 (O_616,N_14875,N_14976);
and UO_617 (O_617,N_14879,N_14932);
nand UO_618 (O_618,N_14975,N_14855);
or UO_619 (O_619,N_14853,N_14876);
or UO_620 (O_620,N_14858,N_14893);
and UO_621 (O_621,N_14905,N_14969);
xor UO_622 (O_622,N_14983,N_14967);
and UO_623 (O_623,N_14946,N_14876);
nand UO_624 (O_624,N_14971,N_14983);
nand UO_625 (O_625,N_14979,N_14930);
or UO_626 (O_626,N_14967,N_14873);
and UO_627 (O_627,N_14964,N_14903);
or UO_628 (O_628,N_14956,N_14972);
or UO_629 (O_629,N_14926,N_14939);
xnor UO_630 (O_630,N_14903,N_14864);
or UO_631 (O_631,N_14938,N_14996);
nor UO_632 (O_632,N_14898,N_14931);
or UO_633 (O_633,N_14874,N_14911);
xor UO_634 (O_634,N_14863,N_14917);
nor UO_635 (O_635,N_14955,N_14857);
nand UO_636 (O_636,N_14913,N_14883);
and UO_637 (O_637,N_14876,N_14898);
nand UO_638 (O_638,N_14923,N_14992);
or UO_639 (O_639,N_14867,N_14897);
nor UO_640 (O_640,N_14911,N_14915);
and UO_641 (O_641,N_14938,N_14981);
xnor UO_642 (O_642,N_14863,N_14922);
or UO_643 (O_643,N_14929,N_14884);
nand UO_644 (O_644,N_14881,N_14985);
or UO_645 (O_645,N_14880,N_14995);
xor UO_646 (O_646,N_14889,N_14982);
xnor UO_647 (O_647,N_14962,N_14925);
and UO_648 (O_648,N_14870,N_14949);
nor UO_649 (O_649,N_14879,N_14888);
or UO_650 (O_650,N_14864,N_14867);
nand UO_651 (O_651,N_14977,N_14931);
nand UO_652 (O_652,N_14947,N_14878);
xor UO_653 (O_653,N_14924,N_14897);
and UO_654 (O_654,N_14893,N_14885);
xnor UO_655 (O_655,N_14991,N_14897);
or UO_656 (O_656,N_14978,N_14988);
nor UO_657 (O_657,N_14894,N_14852);
xnor UO_658 (O_658,N_14947,N_14921);
nand UO_659 (O_659,N_14926,N_14882);
nand UO_660 (O_660,N_14922,N_14996);
nand UO_661 (O_661,N_14910,N_14866);
nor UO_662 (O_662,N_14956,N_14999);
or UO_663 (O_663,N_14920,N_14878);
nor UO_664 (O_664,N_14856,N_14996);
or UO_665 (O_665,N_14983,N_14921);
xnor UO_666 (O_666,N_14885,N_14900);
nor UO_667 (O_667,N_14918,N_14923);
nand UO_668 (O_668,N_14956,N_14946);
and UO_669 (O_669,N_14934,N_14915);
nand UO_670 (O_670,N_14928,N_14967);
xor UO_671 (O_671,N_14902,N_14918);
xor UO_672 (O_672,N_14913,N_14894);
or UO_673 (O_673,N_14946,N_14942);
or UO_674 (O_674,N_14955,N_14944);
nand UO_675 (O_675,N_14978,N_14966);
nor UO_676 (O_676,N_14995,N_14953);
nand UO_677 (O_677,N_14905,N_14902);
or UO_678 (O_678,N_14916,N_14914);
or UO_679 (O_679,N_14918,N_14875);
and UO_680 (O_680,N_14850,N_14949);
nand UO_681 (O_681,N_14916,N_14878);
and UO_682 (O_682,N_14898,N_14851);
nand UO_683 (O_683,N_14997,N_14874);
xnor UO_684 (O_684,N_14932,N_14883);
xnor UO_685 (O_685,N_14876,N_14944);
or UO_686 (O_686,N_14953,N_14960);
xor UO_687 (O_687,N_14860,N_14879);
nor UO_688 (O_688,N_14911,N_14995);
xor UO_689 (O_689,N_14958,N_14898);
nor UO_690 (O_690,N_14999,N_14913);
or UO_691 (O_691,N_14858,N_14975);
or UO_692 (O_692,N_14970,N_14974);
or UO_693 (O_693,N_14965,N_14975);
or UO_694 (O_694,N_14872,N_14972);
nor UO_695 (O_695,N_14884,N_14906);
nand UO_696 (O_696,N_14993,N_14934);
or UO_697 (O_697,N_14960,N_14895);
nand UO_698 (O_698,N_14917,N_14987);
nor UO_699 (O_699,N_14893,N_14921);
xnor UO_700 (O_700,N_14931,N_14899);
or UO_701 (O_701,N_14999,N_14965);
nor UO_702 (O_702,N_14949,N_14951);
or UO_703 (O_703,N_14871,N_14965);
or UO_704 (O_704,N_14907,N_14950);
nand UO_705 (O_705,N_14896,N_14954);
xor UO_706 (O_706,N_14893,N_14926);
nor UO_707 (O_707,N_14993,N_14931);
and UO_708 (O_708,N_14948,N_14939);
and UO_709 (O_709,N_14965,N_14971);
and UO_710 (O_710,N_14906,N_14972);
nor UO_711 (O_711,N_14980,N_14977);
or UO_712 (O_712,N_14910,N_14914);
xor UO_713 (O_713,N_14962,N_14947);
nor UO_714 (O_714,N_14899,N_14871);
or UO_715 (O_715,N_14937,N_14946);
nor UO_716 (O_716,N_14893,N_14883);
and UO_717 (O_717,N_14899,N_14977);
or UO_718 (O_718,N_14934,N_14958);
xnor UO_719 (O_719,N_14925,N_14860);
and UO_720 (O_720,N_14939,N_14892);
and UO_721 (O_721,N_14864,N_14905);
xor UO_722 (O_722,N_14892,N_14954);
or UO_723 (O_723,N_14901,N_14961);
xnor UO_724 (O_724,N_14864,N_14877);
xor UO_725 (O_725,N_14891,N_14978);
or UO_726 (O_726,N_14868,N_14994);
and UO_727 (O_727,N_14868,N_14980);
nand UO_728 (O_728,N_14942,N_14992);
nor UO_729 (O_729,N_14942,N_14969);
and UO_730 (O_730,N_14941,N_14921);
xor UO_731 (O_731,N_14977,N_14884);
or UO_732 (O_732,N_14851,N_14922);
xnor UO_733 (O_733,N_14981,N_14973);
or UO_734 (O_734,N_14925,N_14924);
nand UO_735 (O_735,N_14875,N_14941);
and UO_736 (O_736,N_14949,N_14902);
and UO_737 (O_737,N_14989,N_14962);
or UO_738 (O_738,N_14950,N_14915);
and UO_739 (O_739,N_14880,N_14913);
nor UO_740 (O_740,N_14895,N_14936);
or UO_741 (O_741,N_14856,N_14881);
and UO_742 (O_742,N_14968,N_14993);
nand UO_743 (O_743,N_14943,N_14931);
xor UO_744 (O_744,N_14882,N_14984);
nor UO_745 (O_745,N_14964,N_14895);
nand UO_746 (O_746,N_14875,N_14886);
xnor UO_747 (O_747,N_14933,N_14976);
nor UO_748 (O_748,N_14906,N_14901);
or UO_749 (O_749,N_14872,N_14883);
or UO_750 (O_750,N_14937,N_14938);
nor UO_751 (O_751,N_14947,N_14932);
xnor UO_752 (O_752,N_14917,N_14959);
and UO_753 (O_753,N_14878,N_14907);
and UO_754 (O_754,N_14917,N_14956);
and UO_755 (O_755,N_14938,N_14930);
nor UO_756 (O_756,N_14988,N_14906);
xor UO_757 (O_757,N_14966,N_14863);
and UO_758 (O_758,N_14963,N_14938);
or UO_759 (O_759,N_14889,N_14862);
xor UO_760 (O_760,N_14901,N_14984);
nand UO_761 (O_761,N_14871,N_14985);
xor UO_762 (O_762,N_14850,N_14964);
xnor UO_763 (O_763,N_14989,N_14866);
or UO_764 (O_764,N_14951,N_14970);
nor UO_765 (O_765,N_14999,N_14889);
nand UO_766 (O_766,N_14975,N_14937);
nand UO_767 (O_767,N_14934,N_14875);
nor UO_768 (O_768,N_14908,N_14959);
nor UO_769 (O_769,N_14946,N_14966);
or UO_770 (O_770,N_14891,N_14905);
or UO_771 (O_771,N_14912,N_14889);
or UO_772 (O_772,N_14904,N_14915);
or UO_773 (O_773,N_14873,N_14874);
nand UO_774 (O_774,N_14935,N_14971);
xnor UO_775 (O_775,N_14960,N_14986);
or UO_776 (O_776,N_14968,N_14872);
xor UO_777 (O_777,N_14954,N_14911);
and UO_778 (O_778,N_14976,N_14999);
or UO_779 (O_779,N_14928,N_14895);
nand UO_780 (O_780,N_14927,N_14958);
or UO_781 (O_781,N_14970,N_14927);
or UO_782 (O_782,N_14978,N_14985);
nand UO_783 (O_783,N_14920,N_14981);
nor UO_784 (O_784,N_14907,N_14871);
and UO_785 (O_785,N_14906,N_14950);
nand UO_786 (O_786,N_14996,N_14942);
nand UO_787 (O_787,N_14878,N_14868);
nor UO_788 (O_788,N_14921,N_14931);
nand UO_789 (O_789,N_14938,N_14927);
nand UO_790 (O_790,N_14976,N_14937);
nand UO_791 (O_791,N_14956,N_14973);
and UO_792 (O_792,N_14979,N_14923);
or UO_793 (O_793,N_14964,N_14952);
and UO_794 (O_794,N_14965,N_14912);
or UO_795 (O_795,N_14960,N_14887);
nand UO_796 (O_796,N_14868,N_14974);
nand UO_797 (O_797,N_14912,N_14920);
and UO_798 (O_798,N_14961,N_14913);
xor UO_799 (O_799,N_14875,N_14955);
and UO_800 (O_800,N_14889,N_14899);
nor UO_801 (O_801,N_14875,N_14855);
nand UO_802 (O_802,N_14851,N_14967);
or UO_803 (O_803,N_14855,N_14891);
nor UO_804 (O_804,N_14938,N_14876);
and UO_805 (O_805,N_14897,N_14967);
xnor UO_806 (O_806,N_14937,N_14986);
or UO_807 (O_807,N_14902,N_14956);
or UO_808 (O_808,N_14871,N_14957);
or UO_809 (O_809,N_14968,N_14928);
nand UO_810 (O_810,N_14900,N_14955);
xnor UO_811 (O_811,N_14997,N_14915);
and UO_812 (O_812,N_14970,N_14924);
xnor UO_813 (O_813,N_14897,N_14898);
and UO_814 (O_814,N_14916,N_14939);
or UO_815 (O_815,N_14862,N_14998);
nor UO_816 (O_816,N_14974,N_14927);
and UO_817 (O_817,N_14864,N_14931);
or UO_818 (O_818,N_14901,N_14957);
nor UO_819 (O_819,N_14883,N_14960);
nand UO_820 (O_820,N_14972,N_14886);
and UO_821 (O_821,N_14930,N_14949);
nand UO_822 (O_822,N_14908,N_14976);
xnor UO_823 (O_823,N_14893,N_14945);
nor UO_824 (O_824,N_14851,N_14953);
nor UO_825 (O_825,N_14963,N_14916);
nor UO_826 (O_826,N_14948,N_14981);
and UO_827 (O_827,N_14858,N_14904);
and UO_828 (O_828,N_14996,N_14891);
nor UO_829 (O_829,N_14923,N_14878);
or UO_830 (O_830,N_14916,N_14890);
nor UO_831 (O_831,N_14913,N_14959);
xor UO_832 (O_832,N_14894,N_14927);
nand UO_833 (O_833,N_14928,N_14980);
xor UO_834 (O_834,N_14993,N_14951);
and UO_835 (O_835,N_14919,N_14908);
or UO_836 (O_836,N_14856,N_14961);
nand UO_837 (O_837,N_14935,N_14941);
and UO_838 (O_838,N_14892,N_14963);
nor UO_839 (O_839,N_14902,N_14943);
or UO_840 (O_840,N_14857,N_14994);
and UO_841 (O_841,N_14877,N_14894);
and UO_842 (O_842,N_14913,N_14878);
and UO_843 (O_843,N_14925,N_14940);
or UO_844 (O_844,N_14974,N_14918);
or UO_845 (O_845,N_14867,N_14903);
or UO_846 (O_846,N_14995,N_14975);
nor UO_847 (O_847,N_14915,N_14925);
or UO_848 (O_848,N_14952,N_14973);
nand UO_849 (O_849,N_14922,N_14909);
and UO_850 (O_850,N_14864,N_14884);
and UO_851 (O_851,N_14933,N_14873);
and UO_852 (O_852,N_14921,N_14966);
xor UO_853 (O_853,N_14969,N_14941);
nand UO_854 (O_854,N_14918,N_14916);
nand UO_855 (O_855,N_14895,N_14870);
and UO_856 (O_856,N_14958,N_14858);
nor UO_857 (O_857,N_14914,N_14988);
and UO_858 (O_858,N_14880,N_14962);
nor UO_859 (O_859,N_14872,N_14855);
xor UO_860 (O_860,N_14904,N_14931);
or UO_861 (O_861,N_14924,N_14952);
xor UO_862 (O_862,N_14850,N_14941);
xnor UO_863 (O_863,N_14947,N_14994);
nand UO_864 (O_864,N_14857,N_14970);
nor UO_865 (O_865,N_14924,N_14938);
xor UO_866 (O_866,N_14882,N_14891);
nand UO_867 (O_867,N_14890,N_14980);
xnor UO_868 (O_868,N_14995,N_14987);
nor UO_869 (O_869,N_14898,N_14863);
nand UO_870 (O_870,N_14903,N_14869);
nand UO_871 (O_871,N_14979,N_14961);
nor UO_872 (O_872,N_14917,N_14883);
or UO_873 (O_873,N_14977,N_14862);
nor UO_874 (O_874,N_14926,N_14933);
nor UO_875 (O_875,N_14882,N_14864);
nand UO_876 (O_876,N_14876,N_14884);
or UO_877 (O_877,N_14901,N_14908);
xor UO_878 (O_878,N_14983,N_14986);
nor UO_879 (O_879,N_14907,N_14945);
or UO_880 (O_880,N_14965,N_14988);
and UO_881 (O_881,N_14941,N_14874);
nand UO_882 (O_882,N_14917,N_14886);
nor UO_883 (O_883,N_14850,N_14853);
or UO_884 (O_884,N_14889,N_14891);
nand UO_885 (O_885,N_14938,N_14898);
xnor UO_886 (O_886,N_14915,N_14956);
nor UO_887 (O_887,N_14964,N_14915);
nor UO_888 (O_888,N_14909,N_14994);
xor UO_889 (O_889,N_14924,N_14998);
or UO_890 (O_890,N_14895,N_14990);
nand UO_891 (O_891,N_14991,N_14861);
nor UO_892 (O_892,N_14892,N_14986);
or UO_893 (O_893,N_14943,N_14868);
nand UO_894 (O_894,N_14869,N_14965);
or UO_895 (O_895,N_14943,N_14945);
nor UO_896 (O_896,N_14934,N_14940);
and UO_897 (O_897,N_14855,N_14898);
or UO_898 (O_898,N_14902,N_14876);
nor UO_899 (O_899,N_14903,N_14957);
nand UO_900 (O_900,N_14861,N_14901);
nand UO_901 (O_901,N_14996,N_14964);
nor UO_902 (O_902,N_14865,N_14868);
and UO_903 (O_903,N_14890,N_14926);
nand UO_904 (O_904,N_14987,N_14926);
and UO_905 (O_905,N_14896,N_14903);
and UO_906 (O_906,N_14929,N_14973);
and UO_907 (O_907,N_14981,N_14964);
and UO_908 (O_908,N_14914,N_14984);
xnor UO_909 (O_909,N_14959,N_14957);
nor UO_910 (O_910,N_14915,N_14917);
xor UO_911 (O_911,N_14960,N_14888);
nand UO_912 (O_912,N_14863,N_14902);
xnor UO_913 (O_913,N_14961,N_14953);
nand UO_914 (O_914,N_14912,N_14949);
nor UO_915 (O_915,N_14999,N_14862);
xor UO_916 (O_916,N_14966,N_14995);
or UO_917 (O_917,N_14969,N_14996);
nand UO_918 (O_918,N_14908,N_14958);
nand UO_919 (O_919,N_14921,N_14878);
nor UO_920 (O_920,N_14969,N_14924);
nor UO_921 (O_921,N_14856,N_14861);
and UO_922 (O_922,N_14976,N_14854);
or UO_923 (O_923,N_14893,N_14941);
and UO_924 (O_924,N_14921,N_14970);
xor UO_925 (O_925,N_14944,N_14879);
nor UO_926 (O_926,N_14999,N_14904);
nand UO_927 (O_927,N_14960,N_14920);
nand UO_928 (O_928,N_14888,N_14958);
nand UO_929 (O_929,N_14880,N_14980);
and UO_930 (O_930,N_14972,N_14869);
xnor UO_931 (O_931,N_14906,N_14871);
xnor UO_932 (O_932,N_14993,N_14858);
xnor UO_933 (O_933,N_14872,N_14967);
xor UO_934 (O_934,N_14946,N_14873);
nor UO_935 (O_935,N_14880,N_14872);
or UO_936 (O_936,N_14961,N_14886);
and UO_937 (O_937,N_14902,N_14904);
nand UO_938 (O_938,N_14997,N_14888);
and UO_939 (O_939,N_14900,N_14902);
and UO_940 (O_940,N_14913,N_14911);
nand UO_941 (O_941,N_14990,N_14952);
nor UO_942 (O_942,N_14868,N_14954);
and UO_943 (O_943,N_14979,N_14868);
nor UO_944 (O_944,N_14874,N_14933);
or UO_945 (O_945,N_14962,N_14950);
nor UO_946 (O_946,N_14955,N_14953);
nand UO_947 (O_947,N_14859,N_14982);
and UO_948 (O_948,N_14965,N_14859);
xor UO_949 (O_949,N_14902,N_14853);
nand UO_950 (O_950,N_14936,N_14891);
or UO_951 (O_951,N_14911,N_14851);
nand UO_952 (O_952,N_14889,N_14867);
nor UO_953 (O_953,N_14955,N_14927);
and UO_954 (O_954,N_14923,N_14857);
nand UO_955 (O_955,N_14931,N_14974);
or UO_956 (O_956,N_14886,N_14954);
nor UO_957 (O_957,N_14924,N_14975);
xor UO_958 (O_958,N_14978,N_14936);
nor UO_959 (O_959,N_14922,N_14901);
and UO_960 (O_960,N_14984,N_14956);
xor UO_961 (O_961,N_14901,N_14940);
nand UO_962 (O_962,N_14967,N_14862);
and UO_963 (O_963,N_14928,N_14909);
xnor UO_964 (O_964,N_14854,N_14945);
nand UO_965 (O_965,N_14933,N_14889);
xor UO_966 (O_966,N_14904,N_14956);
nor UO_967 (O_967,N_14989,N_14991);
nor UO_968 (O_968,N_14893,N_14906);
nand UO_969 (O_969,N_14929,N_14960);
or UO_970 (O_970,N_14972,N_14926);
nand UO_971 (O_971,N_14962,N_14905);
and UO_972 (O_972,N_14868,N_14963);
nand UO_973 (O_973,N_14926,N_14896);
or UO_974 (O_974,N_14947,N_14999);
xor UO_975 (O_975,N_14877,N_14971);
xnor UO_976 (O_976,N_14857,N_14952);
xor UO_977 (O_977,N_14910,N_14863);
nand UO_978 (O_978,N_14934,N_14866);
nand UO_979 (O_979,N_14995,N_14881);
or UO_980 (O_980,N_14971,N_14980);
and UO_981 (O_981,N_14955,N_14974);
nor UO_982 (O_982,N_14979,N_14871);
or UO_983 (O_983,N_14929,N_14932);
nor UO_984 (O_984,N_14911,N_14931);
and UO_985 (O_985,N_14964,N_14945);
or UO_986 (O_986,N_14908,N_14873);
and UO_987 (O_987,N_14868,N_14870);
xnor UO_988 (O_988,N_14902,N_14881);
or UO_989 (O_989,N_14955,N_14990);
xor UO_990 (O_990,N_14993,N_14926);
xnor UO_991 (O_991,N_14884,N_14990);
and UO_992 (O_992,N_14887,N_14853);
and UO_993 (O_993,N_14904,N_14968);
nand UO_994 (O_994,N_14885,N_14928);
nand UO_995 (O_995,N_14938,N_14955);
and UO_996 (O_996,N_14957,N_14919);
or UO_997 (O_997,N_14928,N_14853);
nand UO_998 (O_998,N_14911,N_14991);
nor UO_999 (O_999,N_14865,N_14884);
nor UO_1000 (O_1000,N_14949,N_14993);
or UO_1001 (O_1001,N_14917,N_14979);
and UO_1002 (O_1002,N_14914,N_14931);
xor UO_1003 (O_1003,N_14966,N_14895);
and UO_1004 (O_1004,N_14854,N_14903);
xor UO_1005 (O_1005,N_14861,N_14927);
nor UO_1006 (O_1006,N_14853,N_14852);
nand UO_1007 (O_1007,N_14966,N_14905);
or UO_1008 (O_1008,N_14966,N_14856);
nand UO_1009 (O_1009,N_14947,N_14873);
xnor UO_1010 (O_1010,N_14874,N_14876);
nor UO_1011 (O_1011,N_14926,N_14982);
nand UO_1012 (O_1012,N_14972,N_14879);
or UO_1013 (O_1013,N_14901,N_14991);
and UO_1014 (O_1014,N_14875,N_14953);
nand UO_1015 (O_1015,N_14926,N_14915);
or UO_1016 (O_1016,N_14861,N_14977);
nor UO_1017 (O_1017,N_14964,N_14987);
xnor UO_1018 (O_1018,N_14884,N_14858);
nand UO_1019 (O_1019,N_14860,N_14863);
and UO_1020 (O_1020,N_14909,N_14944);
nand UO_1021 (O_1021,N_14931,N_14853);
nor UO_1022 (O_1022,N_14879,N_14864);
and UO_1023 (O_1023,N_14918,N_14862);
nand UO_1024 (O_1024,N_14975,N_14888);
and UO_1025 (O_1025,N_14857,N_14995);
or UO_1026 (O_1026,N_14934,N_14889);
and UO_1027 (O_1027,N_14951,N_14911);
nor UO_1028 (O_1028,N_14854,N_14902);
nor UO_1029 (O_1029,N_14951,N_14891);
xnor UO_1030 (O_1030,N_14983,N_14884);
and UO_1031 (O_1031,N_14974,N_14926);
or UO_1032 (O_1032,N_14882,N_14968);
nand UO_1033 (O_1033,N_14929,N_14864);
nor UO_1034 (O_1034,N_14944,N_14851);
and UO_1035 (O_1035,N_14985,N_14896);
and UO_1036 (O_1036,N_14855,N_14964);
nor UO_1037 (O_1037,N_14864,N_14916);
or UO_1038 (O_1038,N_14961,N_14966);
and UO_1039 (O_1039,N_14916,N_14884);
nor UO_1040 (O_1040,N_14909,N_14926);
or UO_1041 (O_1041,N_14948,N_14952);
or UO_1042 (O_1042,N_14984,N_14932);
or UO_1043 (O_1043,N_14870,N_14880);
nor UO_1044 (O_1044,N_14955,N_14911);
and UO_1045 (O_1045,N_14962,N_14923);
xor UO_1046 (O_1046,N_14950,N_14952);
nor UO_1047 (O_1047,N_14879,N_14880);
xor UO_1048 (O_1048,N_14889,N_14884);
and UO_1049 (O_1049,N_14924,N_14850);
nand UO_1050 (O_1050,N_14959,N_14999);
nor UO_1051 (O_1051,N_14963,N_14953);
nand UO_1052 (O_1052,N_14888,N_14963);
nor UO_1053 (O_1053,N_14995,N_14981);
xor UO_1054 (O_1054,N_14871,N_14961);
or UO_1055 (O_1055,N_14936,N_14981);
xor UO_1056 (O_1056,N_14937,N_14992);
or UO_1057 (O_1057,N_14912,N_14874);
or UO_1058 (O_1058,N_14883,N_14983);
or UO_1059 (O_1059,N_14860,N_14852);
or UO_1060 (O_1060,N_14855,N_14923);
or UO_1061 (O_1061,N_14876,N_14860);
nor UO_1062 (O_1062,N_14957,N_14879);
xor UO_1063 (O_1063,N_14872,N_14943);
nand UO_1064 (O_1064,N_14976,N_14864);
or UO_1065 (O_1065,N_14870,N_14958);
nor UO_1066 (O_1066,N_14955,N_14935);
xor UO_1067 (O_1067,N_14927,N_14922);
nor UO_1068 (O_1068,N_14926,N_14920);
and UO_1069 (O_1069,N_14934,N_14862);
and UO_1070 (O_1070,N_14971,N_14932);
nand UO_1071 (O_1071,N_14893,N_14890);
and UO_1072 (O_1072,N_14875,N_14879);
nor UO_1073 (O_1073,N_14988,N_14897);
xnor UO_1074 (O_1074,N_14954,N_14913);
nand UO_1075 (O_1075,N_14964,N_14927);
nor UO_1076 (O_1076,N_14972,N_14987);
nand UO_1077 (O_1077,N_14901,N_14881);
or UO_1078 (O_1078,N_14888,N_14989);
nor UO_1079 (O_1079,N_14885,N_14854);
xnor UO_1080 (O_1080,N_14926,N_14881);
or UO_1081 (O_1081,N_14944,N_14964);
nand UO_1082 (O_1082,N_14985,N_14954);
or UO_1083 (O_1083,N_14974,N_14938);
xnor UO_1084 (O_1084,N_14969,N_14883);
nor UO_1085 (O_1085,N_14918,N_14949);
nand UO_1086 (O_1086,N_14852,N_14938);
xor UO_1087 (O_1087,N_14899,N_14892);
nor UO_1088 (O_1088,N_14881,N_14945);
nand UO_1089 (O_1089,N_14913,N_14908);
nand UO_1090 (O_1090,N_14890,N_14986);
xor UO_1091 (O_1091,N_14984,N_14992);
nor UO_1092 (O_1092,N_14997,N_14991);
xor UO_1093 (O_1093,N_14858,N_14935);
or UO_1094 (O_1094,N_14918,N_14982);
xnor UO_1095 (O_1095,N_14914,N_14964);
nand UO_1096 (O_1096,N_14954,N_14908);
nor UO_1097 (O_1097,N_14858,N_14887);
nand UO_1098 (O_1098,N_14861,N_14872);
xor UO_1099 (O_1099,N_14977,N_14909);
nor UO_1100 (O_1100,N_14898,N_14987);
or UO_1101 (O_1101,N_14902,N_14894);
or UO_1102 (O_1102,N_14997,N_14935);
xor UO_1103 (O_1103,N_14917,N_14888);
or UO_1104 (O_1104,N_14919,N_14893);
xnor UO_1105 (O_1105,N_14951,N_14880);
xor UO_1106 (O_1106,N_14958,N_14862);
xnor UO_1107 (O_1107,N_14956,N_14876);
or UO_1108 (O_1108,N_14993,N_14916);
xor UO_1109 (O_1109,N_14986,N_14909);
xnor UO_1110 (O_1110,N_14931,N_14915);
nand UO_1111 (O_1111,N_14892,N_14976);
nor UO_1112 (O_1112,N_14940,N_14879);
nand UO_1113 (O_1113,N_14909,N_14947);
and UO_1114 (O_1114,N_14966,N_14949);
nand UO_1115 (O_1115,N_14981,N_14913);
or UO_1116 (O_1116,N_14877,N_14978);
or UO_1117 (O_1117,N_14972,N_14977);
nand UO_1118 (O_1118,N_14953,N_14899);
and UO_1119 (O_1119,N_14870,N_14964);
or UO_1120 (O_1120,N_14899,N_14980);
or UO_1121 (O_1121,N_14886,N_14887);
xnor UO_1122 (O_1122,N_14906,N_14956);
or UO_1123 (O_1123,N_14988,N_14870);
xor UO_1124 (O_1124,N_14961,N_14996);
or UO_1125 (O_1125,N_14899,N_14851);
and UO_1126 (O_1126,N_14992,N_14999);
and UO_1127 (O_1127,N_14880,N_14955);
nor UO_1128 (O_1128,N_14914,N_14867);
nor UO_1129 (O_1129,N_14867,N_14887);
nand UO_1130 (O_1130,N_14950,N_14867);
and UO_1131 (O_1131,N_14914,N_14919);
nor UO_1132 (O_1132,N_14855,N_14874);
nand UO_1133 (O_1133,N_14982,N_14944);
nor UO_1134 (O_1134,N_14996,N_14861);
nand UO_1135 (O_1135,N_14901,N_14928);
nor UO_1136 (O_1136,N_14999,N_14994);
xnor UO_1137 (O_1137,N_14862,N_14936);
nor UO_1138 (O_1138,N_14872,N_14990);
xor UO_1139 (O_1139,N_14857,N_14888);
or UO_1140 (O_1140,N_14939,N_14996);
nand UO_1141 (O_1141,N_14904,N_14916);
xnor UO_1142 (O_1142,N_14897,N_14922);
nand UO_1143 (O_1143,N_14890,N_14957);
nand UO_1144 (O_1144,N_14970,N_14863);
nor UO_1145 (O_1145,N_14937,N_14988);
and UO_1146 (O_1146,N_14997,N_14913);
and UO_1147 (O_1147,N_14940,N_14967);
and UO_1148 (O_1148,N_14996,N_14948);
nand UO_1149 (O_1149,N_14976,N_14987);
and UO_1150 (O_1150,N_14992,N_14912);
or UO_1151 (O_1151,N_14890,N_14907);
or UO_1152 (O_1152,N_14885,N_14851);
nand UO_1153 (O_1153,N_14966,N_14850);
nor UO_1154 (O_1154,N_14851,N_14855);
nand UO_1155 (O_1155,N_14947,N_14853);
and UO_1156 (O_1156,N_14922,N_14867);
or UO_1157 (O_1157,N_14900,N_14963);
nor UO_1158 (O_1158,N_14893,N_14873);
nand UO_1159 (O_1159,N_14964,N_14899);
or UO_1160 (O_1160,N_14875,N_14885);
xor UO_1161 (O_1161,N_14998,N_14928);
nand UO_1162 (O_1162,N_14941,N_14993);
nand UO_1163 (O_1163,N_14900,N_14894);
and UO_1164 (O_1164,N_14978,N_14893);
nand UO_1165 (O_1165,N_14850,N_14875);
nor UO_1166 (O_1166,N_14939,N_14877);
nor UO_1167 (O_1167,N_14859,N_14930);
nand UO_1168 (O_1168,N_14931,N_14964);
nor UO_1169 (O_1169,N_14940,N_14893);
nor UO_1170 (O_1170,N_14993,N_14866);
nor UO_1171 (O_1171,N_14862,N_14914);
nor UO_1172 (O_1172,N_14914,N_14856);
nor UO_1173 (O_1173,N_14884,N_14974);
nor UO_1174 (O_1174,N_14864,N_14919);
nor UO_1175 (O_1175,N_14940,N_14889);
xor UO_1176 (O_1176,N_14854,N_14898);
or UO_1177 (O_1177,N_14929,N_14894);
nor UO_1178 (O_1178,N_14967,N_14955);
xor UO_1179 (O_1179,N_14973,N_14905);
or UO_1180 (O_1180,N_14935,N_14946);
xor UO_1181 (O_1181,N_14886,N_14983);
and UO_1182 (O_1182,N_14975,N_14932);
or UO_1183 (O_1183,N_14942,N_14985);
nand UO_1184 (O_1184,N_14974,N_14893);
nand UO_1185 (O_1185,N_14990,N_14889);
nor UO_1186 (O_1186,N_14858,N_14989);
and UO_1187 (O_1187,N_14864,N_14899);
nand UO_1188 (O_1188,N_14875,N_14902);
nor UO_1189 (O_1189,N_14950,N_14946);
xnor UO_1190 (O_1190,N_14924,N_14976);
xnor UO_1191 (O_1191,N_14860,N_14991);
nand UO_1192 (O_1192,N_14989,N_14961);
nor UO_1193 (O_1193,N_14915,N_14872);
nand UO_1194 (O_1194,N_14915,N_14851);
nand UO_1195 (O_1195,N_14942,N_14979);
and UO_1196 (O_1196,N_14882,N_14901);
nand UO_1197 (O_1197,N_14926,N_14902);
or UO_1198 (O_1198,N_14966,N_14907);
and UO_1199 (O_1199,N_14963,N_14982);
xnor UO_1200 (O_1200,N_14974,N_14998);
nor UO_1201 (O_1201,N_14916,N_14966);
and UO_1202 (O_1202,N_14887,N_14988);
nor UO_1203 (O_1203,N_14942,N_14943);
nand UO_1204 (O_1204,N_14894,N_14963);
and UO_1205 (O_1205,N_14874,N_14927);
and UO_1206 (O_1206,N_14950,N_14919);
nor UO_1207 (O_1207,N_14869,N_14975);
and UO_1208 (O_1208,N_14897,N_14915);
and UO_1209 (O_1209,N_14903,N_14882);
and UO_1210 (O_1210,N_14862,N_14929);
or UO_1211 (O_1211,N_14863,N_14991);
xor UO_1212 (O_1212,N_14867,N_14976);
nand UO_1213 (O_1213,N_14925,N_14884);
and UO_1214 (O_1214,N_14908,N_14876);
nor UO_1215 (O_1215,N_14884,N_14998);
xnor UO_1216 (O_1216,N_14975,N_14940);
nand UO_1217 (O_1217,N_14885,N_14905);
xor UO_1218 (O_1218,N_14976,N_14974);
and UO_1219 (O_1219,N_14965,N_14880);
and UO_1220 (O_1220,N_14984,N_14861);
or UO_1221 (O_1221,N_14946,N_14983);
nand UO_1222 (O_1222,N_14991,N_14878);
and UO_1223 (O_1223,N_14960,N_14857);
and UO_1224 (O_1224,N_14906,N_14913);
nand UO_1225 (O_1225,N_14902,N_14950);
nor UO_1226 (O_1226,N_14920,N_14901);
or UO_1227 (O_1227,N_14967,N_14943);
nand UO_1228 (O_1228,N_14988,N_14912);
nor UO_1229 (O_1229,N_14964,N_14886);
nor UO_1230 (O_1230,N_14883,N_14987);
and UO_1231 (O_1231,N_14870,N_14856);
xor UO_1232 (O_1232,N_14987,N_14960);
nand UO_1233 (O_1233,N_14912,N_14975);
nor UO_1234 (O_1234,N_14871,N_14976);
and UO_1235 (O_1235,N_14988,N_14942);
and UO_1236 (O_1236,N_14973,N_14860);
or UO_1237 (O_1237,N_14864,N_14909);
or UO_1238 (O_1238,N_14912,N_14870);
xnor UO_1239 (O_1239,N_14985,N_14931);
nor UO_1240 (O_1240,N_14885,N_14992);
nor UO_1241 (O_1241,N_14922,N_14920);
nand UO_1242 (O_1242,N_14881,N_14886);
or UO_1243 (O_1243,N_14855,N_14974);
and UO_1244 (O_1244,N_14990,N_14937);
and UO_1245 (O_1245,N_14929,N_14903);
and UO_1246 (O_1246,N_14884,N_14933);
or UO_1247 (O_1247,N_14943,N_14924);
xor UO_1248 (O_1248,N_14921,N_14885);
nor UO_1249 (O_1249,N_14956,N_14925);
nor UO_1250 (O_1250,N_14987,N_14944);
xor UO_1251 (O_1251,N_14921,N_14891);
or UO_1252 (O_1252,N_14907,N_14977);
nand UO_1253 (O_1253,N_14864,N_14963);
xnor UO_1254 (O_1254,N_14869,N_14961);
xnor UO_1255 (O_1255,N_14980,N_14915);
nor UO_1256 (O_1256,N_14850,N_14899);
or UO_1257 (O_1257,N_14929,N_14915);
nor UO_1258 (O_1258,N_14858,N_14914);
nor UO_1259 (O_1259,N_14904,N_14866);
nand UO_1260 (O_1260,N_14858,N_14857);
xor UO_1261 (O_1261,N_14984,N_14925);
or UO_1262 (O_1262,N_14880,N_14998);
and UO_1263 (O_1263,N_14973,N_14853);
nand UO_1264 (O_1264,N_14979,N_14975);
or UO_1265 (O_1265,N_14948,N_14998);
xnor UO_1266 (O_1266,N_14963,N_14941);
and UO_1267 (O_1267,N_14872,N_14890);
nand UO_1268 (O_1268,N_14971,N_14963);
or UO_1269 (O_1269,N_14951,N_14927);
or UO_1270 (O_1270,N_14983,N_14985);
nand UO_1271 (O_1271,N_14885,N_14980);
or UO_1272 (O_1272,N_14958,N_14867);
xnor UO_1273 (O_1273,N_14855,N_14911);
xnor UO_1274 (O_1274,N_14889,N_14935);
and UO_1275 (O_1275,N_14853,N_14908);
or UO_1276 (O_1276,N_14922,N_14978);
and UO_1277 (O_1277,N_14981,N_14855);
and UO_1278 (O_1278,N_14928,N_14878);
nor UO_1279 (O_1279,N_14909,N_14987);
xnor UO_1280 (O_1280,N_14915,N_14892);
nand UO_1281 (O_1281,N_14988,N_14971);
and UO_1282 (O_1282,N_14928,N_14941);
and UO_1283 (O_1283,N_14967,N_14958);
or UO_1284 (O_1284,N_14971,N_14869);
or UO_1285 (O_1285,N_14884,N_14912);
nand UO_1286 (O_1286,N_14859,N_14995);
nor UO_1287 (O_1287,N_14856,N_14941);
nor UO_1288 (O_1288,N_14878,N_14989);
nor UO_1289 (O_1289,N_14969,N_14999);
or UO_1290 (O_1290,N_14968,N_14852);
or UO_1291 (O_1291,N_14882,N_14912);
nand UO_1292 (O_1292,N_14923,N_14866);
nor UO_1293 (O_1293,N_14944,N_14859);
or UO_1294 (O_1294,N_14907,N_14861);
or UO_1295 (O_1295,N_14923,N_14998);
nor UO_1296 (O_1296,N_14879,N_14999);
or UO_1297 (O_1297,N_14929,N_14866);
and UO_1298 (O_1298,N_14962,N_14878);
nand UO_1299 (O_1299,N_14935,N_14970);
and UO_1300 (O_1300,N_14988,N_14922);
and UO_1301 (O_1301,N_14976,N_14865);
xnor UO_1302 (O_1302,N_14894,N_14990);
and UO_1303 (O_1303,N_14982,N_14861);
or UO_1304 (O_1304,N_14966,N_14935);
and UO_1305 (O_1305,N_14892,N_14943);
or UO_1306 (O_1306,N_14987,N_14853);
nor UO_1307 (O_1307,N_14894,N_14940);
nor UO_1308 (O_1308,N_14903,N_14871);
nor UO_1309 (O_1309,N_14875,N_14898);
nand UO_1310 (O_1310,N_14970,N_14980);
nand UO_1311 (O_1311,N_14854,N_14851);
nand UO_1312 (O_1312,N_14938,N_14976);
nor UO_1313 (O_1313,N_14870,N_14942);
and UO_1314 (O_1314,N_14859,N_14916);
nor UO_1315 (O_1315,N_14870,N_14897);
nor UO_1316 (O_1316,N_14973,N_14875);
nand UO_1317 (O_1317,N_14889,N_14938);
xor UO_1318 (O_1318,N_14950,N_14979);
and UO_1319 (O_1319,N_14854,N_14952);
or UO_1320 (O_1320,N_14912,N_14904);
nand UO_1321 (O_1321,N_14992,N_14851);
and UO_1322 (O_1322,N_14939,N_14936);
or UO_1323 (O_1323,N_14885,N_14884);
nor UO_1324 (O_1324,N_14909,N_14897);
nor UO_1325 (O_1325,N_14876,N_14968);
or UO_1326 (O_1326,N_14883,N_14949);
nor UO_1327 (O_1327,N_14908,N_14883);
xor UO_1328 (O_1328,N_14940,N_14927);
nor UO_1329 (O_1329,N_14885,N_14962);
xnor UO_1330 (O_1330,N_14963,N_14883);
or UO_1331 (O_1331,N_14873,N_14903);
or UO_1332 (O_1332,N_14856,N_14864);
xor UO_1333 (O_1333,N_14880,N_14866);
xnor UO_1334 (O_1334,N_14938,N_14944);
and UO_1335 (O_1335,N_14924,N_14944);
or UO_1336 (O_1336,N_14868,N_14993);
or UO_1337 (O_1337,N_14936,N_14914);
or UO_1338 (O_1338,N_14899,N_14933);
or UO_1339 (O_1339,N_14878,N_14965);
and UO_1340 (O_1340,N_14905,N_14938);
and UO_1341 (O_1341,N_14936,N_14962);
xor UO_1342 (O_1342,N_14945,N_14956);
nor UO_1343 (O_1343,N_14971,N_14910);
and UO_1344 (O_1344,N_14863,N_14912);
nand UO_1345 (O_1345,N_14957,N_14881);
nand UO_1346 (O_1346,N_14999,N_14891);
nand UO_1347 (O_1347,N_14929,N_14987);
nor UO_1348 (O_1348,N_14881,N_14906);
nand UO_1349 (O_1349,N_14955,N_14999);
nand UO_1350 (O_1350,N_14951,N_14853);
or UO_1351 (O_1351,N_14928,N_14959);
nor UO_1352 (O_1352,N_14928,N_14969);
nand UO_1353 (O_1353,N_14862,N_14915);
xnor UO_1354 (O_1354,N_14910,N_14873);
nand UO_1355 (O_1355,N_14926,N_14894);
and UO_1356 (O_1356,N_14942,N_14957);
and UO_1357 (O_1357,N_14956,N_14871);
and UO_1358 (O_1358,N_14917,N_14929);
nor UO_1359 (O_1359,N_14903,N_14951);
and UO_1360 (O_1360,N_14933,N_14915);
xor UO_1361 (O_1361,N_14931,N_14854);
or UO_1362 (O_1362,N_14875,N_14963);
xor UO_1363 (O_1363,N_14873,N_14998);
xor UO_1364 (O_1364,N_14897,N_14958);
xor UO_1365 (O_1365,N_14915,N_14896);
xor UO_1366 (O_1366,N_14949,N_14979);
nor UO_1367 (O_1367,N_14882,N_14941);
or UO_1368 (O_1368,N_14980,N_14854);
and UO_1369 (O_1369,N_14865,N_14994);
and UO_1370 (O_1370,N_14966,N_14933);
nand UO_1371 (O_1371,N_14986,N_14942);
and UO_1372 (O_1372,N_14874,N_14994);
nor UO_1373 (O_1373,N_14949,N_14964);
and UO_1374 (O_1374,N_14992,N_14900);
and UO_1375 (O_1375,N_14857,N_14894);
nor UO_1376 (O_1376,N_14979,N_14978);
xor UO_1377 (O_1377,N_14856,N_14981);
and UO_1378 (O_1378,N_14977,N_14988);
nand UO_1379 (O_1379,N_14881,N_14912);
and UO_1380 (O_1380,N_14875,N_14932);
nor UO_1381 (O_1381,N_14919,N_14907);
xor UO_1382 (O_1382,N_14964,N_14897);
or UO_1383 (O_1383,N_14947,N_14899);
xor UO_1384 (O_1384,N_14881,N_14911);
nand UO_1385 (O_1385,N_14977,N_14880);
xnor UO_1386 (O_1386,N_14981,N_14934);
nor UO_1387 (O_1387,N_14974,N_14862);
and UO_1388 (O_1388,N_14904,N_14959);
and UO_1389 (O_1389,N_14990,N_14993);
or UO_1390 (O_1390,N_14871,N_14909);
and UO_1391 (O_1391,N_14910,N_14905);
xnor UO_1392 (O_1392,N_14943,N_14974);
nor UO_1393 (O_1393,N_14874,N_14960);
nor UO_1394 (O_1394,N_14939,N_14974);
nand UO_1395 (O_1395,N_14999,N_14882);
xnor UO_1396 (O_1396,N_14924,N_14993);
xnor UO_1397 (O_1397,N_14924,N_14933);
or UO_1398 (O_1398,N_14968,N_14920);
xnor UO_1399 (O_1399,N_14973,N_14913);
or UO_1400 (O_1400,N_14899,N_14935);
nor UO_1401 (O_1401,N_14959,N_14873);
nand UO_1402 (O_1402,N_14956,N_14884);
xor UO_1403 (O_1403,N_14951,N_14884);
nand UO_1404 (O_1404,N_14933,N_14857);
nor UO_1405 (O_1405,N_14901,N_14941);
or UO_1406 (O_1406,N_14926,N_14951);
and UO_1407 (O_1407,N_14921,N_14863);
and UO_1408 (O_1408,N_14982,N_14956);
and UO_1409 (O_1409,N_14961,N_14922);
xnor UO_1410 (O_1410,N_14958,N_14905);
and UO_1411 (O_1411,N_14886,N_14891);
nor UO_1412 (O_1412,N_14949,N_14955);
nor UO_1413 (O_1413,N_14870,N_14860);
xor UO_1414 (O_1414,N_14994,N_14920);
xnor UO_1415 (O_1415,N_14860,N_14998);
nor UO_1416 (O_1416,N_14907,N_14949);
nand UO_1417 (O_1417,N_14883,N_14887);
xor UO_1418 (O_1418,N_14876,N_14852);
xnor UO_1419 (O_1419,N_14859,N_14876);
xor UO_1420 (O_1420,N_14916,N_14930);
or UO_1421 (O_1421,N_14997,N_14907);
nand UO_1422 (O_1422,N_14903,N_14978);
and UO_1423 (O_1423,N_14879,N_14987);
and UO_1424 (O_1424,N_14919,N_14962);
and UO_1425 (O_1425,N_14909,N_14888);
or UO_1426 (O_1426,N_14947,N_14910);
or UO_1427 (O_1427,N_14955,N_14864);
and UO_1428 (O_1428,N_14908,N_14923);
nand UO_1429 (O_1429,N_14964,N_14858);
and UO_1430 (O_1430,N_14860,N_14993);
nor UO_1431 (O_1431,N_14955,N_14860);
xnor UO_1432 (O_1432,N_14941,N_14983);
xnor UO_1433 (O_1433,N_14929,N_14882);
or UO_1434 (O_1434,N_14949,N_14947);
or UO_1435 (O_1435,N_14942,N_14944);
or UO_1436 (O_1436,N_14995,N_14917);
or UO_1437 (O_1437,N_14933,N_14980);
nor UO_1438 (O_1438,N_14953,N_14968);
or UO_1439 (O_1439,N_14989,N_14956);
nor UO_1440 (O_1440,N_14908,N_14884);
and UO_1441 (O_1441,N_14883,N_14911);
and UO_1442 (O_1442,N_14960,N_14882);
and UO_1443 (O_1443,N_14903,N_14876);
nor UO_1444 (O_1444,N_14873,N_14945);
or UO_1445 (O_1445,N_14860,N_14965);
nand UO_1446 (O_1446,N_14970,N_14969);
and UO_1447 (O_1447,N_14888,N_14911);
nand UO_1448 (O_1448,N_14934,N_14913);
xnor UO_1449 (O_1449,N_14954,N_14942);
nor UO_1450 (O_1450,N_14894,N_14946);
nand UO_1451 (O_1451,N_14927,N_14991);
nand UO_1452 (O_1452,N_14897,N_14954);
and UO_1453 (O_1453,N_14962,N_14870);
and UO_1454 (O_1454,N_14867,N_14893);
nor UO_1455 (O_1455,N_14863,N_14925);
xnor UO_1456 (O_1456,N_14881,N_14976);
and UO_1457 (O_1457,N_14967,N_14874);
nand UO_1458 (O_1458,N_14937,N_14865);
or UO_1459 (O_1459,N_14953,N_14991);
nor UO_1460 (O_1460,N_14959,N_14890);
nor UO_1461 (O_1461,N_14942,N_14983);
and UO_1462 (O_1462,N_14882,N_14978);
nor UO_1463 (O_1463,N_14906,N_14980);
nand UO_1464 (O_1464,N_14888,N_14876);
xor UO_1465 (O_1465,N_14921,N_14998);
nand UO_1466 (O_1466,N_14982,N_14890);
and UO_1467 (O_1467,N_14966,N_14952);
and UO_1468 (O_1468,N_14996,N_14875);
or UO_1469 (O_1469,N_14869,N_14949);
nor UO_1470 (O_1470,N_14906,N_14919);
xnor UO_1471 (O_1471,N_14912,N_14991);
and UO_1472 (O_1472,N_14955,N_14936);
nor UO_1473 (O_1473,N_14866,N_14900);
xnor UO_1474 (O_1474,N_14891,N_14906);
or UO_1475 (O_1475,N_14970,N_14859);
nand UO_1476 (O_1476,N_14893,N_14983);
or UO_1477 (O_1477,N_14997,N_14906);
and UO_1478 (O_1478,N_14929,N_14945);
and UO_1479 (O_1479,N_14939,N_14896);
or UO_1480 (O_1480,N_14904,N_14884);
and UO_1481 (O_1481,N_14974,N_14991);
xor UO_1482 (O_1482,N_14909,N_14861);
or UO_1483 (O_1483,N_14979,N_14908);
nor UO_1484 (O_1484,N_14930,N_14877);
and UO_1485 (O_1485,N_14871,N_14983);
nor UO_1486 (O_1486,N_14989,N_14996);
nor UO_1487 (O_1487,N_14934,N_14942);
xnor UO_1488 (O_1488,N_14982,N_14988);
or UO_1489 (O_1489,N_14874,N_14962);
nor UO_1490 (O_1490,N_14888,N_14943);
nand UO_1491 (O_1491,N_14960,N_14916);
nor UO_1492 (O_1492,N_14937,N_14908);
xor UO_1493 (O_1493,N_14954,N_14984);
xnor UO_1494 (O_1494,N_14966,N_14959);
nand UO_1495 (O_1495,N_14889,N_14925);
or UO_1496 (O_1496,N_14870,N_14981);
or UO_1497 (O_1497,N_14905,N_14945);
nor UO_1498 (O_1498,N_14915,N_14991);
nand UO_1499 (O_1499,N_14859,N_14915);
xnor UO_1500 (O_1500,N_14856,N_14951);
or UO_1501 (O_1501,N_14906,N_14966);
xor UO_1502 (O_1502,N_14982,N_14854);
nor UO_1503 (O_1503,N_14920,N_14990);
nor UO_1504 (O_1504,N_14850,N_14903);
nand UO_1505 (O_1505,N_14878,N_14949);
nand UO_1506 (O_1506,N_14899,N_14916);
or UO_1507 (O_1507,N_14864,N_14983);
nor UO_1508 (O_1508,N_14996,N_14851);
xnor UO_1509 (O_1509,N_14868,N_14856);
xor UO_1510 (O_1510,N_14944,N_14999);
xor UO_1511 (O_1511,N_14864,N_14951);
nor UO_1512 (O_1512,N_14904,N_14950);
or UO_1513 (O_1513,N_14874,N_14887);
nor UO_1514 (O_1514,N_14989,N_14852);
xor UO_1515 (O_1515,N_14937,N_14867);
or UO_1516 (O_1516,N_14929,N_14905);
and UO_1517 (O_1517,N_14851,N_14923);
xnor UO_1518 (O_1518,N_14968,N_14854);
or UO_1519 (O_1519,N_14906,N_14862);
and UO_1520 (O_1520,N_14998,N_14914);
or UO_1521 (O_1521,N_14859,N_14933);
and UO_1522 (O_1522,N_14933,N_14891);
xnor UO_1523 (O_1523,N_14927,N_14935);
or UO_1524 (O_1524,N_14977,N_14942);
and UO_1525 (O_1525,N_14925,N_14972);
and UO_1526 (O_1526,N_14943,N_14954);
nor UO_1527 (O_1527,N_14999,N_14935);
nand UO_1528 (O_1528,N_14908,N_14994);
and UO_1529 (O_1529,N_14869,N_14895);
nor UO_1530 (O_1530,N_14936,N_14917);
and UO_1531 (O_1531,N_14854,N_14910);
nand UO_1532 (O_1532,N_14902,N_14886);
or UO_1533 (O_1533,N_14933,N_14879);
or UO_1534 (O_1534,N_14866,N_14909);
nor UO_1535 (O_1535,N_14861,N_14889);
and UO_1536 (O_1536,N_14939,N_14994);
nor UO_1537 (O_1537,N_14992,N_14852);
xnor UO_1538 (O_1538,N_14960,N_14972);
nor UO_1539 (O_1539,N_14928,N_14861);
nand UO_1540 (O_1540,N_14919,N_14944);
or UO_1541 (O_1541,N_14990,N_14874);
or UO_1542 (O_1542,N_14935,N_14960);
or UO_1543 (O_1543,N_14893,N_14899);
nor UO_1544 (O_1544,N_14927,N_14919);
nand UO_1545 (O_1545,N_14967,N_14865);
or UO_1546 (O_1546,N_14982,N_14911);
xnor UO_1547 (O_1547,N_14990,N_14939);
xor UO_1548 (O_1548,N_14992,N_14983);
or UO_1549 (O_1549,N_14974,N_14910);
or UO_1550 (O_1550,N_14927,N_14957);
nor UO_1551 (O_1551,N_14994,N_14923);
xor UO_1552 (O_1552,N_14975,N_14922);
xnor UO_1553 (O_1553,N_14991,N_14876);
nand UO_1554 (O_1554,N_14959,N_14940);
or UO_1555 (O_1555,N_14936,N_14869);
nand UO_1556 (O_1556,N_14943,N_14972);
and UO_1557 (O_1557,N_14855,N_14929);
nand UO_1558 (O_1558,N_14875,N_14884);
and UO_1559 (O_1559,N_14962,N_14900);
nand UO_1560 (O_1560,N_14970,N_14851);
and UO_1561 (O_1561,N_14888,N_14892);
nand UO_1562 (O_1562,N_14910,N_14909);
nand UO_1563 (O_1563,N_14897,N_14940);
nor UO_1564 (O_1564,N_14860,N_14908);
or UO_1565 (O_1565,N_14917,N_14981);
xnor UO_1566 (O_1566,N_14991,N_14935);
nor UO_1567 (O_1567,N_14909,N_14875);
nor UO_1568 (O_1568,N_14936,N_14889);
nand UO_1569 (O_1569,N_14936,N_14938);
xor UO_1570 (O_1570,N_14875,N_14873);
xor UO_1571 (O_1571,N_14913,N_14852);
or UO_1572 (O_1572,N_14896,N_14964);
nor UO_1573 (O_1573,N_14917,N_14880);
nor UO_1574 (O_1574,N_14958,N_14895);
and UO_1575 (O_1575,N_14905,N_14895);
xor UO_1576 (O_1576,N_14956,N_14863);
nor UO_1577 (O_1577,N_14906,N_14953);
nor UO_1578 (O_1578,N_14871,N_14988);
nand UO_1579 (O_1579,N_14879,N_14927);
and UO_1580 (O_1580,N_14981,N_14852);
xor UO_1581 (O_1581,N_14863,N_14877);
nand UO_1582 (O_1582,N_14932,N_14900);
nand UO_1583 (O_1583,N_14903,N_14930);
nand UO_1584 (O_1584,N_14926,N_14850);
nor UO_1585 (O_1585,N_14996,N_14869);
xnor UO_1586 (O_1586,N_14979,N_14935);
nor UO_1587 (O_1587,N_14994,N_14854);
nand UO_1588 (O_1588,N_14924,N_14931);
xor UO_1589 (O_1589,N_14977,N_14984);
nand UO_1590 (O_1590,N_14926,N_14854);
nor UO_1591 (O_1591,N_14916,N_14983);
nor UO_1592 (O_1592,N_14985,N_14895);
and UO_1593 (O_1593,N_14900,N_14991);
nor UO_1594 (O_1594,N_14876,N_14901);
or UO_1595 (O_1595,N_14945,N_14996);
or UO_1596 (O_1596,N_14861,N_14871);
and UO_1597 (O_1597,N_14949,N_14972);
nand UO_1598 (O_1598,N_14916,N_14928);
nand UO_1599 (O_1599,N_14912,N_14933);
nor UO_1600 (O_1600,N_14963,N_14958);
xor UO_1601 (O_1601,N_14885,N_14932);
nand UO_1602 (O_1602,N_14984,N_14892);
and UO_1603 (O_1603,N_14981,N_14869);
nor UO_1604 (O_1604,N_14918,N_14929);
or UO_1605 (O_1605,N_14937,N_14921);
nor UO_1606 (O_1606,N_14926,N_14988);
nor UO_1607 (O_1607,N_14922,N_14883);
nor UO_1608 (O_1608,N_14994,N_14915);
or UO_1609 (O_1609,N_14888,N_14865);
nor UO_1610 (O_1610,N_14980,N_14893);
or UO_1611 (O_1611,N_14992,N_14978);
and UO_1612 (O_1612,N_14932,N_14949);
or UO_1613 (O_1613,N_14991,N_14919);
nand UO_1614 (O_1614,N_14904,N_14925);
or UO_1615 (O_1615,N_14973,N_14896);
xor UO_1616 (O_1616,N_14894,N_14883);
nor UO_1617 (O_1617,N_14850,N_14883);
nor UO_1618 (O_1618,N_14942,N_14872);
xor UO_1619 (O_1619,N_14852,N_14973);
or UO_1620 (O_1620,N_14901,N_14916);
xor UO_1621 (O_1621,N_14935,N_14900);
or UO_1622 (O_1622,N_14945,N_14914);
or UO_1623 (O_1623,N_14968,N_14910);
nand UO_1624 (O_1624,N_14923,N_14946);
and UO_1625 (O_1625,N_14870,N_14926);
nor UO_1626 (O_1626,N_14947,N_14898);
nand UO_1627 (O_1627,N_14918,N_14998);
nor UO_1628 (O_1628,N_14947,N_14875);
nand UO_1629 (O_1629,N_14871,N_14916);
nand UO_1630 (O_1630,N_14958,N_14889);
or UO_1631 (O_1631,N_14964,N_14937);
and UO_1632 (O_1632,N_14979,N_14861);
or UO_1633 (O_1633,N_14891,N_14939);
and UO_1634 (O_1634,N_14936,N_14984);
or UO_1635 (O_1635,N_14939,N_14853);
xor UO_1636 (O_1636,N_14975,N_14914);
nor UO_1637 (O_1637,N_14852,N_14863);
and UO_1638 (O_1638,N_14874,N_14952);
or UO_1639 (O_1639,N_14921,N_14892);
or UO_1640 (O_1640,N_14956,N_14910);
xnor UO_1641 (O_1641,N_14859,N_14966);
nand UO_1642 (O_1642,N_14969,N_14932);
xnor UO_1643 (O_1643,N_14952,N_14891);
xor UO_1644 (O_1644,N_14977,N_14858);
xnor UO_1645 (O_1645,N_14858,N_14901);
nand UO_1646 (O_1646,N_14890,N_14871);
nor UO_1647 (O_1647,N_14915,N_14852);
nand UO_1648 (O_1648,N_14971,N_14866);
xor UO_1649 (O_1649,N_14926,N_14986);
nand UO_1650 (O_1650,N_14886,N_14923);
and UO_1651 (O_1651,N_14898,N_14921);
or UO_1652 (O_1652,N_14996,N_14977);
and UO_1653 (O_1653,N_14978,N_14909);
or UO_1654 (O_1654,N_14919,N_14885);
and UO_1655 (O_1655,N_14856,N_14985);
nor UO_1656 (O_1656,N_14964,N_14891);
nand UO_1657 (O_1657,N_14953,N_14895);
or UO_1658 (O_1658,N_14889,N_14909);
or UO_1659 (O_1659,N_14974,N_14909);
and UO_1660 (O_1660,N_14924,N_14880);
xor UO_1661 (O_1661,N_14881,N_14875);
nor UO_1662 (O_1662,N_14884,N_14957);
xnor UO_1663 (O_1663,N_14912,N_14877);
nand UO_1664 (O_1664,N_14968,N_14977);
nor UO_1665 (O_1665,N_14926,N_14872);
nor UO_1666 (O_1666,N_14854,N_14881);
or UO_1667 (O_1667,N_14895,N_14994);
or UO_1668 (O_1668,N_14980,N_14990);
and UO_1669 (O_1669,N_14944,N_14878);
xor UO_1670 (O_1670,N_14956,N_14888);
nand UO_1671 (O_1671,N_14931,N_14895);
and UO_1672 (O_1672,N_14921,N_14948);
or UO_1673 (O_1673,N_14911,N_14897);
or UO_1674 (O_1674,N_14861,N_14875);
nor UO_1675 (O_1675,N_14868,N_14951);
nor UO_1676 (O_1676,N_14933,N_14885);
xnor UO_1677 (O_1677,N_14976,N_14876);
and UO_1678 (O_1678,N_14996,N_14966);
nor UO_1679 (O_1679,N_14945,N_14940);
or UO_1680 (O_1680,N_14987,N_14866);
xor UO_1681 (O_1681,N_14934,N_14968);
and UO_1682 (O_1682,N_14869,N_14993);
xnor UO_1683 (O_1683,N_14957,N_14934);
xor UO_1684 (O_1684,N_14896,N_14975);
or UO_1685 (O_1685,N_14896,N_14859);
nand UO_1686 (O_1686,N_14893,N_14962);
or UO_1687 (O_1687,N_14885,N_14855);
or UO_1688 (O_1688,N_14899,N_14926);
or UO_1689 (O_1689,N_14891,N_14919);
nand UO_1690 (O_1690,N_14945,N_14969);
xor UO_1691 (O_1691,N_14974,N_14919);
nand UO_1692 (O_1692,N_14860,N_14855);
or UO_1693 (O_1693,N_14885,N_14991);
and UO_1694 (O_1694,N_14928,N_14881);
nor UO_1695 (O_1695,N_14876,N_14890);
xnor UO_1696 (O_1696,N_14918,N_14888);
nor UO_1697 (O_1697,N_14865,N_14936);
or UO_1698 (O_1698,N_14931,N_14929);
and UO_1699 (O_1699,N_14919,N_14981);
xnor UO_1700 (O_1700,N_14990,N_14873);
nand UO_1701 (O_1701,N_14882,N_14871);
nor UO_1702 (O_1702,N_14869,N_14959);
xnor UO_1703 (O_1703,N_14978,N_14950);
or UO_1704 (O_1704,N_14977,N_14973);
or UO_1705 (O_1705,N_14910,N_14986);
xor UO_1706 (O_1706,N_14952,N_14893);
nor UO_1707 (O_1707,N_14965,N_14921);
nand UO_1708 (O_1708,N_14977,N_14940);
or UO_1709 (O_1709,N_14924,N_14972);
xor UO_1710 (O_1710,N_14921,N_14902);
xor UO_1711 (O_1711,N_14919,N_14966);
and UO_1712 (O_1712,N_14975,N_14952);
nand UO_1713 (O_1713,N_14963,N_14979);
or UO_1714 (O_1714,N_14851,N_14947);
and UO_1715 (O_1715,N_14992,N_14967);
nand UO_1716 (O_1716,N_14894,N_14873);
and UO_1717 (O_1717,N_14920,N_14959);
and UO_1718 (O_1718,N_14915,N_14998);
and UO_1719 (O_1719,N_14890,N_14942);
nor UO_1720 (O_1720,N_14929,N_14980);
nor UO_1721 (O_1721,N_14864,N_14853);
nand UO_1722 (O_1722,N_14907,N_14940);
and UO_1723 (O_1723,N_14975,N_14880);
and UO_1724 (O_1724,N_14933,N_14996);
xor UO_1725 (O_1725,N_14850,N_14948);
or UO_1726 (O_1726,N_14989,N_14880);
nor UO_1727 (O_1727,N_14881,N_14975);
or UO_1728 (O_1728,N_14868,N_14896);
xnor UO_1729 (O_1729,N_14878,N_14983);
and UO_1730 (O_1730,N_14945,N_14872);
nand UO_1731 (O_1731,N_14896,N_14982);
and UO_1732 (O_1732,N_14876,N_14911);
xor UO_1733 (O_1733,N_14943,N_14881);
xor UO_1734 (O_1734,N_14852,N_14950);
or UO_1735 (O_1735,N_14906,N_14907);
nand UO_1736 (O_1736,N_14992,N_14916);
and UO_1737 (O_1737,N_14948,N_14901);
nor UO_1738 (O_1738,N_14988,N_14869);
and UO_1739 (O_1739,N_14932,N_14953);
or UO_1740 (O_1740,N_14922,N_14893);
xor UO_1741 (O_1741,N_14950,N_14995);
nor UO_1742 (O_1742,N_14894,N_14893);
and UO_1743 (O_1743,N_14964,N_14900);
nand UO_1744 (O_1744,N_14983,N_14984);
xor UO_1745 (O_1745,N_14916,N_14851);
or UO_1746 (O_1746,N_14982,N_14970);
or UO_1747 (O_1747,N_14895,N_14974);
xnor UO_1748 (O_1748,N_14894,N_14878);
nand UO_1749 (O_1749,N_14984,N_14887);
nor UO_1750 (O_1750,N_14880,N_14863);
xor UO_1751 (O_1751,N_14982,N_14898);
or UO_1752 (O_1752,N_14992,N_14947);
xnor UO_1753 (O_1753,N_14936,N_14937);
nand UO_1754 (O_1754,N_14947,N_14964);
nor UO_1755 (O_1755,N_14958,N_14938);
nor UO_1756 (O_1756,N_14888,N_14938);
nand UO_1757 (O_1757,N_14900,N_14864);
or UO_1758 (O_1758,N_14903,N_14961);
or UO_1759 (O_1759,N_14998,N_14879);
or UO_1760 (O_1760,N_14863,N_14981);
nor UO_1761 (O_1761,N_14894,N_14915);
or UO_1762 (O_1762,N_14947,N_14990);
or UO_1763 (O_1763,N_14942,N_14982);
or UO_1764 (O_1764,N_14882,N_14953);
nand UO_1765 (O_1765,N_14996,N_14992);
and UO_1766 (O_1766,N_14901,N_14909);
xor UO_1767 (O_1767,N_14988,N_14976);
nand UO_1768 (O_1768,N_14975,N_14929);
or UO_1769 (O_1769,N_14985,N_14917);
nand UO_1770 (O_1770,N_14875,N_14969);
or UO_1771 (O_1771,N_14896,N_14992);
and UO_1772 (O_1772,N_14865,N_14877);
or UO_1773 (O_1773,N_14897,N_14865);
and UO_1774 (O_1774,N_14915,N_14880);
nor UO_1775 (O_1775,N_14878,N_14865);
nor UO_1776 (O_1776,N_14971,N_14891);
nor UO_1777 (O_1777,N_14945,N_14900);
nor UO_1778 (O_1778,N_14865,N_14912);
nor UO_1779 (O_1779,N_14997,N_14879);
nand UO_1780 (O_1780,N_14906,N_14932);
nor UO_1781 (O_1781,N_14937,N_14970);
nor UO_1782 (O_1782,N_14889,N_14921);
xnor UO_1783 (O_1783,N_14893,N_14953);
xnor UO_1784 (O_1784,N_14858,N_14873);
nand UO_1785 (O_1785,N_14941,N_14937);
and UO_1786 (O_1786,N_14972,N_14985);
and UO_1787 (O_1787,N_14942,N_14888);
nor UO_1788 (O_1788,N_14865,N_14982);
nand UO_1789 (O_1789,N_14961,N_14915);
nor UO_1790 (O_1790,N_14908,N_14982);
or UO_1791 (O_1791,N_14976,N_14869);
or UO_1792 (O_1792,N_14864,N_14974);
nand UO_1793 (O_1793,N_14859,N_14877);
and UO_1794 (O_1794,N_14888,N_14944);
and UO_1795 (O_1795,N_14853,N_14870);
nor UO_1796 (O_1796,N_14907,N_14937);
or UO_1797 (O_1797,N_14879,N_14870);
xnor UO_1798 (O_1798,N_14887,N_14890);
xnor UO_1799 (O_1799,N_14929,N_14921);
xor UO_1800 (O_1800,N_14918,N_14997);
nand UO_1801 (O_1801,N_14899,N_14920);
nand UO_1802 (O_1802,N_14858,N_14968);
nand UO_1803 (O_1803,N_14948,N_14975);
nand UO_1804 (O_1804,N_14995,N_14985);
and UO_1805 (O_1805,N_14909,N_14999);
or UO_1806 (O_1806,N_14871,N_14863);
nor UO_1807 (O_1807,N_14882,N_14976);
nand UO_1808 (O_1808,N_14919,N_14873);
xnor UO_1809 (O_1809,N_14884,N_14895);
xor UO_1810 (O_1810,N_14865,N_14918);
and UO_1811 (O_1811,N_14850,N_14984);
and UO_1812 (O_1812,N_14962,N_14879);
or UO_1813 (O_1813,N_14915,N_14975);
xor UO_1814 (O_1814,N_14991,N_14916);
nand UO_1815 (O_1815,N_14930,N_14942);
nand UO_1816 (O_1816,N_14919,N_14973);
or UO_1817 (O_1817,N_14871,N_14886);
xnor UO_1818 (O_1818,N_14995,N_14959);
and UO_1819 (O_1819,N_14990,N_14900);
or UO_1820 (O_1820,N_14995,N_14888);
nor UO_1821 (O_1821,N_14970,N_14938);
and UO_1822 (O_1822,N_14895,N_14911);
or UO_1823 (O_1823,N_14902,N_14973);
or UO_1824 (O_1824,N_14860,N_14919);
nand UO_1825 (O_1825,N_14909,N_14893);
or UO_1826 (O_1826,N_14923,N_14893);
nand UO_1827 (O_1827,N_14937,N_14996);
nor UO_1828 (O_1828,N_14893,N_14966);
or UO_1829 (O_1829,N_14985,N_14868);
and UO_1830 (O_1830,N_14870,N_14871);
and UO_1831 (O_1831,N_14879,N_14925);
or UO_1832 (O_1832,N_14946,N_14891);
nand UO_1833 (O_1833,N_14905,N_14948);
xor UO_1834 (O_1834,N_14978,N_14896);
and UO_1835 (O_1835,N_14937,N_14878);
or UO_1836 (O_1836,N_14921,N_14943);
and UO_1837 (O_1837,N_14896,N_14952);
or UO_1838 (O_1838,N_14959,N_14887);
or UO_1839 (O_1839,N_14971,N_14964);
xnor UO_1840 (O_1840,N_14981,N_14879);
xnor UO_1841 (O_1841,N_14887,N_14899);
nor UO_1842 (O_1842,N_14892,N_14909);
and UO_1843 (O_1843,N_14891,N_14955);
xnor UO_1844 (O_1844,N_14860,N_14953);
nor UO_1845 (O_1845,N_14963,N_14909);
nand UO_1846 (O_1846,N_14969,N_14851);
nor UO_1847 (O_1847,N_14953,N_14856);
nor UO_1848 (O_1848,N_14860,N_14941);
nand UO_1849 (O_1849,N_14875,N_14901);
and UO_1850 (O_1850,N_14950,N_14851);
and UO_1851 (O_1851,N_14869,N_14962);
nor UO_1852 (O_1852,N_14945,N_14920);
nor UO_1853 (O_1853,N_14964,N_14978);
nand UO_1854 (O_1854,N_14995,N_14941);
nand UO_1855 (O_1855,N_14960,N_14914);
nor UO_1856 (O_1856,N_14907,N_14965);
and UO_1857 (O_1857,N_14890,N_14999);
nand UO_1858 (O_1858,N_14906,N_14981);
nor UO_1859 (O_1859,N_14906,N_14872);
nand UO_1860 (O_1860,N_14952,N_14982);
xor UO_1861 (O_1861,N_14952,N_14910);
and UO_1862 (O_1862,N_14985,N_14967);
nand UO_1863 (O_1863,N_14853,N_14979);
xnor UO_1864 (O_1864,N_14888,N_14878);
or UO_1865 (O_1865,N_14852,N_14875);
nand UO_1866 (O_1866,N_14879,N_14899);
nand UO_1867 (O_1867,N_14999,N_14961);
xor UO_1868 (O_1868,N_14875,N_14883);
or UO_1869 (O_1869,N_14905,N_14886);
or UO_1870 (O_1870,N_14992,N_14929);
or UO_1871 (O_1871,N_14993,N_14915);
and UO_1872 (O_1872,N_14861,N_14874);
xor UO_1873 (O_1873,N_14921,N_14975);
nand UO_1874 (O_1874,N_14976,N_14850);
or UO_1875 (O_1875,N_14930,N_14977);
xnor UO_1876 (O_1876,N_14877,N_14958);
nand UO_1877 (O_1877,N_14929,N_14977);
nor UO_1878 (O_1878,N_14945,N_14886);
nand UO_1879 (O_1879,N_14922,N_14874);
nand UO_1880 (O_1880,N_14998,N_14868);
and UO_1881 (O_1881,N_14943,N_14998);
xor UO_1882 (O_1882,N_14989,N_14948);
xor UO_1883 (O_1883,N_14914,N_14878);
or UO_1884 (O_1884,N_14983,N_14857);
and UO_1885 (O_1885,N_14906,N_14929);
nand UO_1886 (O_1886,N_14957,N_14969);
xor UO_1887 (O_1887,N_14876,N_14863);
nand UO_1888 (O_1888,N_14937,N_14920);
nor UO_1889 (O_1889,N_14882,N_14998);
or UO_1890 (O_1890,N_14988,N_14999);
and UO_1891 (O_1891,N_14932,N_14937);
or UO_1892 (O_1892,N_14989,N_14981);
nor UO_1893 (O_1893,N_14892,N_14903);
and UO_1894 (O_1894,N_14985,N_14948);
xnor UO_1895 (O_1895,N_14977,N_14991);
xnor UO_1896 (O_1896,N_14859,N_14867);
nor UO_1897 (O_1897,N_14939,N_14901);
and UO_1898 (O_1898,N_14942,N_14901);
or UO_1899 (O_1899,N_14895,N_14984);
nor UO_1900 (O_1900,N_14871,N_14869);
or UO_1901 (O_1901,N_14876,N_14894);
nor UO_1902 (O_1902,N_14873,N_14935);
and UO_1903 (O_1903,N_14962,N_14865);
or UO_1904 (O_1904,N_14937,N_14968);
or UO_1905 (O_1905,N_14988,N_14939);
nor UO_1906 (O_1906,N_14919,N_14867);
or UO_1907 (O_1907,N_14962,N_14963);
and UO_1908 (O_1908,N_14881,N_14880);
nand UO_1909 (O_1909,N_14937,N_14995);
or UO_1910 (O_1910,N_14881,N_14956);
xnor UO_1911 (O_1911,N_14930,N_14965);
or UO_1912 (O_1912,N_14942,N_14997);
and UO_1913 (O_1913,N_14905,N_14927);
xor UO_1914 (O_1914,N_14947,N_14900);
xor UO_1915 (O_1915,N_14988,N_14885);
or UO_1916 (O_1916,N_14886,N_14948);
and UO_1917 (O_1917,N_14872,N_14970);
or UO_1918 (O_1918,N_14889,N_14900);
nand UO_1919 (O_1919,N_14922,N_14923);
nor UO_1920 (O_1920,N_14960,N_14940);
nand UO_1921 (O_1921,N_14938,N_14908);
xnor UO_1922 (O_1922,N_14995,N_14923);
nand UO_1923 (O_1923,N_14992,N_14963);
nor UO_1924 (O_1924,N_14978,N_14928);
nor UO_1925 (O_1925,N_14899,N_14867);
xnor UO_1926 (O_1926,N_14870,N_14997);
and UO_1927 (O_1927,N_14881,N_14853);
or UO_1928 (O_1928,N_14968,N_14870);
or UO_1929 (O_1929,N_14965,N_14898);
nand UO_1930 (O_1930,N_14939,N_14902);
nand UO_1931 (O_1931,N_14998,N_14981);
and UO_1932 (O_1932,N_14859,N_14919);
and UO_1933 (O_1933,N_14917,N_14885);
xor UO_1934 (O_1934,N_14914,N_14906);
and UO_1935 (O_1935,N_14887,N_14877);
nor UO_1936 (O_1936,N_14888,N_14885);
xnor UO_1937 (O_1937,N_14919,N_14929);
xnor UO_1938 (O_1938,N_14872,N_14879);
nand UO_1939 (O_1939,N_14893,N_14933);
xor UO_1940 (O_1940,N_14977,N_14857);
nand UO_1941 (O_1941,N_14874,N_14975);
or UO_1942 (O_1942,N_14966,N_14861);
xnor UO_1943 (O_1943,N_14921,N_14857);
and UO_1944 (O_1944,N_14978,N_14900);
or UO_1945 (O_1945,N_14886,N_14882);
nor UO_1946 (O_1946,N_14929,N_14954);
or UO_1947 (O_1947,N_14945,N_14941);
nor UO_1948 (O_1948,N_14941,N_14924);
nand UO_1949 (O_1949,N_14902,N_14912);
xnor UO_1950 (O_1950,N_14975,N_14973);
xor UO_1951 (O_1951,N_14999,N_14977);
or UO_1952 (O_1952,N_14869,N_14944);
and UO_1953 (O_1953,N_14872,N_14852);
nand UO_1954 (O_1954,N_14886,N_14874);
nor UO_1955 (O_1955,N_14908,N_14983);
xnor UO_1956 (O_1956,N_14965,N_14868);
and UO_1957 (O_1957,N_14978,N_14960);
nand UO_1958 (O_1958,N_14987,N_14994);
or UO_1959 (O_1959,N_14897,N_14888);
and UO_1960 (O_1960,N_14933,N_14925);
or UO_1961 (O_1961,N_14986,N_14966);
xor UO_1962 (O_1962,N_14916,N_14980);
nor UO_1963 (O_1963,N_14929,N_14950);
or UO_1964 (O_1964,N_14967,N_14889);
nand UO_1965 (O_1965,N_14982,N_14858);
or UO_1966 (O_1966,N_14957,N_14853);
nand UO_1967 (O_1967,N_14936,N_14964);
or UO_1968 (O_1968,N_14962,N_14886);
xor UO_1969 (O_1969,N_14943,N_14856);
nor UO_1970 (O_1970,N_14875,N_14866);
or UO_1971 (O_1971,N_14973,N_14974);
nand UO_1972 (O_1972,N_14977,N_14958);
nand UO_1973 (O_1973,N_14964,N_14882);
and UO_1974 (O_1974,N_14918,N_14925);
and UO_1975 (O_1975,N_14956,N_14986);
or UO_1976 (O_1976,N_14885,N_14852);
or UO_1977 (O_1977,N_14885,N_14864);
or UO_1978 (O_1978,N_14965,N_14876);
or UO_1979 (O_1979,N_14907,N_14868);
and UO_1980 (O_1980,N_14928,N_14906);
or UO_1981 (O_1981,N_14853,N_14915);
nand UO_1982 (O_1982,N_14913,N_14996);
nand UO_1983 (O_1983,N_14904,N_14878);
nand UO_1984 (O_1984,N_14994,N_14898);
xnor UO_1985 (O_1985,N_14874,N_14999);
or UO_1986 (O_1986,N_14913,N_14854);
nand UO_1987 (O_1987,N_14850,N_14858);
xnor UO_1988 (O_1988,N_14901,N_14973);
nand UO_1989 (O_1989,N_14936,N_14878);
xor UO_1990 (O_1990,N_14930,N_14951);
nor UO_1991 (O_1991,N_14934,N_14901);
xor UO_1992 (O_1992,N_14948,N_14931);
or UO_1993 (O_1993,N_14862,N_14939);
nand UO_1994 (O_1994,N_14947,N_14859);
and UO_1995 (O_1995,N_14988,N_14918);
nand UO_1996 (O_1996,N_14925,N_14909);
nor UO_1997 (O_1997,N_14973,N_14895);
xor UO_1998 (O_1998,N_14902,N_14895);
xnor UO_1999 (O_1999,N_14900,N_14948);
endmodule