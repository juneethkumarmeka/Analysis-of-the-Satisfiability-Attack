module basic_5000_50000_5000_25_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
nor U0 (N_0,In_2441,In_1213);
xnor U1 (N_1,In_2879,In_3578);
nand U2 (N_2,In_2596,In_3598);
and U3 (N_3,In_1004,In_706);
nor U4 (N_4,In_1198,In_3269);
and U5 (N_5,In_1534,In_4575);
xor U6 (N_6,In_1728,In_2936);
and U7 (N_7,In_3619,In_1005);
nand U8 (N_8,In_1066,In_673);
or U9 (N_9,In_594,In_1772);
and U10 (N_10,In_2857,In_2248);
xor U11 (N_11,In_875,In_2126);
xnor U12 (N_12,In_480,In_3155);
or U13 (N_13,In_1970,In_783);
nor U14 (N_14,In_2935,In_4828);
nor U15 (N_15,In_2310,In_3464);
xor U16 (N_16,In_3579,In_4767);
and U17 (N_17,In_4077,In_1294);
or U18 (N_18,In_386,In_3709);
and U19 (N_19,In_2353,In_4457);
nand U20 (N_20,In_4768,In_2780);
nor U21 (N_21,In_1469,In_3007);
nand U22 (N_22,In_3382,In_2470);
xnor U23 (N_23,In_1859,In_117);
nand U24 (N_24,In_1172,In_3170);
nand U25 (N_25,In_4059,In_1565);
xnor U26 (N_26,In_1450,In_3980);
nand U27 (N_27,In_205,In_1126);
xnor U28 (N_28,In_541,In_2038);
and U29 (N_29,In_3538,In_2608);
xnor U30 (N_30,In_2678,In_489);
and U31 (N_31,In_4431,In_3359);
nand U32 (N_32,In_2850,In_2401);
xnor U33 (N_33,In_1335,In_4124);
nor U34 (N_34,In_3761,In_3480);
nor U35 (N_35,In_4515,In_746);
nor U36 (N_36,In_2740,In_3953);
nor U37 (N_37,In_2796,In_3584);
nand U38 (N_38,In_3418,In_4119);
nor U39 (N_39,In_4405,In_3190);
or U40 (N_40,In_3985,In_2483);
or U41 (N_41,In_1611,In_1992);
or U42 (N_42,In_2399,In_1443);
and U43 (N_43,In_2753,In_3746);
nand U44 (N_44,In_3315,In_1844);
xnor U45 (N_45,In_4665,In_3930);
or U46 (N_46,In_4011,In_4133);
and U47 (N_47,In_3123,In_1514);
nor U48 (N_48,In_2992,In_3545);
xnor U49 (N_49,In_4425,In_2996);
nor U50 (N_50,In_4784,In_1941);
nor U51 (N_51,In_2061,In_2075);
and U52 (N_52,In_4158,In_2350);
or U53 (N_53,In_4862,In_343);
xnor U54 (N_54,In_140,In_990);
nand U55 (N_55,In_4534,In_935);
nand U56 (N_56,In_2620,In_4184);
nor U57 (N_57,In_845,In_3440);
nand U58 (N_58,In_2865,In_1017);
or U59 (N_59,In_1144,In_1679);
xnor U60 (N_60,In_1850,In_2094);
nand U61 (N_61,In_2934,In_3296);
and U62 (N_62,In_737,In_335);
and U63 (N_63,In_1081,In_4257);
and U64 (N_64,In_4233,In_2484);
nor U65 (N_65,In_1453,In_3271);
and U66 (N_66,In_995,In_330);
nand U67 (N_67,In_2116,In_499);
and U68 (N_68,In_4482,In_2821);
nand U69 (N_69,In_4305,In_2321);
nand U70 (N_70,In_3301,In_692);
and U71 (N_71,In_608,In_3943);
or U72 (N_72,In_3358,In_1794);
or U73 (N_73,In_2172,In_4170);
xor U74 (N_74,In_560,In_1908);
xnor U75 (N_75,In_462,In_4166);
nand U76 (N_76,In_525,In_4302);
nand U77 (N_77,In_2465,In_1252);
nand U78 (N_78,In_2500,In_2);
nand U79 (N_79,In_1865,In_3129);
and U80 (N_80,In_2725,In_4925);
or U81 (N_81,In_1929,In_2820);
nand U82 (N_82,In_1398,In_974);
nor U83 (N_83,In_1113,In_3207);
and U84 (N_84,In_422,In_3940);
xor U85 (N_85,In_2064,In_4404);
nand U86 (N_86,In_2341,In_3154);
or U87 (N_87,In_2463,In_899);
or U88 (N_88,In_4087,In_2811);
or U89 (N_89,In_3230,In_3176);
nor U90 (N_90,In_4114,In_4590);
and U91 (N_91,In_1059,In_4118);
nor U92 (N_92,In_2486,In_2614);
or U93 (N_93,In_4560,In_350);
and U94 (N_94,In_2563,In_1774);
xor U95 (N_95,In_1192,In_790);
xnor U96 (N_96,In_2933,In_3829);
or U97 (N_97,In_4086,In_644);
nor U98 (N_98,In_358,In_2592);
nand U99 (N_99,In_3945,In_2809);
nor U100 (N_100,In_23,In_4888);
nand U101 (N_101,In_3745,In_455);
and U102 (N_102,In_1558,In_471);
nand U103 (N_103,In_3215,In_2642);
nand U104 (N_104,In_3697,In_4081);
xnor U105 (N_105,In_2023,In_482);
or U106 (N_106,In_3703,In_320);
and U107 (N_107,In_333,In_2118);
nor U108 (N_108,In_1617,In_4442);
xor U109 (N_109,In_3887,In_2228);
nor U110 (N_110,In_3281,In_3466);
xnor U111 (N_111,In_4308,In_2425);
and U112 (N_112,In_2730,In_3219);
xor U113 (N_113,In_3775,In_4927);
xor U114 (N_114,In_3729,In_1938);
nand U115 (N_115,In_84,In_2193);
and U116 (N_116,In_4219,In_4702);
xor U117 (N_117,In_1564,In_865);
and U118 (N_118,In_1476,In_4602);
nand U119 (N_119,In_802,In_1354);
or U120 (N_120,In_4183,In_4407);
nand U121 (N_121,In_3222,In_4678);
and U122 (N_122,In_2829,In_3680);
and U123 (N_123,In_2445,In_774);
and U124 (N_124,In_4314,In_3058);
nor U125 (N_125,In_86,In_4584);
nor U126 (N_126,In_2319,In_3556);
or U127 (N_127,In_3467,In_3426);
or U128 (N_128,In_2294,In_689);
and U129 (N_129,In_1542,In_2994);
and U130 (N_130,In_1416,In_3288);
nand U131 (N_131,In_3510,In_33);
or U132 (N_132,In_4418,In_2410);
or U133 (N_133,In_3209,In_240);
and U134 (N_134,In_449,In_2254);
xor U135 (N_135,In_1286,In_714);
or U136 (N_136,In_2090,In_2703);
nand U137 (N_137,In_1226,In_1028);
nor U138 (N_138,In_2339,In_354);
and U139 (N_139,In_3356,In_1588);
or U140 (N_140,In_4452,In_2244);
nor U141 (N_141,In_3122,In_3486);
or U142 (N_142,In_4345,In_3485);
xor U143 (N_143,In_37,In_2259);
nand U144 (N_144,In_2717,In_3182);
and U145 (N_145,In_908,In_2688);
nor U146 (N_146,In_1595,In_2723);
nand U147 (N_147,In_634,In_1472);
xnor U148 (N_148,In_1869,In_1108);
and U149 (N_149,In_2766,In_4631);
and U150 (N_150,In_4089,In_4344);
or U151 (N_151,In_3623,In_1881);
nand U152 (N_152,In_2790,In_4099);
and U153 (N_153,In_940,In_1261);
nand U154 (N_154,In_463,In_2298);
nand U155 (N_155,In_3868,In_1082);
nand U156 (N_156,In_150,In_2777);
nand U157 (N_157,In_2649,In_1615);
nor U158 (N_158,In_3291,In_2531);
nor U159 (N_159,In_4877,In_139);
nand U160 (N_160,In_2057,In_256);
nand U161 (N_161,In_3751,In_667);
and U162 (N_162,In_3353,In_1106);
and U163 (N_163,In_688,In_586);
nand U164 (N_164,In_2546,In_1810);
nor U165 (N_165,In_1698,In_557);
and U166 (N_166,In_633,In_175);
nor U167 (N_167,In_4010,In_4103);
and U168 (N_168,In_3825,In_973);
nor U169 (N_169,In_4147,In_484);
xnor U170 (N_170,In_1667,In_2532);
nor U171 (N_171,In_3397,In_4068);
xnor U172 (N_172,In_4056,In_1227);
xnor U173 (N_173,In_4052,In_1146);
xnor U174 (N_174,In_4821,In_3173);
xnor U175 (N_175,In_3223,In_1829);
or U176 (N_176,In_2424,In_1509);
or U177 (N_177,In_1425,In_1207);
xor U178 (N_178,In_694,In_1918);
nor U179 (N_179,In_4138,In_303);
nor U180 (N_180,In_2887,In_1052);
or U181 (N_181,In_2403,In_475);
nor U182 (N_182,In_1971,In_3616);
nand U183 (N_183,In_2274,In_3691);
and U184 (N_184,In_2151,In_1840);
or U185 (N_185,In_4084,In_411);
xnor U186 (N_186,In_4774,In_3897);
xnor U187 (N_187,In_1018,In_2910);
or U188 (N_188,In_184,In_2683);
or U189 (N_189,In_1737,In_2616);
nand U190 (N_190,In_4146,In_2612);
or U191 (N_191,In_4260,In_2733);
nor U192 (N_192,In_1677,In_614);
and U193 (N_193,In_579,In_3422);
nor U194 (N_194,In_2660,In_3505);
or U195 (N_195,In_1399,In_4758);
and U196 (N_196,In_2835,In_1741);
nand U197 (N_197,In_51,In_2585);
nor U198 (N_198,In_4779,In_1526);
nand U199 (N_199,In_906,In_1742);
nand U200 (N_200,In_4307,In_3807);
nand U201 (N_201,In_4520,In_1733);
or U202 (N_202,In_533,In_2448);
and U203 (N_203,In_705,In_2109);
and U204 (N_204,In_2363,In_69);
and U205 (N_205,In_4243,In_4781);
or U206 (N_206,In_4453,In_38);
and U207 (N_207,In_1937,In_3677);
nor U208 (N_208,In_4972,In_524);
and U209 (N_209,In_4969,In_2591);
nand U210 (N_210,In_2647,In_1201);
nand U211 (N_211,In_724,In_977);
and U212 (N_212,In_3699,In_1795);
nand U213 (N_213,In_1071,In_4738);
and U214 (N_214,In_1999,In_843);
nand U215 (N_215,In_2903,In_1406);
xnor U216 (N_216,In_1051,In_690);
nor U217 (N_217,In_2843,In_3408);
or U218 (N_218,In_4159,In_1490);
nor U219 (N_219,In_2322,In_1298);
or U220 (N_220,In_1403,In_4864);
xor U221 (N_221,In_1641,In_1092);
or U222 (N_222,In_3076,In_4340);
and U223 (N_223,In_2267,In_4533);
xor U224 (N_224,In_1324,In_78);
or U225 (N_225,In_4990,In_3492);
and U226 (N_226,In_2309,In_1727);
nor U227 (N_227,In_2027,In_4065);
nor U228 (N_228,In_3006,In_1358);
nand U229 (N_229,In_1348,In_810);
and U230 (N_230,In_4494,In_3374);
nor U231 (N_231,In_2788,In_4517);
nor U232 (N_232,In_3206,In_1724);
nor U233 (N_233,In_3419,In_3925);
xor U234 (N_234,In_2105,In_4878);
and U235 (N_235,In_4695,In_4708);
nor U236 (N_236,In_71,In_4800);
nand U237 (N_237,In_3029,In_3149);
xor U238 (N_238,In_3895,In_2701);
nand U239 (N_239,In_3479,In_3621);
nor U240 (N_240,In_887,In_3270);
xnor U241 (N_241,In_962,In_1138);
and U242 (N_242,In_266,In_3325);
xor U243 (N_243,In_1921,In_3923);
nand U244 (N_244,In_4450,In_197);
nand U245 (N_245,In_4148,In_4471);
xnor U246 (N_246,In_4920,In_922);
xnor U247 (N_247,In_592,In_1701);
and U248 (N_248,In_3146,In_4540);
nand U249 (N_249,In_1904,In_466);
xnor U250 (N_250,In_1329,In_1410);
nor U251 (N_251,In_4569,In_4291);
and U252 (N_252,In_1699,In_4346);
and U253 (N_253,In_1321,In_3917);
or U254 (N_254,In_4456,In_1911);
xnor U255 (N_255,In_290,In_1731);
or U256 (N_256,In_294,In_3931);
nand U257 (N_257,In_1288,In_132);
or U258 (N_258,In_4055,In_4906);
or U259 (N_259,In_2762,In_1022);
and U260 (N_260,In_3008,In_3617);
and U261 (N_261,In_4994,In_1585);
xnor U262 (N_262,In_3713,In_632);
and U263 (N_263,In_4636,In_701);
or U264 (N_264,In_129,In_3988);
xnor U265 (N_265,In_1898,In_1205);
nand U266 (N_266,In_1356,In_1566);
nor U267 (N_267,In_2641,In_4810);
nand U268 (N_268,In_3760,In_3399);
nor U269 (N_269,In_4217,In_3679);
nand U270 (N_270,In_1740,In_1516);
or U271 (N_271,In_1748,In_1371);
and U272 (N_272,In_3000,In_2412);
xor U273 (N_273,In_2868,In_3794);
nand U274 (N_274,In_4332,In_4213);
and U275 (N_275,In_3112,In_3450);
and U276 (N_276,In_4140,In_555);
nor U277 (N_277,In_1408,In_1713);
nor U278 (N_278,In_4822,In_4619);
nor U279 (N_279,In_2742,In_1189);
and U280 (N_280,In_2986,In_451);
and U281 (N_281,In_3405,In_1002);
and U282 (N_282,In_2231,In_3971);
xor U283 (N_283,In_4171,In_2174);
xnor U284 (N_284,In_3629,In_2139);
or U285 (N_285,In_2051,In_1515);
or U286 (N_286,In_2256,In_4581);
and U287 (N_287,In_1541,In_1610);
nand U288 (N_288,In_2211,In_3625);
nand U289 (N_289,In_1493,In_3753);
xor U290 (N_290,In_3171,In_1843);
nor U291 (N_291,In_4403,In_2908);
or U292 (N_292,In_1427,In_369);
nand U293 (N_293,In_4777,In_3662);
nand U294 (N_294,In_1143,In_3932);
and U295 (N_295,In_1204,In_713);
nor U296 (N_296,In_4751,In_4033);
and U297 (N_297,In_1783,In_1121);
and U298 (N_298,In_2467,In_3782);
nand U299 (N_299,In_2691,In_519);
nand U300 (N_300,In_638,In_4478);
nand U301 (N_301,In_3915,In_3874);
nand U302 (N_302,In_649,In_862);
and U303 (N_303,In_2203,In_1662);
or U304 (N_304,In_1910,In_3871);
and U305 (N_305,In_4428,In_2362);
nand U306 (N_306,In_4977,In_2713);
or U307 (N_307,In_3615,In_1040);
and U308 (N_308,In_2529,In_3258);
xnor U309 (N_309,In_2876,In_170);
nand U310 (N_310,In_3261,In_1323);
or U311 (N_311,In_2805,In_119);
nand U312 (N_312,In_2242,In_4416);
and U313 (N_313,In_4893,In_2594);
or U314 (N_314,In_3049,In_3614);
nand U315 (N_315,In_2358,In_3157);
or U316 (N_316,In_3313,In_376);
nand U317 (N_317,In_133,In_1738);
nand U318 (N_318,In_2624,In_1954);
nor U319 (N_319,In_1796,In_3927);
and U320 (N_320,In_114,In_3557);
nor U321 (N_321,In_274,In_4904);
or U322 (N_322,In_1726,In_3642);
nor U323 (N_323,In_537,In_2750);
nor U324 (N_324,In_4873,In_4288);
or U325 (N_325,In_2106,In_1841);
or U326 (N_326,In_716,In_3855);
nor U327 (N_327,In_1777,In_2001);
nand U328 (N_328,In_2578,In_983);
or U329 (N_329,In_2758,In_3830);
or U330 (N_330,In_1790,In_4211);
or U331 (N_331,In_2571,In_2295);
or U332 (N_332,In_2466,In_1454);
xnor U333 (N_333,In_3150,In_2285);
nor U334 (N_334,In_63,In_4187);
xnor U335 (N_335,In_1225,In_3626);
nor U336 (N_336,In_3078,In_3220);
or U337 (N_337,In_4326,In_585);
nand U338 (N_338,In_1366,In_1957);
nor U339 (N_339,In_2235,In_1468);
and U340 (N_340,In_2002,In_2674);
nor U341 (N_341,In_3067,In_3478);
xor U342 (N_342,In_4891,In_4866);
nand U343 (N_343,In_2157,In_260);
nand U344 (N_344,In_459,In_3824);
or U345 (N_345,In_3267,In_1161);
or U346 (N_346,In_826,In_642);
and U347 (N_347,In_4976,In_2916);
or U348 (N_348,In_4030,In_393);
and U349 (N_349,In_3548,In_611);
nand U350 (N_350,In_1220,In_3816);
nor U351 (N_351,In_4347,In_3959);
and U352 (N_352,In_4577,In_1355);
xnor U353 (N_353,In_4338,In_933);
xor U354 (N_354,In_1787,In_220);
or U355 (N_355,In_4667,In_4120);
or U356 (N_356,In_931,In_1228);
or U357 (N_357,In_2552,In_3095);
nand U358 (N_358,In_1378,In_3221);
and U359 (N_359,In_4348,In_2283);
or U360 (N_360,In_2085,In_4664);
xor U361 (N_361,In_299,In_2468);
and U362 (N_362,In_4773,In_1466);
nor U363 (N_363,In_1925,In_565);
nand U364 (N_364,In_4782,In_2613);
nor U365 (N_365,In_2899,In_1237);
or U366 (N_366,In_4039,In_597);
or U367 (N_367,In_3946,In_3670);
nand U368 (N_368,In_1634,In_1169);
xnor U369 (N_369,In_13,In_222);
nor U370 (N_370,In_2995,In_2034);
xnor U371 (N_371,In_1424,In_3572);
and U372 (N_372,In_1873,In_1722);
and U373 (N_373,In_3728,In_2855);
and U374 (N_374,In_4174,In_4201);
nand U375 (N_375,In_3127,In_1345);
and U376 (N_376,In_3186,In_4251);
nand U377 (N_377,In_2003,In_1353);
or U378 (N_378,In_3063,In_660);
nor U379 (N_379,In_1602,In_3605);
nand U380 (N_380,In_554,In_2830);
nand U381 (N_381,In_4907,In_179);
xnor U382 (N_382,In_3739,In_1589);
xnor U383 (N_383,In_4943,In_203);
nor U384 (N_384,In_4879,In_2891);
and U385 (N_385,In_651,In_3383);
nand U386 (N_386,In_637,In_4648);
nand U387 (N_387,In_2581,In_4377);
xnor U388 (N_388,In_1883,In_3278);
xnor U389 (N_389,In_2333,In_1234);
nor U390 (N_390,In_794,In_656);
nand U391 (N_391,In_2771,In_4769);
or U392 (N_392,In_4916,In_2988);
and U393 (N_393,In_4690,In_1623);
nand U394 (N_394,In_1506,In_4543);
xor U395 (N_395,In_1902,In_4511);
nand U396 (N_396,In_1671,In_1461);
nor U397 (N_397,In_3428,In_226);
xor U398 (N_398,In_876,In_4454);
nor U399 (N_399,In_3237,In_99);
xor U400 (N_400,In_2366,In_1621);
or U401 (N_401,In_894,In_1474);
or U402 (N_402,In_4815,In_2223);
or U403 (N_403,In_262,In_994);
and U404 (N_404,In_1318,In_148);
or U405 (N_405,In_381,In_3570);
nor U406 (N_406,In_733,In_259);
and U407 (N_407,In_104,In_818);
and U408 (N_408,In_2033,In_4018);
or U409 (N_409,In_4381,In_3783);
or U410 (N_410,In_267,In_2927);
xnor U411 (N_411,In_822,In_2694);
and U412 (N_412,In_4670,In_4944);
xnor U413 (N_413,In_483,In_3178);
nand U414 (N_414,In_853,In_485);
nor U415 (N_415,In_4775,In_1072);
nand U416 (N_416,In_3573,In_1899);
nand U417 (N_417,In_4419,In_1124);
nor U418 (N_418,In_4937,In_2956);
nor U419 (N_419,In_2802,In_2566);
nor U420 (N_420,In_4410,In_1160);
nor U421 (N_421,In_1044,In_2914);
nand U422 (N_422,In_1299,In_2328);
nor U423 (N_423,In_4459,In_1782);
nand U424 (N_424,In_1835,In_4355);
or U425 (N_425,In_171,In_2112);
xor U426 (N_426,In_1652,In_2213);
and U427 (N_427,In_275,In_1930);
nand U428 (N_428,In_2508,In_2837);
nand U429 (N_429,In_1823,In_1009);
or U430 (N_430,In_1939,In_112);
nor U431 (N_431,In_4003,In_1441);
or U432 (N_432,In_3410,In_4268);
and U433 (N_433,In_2173,In_4021);
and U434 (N_434,In_3660,In_2711);
and U435 (N_435,In_2707,In_2696);
xor U436 (N_436,In_2798,In_2385);
xnor U437 (N_437,In_4802,In_3159);
nor U438 (N_438,In_893,In_903);
or U439 (N_439,In_3903,In_4046);
xor U440 (N_440,In_4150,In_936);
nor U441 (N_441,In_3803,In_1090);
nand U442 (N_442,In_6,In_4441);
xnor U443 (N_443,In_4761,In_2393);
nand U444 (N_444,In_3866,In_2010);
or U445 (N_445,In_3569,In_3175);
nor U446 (N_446,In_2858,In_2286);
xnor U447 (N_447,In_2562,In_3299);
or U448 (N_448,In_825,In_577);
xnor U449 (N_449,In_3052,In_1940);
nand U450 (N_450,In_2272,In_4541);
or U451 (N_451,In_2110,In_1027);
nor U452 (N_452,In_373,In_2953);
nor U453 (N_453,In_670,In_2431);
and U454 (N_454,In_3878,In_1830);
nor U455 (N_455,In_4278,In_3813);
and U456 (N_456,In_1401,In_2453);
nor U457 (N_457,In_677,In_4144);
and U458 (N_458,In_2923,In_174);
or U459 (N_459,In_2517,In_3036);
and U460 (N_460,In_1451,In_3810);
xor U461 (N_461,In_3968,In_1179);
xor U462 (N_462,In_2030,In_4253);
xnor U463 (N_463,In_1586,In_1364);
and U464 (N_464,In_3608,In_430);
nand U465 (N_465,In_3503,In_4638);
or U466 (N_466,In_4409,In_4884);
and U467 (N_467,In_1665,In_2028);
xor U468 (N_468,In_772,In_4991);
and U469 (N_469,In_3180,In_137);
nor U470 (N_470,In_3520,In_2681);
or U471 (N_471,In_470,In_1868);
xnor U472 (N_472,In_160,In_1637);
or U473 (N_473,In_1297,In_4841);
xnor U474 (N_474,In_1070,In_4279);
xnor U475 (N_475,In_3030,In_199);
nor U476 (N_476,In_719,In_4126);
nor U477 (N_477,In_4681,In_1993);
nor U478 (N_478,In_3708,In_3043);
nand U479 (N_479,In_4490,In_4811);
nor U480 (N_480,In_3516,In_2651);
and U481 (N_481,In_2888,In_1087);
xnor U482 (N_482,In_797,In_1180);
xnor U483 (N_483,In_309,In_2018);
nor U484 (N_484,In_951,In_4128);
nand U485 (N_485,In_4965,In_4548);
nand U486 (N_486,In_254,In_1907);
nand U487 (N_487,In_3607,In_3742);
nand U488 (N_488,In_3453,In_4992);
nand U489 (N_489,In_244,In_4125);
nor U490 (N_490,In_130,In_1923);
nand U491 (N_491,In_4707,In_257);
nand U492 (N_492,In_4161,In_3610);
and U493 (N_493,In_1627,In_2640);
nor U494 (N_494,In_2652,In_4042);
nand U495 (N_495,In_4235,In_4005);
nand U496 (N_496,In_1360,In_2476);
and U497 (N_497,In_2053,In_2506);
nand U498 (N_498,In_1936,In_1870);
nor U499 (N_499,In_113,In_1337);
nor U500 (N_500,In_4890,In_1591);
or U501 (N_501,In_1111,In_2741);
xnor U502 (N_502,In_4280,In_3500);
xor U503 (N_503,In_949,In_1013);
nor U504 (N_504,In_159,In_364);
and U505 (N_505,In_4857,In_4216);
and U506 (N_506,In_4871,In_3748);
nand U507 (N_507,In_2735,In_643);
xor U508 (N_508,In_1876,In_852);
or U509 (N_509,In_4061,In_814);
xnor U510 (N_510,In_2397,In_1449);
and U511 (N_511,In_4637,In_1367);
and U512 (N_512,In_890,In_543);
or U513 (N_513,In_2756,In_2502);
nor U514 (N_514,In_1290,In_2806);
nand U515 (N_515,In_3304,In_4635);
xor U516 (N_516,In_4712,In_2019);
nand U517 (N_517,In_1388,In_2697);
or U518 (N_518,In_4596,In_307);
xnor U519 (N_519,In_2414,In_1685);
nor U520 (N_520,In_762,In_891);
or U521 (N_521,In_2772,In_2443);
nor U522 (N_522,In_4941,In_4266);
xnor U523 (N_523,In_1847,In_1395);
nand U524 (N_524,In_1953,In_4350);
nor U525 (N_525,In_41,In_3494);
nor U526 (N_526,In_3777,In_3239);
xor U527 (N_527,In_1393,In_4919);
nand U528 (N_528,In_3592,In_1177);
and U529 (N_529,In_1706,In_4356);
nand U530 (N_530,In_1926,In_3717);
xor U531 (N_531,In_3024,In_1922);
nor U532 (N_532,In_1001,In_975);
nor U533 (N_533,In_166,In_2783);
xor U534 (N_534,In_1826,In_448);
xor U535 (N_535,In_2559,In_56);
xor U536 (N_536,In_4488,In_4597);
nand U537 (N_537,In_1164,In_3477);
and U538 (N_538,In_4876,In_919);
nand U539 (N_539,In_1268,In_1561);
xnor U540 (N_540,In_3645,In_4655);
and U541 (N_541,In_3297,In_732);
nor U542 (N_542,In_477,In_3553);
nand U543 (N_543,In_3311,In_3880);
nand U544 (N_544,In_1979,In_75);
and U545 (N_545,In_1046,In_200);
nor U546 (N_546,In_4835,In_2207);
xor U547 (N_547,In_102,In_883);
or U548 (N_548,In_3733,In_4143);
nor U549 (N_549,In_2398,In_2885);
xnor U550 (N_550,In_4675,In_626);
nand U551 (N_551,In_4444,In_1149);
nand U552 (N_552,In_4265,In_2898);
or U553 (N_553,In_4093,In_2795);
nand U554 (N_554,In_650,In_3633);
or U555 (N_555,In_787,In_2654);
nor U556 (N_556,In_2070,In_151);
xnor U557 (N_557,In_4491,In_3329);
nor U558 (N_558,In_4275,In_1470);
xnor U559 (N_559,In_2083,In_2519);
xor U560 (N_560,In_2525,In_2631);
nand U561 (N_561,In_408,In_4557);
or U562 (N_562,In_4962,In_2185);
or U563 (N_563,In_3200,In_134);
nor U564 (N_564,In_3151,In_2303);
nand U565 (N_565,In_4749,In_4391);
nor U566 (N_566,In_1533,In_3427);
xnor U567 (N_567,In_3844,In_2017);
nand U568 (N_568,In_628,In_4179);
or U569 (N_569,In_3487,In_2793);
or U570 (N_570,In_2728,In_835);
nor U571 (N_571,In_3391,In_1062);
or U572 (N_572,In_640,In_4020);
or U573 (N_573,In_310,In_4840);
and U574 (N_574,In_3574,In_1504);
xnor U575 (N_575,In_1314,In_3282);
xnor U576 (N_576,In_4911,In_3669);
nand U577 (N_577,In_2524,In_1934);
or U578 (N_578,In_788,In_1411);
nor U579 (N_579,In_341,In_2634);
xor U580 (N_580,In_1556,In_1640);
nand U581 (N_581,In_1102,In_3105);
nor U582 (N_582,In_4863,In_1116);
nor U583 (N_583,In_3766,In_87);
or U584 (N_584,In_601,In_3684);
and U585 (N_585,In_552,In_4809);
nand U586 (N_586,In_3812,In_1088);
nand U587 (N_587,In_3661,In_255);
nand U588 (N_588,In_2883,In_773);
nand U589 (N_589,In_1858,In_2247);
xor U590 (N_590,In_2981,In_2602);
nand U591 (N_591,In_42,In_4113);
nand U592 (N_592,In_1730,In_4561);
nand U593 (N_593,In_4395,In_2812);
xor U594 (N_594,In_2666,In_1293);
nand U595 (N_595,In_3370,In_2794);
and U596 (N_596,In_1346,In_1444);
nor U597 (N_597,In_2396,In_505);
xor U598 (N_598,In_3184,In_3400);
nor U599 (N_599,In_4853,In_340);
nand U600 (N_600,In_1467,In_1745);
nor U601 (N_601,In_204,In_344);
or U602 (N_602,In_3131,In_4339);
nor U603 (N_603,In_1675,In_4360);
and U604 (N_604,In_4653,In_1744);
nor U605 (N_605,In_4228,In_1935);
or U606 (N_606,In_2456,In_4843);
nor U607 (N_607,In_177,In_3263);
and U608 (N_608,In_2915,In_2201);
xor U609 (N_609,In_4477,In_2861);
and U610 (N_610,In_3318,In_1682);
nand U611 (N_611,In_4336,In_4083);
nand U612 (N_612,In_4793,In_2621);
xor U613 (N_613,In_1544,In_2132);
nand U614 (N_614,In_2380,In_1069);
and U615 (N_615,In_1729,In_4050);
xnor U616 (N_616,In_3757,In_311);
nand U617 (N_617,In_4468,In_3640);
or U618 (N_618,In_3065,In_3639);
nand U619 (N_619,In_2357,In_741);
or U620 (N_620,In_2852,In_4510);
and U621 (N_621,In_3901,In_4309);
nand U622 (N_622,In_2224,In_3481);
nand U623 (N_623,In_2949,In_1344);
or U624 (N_624,In_4466,In_3577);
and U625 (N_625,In_2312,In_1141);
nor U626 (N_626,In_196,In_391);
nor U627 (N_627,In_2948,In_968);
nand U628 (N_628,In_4714,In_2549);
or U629 (N_629,In_699,In_3474);
or U630 (N_630,In_1194,In_4718);
and U631 (N_631,In_3412,In_904);
and U632 (N_632,In_4639,In_3750);
and U633 (N_633,In_2273,In_2044);
and U634 (N_634,In_2968,In_1990);
or U635 (N_635,In_2269,In_2297);
nor U636 (N_636,In_2554,In_3309);
nor U637 (N_637,In_4095,In_1576);
nand U638 (N_638,In_3064,In_17);
nor U639 (N_639,In_1158,In_4141);
nor U640 (N_640,In_1739,In_4594);
or U641 (N_641,In_1686,In_1955);
nor U642 (N_642,In_3118,In_3688);
xnor U643 (N_643,In_4763,In_10);
nor U644 (N_644,In_319,In_785);
or U645 (N_645,In_1433,In_3280);
nor U646 (N_646,In_1262,In_3054);
nand U647 (N_647,In_3187,In_3276);
or U648 (N_648,In_2206,In_4);
xnor U649 (N_649,In_971,In_916);
xor U650 (N_650,In_3089,In_1828);
and U651 (N_651,In_2261,In_2428);
and U652 (N_652,In_2799,In_1218);
nand U653 (N_653,In_2589,In_4191);
or U654 (N_654,In_4063,In_2845);
nand U655 (N_655,In_1191,In_1538);
nor U656 (N_656,In_2667,In_3037);
or U657 (N_657,In_1780,In_1901);
and U658 (N_658,In_43,In_4886);
and U659 (N_659,In_1193,In_3051);
nand U660 (N_660,In_1249,In_4736);
xnor U661 (N_661,In_1241,In_3462);
nor U662 (N_662,In_2482,In_3066);
nand U663 (N_663,In_3843,In_2644);
or U664 (N_664,In_2527,In_2073);
xnor U665 (N_665,In_2071,In_4803);
or U666 (N_666,In_4757,In_4207);
nor U667 (N_667,In_245,In_510);
and U668 (N_668,In_4856,In_1505);
or U669 (N_669,In_930,In_915);
and U670 (N_670,In_2225,In_2598);
xor U671 (N_671,In_3380,In_1603);
and U672 (N_672,In_1182,In_999);
nand U673 (N_673,In_3424,In_4283);
or U674 (N_674,In_563,In_1435);
and U675 (N_675,In_115,In_2170);
or U676 (N_676,In_1402,In_4255);
and U677 (N_677,In_4529,In_4669);
and U678 (N_678,In_3292,In_178);
and U679 (N_679,In_4633,In_2127);
or U680 (N_680,In_1700,In_2501);
and U681 (N_681,In_1785,In_1405);
nor U682 (N_682,In_2340,In_1599);
and U683 (N_683,In_4953,In_4624);
xnor U684 (N_684,In_4341,In_1387);
and U685 (N_685,In_3741,In_4498);
or U686 (N_686,In_3197,In_2423);
xnor U687 (N_687,In_4693,In_2943);
xor U688 (N_688,In_2599,In_1372);
xnor U689 (N_689,In_3958,In_2077);
nand U690 (N_690,In_3814,In_3249);
xor U691 (N_691,In_4570,In_3941);
and U692 (N_692,In_1539,In_370);
and U693 (N_693,In_3266,In_1862);
nor U694 (N_694,In_4683,In_218);
xor U695 (N_695,In_4945,In_3804);
nor U696 (N_696,In_3026,In_339);
and U697 (N_697,In_1915,In_4242);
and U698 (N_698,In_3911,In_4220);
nor U699 (N_699,In_3109,In_3056);
xor U700 (N_700,In_1055,In_4957);
nand U701 (N_701,In_4723,In_2146);
or U702 (N_702,In_3165,In_964);
and U703 (N_703,In_4555,In_2277);
or U704 (N_704,In_3681,In_3444);
or U705 (N_705,In_3618,In_316);
xor U706 (N_706,In_4698,In_3929);
nand U707 (N_707,In_2618,In_3140);
nand U708 (N_708,In_4445,In_1996);
or U709 (N_709,In_3341,In_3369);
or U710 (N_710,In_520,In_1646);
nor U711 (N_711,In_145,In_4318);
nor U712 (N_712,In_4578,In_1278);
xor U713 (N_713,In_4009,In_3550);
and U714 (N_714,In_3513,In_2952);
or U715 (N_715,In_1963,In_347);
or U716 (N_716,In_2645,In_2457);
nor U717 (N_717,In_3693,In_776);
nand U718 (N_718,In_454,In_2655);
or U719 (N_719,In_2435,In_495);
nand U720 (N_720,In_827,In_2894);
xor U721 (N_721,In_2816,In_1555);
nand U722 (N_722,In_4954,In_21);
nor U723 (N_723,In_1383,In_4657);
nor U724 (N_724,In_3307,In_1560);
xnor U725 (N_725,In_1651,In_2205);
and U726 (N_726,In_1311,In_135);
nand U727 (N_727,In_3954,In_4163);
and U728 (N_728,In_2054,In_81);
or U729 (N_729,In_1380,In_4506);
and U730 (N_730,In_2048,In_2058);
nand U731 (N_731,In_1648,In_2708);
nand U732 (N_732,In_2005,In_18);
nor U733 (N_733,In_2301,In_2542);
xor U734 (N_734,In_2304,In_3865);
xor U735 (N_735,In_3124,In_1607);
nand U736 (N_736,In_3714,In_1471);
xor U737 (N_737,In_286,In_3549);
or U738 (N_738,In_1392,In_3277);
nand U739 (N_739,In_1168,In_850);
and U740 (N_740,In_97,In_8);
xor U741 (N_741,In_2689,In_336);
and U742 (N_742,In_2997,In_49);
nand U743 (N_743,In_2810,In_1498);
xor U744 (N_744,In_2359,In_2176);
or U745 (N_745,In_4122,In_3108);
xnor U746 (N_746,In_1550,In_778);
xnor U747 (N_747,In_1385,In_3031);
or U748 (N_748,In_4127,In_668);
or U749 (N_749,In_4917,In_2241);
xor U750 (N_750,In_952,In_1570);
and U751 (N_751,In_3965,In_4393);
or U752 (N_752,In_3342,In_763);
xor U753 (N_753,In_4614,In_122);
xor U754 (N_754,In_2253,In_3702);
nor U755 (N_755,In_4984,In_4922);
xor U756 (N_756,In_1230,In_932);
or U757 (N_757,In_395,In_3797);
nor U758 (N_758,In_3704,In_1912);
and U759 (N_759,In_2446,In_549);
or U760 (N_760,In_3885,In_1824);
or U761 (N_761,In_2337,In_780);
nor U762 (N_762,In_1130,In_4493);
and U763 (N_763,In_4023,In_4722);
xor U764 (N_764,In_4959,In_3231);
nand U765 (N_765,In_2325,In_4097);
and U766 (N_766,In_3995,In_2978);
or U767 (N_767,In_421,In_3653);
nor U768 (N_768,In_2405,In_128);
nor U769 (N_769,In_3183,In_4323);
nand U770 (N_770,In_4100,In_4313);
and U771 (N_771,In_1084,In_2495);
nor U772 (N_772,In_4699,In_2983);
nor U773 (N_773,In_3907,In_3033);
nand U774 (N_774,In_4250,In_3599);
or U775 (N_775,In_764,In_3489);
xnor U776 (N_776,In_4396,In_3202);
and U777 (N_777,In_120,In_2014);
nor U778 (N_778,In_101,In_305);
nor U779 (N_779,In_4503,In_1502);
xnor U780 (N_780,In_3846,In_4717);
xor U781 (N_781,In_1962,In_4967);
or U782 (N_782,In_4607,In_4966);
xor U783 (N_783,In_3859,In_45);
or U784 (N_784,In_4236,In_2168);
xor U785 (N_785,In_1678,In_542);
and U786 (N_786,In_4677,In_1303);
or U787 (N_787,In_2814,In_4816);
or U788 (N_788,In_337,In_3451);
nor U789 (N_789,In_717,In_691);
and U790 (N_790,In_4480,In_3659);
xnor U791 (N_791,In_2664,In_1551);
and U792 (N_792,In_3762,In_695);
nor U793 (N_793,In_1797,In_1812);
xnor U794 (N_794,In_2290,In_4458);
or U795 (N_795,In_4933,In_961);
or U796 (N_796,In_4276,In_216);
xor U797 (N_797,In_2976,In_1254);
nor U798 (N_798,In_984,In_530);
nor U799 (N_799,In_239,In_2436);
xnor U800 (N_800,In_3769,In_2893);
xnor U801 (N_801,In_389,In_474);
and U802 (N_802,In_4812,In_3994);
and U803 (N_803,In_1503,In_1222);
nand U804 (N_804,In_3674,In_1209);
nand U805 (N_805,In_4153,In_619);
or U806 (N_806,In_289,In_3432);
or U807 (N_807,In_4006,In_3456);
nor U808 (N_808,In_4131,In_1775);
nand U809 (N_809,In_4975,In_4599);
and U810 (N_810,In_2411,In_90);
or U811 (N_811,In_2999,In_2009);
xnor U812 (N_812,In_3652,In_1831);
xor U813 (N_813,In_3083,In_1914);
or U814 (N_814,In_3863,In_967);
nor U815 (N_815,In_2512,In_901);
nand U816 (N_816,In_3966,In_2437);
nand U817 (N_817,In_1236,In_64);
xor U818 (N_818,In_4043,In_2461);
nor U819 (N_819,In_3395,In_2029);
and U820 (N_820,In_2661,In_89);
or U821 (N_821,In_4497,In_3275);
xnor U822 (N_822,In_2769,In_1527);
xor U823 (N_823,In_509,In_4229);
and U824 (N_824,In_2068,In_3285);
nor U825 (N_825,In_600,In_3678);
nand U826 (N_826,In_683,In_365);
or U827 (N_827,In_2746,In_1577);
or U828 (N_828,In_1167,In_2853);
or U829 (N_829,In_2869,In_2768);
and U830 (N_830,In_3663,In_3381);
and U831 (N_831,In_4603,In_959);
nand U832 (N_832,In_2190,In_3834);
nor U833 (N_833,In_4105,In_4516);
nor U834 (N_834,In_2275,In_209);
xor U835 (N_835,In_1612,In_3028);
nand U836 (N_836,In_2550,In_1846);
and U837 (N_837,In_4580,In_3817);
xnor U838 (N_838,In_3773,In_3594);
nand U839 (N_839,In_2958,In_1043);
and U840 (N_840,In_1887,In_285);
and U841 (N_841,In_2918,In_308);
xor U842 (N_842,In_2402,In_740);
nand U843 (N_843,In_1536,In_4026);
nor U844 (N_844,In_4382,In_2890);
nand U845 (N_845,In_4195,In_2037);
and U846 (N_846,In_1767,In_680);
or U847 (N_847,In_2841,In_2963);
xnor U848 (N_848,In_54,In_2638);
or U849 (N_849,In_74,In_2375);
and U850 (N_850,In_1483,In_4230);
and U851 (N_851,In_4875,In_3820);
or U852 (N_852,In_546,In_194);
xor U853 (N_853,In_435,In_438);
nor U854 (N_854,In_4439,In_2230);
and U855 (N_855,In_803,In_2265);
nor U856 (N_856,In_327,In_3910);
or U857 (N_857,In_4049,In_1208);
nand U858 (N_858,In_4776,In_937);
nor U859 (N_859,In_206,In_2839);
and U860 (N_860,In_2429,In_210);
xnor U861 (N_861,In_3134,In_896);
nand U862 (N_862,In_2015,In_3191);
or U863 (N_863,In_1906,In_1752);
nand U864 (N_864,In_4412,In_2464);
nand U865 (N_865,In_970,In_2234);
and U866 (N_866,In_2973,In_4744);
nand U867 (N_867,In_4421,In_1076);
and U868 (N_868,In_3727,In_131);
or U869 (N_869,In_1557,In_2141);
xnor U870 (N_870,In_1749,In_464);
or U871 (N_871,In_3274,In_1263);
or U872 (N_872,In_2580,In_2663);
xor U873 (N_873,In_2520,In_1872);
xor U874 (N_874,In_4325,In_2849);
or U875 (N_875,In_2942,In_2210);
nor U876 (N_876,In_3604,In_1488);
and U877 (N_877,In_4267,In_4455);
or U878 (N_878,In_3790,In_2434);
xor U879 (N_879,In_528,In_1458);
nand U880 (N_880,In_3446,In_4352);
or U881 (N_881,In_2928,In_2095);
nand U882 (N_882,In_105,In_832);
xor U883 (N_883,In_3268,In_198);
xor U884 (N_884,In_2523,In_2021);
nor U885 (N_885,In_2629,In_2447);
and U886 (N_886,In_3864,In_383);
nor U887 (N_887,In_4551,In_242);
nor U888 (N_888,In_4824,In_4997);
or U889 (N_889,In_2622,In_3540);
and U890 (N_890,In_1991,In_1457);
nand U891 (N_891,In_775,In_2209);
nor U892 (N_892,In_278,In_2833);
nor U893 (N_893,In_1211,In_3247);
nand U894 (N_894,In_1800,In_2006);
nand U895 (N_895,In_738,In_3933);
nand U896 (N_896,In_4641,In_3227);
or U897 (N_897,In_3631,In_3334);
or U898 (N_898,In_4701,In_4057);
xor U899 (N_899,In_4626,In_85);
xor U900 (N_900,In_1688,In_3490);
xor U901 (N_901,In_4234,In_4704);
nand U902 (N_902,In_4642,In_4947);
nand U903 (N_903,In_4008,In_3344);
or U904 (N_904,In_1214,In_3413);
nand U905 (N_905,In_2451,In_3785);
xor U906 (N_906,In_3142,In_3111);
and U907 (N_907,In_12,In_1798);
or U908 (N_908,In_2595,In_3636);
and U909 (N_909,In_3595,In_2087);
and U910 (N_910,In_3876,In_1978);
or U911 (N_911,In_4897,In_3390);
and U912 (N_912,In_3981,In_641);
nand U913 (N_913,In_842,In_4983);
or U914 (N_914,In_4832,In_2196);
xor U915 (N_915,In_4298,In_126);
or U916 (N_916,In_3521,In_4923);
xor U917 (N_917,In_2787,In_3166);
and U918 (N_918,In_1540,In_3720);
nand U919 (N_919,In_4004,In_1495);
nand U920 (N_920,In_2757,In_943);
nor U921 (N_921,In_580,In_1578);
nor U922 (N_922,In_3914,In_3835);
or U923 (N_923,In_3368,In_3587);
nand U924 (N_924,In_767,In_1821);
or U925 (N_925,In_2974,In_1696);
xor U926 (N_926,In_82,In_3744);
nor U927 (N_927,In_3948,In_161);
nor U928 (N_928,In_2218,In_4002);
xnor U929 (N_929,In_757,In_3407);
nand U930 (N_930,In_2198,In_4852);
or U931 (N_931,In_1376,In_3809);
nor U932 (N_932,In_3822,In_442);
nand U933 (N_933,In_4130,In_1235);
xnor U934 (N_934,In_2586,In_3443);
or U935 (N_935,In_666,In_359);
and U936 (N_936,In_3290,In_3764);
nor U937 (N_937,In_3561,In_2395);
xor U938 (N_938,In_3475,In_2284);
nand U939 (N_939,In_460,In_723);
nand U940 (N_940,In_3666,In_494);
xor U941 (N_941,In_1485,In_271);
and U942 (N_942,In_2545,In_2792);
and U943 (N_943,In_1212,In_4770);
nand U944 (N_944,In_3852,In_2197);
and U945 (N_945,In_3331,In_2408);
nand U946 (N_946,In_531,In_3164);
xor U947 (N_947,In_2913,In_4647);
nand U948 (N_948,In_1122,In_2491);
or U949 (N_949,In_1913,In_407);
or U950 (N_950,In_1687,In_1974);
nand U951 (N_951,In_338,In_2767);
nand U952 (N_952,In_4301,In_4185);
xnor U953 (N_953,In_1961,In_1559);
and U954 (N_954,In_3620,In_3624);
nand U955 (N_955,In_3201,In_125);
nand U956 (N_956,In_4795,In_4389);
nand U957 (N_957,In_486,In_1238);
xnor U958 (N_958,In_4363,In_2536);
nand U959 (N_959,In_2705,In_1960);
nand U960 (N_960,In_2611,In_4901);
and U961 (N_961,In_258,In_2163);
or U962 (N_962,In_4854,In_3042);
nand U963 (N_963,In_4710,In_253);
nand U964 (N_964,In_3226,In_264);
nor U965 (N_965,In_2102,In_4589);
xnor U966 (N_966,In_70,In_2966);
nor U967 (N_967,In_1952,In_375);
xor U968 (N_968,In_3488,In_4915);
or U969 (N_969,In_3937,In_3942);
and U970 (N_970,In_3886,In_3833);
or U971 (N_971,In_3463,In_4142);
or U972 (N_972,In_727,In_2365);
nand U973 (N_973,In_1501,In_4640);
xnor U974 (N_974,In_2656,In_1799);
nand U975 (N_975,In_3990,In_806);
nor U976 (N_976,In_4799,In_4842);
and U977 (N_977,In_1101,In_429);
and U978 (N_978,In_3527,In_2957);
nand U979 (N_979,In_2513,In_414);
and U980 (N_980,In_4101,In_236);
xor U981 (N_981,In_121,In_2577);
xor U982 (N_982,In_1683,In_765);
or U983 (N_983,In_2867,In_1430);
xnor U984 (N_984,In_4525,In_2676);
or U985 (N_985,In_1581,In_3650);
xnor U986 (N_986,In_4539,In_3169);
nand U987 (N_987,In_3547,In_4514);
or U988 (N_988,In_4080,In_1513);
xnor U989 (N_989,In_2189,In_2212);
nand U990 (N_990,In_1331,In_182);
xnor U991 (N_991,In_1668,In_48);
and U992 (N_992,In_3459,In_2902);
or U993 (N_993,In_2278,In_3251);
nor U994 (N_994,In_225,In_742);
nor U995 (N_995,In_1919,In_4513);
and U996 (N_996,In_759,In_2148);
xor U997 (N_997,In_1019,In_2658);
nand U998 (N_998,In_2171,In_3414);
nand U999 (N_999,In_3002,In_905);
nor U1000 (N_1000,In_2515,In_4674);
or U1001 (N_1001,In_2020,In_2450);
or U1002 (N_1002,In_2351,In_2088);
nor U1003 (N_1003,In_4709,In_3416);
and U1004 (N_1004,In_2969,In_4500);
or U1005 (N_1005,In_1313,In_4609);
or U1006 (N_1006,In_4819,In_547);
or U1007 (N_1007,In_2137,In_3724);
nor U1008 (N_1008,In_223,In_2937);
nand U1009 (N_1009,In_3340,In_3161);
or U1010 (N_1010,In_4838,In_3630);
and U1011 (N_1011,In_3102,In_4582);
xor U1012 (N_1012,In_1754,In_4989);
or U1013 (N_1013,In_4627,In_3319);
or U1014 (N_1014,In_830,In_1155);
or U1015 (N_1015,In_1771,In_1033);
nand U1016 (N_1016,In_631,In_2832);
and U1017 (N_1017,In_2938,In_3759);
nor U1018 (N_1018,In_2895,In_963);
nand U1019 (N_1019,In_4939,In_1379);
xor U1020 (N_1020,In_4844,In_2123);
xnor U1021 (N_1021,In_2091,In_3185);
and U1022 (N_1022,In_2889,In_582);
xor U1023 (N_1023,In_2169,In_2188);
or U1024 (N_1024,In_3203,In_1592);
or U1025 (N_1025,In_2568,In_4223);
nor U1026 (N_1026,In_4960,In_192);
nor U1027 (N_1027,In_3144,In_28);
nand U1028 (N_1028,In_2114,In_345);
or U1029 (N_1029,In_3867,In_4522);
and U1030 (N_1030,In_2504,In_3779);
xnor U1031 (N_1031,In_1049,In_2670);
and U1032 (N_1032,In_750,In_4051);
nand U1033 (N_1033,In_3772,In_4711);
or U1034 (N_1034,In_1692,In_841);
nor U1035 (N_1035,In_4887,In_1766);
or U1036 (N_1036,In_3046,In_3924);
nor U1037 (N_1037,In_4139,In_4662);
nor U1038 (N_1038,In_880,In_3632);
nor U1039 (N_1039,In_1848,In_507);
nand U1040 (N_1040,In_4559,In_2252);
and U1041 (N_1041,In_3951,In_2152);
xor U1042 (N_1042,In_3593,In_4566);
xor U1043 (N_1043,In_4286,In_4869);
nor U1044 (N_1044,In_2971,In_2659);
nor U1045 (N_1045,In_1891,In_1245);
nand U1046 (N_1046,In_954,In_3672);
nand U1047 (N_1047,In_4437,In_2154);
xnor U1048 (N_1048,In_831,In_3447);
and U1049 (N_1049,In_2329,In_4579);
and U1050 (N_1050,In_2760,In_2067);
nor U1051 (N_1051,In_111,In_1670);
xor U1052 (N_1052,In_1357,In_2860);
or U1053 (N_1053,In_946,In_4505);
and U1054 (N_1054,In_2646,In_1163);
nor U1055 (N_1055,In_1422,In_1573);
xnor U1056 (N_1056,In_1375,In_1041);
xnor U1057 (N_1057,In_2308,In_3671);
xnor U1058 (N_1058,In_1362,In_4546);
xnor U1059 (N_1059,In_2896,In_912);
and U1060 (N_1060,In_2348,In_2604);
nand U1061 (N_1061,In_3070,In_4894);
and U1062 (N_1062,In_3384,In_4747);
xnor U1063 (N_1063,In_3255,In_1804);
nor U1064 (N_1064,In_3177,In_3972);
nor U1065 (N_1065,In_2317,In_155);
nand U1066 (N_1066,In_1056,In_4820);
xnor U1067 (N_1067,In_636,In_715);
and U1068 (N_1068,In_1296,In_1279);
xnor U1069 (N_1069,In_3236,In_2615);
nand U1070 (N_1070,In_4849,In_4630);
and U1071 (N_1071,In_4615,In_1644);
and U1072 (N_1072,In_394,In_3894);
nor U1073 (N_1073,In_207,In_1091);
and U1074 (N_1074,In_3740,In_2838);
xor U1075 (N_1075,In_4406,In_3252);
nor U1076 (N_1076,In_1507,In_1445);
and U1077 (N_1077,In_4750,In_3121);
nand U1078 (N_1078,In_1900,In_3706);
and U1079 (N_1079,In_1875,In_3606);
or U1080 (N_1080,In_3551,In_4899);
or U1081 (N_1081,In_3542,In_1010);
nor U1082 (N_1082,In_1413,In_2452);
nand U1083 (N_1083,In_1036,In_838);
or U1084 (N_1084,In_1743,In_473);
or U1085 (N_1085,In_2582,In_406);
nor U1086 (N_1086,In_2623,In_534);
or U1087 (N_1087,In_60,In_2314);
and U1088 (N_1088,In_4608,In_2906);
and U1089 (N_1089,In_3193,In_4946);
xor U1090 (N_1090,In_4860,In_4706);
or U1091 (N_1091,In_2985,In_3326);
nor U1092 (N_1092,In_2801,In_4805);
or U1093 (N_1093,In_4721,In_2318);
and U1094 (N_1094,In_944,In_1058);
xnor U1095 (N_1095,In_4337,In_3634);
or U1096 (N_1096,In_3071,In_2345);
xor U1097 (N_1097,In_819,In_4423);
xnor U1098 (N_1098,In_921,In_3712);
and U1099 (N_1099,In_2778,In_1137);
nand U1100 (N_1100,In_2200,In_1598);
and U1101 (N_1101,In_2866,In_1223);
and U1102 (N_1102,In_3308,In_3612);
or U1103 (N_1103,In_3125,In_4586);
xor U1104 (N_1104,In_2103,In_4394);
nor U1105 (N_1105,In_4263,In_3791);
or U1106 (N_1106,In_3022,In_431);
and U1107 (N_1107,In_443,In_589);
or U1108 (N_1108,In_4481,In_426);
and U1109 (N_1109,In_3181,In_2726);
nor U1110 (N_1110,In_4072,In_4955);
nor U1111 (N_1111,In_3320,In_2342);
nor U1112 (N_1112,In_1535,In_169);
and U1113 (N_1113,In_4924,In_2687);
nand U1114 (N_1114,In_2871,In_2072);
or U1115 (N_1115,In_4553,In_2807);
xor U1116 (N_1116,In_2917,In_4935);
or U1117 (N_1117,In_4064,In_2022);
nor U1118 (N_1118,In_1135,In_1026);
or U1119 (N_1119,In_1153,In_55);
nand U1120 (N_1120,In_3723,In_704);
nor U1121 (N_1121,In_858,In_3347);
nor U1122 (N_1122,In_4422,In_4387);
nor U1123 (N_1123,In_4889,In_1590);
nor U1124 (N_1124,In_424,In_4524);
or U1125 (N_1125,In_1897,In_4304);
nor U1126 (N_1126,In_2911,In_2391);
nor U1127 (N_1127,In_7,In_1746);
nor U1128 (N_1128,In_3949,In_4071);
xnor U1129 (N_1129,In_3294,In_1768);
and U1130 (N_1130,In_4293,In_4277);
and U1131 (N_1131,In_1657,In_4366);
nor U1132 (N_1132,In_2181,In_1751);
xor U1133 (N_1133,In_2747,In_3448);
xor U1134 (N_1134,In_2270,In_2555);
or U1135 (N_1135,In_1977,In_1769);
or U1136 (N_1136,In_1863,In_569);
xnor U1137 (N_1137,In_4426,In_868);
nor U1138 (N_1138,In_1763,In_3575);
nand U1139 (N_1139,In_1139,In_3836);
or U1140 (N_1140,In_1125,In_3850);
and U1141 (N_1141,In_1428,In_2781);
xor U1142 (N_1142,In_2862,In_4909);
xnor U1143 (N_1143,In_4502,In_567);
or U1144 (N_1144,In_3345,In_969);
xnor U1145 (N_1145,In_2257,In_3138);
xnor U1146 (N_1146,In_979,In_3483);
or U1147 (N_1147,In_1302,In_1455);
nor U1148 (N_1148,In_1031,In_781);
xnor U1149 (N_1149,In_4285,In_2836);
or U1150 (N_1150,In_2700,In_4519);
nor U1151 (N_1151,In_3826,In_4913);
xnor U1152 (N_1152,In_2150,In_659);
nor U1153 (N_1153,In_2490,In_1359);
and U1154 (N_1154,In_2712,In_4436);
and U1155 (N_1155,In_1301,In_1548);
nand U1156 (N_1156,In_107,In_1446);
nor U1157 (N_1157,In_3992,In_3195);
or U1158 (N_1158,In_2459,In_2422);
nor U1159 (N_1159,In_2743,In_513);
nand U1160 (N_1160,In_986,In_2415);
xnor U1161 (N_1161,In_1475,In_1809);
nand U1162 (N_1162,In_2097,In_2657);
nand U1163 (N_1163,In_1714,In_149);
xnor U1164 (N_1164,In_1833,In_1703);
xnor U1165 (N_1165,In_2130,In_265);
nor U1166 (N_1166,In_3675,In_4383);
xor U1167 (N_1167,In_708,In_3718);
or U1168 (N_1168,In_2016,In_3364);
xnor U1169 (N_1169,In_1107,In_3899);
nand U1170 (N_1170,In_368,In_859);
or U1171 (N_1171,In_1497,In_4446);
nand U1172 (N_1172,In_1452,In_4644);
xnor U1173 (N_1173,In_4613,In_183);
and U1174 (N_1174,In_1691,In_4310);
nor U1175 (N_1175,In_3947,In_374);
xnor U1176 (N_1176,In_4349,In_1707);
or U1177 (N_1177,In_116,In_3017);
nand U1178 (N_1178,In_4523,In_808);
nor U1179 (N_1179,In_1958,In_1669);
nor U1180 (N_1180,In_4826,In_1370);
and U1181 (N_1181,In_1986,In_4585);
xnor U1182 (N_1182,In_4620,In_3113);
or U1183 (N_1183,In_2041,In_4364);
nor U1184 (N_1184,In_3199,In_2878);
and U1185 (N_1185,In_62,In_353);
nor U1186 (N_1186,In_230,In_4688);
xnor U1187 (N_1187,In_1547,In_1284);
xor U1188 (N_1188,In_4908,In_3586);
nand U1189 (N_1189,In_2607,In_1802);
xor U1190 (N_1190,In_3114,In_3687);
or U1191 (N_1191,In_4329,In_2059);
xor U1192 (N_1192,In_2548,In_3583);
nand U1193 (N_1193,In_420,In_4562);
or U1194 (N_1194,In_4152,In_4660);
nor U1195 (N_1195,In_1054,In_3838);
or U1196 (N_1196,In_4145,In_1407);
and U1197 (N_1197,In_3194,In_4645);
or U1198 (N_1198,In_4102,In_3770);
and U1199 (N_1199,In_4365,In_4588);
xnor U1200 (N_1200,In_4132,In_3393);
nor U1201 (N_1201,In_304,In_180);
xor U1202 (N_1202,In_4287,In_3204);
xnor U1203 (N_1203,In_100,In_3546);
xor U1204 (N_1204,In_1956,In_2082);
nand U1205 (N_1205,In_4549,In_4786);
and U1206 (N_1206,In_3872,In_1884);
and U1207 (N_1207,In_3229,In_4846);
nand U1208 (N_1208,In_39,In_3567);
nor U1209 (N_1209,In_2477,In_1866);
xor U1210 (N_1210,In_472,In_1666);
nand U1211 (N_1211,In_3366,In_1702);
xnor U1212 (N_1212,In_2360,In_4729);
or U1213 (N_1213,In_2281,In_4289);
nand U1214 (N_1214,In_3978,In_3069);
nor U1215 (N_1215,In_3163,In_2050);
xor U1216 (N_1216,In_2099,In_1521);
and U1217 (N_1217,In_32,In_1257);
nor U1218 (N_1218,In_1878,In_753);
and U1219 (N_1219,In_4384,In_1849);
or U1220 (N_1220,In_366,In_953);
nor U1221 (N_1221,In_1240,In_1008);
or U1222 (N_1222,In_457,In_3132);
nand U1223 (N_1223,In_2900,In_3906);
xnor U1224 (N_1224,In_2356,In_3473);
xnor U1225 (N_1225,In_413,In_2335);
nor U1226 (N_1226,In_1807,In_4066);
and U1227 (N_1227,In_1969,In_1042);
nor U1228 (N_1228,In_1145,In_4948);
and U1229 (N_1229,In_2404,In_176);
and U1230 (N_1230,In_4299,In_833);
nand U1231 (N_1231,In_625,In_3233);
xnor U1232 (N_1232,In_1014,In_950);
or U1233 (N_1233,In_4804,In_1608);
nor U1234 (N_1234,In_2630,In_4073);
nor U1235 (N_1235,In_3,In_2480);
or U1236 (N_1236,In_726,In_925);
or U1237 (N_1237,In_1597,In_4628);
nand U1238 (N_1238,In_2739,In_2187);
nand U1239 (N_1239,In_2987,In_4547);
nand U1240 (N_1240,In_3896,In_888);
nor U1241 (N_1241,In_2240,In_3683);
nor U1242 (N_1242,In_1187,In_988);
xnor U1243 (N_1243,In_718,In_1186);
nand U1244 (N_1244,In_1373,In_173);
and U1245 (N_1245,In_751,In_3350);
and U1246 (N_1246,In_283,In_2716);
nor U1247 (N_1247,In_2920,In_501);
xnor U1248 (N_1248,In_2579,In_2098);
and U1249 (N_1249,In_3765,In_1037);
nor U1250 (N_1250,In_3649,In_3158);
nand U1251 (N_1251,In_1496,In_2751);
nand U1252 (N_1252,In_4753,In_1050);
xor U1253 (N_1253,In_2372,In_4870);
nand U1254 (N_1254,In_4475,In_1269);
and U1255 (N_1255,In_4996,In_1709);
xor U1256 (N_1256,In_3388,In_1568);
or U1257 (N_1257,In_871,In_94);
xor U1258 (N_1258,In_985,In_3406);
xor U1259 (N_1259,In_863,In_529);
and U1260 (N_1260,In_1190,In_1642);
or U1261 (N_1261,In_4850,In_1489);
xnor U1262 (N_1262,In_2856,In_156);
and U1263 (N_1263,In_1280,In_444);
nor U1264 (N_1264,In_4663,In_4032);
nor U1265 (N_1265,In_3667,In_4269);
nor U1266 (N_1266,In_1307,In_4380);
or U1267 (N_1267,In_1855,In_4526);
or U1268 (N_1268,In_4940,In_4652);
xor U1269 (N_1269,In_1282,In_4634);
or U1270 (N_1270,In_2191,In_4831);
or U1271 (N_1271,In_73,In_1575);
xnor U1272 (N_1272,In_3831,In_404);
nor U1273 (N_1273,In_1928,In_3068);
xor U1274 (N_1274,In_2161,In_3167);
and U1275 (N_1275,In_40,In_873);
xor U1276 (N_1276,In_2249,In_3098);
nand U1277 (N_1277,In_1024,In_3023);
nand U1278 (N_1278,In_604,In_1674);
or U1279 (N_1279,In_934,In_4797);
nor U1280 (N_1280,In_796,In_3234);
nor U1281 (N_1281,In_1491,In_612);
nor U1282 (N_1282,In_2961,In_2262);
nand U1283 (N_1283,In_1755,In_2886);
xor U1284 (N_1284,In_3305,In_298);
nor U1285 (N_1285,In_3110,In_1500);
nor U1286 (N_1286,In_1332,In_3355);
nor U1287 (N_1287,In_3365,In_2327);
xor U1288 (N_1288,In_4254,In_2031);
nor U1289 (N_1289,In_4914,In_4177);
or U1290 (N_1290,In_329,In_2379);
xor U1291 (N_1291,In_1628,In_168);
or U1292 (N_1292,In_2076,In_4117);
nor U1293 (N_1293,In_1029,In_4895);
xor U1294 (N_1294,In_4684,In_4572);
nor U1295 (N_1295,In_16,In_57);
or U1296 (N_1296,In_1003,In_1060);
and U1297 (N_1297,In_606,In_2478);
xor U1298 (N_1298,In_3732,In_3482);
and U1299 (N_1299,In_4035,In_3771);
nor U1300 (N_1300,In_1386,In_1292);
and U1301 (N_1301,In_3339,In_878);
and U1302 (N_1302,In_30,In_756);
nand U1303 (N_1303,In_229,In_103);
or U1304 (N_1304,In_1860,In_4330);
xor U1305 (N_1305,In_4202,In_1654);
and U1306 (N_1306,In_558,In_3302);
and U1307 (N_1307,In_3208,In_1068);
and U1308 (N_1308,In_3888,In_118);
xor U1309 (N_1309,In_2653,In_4112);
or U1310 (N_1310,In_4479,In_1006);
nand U1311 (N_1311,In_2079,In_25);
nand U1312 (N_1312,In_3079,In_3970);
and U1313 (N_1313,In_109,In_574);
nand U1314 (N_1314,In_3788,In_924);
and U1315 (N_1315,In_4601,In_3332);
xor U1316 (N_1316,In_1417,In_621);
or U1317 (N_1317,In_2011,In_3295);
or U1318 (N_1318,In_1690,In_2389);
nand U1319 (N_1319,In_2946,In_1305);
nand U1320 (N_1320,In_3798,In_4780);
nand U1321 (N_1321,In_1776,In_2679);
xor U1322 (N_1322,In_4896,In_1717);
nand U1323 (N_1323,In_4833,In_1672);
nand U1324 (N_1324,In_95,In_669);
or U1325 (N_1325,In_4725,In_4958);
xnor U1326 (N_1326,In_2039,In_2732);
and U1327 (N_1327,In_1917,In_4461);
nor U1328 (N_1328,In_19,In_1511);
xor U1329 (N_1329,In_1333,In_2715);
nand U1330 (N_1330,In_2975,In_2202);
nand U1331 (N_1331,In_3225,In_2156);
xnor U1332 (N_1332,In_3890,In_545);
xnor U1333 (N_1333,In_1814,In_1285);
nor U1334 (N_1334,In_662,In_861);
or U1335 (N_1335,In_1757,In_2718);
nand U1336 (N_1336,In_1664,In_469);
xnor U1337 (N_1337,In_3889,In_3944);
nand U1338 (N_1338,In_2754,In_2336);
nand U1339 (N_1339,In_215,In_1229);
and U1340 (N_1340,In_4928,In_902);
nor U1341 (N_1341,In_3767,In_3103);
xor U1342 (N_1342,In_423,In_4295);
and U1343 (N_1343,In_4270,In_1063);
nor U1344 (N_1344,In_263,In_2925);
nand U1345 (N_1345,In_193,In_400);
xor U1346 (N_1346,In_141,In_3543);
nor U1347 (N_1347,In_3335,In_3338);
nand U1348 (N_1348,In_4186,In_3352);
nand U1349 (N_1349,In_3210,In_599);
nand U1350 (N_1350,In_3116,In_798);
and U1351 (N_1351,In_3588,In_4169);
or U1352 (N_1352,In_3003,In_1325);
xnor U1353 (N_1353,In_945,In_2131);
nor U1354 (N_1354,In_4680,In_870);
nand U1355 (N_1355,In_1964,In_1258);
and U1356 (N_1356,In_3909,In_1633);
xor U1357 (N_1357,In_2534,In_4760);
nand U1358 (N_1358,In_4632,In_2493);
and U1359 (N_1359,In_3248,In_3435);
or U1360 (N_1360,In_1528,In_2574);
nand U1361 (N_1361,In_4496,In_3722);
nand U1362 (N_1362,In_1377,In_328);
or U1363 (N_1363,In_3983,In_4247);
or U1364 (N_1364,In_2409,In_3849);
xor U1365 (N_1365,In_3119,In_4772);
nor U1366 (N_1366,In_2177,In_2872);
or U1367 (N_1367,In_3690,In_34);
nand U1368 (N_1368,In_2208,In_1818);
and U1369 (N_1369,In_1419,In_4936);
xnor U1370 (N_1370,In_3789,In_895);
and U1371 (N_1371,In_707,In_3504);
and U1372 (N_1372,In_1927,In_2625);
and U1373 (N_1373,In_2540,In_1892);
nand U1374 (N_1374,In_1173,In_2964);
and U1375 (N_1375,In_1635,In_4351);
xnor U1376 (N_1376,In_3977,In_1244);
or U1377 (N_1377,In_1479,In_1275);
or U1378 (N_1378,In_3465,In_1085);
and U1379 (N_1379,In_3107,In_2232);
nand U1380 (N_1380,In_539,In_4705);
xnor U1381 (N_1381,In_947,In_2136);
or U1382 (N_1382,In_3515,In_2573);
and U1383 (N_1383,In_4264,In_562);
and U1384 (N_1384,In_4495,In_276);
or U1385 (N_1385,In_217,In_3715);
or U1386 (N_1386,In_1478,In_4713);
xnor U1387 (N_1387,In_3851,In_926);
and U1388 (N_1388,In_4196,In_3379);
nor U1389 (N_1389,In_224,In_1994);
xnor U1390 (N_1390,In_2074,In_1350);
or U1391 (N_1391,In_2347,In_3472);
and U1392 (N_1392,In_3571,In_419);
nor U1393 (N_1393,In_4376,In_2556);
xnor U1394 (N_1394,In_3316,In_2848);
and U1395 (N_1395,In_3781,In_2047);
xor U1396 (N_1396,In_4085,In_2255);
and U1397 (N_1397,In_380,In_3665);
and U1398 (N_1398,In_4300,In_2107);
and U1399 (N_1399,In_3801,In_3117);
nor U1400 (N_1400,In_4938,In_3627);
and U1401 (N_1401,In_1080,In_1384);
and U1402 (N_1402,In_2765,In_1057);
or U1403 (N_1403,In_2260,In_2236);
or U1404 (N_1404,In_4567,In_3796);
or U1405 (N_1405,In_2258,In_684);
xnor U1406 (N_1406,In_146,In_4950);
xnor U1407 (N_1407,In_657,In_1480);
or U1408 (N_1408,In_4321,In_3496);
nor U1409 (N_1409,In_3918,In_4226);
nand U1410 (N_1410,In_46,In_624);
nand U1411 (N_1411,In_511,In_678);
nand U1412 (N_1412,In_3198,In_527);
and U1413 (N_1413,In_1987,In_219);
or U1414 (N_1414,In_4968,In_4244);
nor U1415 (N_1415,In_581,In_4424);
nand U1416 (N_1416,In_3514,In_2510);
xnor U1417 (N_1417,In_3404,In_2709);
xnor U1418 (N_1418,In_4910,In_382);
and U1419 (N_1419,In_2046,In_992);
and U1420 (N_1420,In_4194,In_3040);
xnor U1421 (N_1421,In_2984,In_4483);
and U1422 (N_1422,In_652,In_1982);
nand U1423 (N_1423,In_2704,In_3881);
xnor U1424 (N_1424,In_3576,In_3544);
nand U1425 (N_1425,In_437,In_4813);
xor U1426 (N_1426,In_2195,In_664);
nor U1427 (N_1427,In_4180,In_2332);
nand U1428 (N_1428,In_2609,In_4982);
nand U1429 (N_1429,In_1260,In_623);
nand U1430 (N_1430,In_4334,In_2462);
nand U1431 (N_1431,In_3862,In_3498);
and U1432 (N_1432,In_461,In_1600);
xor U1433 (N_1433,In_2138,In_2680);
or U1434 (N_1434,In_2419,In_2970);
nor U1435 (N_1435,In_1115,In_3590);
and U1436 (N_1436,In_1391,In_2313);
nand U1437 (N_1437,In_1185,In_2764);
nand U1438 (N_1438,In_3555,In_2135);
xor U1439 (N_1439,In_3378,In_720);
or U1440 (N_1440,In_4189,In_3211);
or U1441 (N_1441,In_2035,In_4292);
nor U1442 (N_1442,In_1546,In_4592);
nor U1443 (N_1443,In_4818,In_1338);
nor U1444 (N_1444,In_4390,In_4238);
and U1445 (N_1445,In_544,In_4206);
and U1446 (N_1446,In_1224,In_3499);
nor U1447 (N_1447,In_3192,In_823);
and U1448 (N_1448,In_1708,In_356);
nand U1449 (N_1449,In_491,In_4115);
nand U1450 (N_1450,In_1583,In_1756);
xnor U1451 (N_1451,In_4742,In_1625);
or U1452 (N_1452,In_2373,In_686);
nor U1453 (N_1453,In_4025,In_108);
and U1454 (N_1454,In_4354,In_268);
xor U1455 (N_1455,In_2492,In_4465);
nand U1456 (N_1456,In_3265,In_3445);
nor U1457 (N_1457,In_2880,In_1924);
nand U1458 (N_1458,In_3476,In_3705);
or U1459 (N_1459,In_2438,In_789);
nor U1460 (N_1460,In_2932,In_2972);
nand U1461 (N_1461,In_4091,In_2706);
or U1462 (N_1462,In_2693,In_793);
nor U1463 (N_1463,In_3174,In_4766);
nand U1464 (N_1464,In_3135,In_4979);
xor U1465 (N_1465,In_553,In_2226);
nand U1466 (N_1466,In_1105,In_1499);
nor U1467 (N_1467,In_4104,In_3698);
and U1468 (N_1468,In_849,In_1734);
xor U1469 (N_1469,In_3321,In_2246);
or U1470 (N_1470,In_942,In_2572);
nor U1471 (N_1471,In_2749,In_2773);
nor U1472 (N_1472,In_251,In_3403);
nor U1473 (N_1473,In_2499,In_3986);
and U1474 (N_1474,In_67,In_3735);
or U1475 (N_1475,In_4600,In_879);
nand U1476 (N_1476,In_2776,In_1053);
or U1477 (N_1477,In_3784,In_2979);
xor U1478 (N_1478,In_2675,In_1347);
xor U1479 (N_1479,In_4518,In_654);
or U1480 (N_1480,In_3343,In_2078);
xnor U1481 (N_1481,In_3982,In_4168);
xor U1482 (N_1482,In_3854,In_1312);
xor U1483 (N_1483,In_1735,In_1349);
xor U1484 (N_1484,In_3747,In_1647);
nand U1485 (N_1485,In_4090,In_2692);
and U1486 (N_1486,In_3035,In_564);
xor U1487 (N_1487,In_4016,In_3293);
nand U1488 (N_1488,In_1966,In_1271);
and U1489 (N_1489,In_3509,In_2564);
or U1490 (N_1490,In_1983,In_476);
or U1491 (N_1491,In_2819,In_2940);
nand U1492 (N_1492,In_1531,In_729);
nand U1493 (N_1493,In_815,In_500);
nor U1494 (N_1494,In_300,In_2738);
nand U1495 (N_1495,In_1933,In_3238);
or U1496 (N_1496,In_855,In_1832);
xor U1497 (N_1497,In_284,In_4912);
or U1498 (N_1498,In_3314,In_2669);
nand U1499 (N_1499,In_2115,In_1562);
xnor U1500 (N_1500,In_4827,In_595);
and U1501 (N_1501,In_2628,In_4654);
and U1502 (N_1502,In_856,In_1889);
or U1503 (N_1503,In_2789,In_3493);
and U1504 (N_1504,In_1110,In_3646);
nand U1505 (N_1505,In_739,In_1659);
xor U1506 (N_1506,In_1459,In_3470);
xor U1507 (N_1507,In_1626,In_3875);
nor U1508 (N_1508,In_4598,In_2417);
or U1509 (N_1509,In_4883,In_3893);
and U1510 (N_1510,In_4611,In_3015);
nor U1511 (N_1511,In_2125,In_4415);
nor U1512 (N_1512,In_602,In_1320);
and U1513 (N_1513,In_228,In_811);
or U1514 (N_1514,In_4764,In_2698);
and U1515 (N_1515,In_4106,In_1326);
or U1516 (N_1516,In_3073,In_318);
nand U1517 (N_1517,In_234,In_2551);
xor U1518 (N_1518,In_2877,In_914);
nor U1519 (N_1519,In_3420,In_730);
nor U1520 (N_1520,In_2460,In_889);
xnor U1521 (N_1521,In_2149,In_1287);
nor U1522 (N_1522,In_4501,In_249);
or U1523 (N_1523,In_3349,In_3439);
xnor U1524 (N_1524,In_3093,In_1813);
nor U1525 (N_1525,In_2965,In_2320);
or U1526 (N_1526,In_1203,In_2324);
nand U1527 (N_1527,In_645,In_1015);
and U1528 (N_1528,In_2731,In_1083);
and U1529 (N_1529,In_4261,In_1246);
xnor U1530 (N_1530,In_2626,In_2338);
nand U1531 (N_1531,In_3559,In_302);
and U1532 (N_1532,In_4564,In_3431);
nor U1533 (N_1533,In_2892,In_1817);
and U1534 (N_1534,In_2496,In_4792);
or U1535 (N_1535,In_860,In_4109);
nand U1536 (N_1536,In_817,In_1643);
nor U1537 (N_1537,In_1412,In_153);
nand U1538 (N_1538,In_3756,In_570);
and U1539 (N_1539,In_409,In_65);
nand U1540 (N_1540,In_2847,In_3996);
and U1541 (N_1541,In_2962,In_3832);
xnor U1542 (N_1542,In_2668,In_2370);
and U1543 (N_1543,In_4521,In_3786);
nor U1544 (N_1544,In_616,In_4778);
nor U1545 (N_1545,In_4730,In_3011);
or U1546 (N_1546,In_1093,In_3087);
and U1547 (N_1547,In_1851,In_618);
and U1548 (N_1548,In_514,In_2287);
nand U1549 (N_1549,In_235,In_1903);
or U1550 (N_1550,In_1482,In_3934);
or U1551 (N_1551,In_4661,In_2584);
nand U1552 (N_1552,In_355,In_1100);
nor U1553 (N_1553,In_752,In_4231);
xor U1554 (N_1554,In_3839,In_4136);
nor U1555 (N_1555,In_4214,In_1520);
nor U1556 (N_1556,In_2143,In_4531);
nand U1557 (N_1557,In_314,In_3993);
and U1558 (N_1558,In_3898,In_3059);
xor U1559 (N_1559,In_1976,In_4855);
nor U1560 (N_1560,In_27,In_4224);
and U1561 (N_1561,In_4796,In_3452);
nor U1562 (N_1562,In_568,In_4069);
or U1563 (N_1563,In_846,In_4303);
nand U1564 (N_1564,In_2734,In_3969);
nand U1565 (N_1565,In_3362,In_3508);
nor U1566 (N_1566,In_4964,In_4053);
nand U1567 (N_1567,In_3104,In_3401);
xnor U1568 (N_1568,In_1549,In_4031);
xor U1569 (N_1569,In_2280,In_456);
nand U1570 (N_1570,In_3433,In_4252);
nor U1571 (N_1571,In_1281,In_3377);
or U1572 (N_1572,In_2518,In_2479);
and U1573 (N_1573,In_877,In_3273);
or U1574 (N_1574,In_4019,In_2488);
nor U1575 (N_1575,In_884,In_939);
nand U1576 (N_1576,In_2785,In_2565);
nand U1577 (N_1577,In_3050,In_3014);
nor U1578 (N_1578,In_3979,In_3436);
and U1579 (N_1579,In_2394,In_4961);
or U1580 (N_1580,In_4149,In_1594);
and U1581 (N_1581,In_2931,In_1394);
nand U1582 (N_1582,In_2063,In_4929);
nor U1583 (N_1583,In_3780,In_3228);
and U1584 (N_1584,In_3136,In_2722);
nand U1585 (N_1585,In_4027,In_5);
and U1586 (N_1586,In_4385,In_445);
and U1587 (N_1587,In_4028,In_4974);
or U1588 (N_1588,In_648,In_3438);
or U1589 (N_1589,In_609,In_3336);
and U1590 (N_1590,In_829,In_2239);
nand U1591 (N_1591,In_2671,In_2511);
nor U1592 (N_1592,In_4397,In_1369);
xor U1593 (N_1593,In_496,In_2473);
xor U1594 (N_1594,In_4552,In_144);
xor U1595 (N_1595,In_2784,In_2100);
nand U1596 (N_1596,In_3141,In_3284);
nor U1597 (N_1597,In_4489,In_4987);
nor U1598 (N_1598,In_676,In_4550);
xnor U1599 (N_1599,In_1016,In_1174);
and U1600 (N_1600,In_315,In_4282);
or U1601 (N_1601,In_247,In_2007);
nand U1602 (N_1602,In_396,In_2603);
or U1603 (N_1603,In_15,In_1272);
xor U1604 (N_1604,In_4861,In_317);
or U1605 (N_1605,In_4656,In_548);
nor U1606 (N_1606,In_4240,In_291);
or U1607 (N_1607,In_2268,In_1104);
or U1608 (N_1608,In_172,In_415);
nand U1609 (N_1609,In_1098,In_2276);
or U1610 (N_1610,In_809,In_834);
or U1611 (N_1611,In_1985,In_4205);
nand U1612 (N_1612,In_4787,In_996);
and U1613 (N_1613,In_452,In_1765);
xor U1614 (N_1614,In_2522,In_1805);
nand U1615 (N_1615,In_3806,In_3818);
nor U1616 (N_1616,In_1552,In_3920);
xor U1617 (N_1617,In_538,In_2433);
and U1618 (N_1618,In_4898,In_3568);
nor U1619 (N_1619,In_4735,In_2392);
nor U1620 (N_1620,In_2544,In_3469);
nor U1621 (N_1621,In_2695,In_1931);
and U1622 (N_1622,In_4865,In_3664);
xnor U1623 (N_1623,In_1086,In_4451);
or U1624 (N_1624,In_2111,In_387);
and U1625 (N_1625,In_2977,In_2617);
or U1626 (N_1626,In_2561,In_4507);
or U1627 (N_1627,In_187,In_361);
or U1628 (N_1628,In_566,In_2454);
or U1629 (N_1629,In_2497,In_398);
xor U1630 (N_1630,In_3009,In_2243);
xnor U1631 (N_1631,In_434,In_3371);
or U1632 (N_1632,In_2155,In_2516);
or U1633 (N_1633,In_2632,In_3554);
nand U1634 (N_1634,In_3754,In_2567);
xor U1635 (N_1635,In_745,In_4574);
nand U1636 (N_1636,In_2557,In_1165);
and U1637 (N_1637,In_2939,In_2558);
nor U1638 (N_1638,In_4536,In_3530);
nor U1639 (N_1639,In_4044,In_4342);
xnor U1640 (N_1640,In_3264,In_3262);
or U1641 (N_1641,In_1032,In_4839);
nor U1642 (N_1642,In_1762,In_1255);
xor U1643 (N_1643,In_2947,In_1464);
xnor U1644 (N_1644,In_2690,In_4320);
or U1645 (N_1645,In_3602,In_250);
nand U1646 (N_1646,In_3153,In_1316);
nand U1647 (N_1647,In_2160,In_2220);
and U1648 (N_1648,In_3891,In_1545);
nor U1649 (N_1649,In_1619,In_3324);
or U1650 (N_1650,In_4038,In_1997);
xnor U1651 (N_1651,In_3758,In_20);
nand U1652 (N_1652,In_2533,In_989);
xnor U1653 (N_1653,In_2539,In_2060);
and U1654 (N_1654,In_1327,In_3710);
nand U1655 (N_1655,In_2056,In_4188);
and U1656 (N_1656,In_744,In_4783);
nor U1657 (N_1657,In_1584,In_4858);
nor U1658 (N_1658,In_2052,In_2677);
and U1659 (N_1659,In_3955,In_1020);
or U1660 (N_1660,In_4571,In_3497);
xor U1661 (N_1661,In_1822,In_59);
and U1662 (N_1662,In_3736,In_3963);
xnor U1663 (N_1663,In_4733,In_2418);
nand U1664 (N_1664,In_3430,In_2354);
or U1665 (N_1665,In_4762,In_2384);
or U1666 (N_1666,In_1523,In_3461);
or U1667 (N_1667,In_1132,In_1947);
nor U1668 (N_1668,In_2245,In_4129);
nand U1669 (N_1669,In_743,In_1596);
nor U1670 (N_1670,In_4825,In_1352);
nand U1671 (N_1671,In_3244,In_1159);
nor U1672 (N_1672,In_3012,In_4060);
nand U1673 (N_1673,In_3005,In_1064);
xnor U1674 (N_1674,In_2474,In_2214);
nand U1675 (N_1675,In_1720,In_2390);
nor U1676 (N_1676,In_2065,In_2803);
and U1677 (N_1677,In_1023,In_4499);
nand U1678 (N_1678,In_186,In_1199);
nor U1679 (N_1679,In_1705,In_4867);
and U1680 (N_1680,In_4808,In_3032);
nand U1681 (N_1681,In_2684,In_1409);
or U1682 (N_1682,In_2844,In_1251);
or U1683 (N_1683,In_2229,In_575);
and U1684 (N_1684,In_965,In_3074);
and U1685 (N_1685,In_1695,In_1151);
nor U1686 (N_1686,In_3246,In_326);
nor U1687 (N_1687,In_2042,In_3523);
xnor U1688 (N_1688,In_4098,In_1689);
nor U1689 (N_1689,In_2627,In_1711);
nand U1690 (N_1690,In_2993,In_4190);
nand U1691 (N_1691,In_47,In_1793);
nand U1692 (N_1692,In_1693,In_3232);
nor U1693 (N_1693,In_1365,In_685);
nand U1694 (N_1694,In_2901,In_1718);
or U1695 (N_1695,In_3097,In_702);
nor U1696 (N_1696,In_96,In_679);
nor U1697 (N_1697,In_3774,In_1477);
nor U1698 (N_1698,In_4199,In_2547);
or U1699 (N_1699,In_2637,In_313);
or U1700 (N_1700,In_3460,In_4362);
or U1701 (N_1701,In_3695,In_1571);
xor U1702 (N_1702,In_497,In_2407);
and U1703 (N_1703,In_998,In_3628);
and U1704 (N_1704,In_3322,In_3101);
and U1705 (N_1705,In_779,In_2639);
xor U1706 (N_1706,In_2439,In_3044);
xor U1707 (N_1707,In_202,In_2180);
nand U1708 (N_1708,In_3115,In_1871);
xnor U1709 (N_1709,In_722,In_9);
nand U1710 (N_1710,In_2427,In_3860);
nand U1711 (N_1711,In_1196,In_221);
or U1712 (N_1712,In_3004,In_1886);
or U1713 (N_1713,In_2144,In_4297);
nor U1714 (N_1714,In_3658,In_2605);
or U1715 (N_1715,In_3287,In_2449);
and U1716 (N_1716,In_2167,In_3168);
and U1717 (N_1717,In_2326,In_2388);
and U1718 (N_1718,In_3676,In_348);
xnor U1719 (N_1719,In_3976,In_4998);
xor U1720 (N_1720,In_766,In_325);
nand U1721 (N_1721,In_4740,In_371);
and U1722 (N_1722,In_4563,In_3692);
nor U1723 (N_1723,In_3310,In_957);
xnor U1724 (N_1724,In_106,In_770);
or U1725 (N_1725,In_1351,In_4210);
xor U1726 (N_1726,In_4484,In_3957);
and U1727 (N_1727,In_2727,In_2331);
or U1728 (N_1728,In_4486,In_3638);
or U1729 (N_1729,In_3458,In_450);
or U1730 (N_1730,In_4673,In_3950);
and U1731 (N_1731,In_4463,In_3635);
nand U1732 (N_1732,In_3100,In_2721);
and U1733 (N_1733,In_288,In_2543);
and U1734 (N_1734,In_279,In_4921);
xnor U1735 (N_1735,In_3001,In_721);
and U1736 (N_1736,In_4249,In_4830);
nor U1737 (N_1737,In_4942,In_864);
nand U1738 (N_1738,In_4322,In_2183);
or U1739 (N_1739,In_3961,In_3536);
nor U1740 (N_1740,In_980,In_4245);
xnor U1741 (N_1741,In_2930,In_3363);
xnor U1742 (N_1742,In_4272,In_1681);
xor U1743 (N_1743,In_1788,In_572);
xnor U1744 (N_1744,In_1486,In_2420);
xor U1745 (N_1745,In_3752,In_50);
xnor U1746 (N_1746,In_4368,In_1077);
nand U1747 (N_1747,In_4306,In_3286);
nor U1748 (N_1748,In_2494,In_4107);
and U1749 (N_1749,In_3027,In_1563);
nand U1750 (N_1750,In_551,In_2346);
nand U1751 (N_1751,In_3541,In_1128);
xor U1752 (N_1752,In_1215,In_3172);
nor U1753 (N_1753,In_854,In_4013);
nor U1754 (N_1754,In_3738,In_1710);
nor U1755 (N_1755,In_2980,In_3637);
and U1756 (N_1756,In_504,In_2271);
or U1757 (N_1757,In_4903,In_2192);
and U1758 (N_1758,In_293,In_124);
or U1759 (N_1759,In_2013,In_4096);
nor U1760 (N_1760,In_4449,In_1243);
nor U1761 (N_1761,In_3096,In_3847);
xnor U1762 (N_1762,In_1421,In_416);
or U1763 (N_1763,In_4791,In_2475);
nor U1764 (N_1764,In_851,In_1021);
or U1765 (N_1765,In_3585,In_3337);
or U1766 (N_1766,In_2008,In_4440);
and U1767 (N_1767,In_2400,In_468);
xnor U1768 (N_1768,In_3840,In_4092);
and U1769 (N_1769,In_1684,In_508);
nor U1770 (N_1770,In_1861,In_4319);
nor U1771 (N_1771,In_4554,In_674);
nand U1772 (N_1772,In_3613,In_596);
xnor U1773 (N_1773,In_467,In_3259);
nor U1774 (N_1774,In_3755,In_1134);
and U1775 (N_1775,In_2826,In_4328);
or U1776 (N_1776,In_1120,In_1437);
and U1777 (N_1777,In_3196,In_3212);
xor U1778 (N_1778,In_866,In_2636);
or U1779 (N_1779,In_4952,In_4798);
or U1780 (N_1780,In_3648,In_3333);
nand U1781 (N_1781,In_3126,In_526);
and U1782 (N_1782,In_3919,In_3279);
nor U1783 (N_1783,In_607,In_2406);
nand U1784 (N_1784,In_3162,In_227);
nand U1785 (N_1785,In_4271,In_4155);
nor U1786 (N_1786,In_1197,In_1893);
nor U1787 (N_1787,In_2685,In_4606);
and U1788 (N_1788,In_4692,In_1140);
nor U1789 (N_1789,In_2311,In_3795);
xnor U1790 (N_1790,In_2828,In_2960);
and U1791 (N_1791,In_4173,In_3160);
xnor U1792 (N_1792,In_2633,In_2166);
nor U1793 (N_1793,In_4676,In_1880);
nor U1794 (N_1794,In_540,In_2343);
nand U1795 (N_1795,In_1148,In_79);
nand U1796 (N_1796,In_3082,In_3711);
xor U1797 (N_1797,In_2530,In_4165);
nand U1798 (N_1798,In_2043,In_4727);
and U1799 (N_1799,In_213,In_1397);
nand U1800 (N_1800,In_1300,In_158);
or U1801 (N_1801,In_1510,In_4544);
nor U1802 (N_1802,In_3837,In_1114);
xor U1803 (N_1803,In_1770,In_154);
xnor U1804 (N_1804,In_4686,In_1075);
and U1805 (N_1805,In_4617,In_681);
xnor U1806 (N_1806,In_3021,In_844);
nor U1807 (N_1807,In_4232,In_1825);
nand U1808 (N_1808,In_3506,In_3998);
and U1809 (N_1809,In_928,In_2413);
nand U1810 (N_1810,In_3792,In_4470);
nand U1811 (N_1811,In_4435,In_1864);
nor U1812 (N_1812,In_3147,In_1487);
nor U1813 (N_1813,In_3823,In_4745);
and U1814 (N_1814,In_3730,In_4034);
nor U1815 (N_1815,In_1781,In_731);
or U1816 (N_1816,In_991,In_1231);
xnor U1817 (N_1817,In_4041,In_2092);
nor U1818 (N_1818,In_465,In_2870);
nor U1819 (N_1819,In_4687,In_897);
nand U1820 (N_1820,In_2813,In_4473);
nor U1821 (N_1821,In_3072,In_675);
nor U1822 (N_1822,In_2509,In_3152);
and U1823 (N_1823,In_4123,In_4259);
xor U1824 (N_1824,In_458,In_4934);
or U1825 (N_1825,In_4743,In_4931);
nor U1826 (N_1826,In_3533,In_1109);
xnor U1827 (N_1827,In_4973,In_703);
xnor U1828 (N_1828,In_4771,In_4209);
and U1829 (N_1829,In_428,In_4682);
nor U1830 (N_1830,In_2597,In_2182);
and U1831 (N_1831,In_231,In_1065);
and U1832 (N_1832,In_2954,In_1206);
or U1833 (N_1833,In_3512,In_4535);
or U1834 (N_1834,In_1283,In_1012);
nor U1835 (N_1835,In_1948,In_4836);
or U1836 (N_1836,In_4658,In_613);
nor U1837 (N_1837,In_403,In_4847);
nand U1838 (N_1838,In_1447,In_918);
or U1839 (N_1839,In_4315,In_1038);
nor U1840 (N_1840,In_2299,In_2472);
nor U1841 (N_1841,In_1219,In_3622);
or U1842 (N_1842,In_1601,In_1645);
nand U1843 (N_1843,In_639,In_4837);
or U1844 (N_1844,In_2282,In_1273);
xnor U1845 (N_1845,In_2521,In_1773);
and U1846 (N_1846,In_2323,In_4427);
nor U1847 (N_1847,In_1553,In_3099);
nand U1848 (N_1848,In_4413,In_1758);
and U1849 (N_1849,In_4014,In_3243);
nor U1850 (N_1850,In_3564,In_1697);
xnor U1851 (N_1851,In_3442,In_1827);
nand U1852 (N_1852,In_3987,In_2665);
nand U1853 (N_1853,In_4359,In_1176);
and U1854 (N_1854,In_2355,In_1340);
xor U1855 (N_1855,In_2184,In_2024);
xor U1856 (N_1856,In_2822,In_3725);
or U1857 (N_1857,In_273,In_2736);
nand U1858 (N_1858,In_1073,In_522);
nand U1859 (N_1859,In_4679,In_2840);
or U1860 (N_1860,In_321,In_446);
nand U1861 (N_1861,In_1432,In_447);
or U1862 (N_1862,In_1363,In_3913);
xnor U1863 (N_1863,In_1616,In_1786);
nand U1864 (N_1864,In_2541,In_4246);
nor U1865 (N_1865,In_2643,In_1613);
xor U1866 (N_1866,In_1119,In_3303);
or U1867 (N_1867,In_29,In_1291);
and U1868 (N_1868,In_2797,In_2292);
nand U1869 (N_1869,In_1308,In_185);
nand U1870 (N_1870,In_761,In_4949);
nor U1871 (N_1871,In_3289,In_3257);
nor U1872 (N_1872,In_1460,In_4504);
or U1873 (N_1873,In_4988,In_3468);
nand U1874 (N_1874,In_2194,In_3454);
nor U1875 (N_1875,In_3529,In_3188);
or U1876 (N_1876,In_2217,In_2827);
and U1877 (N_1877,In_3989,In_1097);
xnor U1878 (N_1878,In_892,In_777);
nand U1879 (N_1879,In_503,In_297);
xnor U1880 (N_1880,In_208,In_4040);
nand U1881 (N_1881,In_1895,In_4715);
and U1882 (N_1882,In_2779,In_4741);
or U1883 (N_1883,In_2808,In_4467);
nand U1884 (N_1884,In_147,In_1951);
or U1885 (N_1885,In_672,In_1661);
xnor U1886 (N_1886,In_4237,In_1820);
nand U1887 (N_1887,In_3900,In_966);
nor U1888 (N_1888,In_2922,In_1216);
xnor U1889 (N_1889,In_277,In_2682);
nand U1890 (N_1890,In_816,In_682);
or U1891 (N_1891,In_2761,In_3501);
and U1892 (N_1892,In_3128,In_362);
or U1893 (N_1893,In_4963,In_1039);
and U1894 (N_1894,In_3562,In_1944);
xor U1895 (N_1895,In_3597,In_481);
nor U1896 (N_1896,In_2635,In_1629);
or U1897 (N_1897,In_3563,In_587);
nor U1898 (N_1898,In_2882,In_2089);
nor U1899 (N_1899,In_2955,In_687);
or U1900 (N_1900,In_1309,In_2266);
nor U1901 (N_1901,In_4732,In_4918);
and U1902 (N_1902,In_4788,In_1942);
and U1903 (N_1903,In_4487,In_917);
xor U1904 (N_1904,In_2119,In_3734);
or U1905 (N_1905,In_4273,In_2471);
nor U1906 (N_1906,In_4981,In_312);
xnor U1907 (N_1907,In_4045,In_2383);
or U1908 (N_1908,In_1095,In_4121);
or U1909 (N_1909,In_2134,In_4022);
xnor U1910 (N_1910,In_4868,In_2307);
nor U1911 (N_1911,In_3048,In_1334);
and U1912 (N_1912,In_1418,In_4986);
or U1913 (N_1913,In_1414,In_4402);
nand U1914 (N_1914,In_2842,In_2369);
nand U1915 (N_1915,In_1732,In_1289);
nand U1916 (N_1916,In_4239,In_4429);
or U1917 (N_1917,In_1250,In_3061);
xnor U1918 (N_1918,In_2036,In_4399);
and U1919 (N_1919,In_1396,In_58);
xnor U1920 (N_1920,In_4650,In_2251);
xnor U1921 (N_1921,In_1721,In_2368);
and U1922 (N_1922,In_357,In_1274);
nor U1923 (N_1923,In_1764,In_3441);
or U1924 (N_1924,In_4192,In_3392);
and U1925 (N_1925,In_3019,In_3926);
and U1926 (N_1926,In_246,In_4218);
nand U1927 (N_1927,In_1867,In_2264);
nor U1928 (N_1928,In_4411,In_143);
xor U1929 (N_1929,In_2755,In_417);
nor U1930 (N_1930,In_3205,In_4222);
nor U1931 (N_1931,In_769,In_4448);
or U1932 (N_1932,In_2133,In_3534);
and U1933 (N_1933,In_2873,In_4537);
nor U1934 (N_1934,In_2587,In_578);
xor U1935 (N_1935,In_360,In_1984);
nor U1936 (N_1936,In_2673,In_4017);
nand U1937 (N_1937,In_2279,In_747);
or U1938 (N_1938,In_385,In_828);
xnor U1939 (N_1939,In_3283,In_4176);
xnor U1940 (N_1940,In_261,In_3912);
nand U1941 (N_1941,In_1147,In_2237);
xnor U1942 (N_1942,In_2859,In_929);
xnor U1943 (N_1943,In_4438,In_110);
nor U1944 (N_1944,In_4545,In_2909);
nand U1945 (N_1945,In_3763,In_397);
and U1946 (N_1946,In_2719,In_1431);
or U1947 (N_1947,In_1609,In_3372);
and U1948 (N_1948,In_4371,In_3421);
xnor U1949 (N_1949,In_377,In_93);
nor U1950 (N_1950,In_3938,In_1656);
xor U1951 (N_1951,In_3327,In_4262);
xnor U1952 (N_1952,In_710,In_4573);
and U1953 (N_1953,In_4434,In_3402);
or U1954 (N_1954,In_872,In_847);
or U1955 (N_1955,In_2576,In_1089);
or U1956 (N_1956,In_1175,In_3423);
or U1957 (N_1957,In_1856,In_1328);
or U1958 (N_1958,In_1518,In_655);
nand U1959 (N_1959,In_1981,In_2444);
xor U1960 (N_1960,In_2919,In_1658);
or U1961 (N_1961,In_1319,In_1336);
xor U1962 (N_1962,In_4047,In_1845);
nor U1963 (N_1963,In_66,In_840);
xor U1964 (N_1964,In_2526,In_1389);
nor U1965 (N_1965,In_1035,In_26);
nand U1966 (N_1966,In_948,In_4373);
or U1967 (N_1967,In_4508,In_725);
or U1968 (N_1968,In_195,In_4932);
and U1969 (N_1969,In_2421,In_799);
and U1970 (N_1970,In_3517,In_1620);
and U1971 (N_1971,In_4971,In_433);
and U1972 (N_1972,In_3719,In_4834);
and U1973 (N_1973,In_4369,In_36);
nor U1974 (N_1974,In_1202,In_4116);
xor U1975 (N_1975,In_3354,In_4361);
xor U1976 (N_1976,In_4172,In_784);
nand U1977 (N_1977,In_4353,In_123);
nand U1978 (N_1978,In_378,In_2897);
xnor U1979 (N_1979,In_157,In_1916);
nor U1980 (N_1980,In_3668,In_4469);
or U1981 (N_1981,In_4432,In_324);
or U1982 (N_1982,In_2982,In_1572);
and U1983 (N_1983,In_2084,In_4343);
nand U1984 (N_1984,In_2991,In_4646);
xnor U1985 (N_1985,In_3999,In_2583);
nand U1986 (N_1986,In_1456,In_502);
or U1987 (N_1987,In_2782,In_3020);
or U1988 (N_1988,In_665,In_3800);
or U1989 (N_1989,In_2426,In_3088);
nor U1990 (N_1990,In_1436,In_2025);
or U1991 (N_1991,In_3997,In_405);
or U1992 (N_1992,In_512,In_3396);
nand U1993 (N_1993,In_2145,In_488);
nand U1994 (N_1994,In_1448,In_2222);
xnor U1995 (N_1995,In_4625,In_243);
or U1996 (N_1996,In_3811,In_2823);
nor U1997 (N_1997,In_61,In_972);
or U1998 (N_1998,In_3883,In_1704);
and U1999 (N_1999,In_2069,In_4872);
nor U2000 (N_2000,N_1610,N_1308);
nor U2001 (N_2001,N_355,N_1099);
and U2002 (N_2002,N_922,N_1433);
or U2003 (N_2003,N_92,In_4430);
nand U2004 (N_2004,N_1932,N_370);
and U2005 (N_2005,N_1909,N_91);
and U2006 (N_2006,In_2710,In_1842);
nand U2007 (N_2007,N_1561,N_477);
xnor U2008 (N_2008,In_3041,N_665);
or U2009 (N_2009,N_909,N_894);
or U2010 (N_2010,N_845,N_1739);
nor U2011 (N_2011,N_1876,N_867);
and U2012 (N_2012,N_1089,N_997);
nand U2013 (N_2013,N_1450,N_825);
nor U2014 (N_2014,In_630,N_1382);
and U2015 (N_2015,In_342,N_490);
or U2016 (N_2016,N_1197,N_262);
and U2017 (N_2017,N_1741,In_2382);
xnor U2018 (N_2018,N_958,N_624);
or U2019 (N_2019,In_1932,N_175);
nand U2020 (N_2020,N_139,N_1816);
xor U2021 (N_2021,In_292,N_1032);
nor U2022 (N_2022,N_1481,N_809);
and U2023 (N_2023,In_4157,In_4874);
xnor U2024 (N_2024,In_4197,N_851);
xnor U2025 (N_2025,N_837,N_555);
and U2026 (N_2026,In_4859,N_171);
and U2027 (N_2027,N_1596,N_1408);
or U2028 (N_2028,N_94,In_3217);
nor U2029 (N_2029,N_783,N_674);
xor U2030 (N_2030,N_1149,N_1779);
and U2031 (N_2031,N_944,N_1146);
nor U2032 (N_2032,N_518,N_79);
xor U2033 (N_2033,In_622,N_1040);
nor U2034 (N_2034,N_300,N_1363);
nor U2035 (N_2035,In_2570,N_236);
or U2036 (N_2036,N_1436,N_1035);
nand U2037 (N_2037,N_1843,N_733);
nor U2038 (N_2038,N_1728,N_1860);
or U2039 (N_2039,In_3429,N_1888);
nor U2040 (N_2040,N_141,N_609);
xor U2041 (N_2041,N_738,N_1716);
or U2042 (N_2042,N_245,In_2907);
or U2043 (N_2043,N_956,In_4258);
and U2044 (N_2044,N_1396,N_663);
nand U2045 (N_2045,N_905,In_4015);
or U2046 (N_2046,In_4565,N_88);
or U2047 (N_2047,N_563,N_912);
or U2048 (N_2048,N_1713,In_4587);
nor U2049 (N_2049,N_266,In_280);
and U2050 (N_2050,In_1265,N_1462);
nor U2051 (N_2051,N_725,N_869);
xor U2052 (N_2052,N_1364,In_3686);
nand U2053 (N_2053,N_240,N_1542);
nand U2054 (N_2054,N_1067,In_498);
xnor U2055 (N_2055,N_1361,N_577);
or U2056 (N_2056,N_618,In_523);
nand U2057 (N_2057,N_312,In_4162);
nand U2058 (N_2058,N_1847,In_3437);
nor U2059 (N_2059,N_93,In_164);
nor U2060 (N_2060,N_1114,In_3858);
nor U2061 (N_2061,N_425,N_1689);
nor U2062 (N_2062,N_1045,N_5);
xnor U2063 (N_2063,N_1420,N_1650);
nand U2064 (N_2064,In_1310,N_964);
or U2065 (N_2065,N_1482,In_1341);
nor U2066 (N_2066,N_433,N_162);
or U2067 (N_2067,In_4700,N_1511);
nor U2068 (N_2068,N_1016,N_1472);
nor U2069 (N_2069,N_1071,N_1072);
nor U2070 (N_2070,In_1374,N_1572);
nand U2071 (N_2071,In_2432,N_1271);
nor U2072 (N_2072,In_3902,N_197);
nor U2073 (N_2073,N_1260,N_234);
or U2074 (N_2074,In_3213,N_1512);
and U2075 (N_2075,In_4621,In_1998);
and U2076 (N_2076,N_1231,N_1729);
xor U2077 (N_2077,N_1671,In_910);
nor U2078 (N_2078,In_2535,N_1185);
and U2079 (N_2079,In_3960,N_318);
nor U2080 (N_2080,N_168,N_1520);
nand U2081 (N_2081,In_4076,N_826);
and U2082 (N_2082,In_3471,N_726);
nand U2083 (N_2083,N_499,N_1905);
xor U2084 (N_2084,In_334,N_692);
or U2085 (N_2085,N_1452,N_1645);
or U2086 (N_2086,In_4290,N_34);
and U2087 (N_2087,In_1836,N_1960);
xor U2088 (N_2088,In_2737,N_254);
nor U2089 (N_2089,N_1992,N_1080);
and U2090 (N_2090,N_975,N_852);
nor U2091 (N_2091,N_1014,In_1481);
or U2092 (N_2092,N_1873,N_879);
nand U2093 (N_2093,N_1201,N_1144);
and U2094 (N_2094,In_2672,N_1269);
xnor U2095 (N_2095,In_4193,N_523);
and U2096 (N_2096,N_46,N_1344);
xnor U2097 (N_2097,In_1888,In_3357);
nand U2098 (N_2098,In_4164,In_591);
or U2099 (N_2099,N_1299,N_229);
nand U2100 (N_2100,In_2745,N_1367);
and U2101 (N_2101,In_4746,N_1176);
and U2102 (N_2102,N_410,N_1754);
nor U2103 (N_2103,In_1217,N_562);
and U2104 (N_2104,N_1188,In_2000);
or U2105 (N_2105,N_1621,N_1827);
xor U2106 (N_2106,N_1012,N_329);
and U2107 (N_2107,N_1912,N_828);
xnor U2108 (N_2108,N_675,N_259);
xor U2109 (N_2109,N_1219,N_730);
nor U2110 (N_2110,N_1976,N_315);
or U2111 (N_2111,N_1653,In_3306);
and U2112 (N_2112,N_80,N_704);
nor U2113 (N_2113,In_2662,N_1846);
or U2114 (N_2114,N_1319,N_1604);
nor U2115 (N_2115,In_941,N_1127);
nand U2116 (N_2116,In_1525,N_1745);
and U2117 (N_2117,In_379,N_19);
nand U2118 (N_2118,In_3060,N_1163);
xor U2119 (N_2119,N_981,In_4281);
nand U2120 (N_2120,N_1421,In_3921);
xor U2121 (N_2121,N_641,In_1778);
xnor U2122 (N_2122,N_270,N_566);
and U2123 (N_2123,In_4659,N_779);
xnor U2124 (N_2124,N_1444,In_269);
nor U2125 (N_2125,N_586,In_3298);
nand U2126 (N_2126,In_760,In_2825);
and U2127 (N_2127,N_1692,N_1614);
nor U2128 (N_2128,N_1765,N_1000);
nor U2129 (N_2129,In_3701,N_1737);
or U2130 (N_2130,N_1812,In_4576);
and U2131 (N_2131,N_653,N_953);
and U2132 (N_2132,In_4317,N_1335);
and U2133 (N_2133,N_1486,N_973);
or U2134 (N_2134,In_2215,N_1286);
or U2135 (N_2135,N_695,In_1943);
nand U2136 (N_2136,N_1661,N_1649);
nand U2137 (N_2137,N_903,N_858);
and U2138 (N_2138,N_1439,N_1525);
nor U2139 (N_2139,N_1730,N_1130);
and U2140 (N_2140,In_3778,N_272);
xor U2141 (N_2141,N_1505,N_1908);
nor U2142 (N_2142,In_35,N_743);
or U2143 (N_2143,N_574,N_821);
xor U2144 (N_2144,In_1253,N_1921);
xor U2145 (N_2145,N_448,N_1025);
or U2146 (N_2146,N_1063,In_1429);
or U2147 (N_2147,In_4716,N_600);
nand U2148 (N_2148,N_1404,N_1585);
xnor U2149 (N_2149,N_1077,N_1118);
nor U2150 (N_2150,In_791,N_787);
nor U2151 (N_2151,N_1097,N_750);
or U2152 (N_2152,In_1614,N_1441);
nand U2153 (N_2153,N_1519,N_933);
or U2154 (N_2154,N_1178,N_1143);
xor U2155 (N_2155,N_45,N_1759);
or U2156 (N_2156,N_47,N_1372);
xnor U2157 (N_2157,In_3737,In_881);
or U2158 (N_2158,In_1267,N_1959);
nand U2159 (N_2159,N_1915,In_88);
or U2160 (N_2160,N_1801,N_282);
nor U2161 (N_2161,N_521,N_1457);
xor U2162 (N_2162,N_406,N_934);
or U2163 (N_2163,In_1995,In_4200);
xor U2164 (N_2164,N_948,N_123);
or U2165 (N_2165,N_28,N_651);
and U2166 (N_2166,N_220,In_1593);
or U2167 (N_2167,In_3877,In_4048);
nor U2168 (N_2168,In_697,N_44);
nor U2169 (N_2169,N_812,In_920);
or U2170 (N_2170,N_1786,N_372);
and U2171 (N_2171,In_4726,N_900);
nand U2172 (N_2172,N_250,In_138);
or U2173 (N_2173,N_584,N_9);
or U2174 (N_2174,N_51,N_987);
xor U2175 (N_2175,In_1837,In_3398);
or U2176 (N_2176,N_1562,N_676);
or U2177 (N_2177,In_1094,In_127);
or U2178 (N_2178,N_540,In_807);
or U2179 (N_2179,In_1156,In_2330);
and U2180 (N_2180,N_1503,N_712);
xor U2181 (N_2181,N_1546,N_817);
and U2182 (N_2182,N_1894,N_429);
or U2183 (N_2183,N_1760,N_1315);
nand U2184 (N_2184,N_160,N_132);
nor U2185 (N_2185,In_3808,N_896);
or U2186 (N_2186,N_842,N_1615);
and U2187 (N_2187,In_1304,N_488);
and U2188 (N_2188,N_1936,N_531);
nand U2189 (N_2189,N_14,N_1620);
xnor U2190 (N_2190,N_633,N_1011);
xnor U2191 (N_2191,N_1670,N_1028);
or U2192 (N_2192,In_212,In_1606);
nor U2193 (N_2193,N_892,N_1631);
or U2194 (N_2194,N_1200,N_669);
nand U2195 (N_2195,N_369,N_590);
nand U2196 (N_2196,N_645,N_25);
nand U2197 (N_2197,In_3975,N_847);
nor U2198 (N_2198,In_3525,N_967);
nand U2199 (N_2199,N_115,N_696);
and U2200 (N_2200,In_3367,In_4388);
or U2201 (N_2201,In_3952,In_2863);
and U2202 (N_2202,N_289,N_85);
xor U2203 (N_2203,N_1076,N_1547);
and U2204 (N_2204,N_434,N_1613);
nor U2205 (N_2205,N_242,N_398);
nor U2206 (N_2206,N_959,N_1424);
nor U2207 (N_2207,N_1468,N_595);
or U2208 (N_2208,N_1339,N_1567);
nand U2209 (N_2209,N_349,N_153);
xor U2210 (N_2210,N_947,In_782);
nor U2211 (N_2211,In_4012,N_1236);
or U2212 (N_2212,N_1663,N_1373);
nand U2213 (N_2213,In_2505,N_1533);
or U2214 (N_2214,In_735,N_1586);
xnor U2215 (N_2215,N_1500,N_1872);
and U2216 (N_2216,N_542,N_769);
or U2217 (N_2217,In_792,N_1029);
or U2218 (N_2218,N_1640,N_1453);
nor U2219 (N_2219,In_3254,N_1541);
or U2220 (N_2220,N_1923,N_592);
nor U2221 (N_2221,N_1206,N_1151);
xnor U2222 (N_2222,In_4765,In_3856);
and U2223 (N_2223,In_4151,N_249);
or U2224 (N_2224,In_536,In_4814);
or U2225 (N_2225,In_2104,N_1731);
and U2226 (N_2226,N_1857,N_758);
nand U2227 (N_2227,N_1916,N_557);
nand U2228 (N_2228,In_1233,In_2553);
and U2229 (N_2229,N_844,N_951);
xnor U2230 (N_2230,N_1487,In_4335);
and U2231 (N_2231,In_4324,In_4203);
or U2232 (N_2232,N_932,N_1036);
nor U2233 (N_2233,N_883,N_2);
nand U2234 (N_2234,In_1949,In_4643);
nor U2235 (N_2235,N_1679,In_3768);
nor U2236 (N_2236,N_766,N_1991);
and U2237 (N_2237,N_679,N_1414);
nand U2238 (N_2238,In_2263,In_3415);
or U2239 (N_2239,N_49,N_1125);
and U2240 (N_2240,In_3245,N_1177);
xor U2241 (N_2241,N_381,N_1556);
and U2242 (N_2242,In_191,N_1117);
nand U2243 (N_2243,N_1557,N_1719);
nand U2244 (N_2244,In_4956,N_536);
and U2245 (N_2245,N_474,N_1289);
xor U2246 (N_2246,N_1884,In_2129);
xor U2247 (N_2247,N_100,N_1265);
nor U2248 (N_2248,In_4372,N_720);
or U2249 (N_2249,N_805,N_180);
nor U2250 (N_2250,N_1840,N_1774);
or U2251 (N_2251,N_646,In_2049);
xnor U2252 (N_2252,N_737,In_1712);
nand U2253 (N_2253,In_1462,N_227);
nand U2254 (N_2254,N_1173,N_1580);
and U2255 (N_2255,In_3552,N_1982);
nor U2256 (N_2256,N_331,N_1849);
and U2257 (N_2257,N_105,N_316);
or U2258 (N_2258,N_880,In_3643);
nor U2259 (N_2259,N_1961,N_90);
nand U2260 (N_2260,N_1135,N_1901);
or U2261 (N_2261,N_319,N_864);
xor U2262 (N_2262,N_111,N_1523);
or U2263 (N_2263,N_489,N_287);
nand U2264 (N_2264,N_917,N_252);
nor U2265 (N_2265,N_1672,In_588);
nand U2266 (N_2266,N_517,N_278);
nor U2267 (N_2267,N_647,N_591);
xor U2268 (N_2268,N_211,N_1554);
nor U2269 (N_2269,N_1013,N_1418);
nand U2270 (N_2270,N_1646,N_337);
nand U2271 (N_2271,N_1307,In_3532);
nor U2272 (N_2272,N_506,In_1920);
nor U2273 (N_2273,In_561,In_4182);
xor U2274 (N_2274,In_4829,N_1355);
and U2275 (N_2275,N_1049,In_346);
xor U2276 (N_2276,In_709,In_2752);
nor U2277 (N_2277,N_537,N_1515);
and U2278 (N_2278,N_1968,N_534);
nand U2279 (N_2279,N_1589,N_1132);
nor U2280 (N_2280,N_419,N_715);
nand U2281 (N_2281,N_1891,N_1855);
or U2282 (N_2282,N_1270,N_1978);
nand U2283 (N_2283,N_838,In_1632);
nor U2284 (N_2284,N_151,N_177);
nand U2285 (N_2285,N_1601,N_1226);
nand U2286 (N_2286,N_20,N_297);
and U2287 (N_2287,In_3081,In_4062);
xor U2288 (N_2288,N_441,In_4294);
and U2289 (N_2289,N_974,N_1509);
nand U2290 (N_2290,N_1255,N_1395);
and U2291 (N_2291,In_4759,In_3611);
and U2292 (N_2292,In_2503,In_1723);
or U2293 (N_2293,In_162,In_3387);
xor U2294 (N_2294,N_1350,In_1188);
and U2295 (N_2295,N_1600,N_232);
nand U2296 (N_2296,N_1458,In_3842);
or U2297 (N_2297,N_795,N_1819);
xor U2298 (N_2298,N_1538,N_24);
and U2299 (N_2299,In_3080,N_465);
xor U2300 (N_2300,N_1788,In_4629);
or U2301 (N_2301,In_432,N_13);
nor U2302 (N_2302,In_1047,In_2121);
nor U2303 (N_2303,N_320,In_4527);
or U2304 (N_2304,N_362,N_1369);
nor U2305 (N_2305,N_1701,N_672);
nand U2306 (N_2306,N_1093,N_1794);
nand U2307 (N_2307,N_544,N_1638);
or U2308 (N_2308,In_2786,N_1342);
xnor U2309 (N_2309,In_4542,N_1241);
nor U2310 (N_2310,In_3053,N_1243);
nand U2311 (N_2311,N_1340,N_597);
nand U2312 (N_2312,N_1278,N_357);
and U2313 (N_2313,In_3300,In_76);
nand U2314 (N_2314,N_273,In_1519);
or U2315 (N_2315,In_2227,N_1041);
xor U2316 (N_2316,N_206,N_222);
and U2317 (N_2317,N_859,N_1950);
or U2318 (N_2318,In_296,N_1537);
and U2319 (N_2319,In_3879,N_1321);
xnor U2320 (N_2320,In_487,N_1558);
nand U2321 (N_2321,In_4001,In_4902);
and U2322 (N_2322,N_1514,N_281);
or U2323 (N_2323,N_889,In_3143);
or U2324 (N_2324,In_4980,N_765);
xor U2325 (N_2325,N_545,In_1854);
or U2326 (N_2326,N_1881,In_1440);
or U2327 (N_2327,In_2374,N_12);
nor U2328 (N_2328,N_553,N_1101);
and U2329 (N_2329,In_3696,N_1285);
nor U2330 (N_2330,N_209,N_830);
and U2331 (N_2331,N_1836,N_1858);
or U2332 (N_2332,In_1580,In_813);
xnor U2333 (N_2333,N_1680,In_4970);
nand U2334 (N_2334,N_1612,N_1136);
xor U2335 (N_2335,N_1682,N_137);
and U2336 (N_2336,N_1817,N_446);
xnor U2337 (N_2337,In_4734,In_938);
or U2338 (N_2338,N_1919,N_1274);
and U2339 (N_2339,N_1979,N_1187);
xnor U2340 (N_2340,N_217,N_313);
xnor U2341 (N_2341,N_1980,In_3776);
xnor U2342 (N_2342,N_1814,N_244);
nor U2343 (N_2343,N_391,In_712);
and U2344 (N_2344,N_886,N_1242);
nand U2345 (N_2345,N_1530,In_1896);
nor U2346 (N_2346,In_3409,N_854);
nor U2347 (N_2347,In_1306,N_1681);
or U2348 (N_2348,N_69,In_4460);
or U2349 (N_2349,N_1575,N_925);
nand U2350 (N_2350,N_67,In_1045);
nand U2351 (N_2351,N_1153,N_364);
or U2352 (N_2352,N_221,In_1676);
nand U2353 (N_2353,N_882,N_1727);
xor U2354 (N_2354,In_913,N_794);
and U2355 (N_2355,N_1685,N_526);
nor U2356 (N_2356,N_1059,N_1448);
and U2357 (N_2357,N_60,N_705);
and U2358 (N_2358,N_700,In_2929);
xor U2359 (N_2359,N_1075,In_620);
nor U2360 (N_2360,N_1655,In_3644);
nand U2361 (N_2361,In_573,N_279);
xor U2362 (N_2362,N_1875,N_1922);
or U2363 (N_2363,N_1008,N_797);
nand U2364 (N_2364,In_4485,N_875);
or U2365 (N_2365,N_1989,In_1259);
or U2366 (N_2366,In_2165,N_1513);
nor U2367 (N_2367,In_3743,N_1704);
xor U2368 (N_2368,N_1632,In_2864);
and U2369 (N_2369,In_4756,In_402);
xnor U2370 (N_2370,N_921,N_1599);
and U2371 (N_2371,N_1676,In_2080);
xnor U2372 (N_2372,In_2293,N_400);
nor U2373 (N_2373,N_1693,In_4930);
nor U2374 (N_2374,N_1570,N_1956);
nor U2375 (N_2375,N_1733,N_611);
xnor U2376 (N_2376,In_909,In_1815);
or U2377 (N_2377,In_53,In_1806);
and U2378 (N_2378,In_4794,N_485);
nand U2379 (N_2379,N_322,In_3139);
and U2380 (N_2380,In_1048,In_1965);
or U2381 (N_2381,N_1262,N_761);
xnor U2382 (N_2382,N_1221,In_4447);
xnor U2383 (N_2383,In_1747,N_1643);
nor U2384 (N_2384,N_1399,In_4926);
xor U2385 (N_2385,N_7,In_399);
and U2386 (N_2386,N_1381,N_345);
or U2387 (N_2387,N_814,In_1434);
xor U2388 (N_2388,In_24,N_23);
and U2389 (N_2389,N_407,N_1290);
or U2390 (N_2390,N_1210,In_3802);
and U2391 (N_2391,N_1810,N_942);
and U2392 (N_2392,N_409,N_1882);
or U2393 (N_2393,In_3075,N_1057);
nand U2394 (N_2394,In_4985,N_112);
xor U2395 (N_2395,N_570,N_656);
xnor U2396 (N_2396,N_114,In_4408);
xor U2397 (N_2397,In_1801,N_1944);
or U2398 (N_2398,N_585,In_4327);
and U2399 (N_2399,In_4593,In_4719);
nand U2400 (N_2400,N_1972,N_1303);
and U2401 (N_2401,In_4755,In_3967);
nand U2402 (N_2402,N_1256,In_2924);
and U2403 (N_2403,N_1345,N_1471);
and U2404 (N_2404,N_694,In_188);
or U2405 (N_2405,In_1753,N_1393);
nand U2406 (N_2406,N_1109,N_1707);
xnor U2407 (N_2407,In_4666,N_200);
nor U2408 (N_2408,N_40,N_1432);
xor U2409 (N_2409,N_129,N_1506);
xnor U2410 (N_2410,N_1272,In_281);
xnor U2411 (N_2411,In_4331,N_832);
xnor U2412 (N_2412,In_4703,In_3084);
and U2413 (N_2413,N_1337,In_2458);
xnor U2414 (N_2414,N_1394,N_378);
or U2415 (N_2415,N_147,N_1995);
xnor U2416 (N_2416,In_2593,In_3657);
nor U2417 (N_2417,In_2081,In_427);
nor U2418 (N_2418,In_2291,In_3848);
nand U2419 (N_2419,N_140,N_443);
and U2420 (N_2420,N_1983,In_1210);
nor U2421 (N_2421,N_1060,In_3916);
and U2422 (N_2422,N_251,In_2221);
nand U2423 (N_2423,N_1238,N_698);
xnor U2424 (N_2424,N_1223,N_1357);
nor U2425 (N_2425,N_1440,In_3156);
or U2426 (N_2426,N_1683,N_226);
xnor U2427 (N_2427,N_872,In_4728);
nand U2428 (N_2428,In_68,In_1170);
nand U2429 (N_2429,In_2774,N_1435);
nand U2430 (N_2430,In_349,In_3700);
nand U2431 (N_2431,N_1662,In_425);
nand U2432 (N_2432,N_1973,In_3010);
nand U2433 (N_2433,N_344,N_955);
or U2434 (N_2434,In_1636,N_1110);
nand U2435 (N_2435,N_431,In_2055);
nor U2436 (N_2436,N_166,N_418);
or U2437 (N_2437,N_1098,In_1882);
nand U2438 (N_2438,In_4036,N_1085);
nor U2439 (N_2439,N_420,N_874);
nand U2440 (N_2440,In_556,N_210);
nor U2441 (N_2441,N_615,N_648);
or U2442 (N_2442,N_1634,In_4094);
or U2443 (N_2443,N_1196,In_2045);
or U2444 (N_2444,In_1127,N_1220);
nand U2445 (N_2445,N_789,In_142);
or U2446 (N_2446,In_2387,N_76);
or U2447 (N_2447,N_736,N_995);
nor U2448 (N_2448,N_269,N_1492);
nand U2449 (N_2449,N_1061,In_3034);
nor U2450 (N_2450,In_1649,N_1447);
or U2451 (N_2451,N_793,In_2302);
or U2452 (N_2452,In_2352,N_1082);
nor U2453 (N_2453,N_1442,In_2619);
nor U2454 (N_2454,N_1493,N_174);
or U2455 (N_2455,N_962,In_982);
and U2456 (N_2456,In_2874,In_3495);
xor U2457 (N_2457,N_1284,N_1212);
xor U2458 (N_2458,In_3882,In_1096);
xnor U2459 (N_2459,N_841,In_1195);
nor U2460 (N_2460,In_2296,In_4612);
nand U2461 (N_2461,In_2316,In_1638);
nor U2462 (N_2462,N_1611,N_486);
and U2463 (N_2463,N_1474,In_3841);
or U2464 (N_2464,N_503,In_2250);
nand U2465 (N_2465,N_1656,N_831);
or U2466 (N_2466,N_1711,N_1087);
nand U2467 (N_2467,N_1233,In_2590);
and U2468 (N_2468,N_502,In_2238);
xnor U2469 (N_2469,N_576,N_701);
and U2470 (N_2470,In_363,N_26);
and U2471 (N_2471,N_901,N_351);
and U2472 (N_2472,N_1006,N_1423);
or U2473 (N_2473,In_2289,N_1673);
and U2474 (N_2474,In_800,N_361);
nand U2475 (N_2475,In_1543,N_1287);
nor U2476 (N_2476,N_191,In_4378);
nor U2477 (N_2477,N_10,N_790);
nand U2478 (N_2478,N_1866,N_1895);
or U2479 (N_2479,N_1898,In_163);
nor U2480 (N_2480,In_1404,N_204);
nand U2481 (N_2481,In_4208,In_2990);
or U2482 (N_2482,N_1066,N_238);
and U2483 (N_2483,N_1002,In_1784);
or U2484 (N_2484,N_1166,N_816);
or U2485 (N_2485,N_1247,N_1155);
and U2486 (N_2486,In_2514,N_1485);
and U2487 (N_2487,In_1025,In_3892);
or U2488 (N_2488,N_1838,N_753);
or U2489 (N_2489,N_1422,In_3039);
nor U2490 (N_2490,In_2851,N_159);
xnor U2491 (N_2491,In_3805,In_287);
or U2492 (N_2492,N_1490,In_4905);
xnor U2493 (N_2493,N_1581,In_190);
nand U2494 (N_2494,N_1124,N_1325);
nand U2495 (N_2495,In_2875,N_888);
xnor U2496 (N_2496,N_1784,In_4358);
or U2497 (N_2497,In_1760,In_3449);
or U2498 (N_2498,N_195,In_1663);
xnor U2499 (N_2499,In_189,N_1438);
xor U2500 (N_2500,In_2164,N_1336);
or U2501 (N_2501,N_1744,In_3853);
xnor U2502 (N_2502,N_1924,In_771);
and U2503 (N_2503,N_1687,In_4386);
xnor U2504 (N_2504,N_1354,In_1361);
xnor U2505 (N_2505,N_1853,N_949);
xor U2506 (N_2506,N_760,In_1400);
and U2507 (N_2507,In_4156,N_887);
nand U2508 (N_2508,N_380,In_886);
xnor U2509 (N_2509,In_4694,In_517);
xnor U2510 (N_2510,N_619,N_1669);
and U2511 (N_2511,N_53,N_325);
nor U2512 (N_2512,N_1736,N_1815);
xor U2513 (N_2513,N_1773,N_1918);
nand U2514 (N_2514,N_1769,In_4007);
xnor U2515 (N_2515,In_2219,In_3502);
nand U2516 (N_2516,N_667,N_1494);
and U2517 (N_2517,N_157,N_1778);
nand U2518 (N_2518,N_1867,In_981);
nor U2519 (N_2519,N_212,N_1746);
nor U2520 (N_2520,N_117,N_920);
nor U2521 (N_2521,In_836,N_1618);
xnor U2522 (N_2522,N_1931,In_4790);
and U2523 (N_2523,N_478,N_1552);
nor U2524 (N_2524,N_757,In_1567);
or U2525 (N_2525,N_1616,N_643);
or U2526 (N_2526,N_777,N_218);
nor U2527 (N_2527,N_1772,In_821);
nor U2528 (N_2528,In_1660,N_1675);
or U2529 (N_2529,N_1584,In_3250);
xor U2530 (N_2530,In_1103,N_1642);
nor U2531 (N_2531,N_1688,N_1334);
nand U2532 (N_2532,In_2724,In_1819);
xnor U2533 (N_2533,N_686,N_1138);
nand U2534 (N_2534,N_1560,N_551);
xor U2535 (N_2535,In_4160,N_1822);
or U2536 (N_2536,In_795,N_469);
nand U2537 (N_2537,N_1052,N_910);
or U2538 (N_2538,N_620,N_101);
xnor U2539 (N_2539,N_746,N_1539);
xor U2540 (N_2540,N_1949,N_596);
or U2541 (N_2541,N_762,N_1167);
or U2542 (N_2542,N_1780,N_1351);
xor U2543 (N_2543,In_3511,N_1306);
nand U2544 (N_2544,N_454,N_1412);
nor U2545 (N_2545,N_309,N_1195);
nand U2546 (N_2546,N_161,N_1465);
nand U2547 (N_2547,N_417,N_865);
nand U2548 (N_2548,In_2386,In_4181);
xnor U2549 (N_2549,N_348,N_533);
nand U2550 (N_2550,N_1083,N_308);
and U2551 (N_2551,In_1099,N_224);
or U2552 (N_2552,N_1017,N_136);
or U2553 (N_2553,N_843,N_386);
nand U2554 (N_2554,N_929,N_317);
nand U2555 (N_2555,In_3148,N_870);
or U2556 (N_2556,N_267,In_4672);
or U2557 (N_2557,N_1808,N_603);
or U2558 (N_2558,N_198,In_4556);
xnor U2559 (N_2559,In_3106,N_1841);
nor U2560 (N_2560,In_270,N_1799);
xnor U2561 (N_2561,In_3870,In_4067);
xnor U2562 (N_2562,N_1276,In_1653);
nand U2563 (N_2563,N_754,N_1217);
nand U2564 (N_2564,N_1548,In_3389);
nor U2565 (N_2565,N_1892,In_3857);
nor U2566 (N_2566,N_670,In_211);
nor U2567 (N_2567,In_3539,N_1883);
xnor U2568 (N_2568,N_172,N_890);
nor U2569 (N_2569,N_1437,In_3038);
and U2570 (N_2570,In_1857,N_208);
or U2571 (N_2571,N_48,N_65);
nand U2572 (N_2572,In_1967,N_840);
or U2573 (N_2573,N_1079,N_35);
nor U2574 (N_2574,N_1844,In_598);
xor U2575 (N_2575,N_1696,N_628);
nor U2576 (N_2576,In_1390,In_3094);
and U2577 (N_2577,N_497,N_511);
nand U2578 (N_2578,N_1756,In_3240);
xnor U2579 (N_2579,N_1700,N_125);
and U2580 (N_2580,N_1461,N_1317);
nand U2581 (N_2581,N_1463,N_1768);
xnor U2582 (N_2582,N_1326,N_464);
and U2583 (N_2583,N_440,N_467);
or U2584 (N_2584,In_4111,N_810);
or U2585 (N_2585,N_1578,N_1283);
nor U2586 (N_2586,N_187,In_4379);
nor U2587 (N_2587,N_1062,N_298);
nand U2588 (N_2588,In_4731,In_4685);
xor U2589 (N_2589,In_4204,In_4375);
nor U2590 (N_2590,N_1070,N_731);
nand U2591 (N_2591,In_3589,In_233);
or U2592 (N_2592,N_1054,In_2440);
or U2593 (N_2593,N_415,N_579);
or U2594 (N_2594,N_1009,N_190);
nor U2595 (N_2595,N_512,In_1011);
nand U2596 (N_2596,N_1796,N_1129);
xor U2597 (N_2597,N_1409,N_515);
nand U2598 (N_2598,N_1859,In_2142);
nand U2599 (N_2599,N_148,N_1787);
or U2600 (N_2600,In_3260,N_788);
and U2601 (N_2601,N_685,N_461);
nor U2602 (N_2602,In_3819,N_575);
xnor U2603 (N_2603,In_3137,N_1467);
nor U2604 (N_2604,In_4154,N_1879);
nor U2605 (N_2605,N_1821,In_647);
or U2606 (N_2606,N_993,In_3057);
and U2607 (N_2607,N_265,In_1791);
and U2608 (N_2608,N_1835,N_1376);
or U2609 (N_2609,N_1431,N_721);
or U2610 (N_2610,In_4178,N_1885);
nand U2611 (N_2611,In_4851,N_1434);
or U2612 (N_2612,N_1365,In_1342);
nor U2613 (N_2613,N_1268,In_4671);
or U2614 (N_2614,In_1382,N_327);
nand U2615 (N_2615,N_848,In_1256);
xor U2616 (N_2616,N_449,N_1312);
or U2617 (N_2617,In_1152,N_751);
nor U2618 (N_2618,N_31,N_1863);
nor U2619 (N_2619,N_377,In_3535);
nor U2620 (N_2620,In_4528,In_960);
and U2621 (N_2621,In_1532,N_1425);
and U2622 (N_2622,In_4885,N_1443);
nor U2623 (N_2623,N_1449,N_1551);
or U2624 (N_2624,N_201,In_2600);
and U2625 (N_2625,N_154,N_1031);
nand U2626 (N_2626,N_1628,N_1103);
nor U2627 (N_2627,In_3707,N_1104);
xnor U2628 (N_2628,N_307,N_936);
nor U2629 (N_2629,N_520,N_367);
nor U2630 (N_2630,In_4754,In_1630);
nor U2631 (N_2631,N_1046,N_1917);
nand U2632 (N_2632,N_1933,In_2032);
xnor U2633 (N_2633,N_1343,N_285);
or U2634 (N_2634,In_1736,In_4070);
nor U2635 (N_2635,In_3224,In_1517);
nor U2636 (N_2636,N_1998,N_614);
xor U2637 (N_2637,In_3086,N_1192);
or U2638 (N_2638,In_1811,N_1824);
xor U2639 (N_2639,N_748,N_941);
nand U2640 (N_2640,In_907,In_4433);
xor U2641 (N_2641,In_2884,N_1495);
or U2642 (N_2642,In_4311,N_1588);
xnor U2643 (N_2643,N_1460,N_1893);
xnor U2644 (N_2644,N_1842,In_4108);
nand U2645 (N_2645,N_739,In_4134);
nor U2646 (N_2646,N_1630,N_1022);
or U2647 (N_2647,N_1090,N_565);
and U2648 (N_2648,N_1761,N_1451);
or U2649 (N_2649,N_1108,N_718);
nand U2650 (N_2650,In_3991,N_713);
xor U2651 (N_2651,In_3522,N_804);
or U2652 (N_2652,In_882,N_784);
xor U2653 (N_2653,In_3373,N_877);
and U2654 (N_2654,N_184,In_2729);
xnor U2655 (N_2655,N_1405,In_392);
or U2656 (N_2656,N_1510,N_124);
and U2657 (N_2657,N_1906,N_401);
or U2658 (N_2658,N_1954,In_2941);
or U2659 (N_2659,N_602,In_2989);
nor U2660 (N_2660,N_326,N_263);
xnor U2661 (N_2661,N_142,In_3558);
xor U2662 (N_2662,N_535,N_836);
and U2663 (N_2663,In_4284,N_1183);
xor U2664 (N_2664,N_1743,N_1785);
xnor U2665 (N_2665,N_928,N_798);
and U2666 (N_2666,N_1251,N_1341);
xnor U2667 (N_2667,N_1261,In_1622);
and U2668 (N_2668,N_1941,In_4212);
and U2669 (N_2669,In_1909,In_755);
nand U2670 (N_2670,In_3253,N_1988);
nand U2671 (N_2671,In_1894,In_92);
or U2672 (N_2672,N_1058,N_1811);
and U2673 (N_2673,N_1996,N_430);
and U2674 (N_2674,N_759,N_52);
or U2675 (N_2675,N_1762,N_811);
and U2676 (N_2676,N_223,N_1782);
nand U2677 (N_2677,N_1684,N_253);
xnor U2678 (N_2678,N_1047,In_2945);
and U2679 (N_2679,N_1021,N_284);
and U2680 (N_2680,N_1368,In_2481);
nand U2681 (N_2681,N_1302,N_857);
or U2682 (N_2682,N_741,N_539);
nor U2683 (N_2683,In_3566,N_32);
nor U2684 (N_2684,In_532,In_2686);
nand U2685 (N_2685,N_1305,N_1579);
xor U2686 (N_2686,In_2288,In_2364);
xnor U2687 (N_2687,N_182,N_671);
and U2688 (N_2688,N_749,N_1636);
xnor U2689 (N_2689,N_1100,N_1020);
nor U2690 (N_2690,In_3045,In_4848);
nand U2691 (N_2691,N_1721,N_4);
and U2692 (N_2692,In_1808,N_1791);
xor U2693 (N_2693,N_689,N_1426);
nor U2694 (N_2694,In_1508,N_1323);
nand U2695 (N_2695,In_4622,N_413);
and U2696 (N_2696,N_1940,N_243);
and U2697 (N_2697,N_1383,N_1055);
and U2698 (N_2698,N_1131,In_3609);
nor U2699 (N_2699,N_1288,In_91);
or U2700 (N_2700,In_490,In_3601);
xnor U2701 (N_2701,N_571,N_1213);
nor U2702 (N_2702,N_1569,N_1914);
xor U2703 (N_2703,In_857,In_1242);
and U2704 (N_2704,N_1327,N_1828);
and U2705 (N_2705,N_1179,N_1489);
or U2706 (N_2706,In_1680,In_1582);
xor U2707 (N_2707,N_472,N_1162);
or U2708 (N_2708,N_56,N_82);
nor U2709 (N_2709,N_70,N_414);
or U2710 (N_2710,N_1199,N_1478);
xor U2711 (N_2711,N_1480,N_442);
or U2712 (N_2712,In_3560,N_1388);
xnor U2713 (N_2713,N_411,N_296);
or U2714 (N_2714,N_452,In_412);
xor U2715 (N_2715,N_636,N_1592);
and U2716 (N_2716,N_806,N_1184);
nor U2717 (N_2717,N_36,In_4649);
nor U2718 (N_2718,N_1877,N_1475);
or U2719 (N_2719,N_549,N_122);
or U2720 (N_2720,N_907,N_213);
nor U2721 (N_2721,N_654,In_152);
and U2722 (N_2722,N_1839,In_4568);
or U2723 (N_2723,N_384,In_2791);
or U2724 (N_2724,N_587,In_4398);
xor U2725 (N_2725,In_3936,In_3330);
or U2726 (N_2726,N_1298,N_1524);
or U2727 (N_2727,N_1971,N_1823);
nand U2728 (N_2728,N_637,In_711);
xnor U2729 (N_2729,N_969,N_15);
nand U2730 (N_2730,In_4691,N_1720);
xor U2731 (N_2731,N_393,N_1800);
nand U2732 (N_2732,N_1378,N_189);
nor U2733 (N_2733,N_1137,N_1228);
xor U2734 (N_2734,In_2216,N_1264);
or U2735 (N_2735,N_1497,In_1879);
nand U2736 (N_2736,In_252,In_3241);
or U2737 (N_2737,N_776,N_650);
nand U2738 (N_2738,N_895,In_3928);
xnor U2739 (N_2739,In_993,N_231);
nand U2740 (N_2740,In_3694,N_192);
nor U2741 (N_2741,N_1254,In_1343);
nand U2742 (N_2742,In_2367,N_1587);
or U2743 (N_2743,N_481,In_31);
or U2744 (N_2744,N_1419,In_734);
and U2745 (N_2745,In_1885,N_1456);
and U2746 (N_2746,N_109,N_1939);
xnor U2747 (N_2747,N_822,N_1123);
nor U2748 (N_2748,In_754,N_1348);
and U2749 (N_2749,In_2469,In_3457);
and U2750 (N_2750,N_594,In_1522);
nand U2751 (N_2751,N_717,In_3565);
nand U2752 (N_2752,In_3600,In_4417);
nor U2753 (N_2753,In_2834,In_4616);
nand U2754 (N_2754,N_658,In_1874);
or U2755 (N_2755,N_476,N_203);
xor U2756 (N_2756,N_1191,N_426);
or U2757 (N_2757,In_372,N_979);
xor U2758 (N_2758,In_3531,In_801);
xnor U2759 (N_2759,In_820,N_1091);
and U2760 (N_2760,In_3861,N_913);
nand U2761 (N_2761,N_742,N_773);
nand U2762 (N_2762,N_169,N_756);
nand U2763 (N_2763,N_74,N_1112);
or U2764 (N_2764,In_1877,N_1657);
and U2765 (N_2765,In_1473,N_1322);
or U2766 (N_2766,N_1577,N_1726);
nor U2767 (N_2767,N_1802,N_677);
nor U2768 (N_2768,In_3120,In_4618);
xor U2769 (N_2769,N_1776,N_876);
nor U2770 (N_2770,In_1423,N_295);
nor U2771 (N_2771,N_601,In_4880);
or U2772 (N_2772,In_3062,N_1156);
nand U2773 (N_2773,N_1147,N_383);
nand U2774 (N_2774,N_1349,N_1139);
or U2775 (N_2775,N_1234,N_186);
and U2776 (N_2776,N_916,N_629);
and U2777 (N_2777,In_2430,N_1064);
and U2778 (N_2778,N_333,In_3655);
nor U2779 (N_2779,N_800,In_956);
nand U2780 (N_2780,N_1428,N_64);
xor U2781 (N_2781,N_1120,In_2817);
nand U2782 (N_2782,N_1211,N_1518);
or U2783 (N_2783,N_626,In_4227);
and U2784 (N_2784,N_373,N_1332);
and U2785 (N_2785,In_3973,In_635);
nor U2786 (N_2786,N_524,In_1852);
and U2787 (N_2787,N_301,In_1074);
nor U2788 (N_2788,In_1171,N_740);
nor U2789 (N_2789,N_310,N_128);
and U2790 (N_2790,N_1740,N_926);
or U2791 (N_2791,N_423,N_97);
nor U2792 (N_2792,N_908,N_1582);
xor U2793 (N_2793,N_1225,N_1275);
and U2794 (N_2794,N_395,N_1488);
nand U2795 (N_2795,N_850,N_444);
nor U2796 (N_2796,In_4785,N_1999);
xnor U2797 (N_2797,N_1735,In_1945);
nor U2798 (N_2798,N_314,In_3375);
and U2799 (N_2799,N_299,In_2944);
nor U2800 (N_2800,N_984,In_1492);
nand U2801 (N_2801,In_1529,N_1074);
nand U2802 (N_2802,N_707,N_102);
nand U2803 (N_2803,In_2998,In_1118);
and U2804 (N_2804,In_1946,N_87);
and U2805 (N_2805,N_1623,N_1690);
or U2806 (N_2806,N_1896,N_1591);
and U2807 (N_2807,N_127,N_661);
or U2808 (N_2808,N_541,N_149);
and U2809 (N_2809,N_1622,N_194);
nand U2810 (N_2810,In_1512,In_824);
nor U2811 (N_2811,In_2004,N_1502);
nand U2812 (N_2812,N_42,In_1604);
or U2813 (N_2813,In_629,N_655);
nand U2814 (N_2814,N_324,N_513);
or U2815 (N_2815,N_1446,In_1988);
xnor U2816 (N_2816,In_2759,In_3673);
xor U2817 (N_2817,N_1042,N_778);
or U2818 (N_2818,In_3828,N_1466);
or U2819 (N_2819,In_11,N_1205);
and U2820 (N_2820,N_1263,N_786);
or U2821 (N_2821,In_3845,In_4999);
and U2822 (N_2822,N_1331,N_630);
or U2823 (N_2823,N_546,N_342);
and U2824 (N_2824,N_930,N_1911);
nor U2825 (N_2825,In_839,In_3651);
xnor U2826 (N_2826,N_103,N_1086);
or U2827 (N_2827,N_1603,N_977);
xnor U2828 (N_2828,N_943,N_1347);
xor U2829 (N_2829,N_1385,In_2967);
nor U2830 (N_2830,N_1660,N_1281);
and U2831 (N_2831,N_938,In_3242);
xor U2832 (N_2832,N_1813,N_871);
and U2833 (N_2833,In_1789,N_468);
nand U2834 (N_2834,N_33,N_1658);
xnor U2835 (N_2835,In_2881,N_0);
nor U2836 (N_2836,In_436,In_4538);
nand U2837 (N_2837,N_358,In_661);
or U2838 (N_2838,N_1389,In_1438);
nand U2839 (N_2839,In_653,In_3133);
and U2840 (N_2840,N_1806,In_837);
or U2841 (N_2841,N_1253,N_341);
or U2842 (N_2842,N_134,N_99);
nand U2843 (N_2843,In_4806,N_1479);
or U2844 (N_2844,N_379,N_1445);
nand U2845 (N_2845,In_2560,N_568);
nand U2846 (N_2846,N_462,N_1154);
nor U2847 (N_2847,In_927,N_389);
xor U2848 (N_2848,N_1065,N_1415);
and U2849 (N_2849,In_3984,N_1403);
and U2850 (N_2850,N_258,N_1249);
and U2851 (N_2851,In_2831,In_4993);
or U2852 (N_2852,N_994,In_3491);
nor U2853 (N_2853,N_904,N_1504);
nor U2854 (N_2854,N_724,In_3312);
nand U2855 (N_2855,N_1818,N_1304);
nand U2856 (N_2856,In_14,In_4167);
nor U2857 (N_2857,In_1381,In_1554);
nand U2858 (N_2858,In_3361,N_483);
xor U2859 (N_2859,N_891,N_494);
and U2860 (N_2860,In_214,N_1018);
nand U2861 (N_2861,In_2650,N_1170);
nor U2862 (N_2862,In_848,In_388);
nor U2863 (N_2863,In_3935,N_957);
or U2864 (N_2864,In_237,N_1145);
nor U2865 (N_2865,In_671,N_983);
nand U2866 (N_2866,In_295,In_1200);
or U2867 (N_2867,N_1927,N_457);
and U2868 (N_2868,N_1416,In_3526);
xnor U2869 (N_2869,N_582,N_1360);
xnor U2870 (N_2870,N_396,N_1757);
nor U2871 (N_2871,In_987,N_1535);
nor U2872 (N_2872,N_982,N_1427);
nand U2873 (N_2873,N_18,In_2349);
nand U2874 (N_2874,N_732,N_1804);
xnor U2875 (N_2875,N_439,In_4604);
or U2876 (N_2876,N_1869,N_1088);
and U2877 (N_2877,In_3964,N_923);
or U2878 (N_2878,N_1837,N_277);
and U2879 (N_2879,In_3904,N_1609);
nand U2880 (N_2880,N_1874,N_1970);
nand U2881 (N_2881,In_1183,N_1742);
or U2882 (N_2882,N_1273,N_593);
xnor U2883 (N_2883,In_3216,In_2062);
xor U2884 (N_2884,N_1595,N_1809);
nand U2885 (N_2885,N_50,N_1374);
xor U2886 (N_2886,N_1126,In_4623);
nand U2887 (N_2887,In_3905,In_3581);
and U2888 (N_2888,N_1697,N_1406);
or U2889 (N_2889,In_3731,In_1639);
or U2890 (N_2890,N_1499,N_1717);
nand U2891 (N_2891,N_447,N_156);
nand U2892 (N_2892,N_185,N_1115);
nand U2893 (N_2893,In_2537,N_416);
nor U2894 (N_2894,N_1227,In_4951);
xor U2895 (N_2895,In_4605,N_752);
or U2896 (N_2896,N_1266,N_885);
nand U2897 (N_2897,N_1948,N_104);
xor U2898 (N_2898,N_727,In_1650);
or U2899 (N_2899,N_1318,N_1534);
nor U2900 (N_2900,N_63,In_2300);
or U2901 (N_2901,In_77,In_4724);
nand U2902 (N_2902,N_613,In_232);
xor U2903 (N_2903,N_196,N_1208);
nor U2904 (N_2904,N_1330,N_1068);
xor U2905 (N_2905,In_1989,N_1686);
or U2906 (N_2906,N_968,N_62);
and U2907 (N_2907,N_1454,N_1379);
xor U2908 (N_2908,N_1920,N_853);
nand U2909 (N_2909,N_1648,N_824);
nand U2910 (N_2910,In_4472,In_550);
or U2911 (N_2911,In_4978,N_573);
or U2912 (N_2912,N_1937,In_453);
xor U2913 (N_2913,N_1749,N_1635);
or U2914 (N_2914,N_89,N_1722);
or U2915 (N_2915,N_1529,In_2818);
nand U2916 (N_2916,In_4464,N_207);
or U2917 (N_2917,In_1618,In_181);
xor U2918 (N_2918,N_1043,N_1890);
or U2919 (N_2919,N_1644,In_3016);
and U2920 (N_2920,N_1398,N_559);
or U2921 (N_2921,N_1498,In_1339);
or U2922 (N_2922,N_1832,In_1123);
and U2923 (N_2923,N_387,In_4697);
nor U2924 (N_2924,N_343,N_782);
nand U2925 (N_2925,N_292,In_646);
and U2926 (N_2926,In_1368,N_507);
and U2927 (N_2927,N_1301,N_1168);
xnor U2928 (N_2928,In_3596,N_390);
nand U2929 (N_2929,In_241,In_4668);
or U2930 (N_2930,N_121,In_610);
nand U2931 (N_2931,N_363,In_1150);
xor U2932 (N_2932,In_401,N_605);
and U2933 (N_2933,N_1164,N_911);
or U2934 (N_2934,N_388,N_1624);
and U2935 (N_2935,N_1871,N_1084);
xnor U2936 (N_2936,In_2026,In_804);
xnor U2937 (N_2937,N_768,N_899);
and U2938 (N_2938,N_1654,N_719);
or U2939 (N_2939,In_2096,In_4374);
and U2940 (N_2940,In_2846,N_330);
and U2941 (N_2941,N_1371,N_404);
and U2942 (N_2942,N_989,In_2120);
xor U2943 (N_2943,N_829,N_1484);
nand U2944 (N_2944,N_1709,In_3873);
and U2945 (N_2945,N_1232,N_914);
nand U2946 (N_2946,In_2569,N_120);
or U2947 (N_2947,In_2720,In_590);
xor U2948 (N_2948,N_532,N_1171);
xor U2949 (N_2949,N_1829,N_41);
xnor U2950 (N_2950,N_1430,N_1157);
nand U2951 (N_2951,In_2162,In_4558);
or U2952 (N_2952,In_1673,In_2371);
xnor U2953 (N_2953,N_1113,N_30);
nor U2954 (N_2954,N_1159,In_3025);
nor U2955 (N_2955,N_424,N_81);
xor U2956 (N_2956,N_1753,N_290);
nand U2957 (N_2957,N_408,N_451);
or U2958 (N_2958,N_1033,In_3685);
and U2959 (N_2959,N_1282,In_3091);
nand U2960 (N_2960,N_246,N_1555);
nand U2961 (N_2961,In_2186,In_900);
xnor U2962 (N_2962,N_1990,N_525);
nand U2963 (N_2963,In_4078,N_1161);
nand U2964 (N_2964,N_1280,N_1723);
xnor U2965 (N_2965,N_1142,In_3580);
and U2966 (N_2966,N_710,In_4075);
nand U2967 (N_2967,N_1699,N_1128);
nor U2968 (N_2968,N_436,In_2905);
or U2969 (N_2969,In_4817,N_1607);
or U2970 (N_2970,N_1750,N_550);
or U2971 (N_2971,In_1761,N_862);
nor U2972 (N_2972,N_1250,In_4737);
nor U2973 (N_2973,N_530,N_306);
and U2974 (N_2974,In_1968,In_615);
nand U2975 (N_2975,N_427,N_1222);
xor U2976 (N_2976,N_1710,N_1380);
or U2977 (N_2977,In_1112,N_1324);
and U2978 (N_2978,N_1291,N_366);
or U2979 (N_2979,N_1034,In_331);
or U2980 (N_2980,N_813,N_1594);
or U2981 (N_2981,In_3394,N_347);
or U2982 (N_2982,In_1442,N_558);
nand U2983 (N_2983,N_1230,N_1708);
nand U2984 (N_2984,N_6,N_1652);
nor U2985 (N_2985,N_412,In_2926);
and U2986 (N_2986,N_924,N_1943);
and U2987 (N_2987,In_2455,N_1407);
and U2988 (N_2988,In_2804,N_1963);
nand U2989 (N_2989,N_86,N_728);
xnor U2990 (N_2990,N_1279,In_3682);
nor U2991 (N_2991,In_2606,In_4509);
and U2992 (N_2992,N_1216,N_1390);
and U2993 (N_2993,In_4512,In_2800);
xor U2994 (N_2994,N_785,N_1309);
nor U2995 (N_2995,In_2744,In_603);
and U2996 (N_2996,N_150,N_1248);
or U2997 (N_2997,N_77,N_170);
xnor U2998 (N_2998,N_1803,In_1750);
or U2999 (N_2999,In_2153,In_2377);
and U3000 (N_3000,N_1864,N_256);
nor U3001 (N_3001,In_1494,N_1783);
nor U3002 (N_3002,N_516,In_3317);
or U3003 (N_3003,N_1549,In_786);
xor U3004 (N_3004,In_4256,N_683);
and U3005 (N_3005,In_1142,In_4082);
or U3006 (N_3006,N_1665,N_275);
xnor U3007 (N_3007,N_455,N_919);
nand U3008 (N_3008,N_1792,In_201);
xnor U3009 (N_3009,In_1905,In_3360);
or U3010 (N_3010,N_1593,In_1295);
or U3011 (N_3011,N_328,N_827);
and U3012 (N_3012,In_4748,In_1719);
or U3013 (N_3013,N_286,N_961);
nor U3014 (N_3014,In_2124,N_54);
nand U3015 (N_3015,N_684,N_1573);
and U3016 (N_3016,N_450,N_1193);
or U3017 (N_3017,N_527,N_1338);
or U3018 (N_3018,N_893,In_1007);
or U3019 (N_3019,N_1094,N_458);
nor U3020 (N_3020,In_1330,N_1352);
and U3021 (N_3021,In_384,N_640);
xor U3022 (N_3022,N_1926,N_233);
xor U3023 (N_3023,In_2086,N_878);
xnor U3024 (N_3024,N_744,N_421);
or U3025 (N_3025,N_216,N_729);
xnor U3026 (N_3026,N_1674,In_1079);
and U3027 (N_3027,N_1134,N_1001);
or U3028 (N_3028,N_71,N_1747);
or U3029 (N_3029,In_3507,N_59);
nor U3030 (N_3030,In_2416,In_1725);
nand U3031 (N_3031,N_1258,In_165);
xnor U3032 (N_3032,In_1524,N_723);
or U3033 (N_3033,N_660,N_1583);
nor U3034 (N_3034,N_1748,N_1712);
xor U3035 (N_3035,N_498,N_985);
nor U3036 (N_3036,In_2012,N_84);
or U3037 (N_3037,N_818,N_1527);
nor U3038 (N_3038,In_1716,N_1627);
and U3039 (N_3039,In_4248,In_4333);
xnor U3040 (N_3040,N_1850,In_4807);
and U3041 (N_3041,N_1218,N_1559);
nand U3042 (N_3042,In_2699,In_3689);
xor U3043 (N_3043,N_1543,N_460);
nor U3044 (N_3044,N_808,In_167);
nand U3045 (N_3045,N_510,N_1987);
nand U3046 (N_3046,N_214,N_1391);
nand U3047 (N_3047,N_1158,N_1507);
or U3048 (N_3048,N_1910,N_1767);
or U3049 (N_3049,In_748,N_1150);
and U3050 (N_3050,In_978,N_965);
or U3051 (N_3051,N_1358,In_2334);
or U3052 (N_3052,In_3047,In_1959);
nor U3053 (N_3053,N_1295,N_638);
xnor U3054 (N_3054,N_548,N_1160);
and U3055 (N_3055,N_1190,N_702);
or U3056 (N_3056,In_3974,In_2702);
or U3057 (N_3057,N_1725,In_418);
and U3058 (N_3058,N_22,N_1777);
nor U3059 (N_3059,In_2824,N_781);
nand U3060 (N_3060,In_2093,In_4414);
and U3061 (N_3061,N_1606,N_1386);
and U3062 (N_3062,In_4221,N_1732);
or U3063 (N_3063,N_1292,In_583);
nand U3064 (N_3064,In_4443,In_4000);
nor U3065 (N_3065,In_4058,N_1528);
or U3066 (N_3066,N_1678,In_1574);
and U3067 (N_3067,In_1131,N_1706);
or U3068 (N_3068,N_1402,N_336);
nand U3069 (N_3069,N_135,In_1624);
nor U3070 (N_3070,In_351,In_584);
or U3071 (N_3071,N_1257,N_106);
nor U3072 (N_3072,In_4801,N_271);
nand U3073 (N_3073,In_2122,In_3092);
xnor U3074 (N_3074,In_4110,In_2108);
nor U3075 (N_3075,In_1853,N_1574);
or U3076 (N_3076,N_1392,N_693);
nor U3077 (N_3077,In_867,In_1);
nand U3078 (N_3078,N_1522,In_72);
nor U3079 (N_3079,N_1974,In_2315);
or U3080 (N_3080,N_706,N_493);
nor U3081 (N_3081,N_569,N_866);
nand U3082 (N_3082,In_1166,N_1048);
and U3083 (N_3083,N_181,In_3656);
xor U3084 (N_3084,In_1569,N_260);
or U3085 (N_3085,In_2507,In_4054);
nand U3086 (N_3086,N_774,In_1579);
xnor U3087 (N_3087,In_2538,N_1455);
and U3088 (N_3088,N_1900,N_475);
nand U3089 (N_3089,In_3090,In_1631);
xor U3090 (N_3090,N_1886,N_1964);
nand U3091 (N_3091,N_803,In_410);
nor U3092 (N_3092,In_4420,In_4881);
nor U3093 (N_3093,N_976,N_543);
and U3094 (N_3094,N_986,N_1526);
xnor U3095 (N_3095,In_3799,N_143);
and U3096 (N_3096,N_1958,N_1605);
xor U3097 (N_3097,In_1715,In_885);
nand U3098 (N_3098,N_1938,N_522);
or U3099 (N_3099,In_518,N_1152);
nand U3100 (N_3100,N_1224,In_3077);
xor U3101 (N_3101,In_2147,N_248);
nand U3102 (N_3102,In_4823,N_16);
nand U3103 (N_3103,N_1625,N_1564);
nor U3104 (N_3104,In_1129,N_980);
nand U3105 (N_3105,In_238,In_22);
nand U3106 (N_3106,N_1985,In_1162);
nand U3107 (N_3107,N_375,In_4296);
nor U3108 (N_3108,In_1067,N_931);
nand U3109 (N_3109,In_2361,N_1198);
or U3110 (N_3110,N_1078,N_178);
and U3111 (N_3111,In_1890,N_1969);
nand U3112 (N_3112,In_2489,N_1244);
nor U3113 (N_3113,N_714,N_1962);
or U3114 (N_3114,N_988,N_255);
xor U3115 (N_3115,N_1328,N_167);
or U3116 (N_3116,N_1477,In_2158);
nand U3117 (N_3117,N_1880,N_1805);
nand U3118 (N_3118,N_8,N_1346);
or U3119 (N_3119,N_193,In_352);
xnor U3120 (N_3120,N_622,N_1375);
or U3121 (N_3121,N_1563,In_332);
nand U3122 (N_3122,N_435,In_3591);
nand U3123 (N_3123,In_1239,N_697);
xnor U3124 (N_3124,In_4367,N_276);
nand U3125 (N_3125,In_3815,N_1053);
nor U3126 (N_3126,N_1986,N_1069);
xor U3127 (N_3127,In_4370,In_272);
xnor U3128 (N_3128,N_1015,N_1536);
and U3129 (N_3129,N_897,In_758);
or U3130 (N_3130,N_1310,N_1997);
xor U3131 (N_3131,N_1366,In_3376);
and U3132 (N_3132,In_441,N_39);
or U3133 (N_3133,N_332,N_1202);
nor U3134 (N_3134,N_228,In_1975);
xor U3135 (N_3135,In_1322,N_1807);
xor U3136 (N_3136,N_561,N_1617);
nor U3137 (N_3137,N_1102,N_915);
xor U3138 (N_3138,In_3351,N_1172);
xor U3139 (N_3139,In_80,N_1629);
or U3140 (N_3140,N_73,N_501);
nand U3141 (N_3141,N_560,N_1532);
nor U3142 (N_3142,N_1677,N_1826);
xnor U3143 (N_3143,N_1106,N_268);
and U3144 (N_3144,N_482,N_604);
nand U3145 (N_3145,N_937,In_3055);
and U3146 (N_3146,N_722,In_2442);
xnor U3147 (N_3147,N_770,N_687);
or U3148 (N_3148,N_1239,In_2950);
xor U3149 (N_3149,N_792,N_356);
nor U3150 (N_3150,N_1568,N_1353);
nor U3151 (N_3151,In_1061,In_2770);
xnor U3152 (N_3152,In_576,N_863);
or U3153 (N_3153,In_4137,In_605);
or U3154 (N_3154,In_559,N_399);
xor U3155 (N_3155,N_428,N_775);
xnor U3156 (N_3156,In_2748,N_1476);
or U3157 (N_3157,N_1957,In_3346);
nor U3158 (N_3158,In_1465,N_155);
nor U3159 (N_3159,N_1121,In_1317);
nor U3160 (N_3160,N_939,In_3328);
or U3161 (N_3161,N_1483,In_805);
xor U3162 (N_3162,N_1095,N_991);
and U3163 (N_3163,In_478,N_1207);
nand U3164 (N_3164,N_635,In_4400);
xor U3165 (N_3165,N_1039,N_1501);
nor U3166 (N_3166,N_508,N_711);
xor U3167 (N_3167,N_1521,In_1439);
nor U3168 (N_3168,N_491,N_839);
nor U3169 (N_3169,In_3524,In_2066);
or U3170 (N_3170,In_3256,N_1865);
and U3171 (N_3171,N_617,In_1248);
nand U3172 (N_3172,In_3647,In_3939);
and U3173 (N_3173,In_4241,N_1027);
nand U3174 (N_3174,N_1928,N_432);
nand U3175 (N_3175,N_339,In_2199);
xnor U3176 (N_3176,N_1470,In_2305);
xnor U3177 (N_3177,In_2175,N_1245);
nand U3178 (N_3178,In_1779,N_680);
xor U3179 (N_3179,N_1781,N_1370);
and U3180 (N_3180,N_1429,N_1056);
nor U3181 (N_3181,N_1639,N_868);
nor U3182 (N_3182,N_990,In_3726);
xor U3183 (N_3183,In_4225,N_247);
nand U3184 (N_3184,N_1377,N_130);
nor U3185 (N_3185,N_11,In_3821);
xnor U3186 (N_3186,In_1078,N_1464);
nand U3187 (N_3187,N_846,In_4024);
or U3188 (N_3188,N_95,In_4900);
xnor U3189 (N_3189,N_288,In_3654);
or U3190 (N_3190,In_1530,N_552);
nand U3191 (N_3191,N_1861,N_1296);
or U3192 (N_3192,N_340,N_1770);
nor U3193 (N_3193,N_487,In_1136);
nand U3194 (N_3194,In_83,In_4037);
or U3195 (N_3195,N_1946,N_371);
or U3196 (N_3196,N_1668,N_538);
nor U3197 (N_3197,N_1664,N_1297);
and U3198 (N_3198,N_801,N_902);
xor U3199 (N_3199,In_2128,In_2344);
nor U3200 (N_3200,N_583,In_1426);
and U3201 (N_3201,N_1825,N_978);
and U3202 (N_3202,In_911,N_819);
nor U3203 (N_3203,N_1887,In_2648);
and U3204 (N_3204,N_1831,N_225);
xnor U3205 (N_3205,In_4595,N_644);
nand U3206 (N_3206,N_763,N_1945);
and U3207 (N_3207,In_2815,N_1214);
nor U3208 (N_3208,N_113,N_849);
nand U3209 (N_3209,In_535,N_1868);
nand U3210 (N_3210,N_1602,In_2959);
and U3211 (N_3211,N_1252,N_567);
xor U3212 (N_3212,N_1590,N_1695);
or U3213 (N_3213,In_4882,In_3827);
xor U3214 (N_3214,N_1329,N_261);
or U3215 (N_3215,N_682,N_906);
and U3216 (N_3216,N_199,In_2904);
nand U3217 (N_3217,In_898,In_3348);
or U3218 (N_3218,N_927,In_1655);
nor U3219 (N_3219,In_322,N_681);
and U3220 (N_3220,N_1718,N_504);
xor U3221 (N_3221,In_976,In_1972);
and U3222 (N_3222,N_1793,N_1019);
nor U3223 (N_3223,N_556,N_1598);
and U3224 (N_3224,N_305,N_291);
nor U3225 (N_3225,N_3,N_1597);
and U3226 (N_3226,In_3641,N_437);
or U3227 (N_3227,N_642,N_1771);
nor U3228 (N_3228,N_133,N_1267);
nor U3229 (N_3229,In_2951,N_627);
and U3230 (N_3230,N_83,In_2179);
nand U3231 (N_3231,N_1897,N_1930);
nor U3232 (N_3232,N_1975,In_3962);
and U3233 (N_3233,N_1966,N_96);
nand U3234 (N_3234,In_617,N_146);
nand U3235 (N_3235,N_29,N_116);
xnor U3236 (N_3236,N_935,N_621);
nor U3237 (N_3237,N_1037,In_4198);
nor U3238 (N_3238,N_496,N_202);
xor U3239 (N_3239,N_1715,N_1203);
nand U3240 (N_3240,In_3484,N_1141);
nor U3241 (N_3241,N_1608,N_479);
xnor U3242 (N_3242,N_1913,N_1387);
or U3243 (N_3243,In_4610,In_301);
nor U3244 (N_3244,N_1050,N_402);
or U3245 (N_3245,N_1105,In_1759);
xor U3246 (N_3246,In_2306,In_700);
xor U3247 (N_3247,In_4215,In_3749);
and U3248 (N_3248,In_0,In_515);
nor U3249 (N_3249,N_1659,In_2498);
nand U3250 (N_3250,N_405,N_183);
xor U3251 (N_3251,N_861,In_3130);
xor U3252 (N_3252,In_4591,In_1247);
nor U3253 (N_3253,N_1764,N_1174);
nand U3254 (N_3254,N_98,N_492);
or U3255 (N_3255,In_4689,In_1605);
nor U3256 (N_3256,In_248,N_176);
or U3257 (N_3257,N_554,N_657);
or U3258 (N_3258,In_2775,N_131);
and U3259 (N_3259,In_493,In_1834);
and U3260 (N_3260,N_500,N_283);
or U3261 (N_3261,N_27,In_1420);
nor U3262 (N_3262,N_353,N_1181);
or U3263 (N_3263,N_1314,N_971);
xor U3264 (N_3264,N_179,In_3787);
xor U3265 (N_3265,N_119,N_1165);
and U3266 (N_3266,N_1508,In_663);
or U3267 (N_3267,N_163,N_1751);
nand U3268 (N_3268,N_58,In_3179);
nand U3269 (N_3269,In_923,N_1359);
nand U3270 (N_3270,N_138,N_1004);
xnor U3271 (N_3271,N_1119,In_2714);
nor U3272 (N_3272,N_1459,N_1981);
xnor U3273 (N_3273,N_771,N_118);
xor U3274 (N_3274,N_1889,N_547);
nand U3275 (N_3275,N_666,In_3528);
nand U3276 (N_3276,N_1576,N_625);
nor U3277 (N_3277,N_519,N_360);
or U3278 (N_3278,N_509,N_1026);
nand U3279 (N_3279,In_1030,In_4274);
and U3280 (N_3280,In_521,N_463);
and U3281 (N_3281,N_881,N_422);
nand U3282 (N_3282,N_1925,In_1266);
nand U3283 (N_3283,N_1798,In_3884);
xnor U3284 (N_3284,N_235,N_335);
and U3285 (N_3285,N_1903,N_992);
or U3286 (N_3286,In_2381,In_658);
and U3287 (N_3287,In_98,In_323);
and U3288 (N_3288,N_1854,In_506);
and U3289 (N_3289,N_374,N_581);
nor U3290 (N_3290,N_75,N_1984);
nand U3291 (N_3291,In_3956,N_352);
or U3292 (N_3292,N_1293,N_612);
nand U3293 (N_3293,N_1856,N_652);
nor U3294 (N_3294,In_1463,In_4462);
or U3295 (N_3295,N_334,N_649);
and U3296 (N_3296,N_368,N_1967);
nor U3297 (N_3297,N_780,N_1904);
and U3298 (N_3298,In_1133,N_1651);
nand U3299 (N_3299,N_311,N_1356);
nand U3300 (N_3300,N_21,In_439);
nand U3301 (N_3301,N_945,In_1315);
nand U3302 (N_3302,In_997,N_673);
nor U3303 (N_3303,In_1587,N_144);
nand U3304 (N_3304,N_529,N_37);
nor U3305 (N_3305,N_940,N_1316);
nor U3306 (N_3306,In_4530,In_479);
or U3307 (N_3307,In_874,N_1703);
xnor U3308 (N_3308,In_2140,In_768);
and U3309 (N_3309,N_606,In_1154);
or U3310 (N_3310,N_1641,N_946);
or U3311 (N_3311,N_1194,N_484);
or U3312 (N_3312,In_1839,N_699);
nor U3313 (N_3313,In_2376,N_688);
and U3314 (N_3314,In_1792,N_403);
nand U3315 (N_3315,N_480,N_385);
nor U3316 (N_3316,In_955,N_1294);
xnor U3317 (N_3317,N_1397,In_4175);
nand U3318 (N_3318,N_239,In_4789);
xnor U3319 (N_3319,In_44,In_4392);
xnor U3320 (N_3320,N_1362,In_3519);
nor U3321 (N_3321,In_367,In_1415);
xnor U3322 (N_3322,In_2233,N_1929);
nand U3323 (N_3323,In_136,N_257);
or U3324 (N_3324,N_158,N_918);
nor U3325 (N_3325,N_1758,In_4651);
and U3326 (N_3326,N_1571,N_796);
nor U3327 (N_3327,N_466,N_1565);
nor U3328 (N_3328,N_1766,N_1852);
nor U3329 (N_3329,In_4532,N_1965);
nand U3330 (N_3330,N_599,N_1148);
or U3331 (N_3331,In_3869,In_2159);
nor U3332 (N_3332,In_2588,In_2854);
nor U3333 (N_3333,In_1816,In_4088);
nor U3334 (N_3334,N_376,In_1264);
nor U3335 (N_3335,N_1400,N_1952);
and U3336 (N_3336,N_1473,In_3018);
and U3337 (N_3337,N_108,In_2528);
xor U3338 (N_3338,In_1537,In_1803);
or U3339 (N_3339,N_471,N_293);
nor U3340 (N_3340,N_564,N_1878);
or U3341 (N_3341,N_1410,N_1833);
and U3342 (N_3342,In_2763,N_1942);
or U3343 (N_3343,N_1775,In_3386);
nand U3344 (N_3344,N_598,N_1411);
nor U3345 (N_3345,N_1834,N_188);
xnor U3346 (N_3346,In_627,N_1694);
and U3347 (N_3347,N_294,N_1666);
or U3348 (N_3348,N_860,N_799);
and U3349 (N_3349,N_1003,N_1030);
xor U3350 (N_3350,In_1184,N_1023);
xnor U3351 (N_3351,In_2178,N_1553);
nor U3352 (N_3352,N_1705,N_17);
xnor U3353 (N_3353,N_1795,N_1820);
nor U3354 (N_3354,In_3603,In_3417);
xnor U3355 (N_3355,N_354,In_2040);
or U3356 (N_3356,N_1907,N_438);
and U3357 (N_3357,N_954,N_1698);
nand U3358 (N_3358,N_960,N_230);
and U3359 (N_3359,In_1178,N_802);
nor U3360 (N_3360,N_1133,In_3716);
or U3361 (N_3361,N_963,N_514);
and U3362 (N_3362,In_2601,N_323);
xor U3363 (N_3363,In_1277,N_165);
nor U3364 (N_3364,In_2117,N_346);
or U3365 (N_3365,N_215,N_264);
xnor U3366 (N_3366,N_528,In_1000);
nor U3367 (N_3367,In_4583,In_3908);
xor U3368 (N_3368,N_66,N_241);
xor U3369 (N_3369,In_3085,In_4696);
xor U3370 (N_3370,In_1270,N_107);
or U3371 (N_3371,N_280,N_473);
xor U3372 (N_3372,N_173,N_470);
or U3373 (N_3373,In_4079,In_2485);
or U3374 (N_3374,N_1229,N_1175);
nor U3375 (N_3375,In_3411,In_4312);
and U3376 (N_3376,In_3518,N_1116);
nor U3377 (N_3377,In_1221,In_492);
xnor U3378 (N_3378,N_1333,N_1845);
nand U3379 (N_3379,N_807,N_1516);
nor U3380 (N_3380,N_359,N_445);
xnor U3381 (N_3381,N_835,In_593);
xor U3382 (N_3382,N_678,N_734);
and U3383 (N_3383,N_152,In_440);
nor U3384 (N_3384,N_1848,N_1384);
nand U3385 (N_3385,N_616,N_1947);
nor U3386 (N_3386,In_4135,N_1189);
nor U3387 (N_3387,N_1763,N_1320);
nor U3388 (N_3388,In_3582,N_1038);
or U3389 (N_3389,N_1955,N_392);
nor U3390 (N_3390,N_1417,N_1790);
or U3391 (N_3391,N_1122,N_1186);
or U3392 (N_3392,In_1034,In_869);
xor U3393 (N_3393,N_970,N_709);
and U3394 (N_3394,In_728,N_589);
nand U3395 (N_3395,N_772,N_505);
and U3396 (N_3396,In_3721,N_382);
xnor U3397 (N_3397,N_1862,In_2921);
xnor U3398 (N_3398,N_1789,N_659);
and U3399 (N_3399,N_1714,N_855);
and U3400 (N_3400,In_1157,N_767);
nor U3401 (N_3401,N_764,N_623);
and U3402 (N_3402,N_610,N_1566);
xor U3403 (N_3403,N_703,N_1313);
or U3404 (N_3404,In_306,In_1181);
nor U3405 (N_3405,N_1073,N_38);
and U3406 (N_3406,N_1934,N_274);
and U3407 (N_3407,N_745,N_456);
nand U3408 (N_3408,N_668,In_2487);
or U3409 (N_3409,In_2204,N_634);
nor U3410 (N_3410,N_1081,In_1838);
or U3411 (N_3411,N_1246,N_495);
nand U3412 (N_3412,N_820,N_126);
nand U3413 (N_3413,In_3425,N_1107);
or U3414 (N_3414,N_1619,N_1);
nand U3415 (N_3415,In_3189,N_205);
xnor U3416 (N_3416,N_1830,N_966);
and U3417 (N_3417,In_2575,In_390);
nor U3418 (N_3418,N_1111,In_3434);
nor U3419 (N_3419,N_834,In_4474);
nor U3420 (N_3420,In_1276,In_4074);
or U3421 (N_3421,In_52,N_321);
nand U3422 (N_3422,N_1140,N_1637);
nor U3423 (N_3423,N_453,N_55);
and U3424 (N_3424,N_1724,In_4476);
nand U3425 (N_3425,N_365,In_282);
and U3426 (N_3426,N_1024,N_873);
nor U3427 (N_3427,N_43,In_3272);
nand U3428 (N_3428,N_110,In_4029);
xor U3429 (N_3429,N_588,N_998);
nor U3430 (N_3430,N_1734,N_1401);
nor U3431 (N_3431,N_735,N_791);
xor U3432 (N_3432,N_57,In_3537);
xnor U3433 (N_3433,In_958,N_691);
nor U3434 (N_3434,In_3145,N_1413);
and U3435 (N_3435,In_3922,In_2101);
or U3436 (N_3436,N_662,N_397);
nor U3437 (N_3437,N_1755,N_1259);
or U3438 (N_3438,In_4845,N_578);
nand U3439 (N_3439,N_690,In_3235);
xnor U3440 (N_3440,N_708,N_237);
nor U3441 (N_3441,In_571,In_3455);
nand U3442 (N_3442,In_1694,N_1994);
xnor U3443 (N_3443,N_78,N_1550);
xnor U3444 (N_3444,N_1051,N_1496);
nor U3445 (N_3445,N_823,In_1232);
and U3446 (N_3446,In_693,N_952);
and U3447 (N_3447,N_1545,N_61);
or U3448 (N_3448,In_698,In_1980);
nor U3449 (N_3449,N_1953,In_2912);
nor U3450 (N_3450,In_4892,N_1007);
nand U3451 (N_3451,N_1902,N_1180);
nor U3452 (N_3452,N_1005,In_2113);
or U3453 (N_3453,N_1240,N_338);
nor U3454 (N_3454,In_736,In_3214);
nand U3455 (N_3455,In_3323,N_631);
and U3456 (N_3456,N_164,N_815);
nand U3457 (N_3457,N_632,In_4752);
nor U3458 (N_3458,N_1096,N_747);
nand U3459 (N_3459,N_607,N_1182);
or U3460 (N_3460,N_1517,N_1209);
nand U3461 (N_3461,N_304,N_1092);
nand U3462 (N_3462,In_3218,N_755);
and U3463 (N_3463,N_1977,N_1935);
xnor U3464 (N_3464,N_716,In_1484);
and U3465 (N_3465,N_1993,N_145);
and U3466 (N_3466,N_1277,In_1117);
xnor U3467 (N_3467,N_1851,N_1544);
or U3468 (N_3468,N_639,N_1531);
nand U3469 (N_3469,N_459,In_749);
and U3470 (N_3470,N_1951,In_2610);
and U3471 (N_3471,In_3793,N_1633);
and U3472 (N_3472,N_1738,In_3013);
nor U3473 (N_3473,In_3385,N_1300);
nor U3474 (N_3474,N_1540,N_219);
xor U3475 (N_3475,N_1237,In_1950);
xnor U3476 (N_3476,N_1702,N_72);
nand U3477 (N_3477,N_394,N_1215);
nor U3478 (N_3478,N_1169,N_950);
xor U3479 (N_3479,N_1044,In_4739);
and U3480 (N_3480,N_1491,N_1752);
nor U3481 (N_3481,N_1691,N_350);
nor U3482 (N_3482,N_833,N_302);
nor U3483 (N_3483,N_303,N_1899);
and U3484 (N_3484,In_1973,N_884);
nand U3485 (N_3485,In_4316,N_1626);
or U3486 (N_3486,N_1204,N_1235);
nor U3487 (N_3487,In_516,N_1647);
nand U3488 (N_3488,N_1870,N_856);
xor U3489 (N_3489,In_812,N_1667);
and U3490 (N_3490,N_572,In_4401);
xor U3491 (N_3491,In_4720,N_1311);
nand U3492 (N_3492,In_2378,In_696);
and U3493 (N_3493,In_4995,N_68);
and U3494 (N_3494,N_1797,In_4492);
xor U3495 (N_3495,N_996,In_4357);
or U3496 (N_3496,N_1010,N_1469);
and U3497 (N_3497,N_972,N_664);
or U3498 (N_3498,N_580,N_608);
nand U3499 (N_3499,N_999,N_898);
and U3500 (N_3500,In_920,In_4357);
xor U3501 (N_3501,N_1406,N_30);
nor U3502 (N_3502,In_2204,In_233);
xor U3503 (N_3503,In_2117,In_3560);
xor U3504 (N_3504,N_430,N_94);
and U3505 (N_3505,N_57,N_1328);
or U3506 (N_3506,N_1315,N_737);
and U3507 (N_3507,N_588,N_1132);
or U3508 (N_3508,N_856,N_123);
nand U3509 (N_3509,N_618,In_92);
nor U3510 (N_3510,N_781,In_3964);
and U3511 (N_3511,In_2117,N_1177);
nand U3512 (N_3512,In_593,N_224);
nor U3513 (N_3513,In_4558,In_1000);
and U3514 (N_3514,In_1631,N_604);
nand U3515 (N_3515,N_1956,In_1650);
and U3516 (N_3516,N_1706,N_148);
nor U3517 (N_3517,N_1586,N_1716);
or U3518 (N_3518,In_4746,N_1876);
nor U3519 (N_3519,N_309,N_22);
and U3520 (N_3520,N_861,N_1328);
xnor U3521 (N_3521,N_1336,In_3519);
xnor U3522 (N_3522,In_4110,N_1189);
nor U3523 (N_3523,In_3651,In_3737);
or U3524 (N_3524,N_1140,N_1418);
nand U3525 (N_3525,N_64,N_1245);
or U3526 (N_3526,N_1829,N_1501);
xor U3527 (N_3527,N_408,N_721);
xnor U3528 (N_3528,N_1264,In_1221);
and U3529 (N_3529,N_886,N_767);
nor U3530 (N_3530,In_837,In_4605);
nor U3531 (N_3531,N_443,N_1211);
and U3532 (N_3532,N_1660,In_4724);
nand U3533 (N_3533,N_1550,In_1248);
nand U3534 (N_3534,In_2129,In_2528);
and U3535 (N_3535,In_3045,N_1706);
xnor U3536 (N_3536,In_4823,In_4671);
and U3537 (N_3537,N_973,N_13);
or U3538 (N_3538,N_269,In_3047);
nor U3539 (N_3539,N_647,In_3235);
xor U3540 (N_3540,N_1557,N_1024);
or U3541 (N_3541,N_1288,N_1696);
nor U3542 (N_3542,N_1572,In_1492);
nor U3543 (N_3543,In_4649,In_2998);
nand U3544 (N_3544,In_1195,In_3962);
nor U3545 (N_3545,In_4785,N_74);
nor U3546 (N_3546,N_212,In_2710);
xor U3547 (N_3547,In_4388,In_306);
or U3548 (N_3548,N_747,In_2062);
xor U3549 (N_3549,N_588,N_31);
nor U3550 (N_3550,N_1925,N_267);
nor U3551 (N_3551,N_1033,N_1244);
and U3552 (N_3552,In_372,N_817);
and U3553 (N_3553,N_1438,N_1593);
or U3554 (N_3554,In_410,In_3870);
nand U3555 (N_3555,In_1882,N_1058);
nor U3556 (N_3556,In_1725,N_1928);
nor U3557 (N_3557,N_1618,In_3148);
nand U3558 (N_3558,In_2124,N_1973);
xor U3559 (N_3559,N_569,N_1567);
or U3560 (N_3560,N_957,In_2377);
and U3561 (N_3561,N_1108,N_1191);
or U3562 (N_3562,In_4807,N_55);
and U3563 (N_3563,In_4135,In_711);
or U3564 (N_3564,N_1856,N_592);
nor U3565 (N_3565,In_1481,N_515);
nor U3566 (N_3566,N_1794,N_751);
nand U3567 (N_3567,N_964,In_4565);
xnor U3568 (N_3568,N_1337,In_3386);
and U3569 (N_3569,N_1157,N_853);
nand U3570 (N_3570,N_1264,In_516);
xnor U3571 (N_3571,In_2775,N_147);
nor U3572 (N_3572,N_989,N_184);
or U3573 (N_3573,In_3060,In_4000);
xor U3574 (N_3574,In_3013,N_152);
and U3575 (N_3575,N_275,N_1606);
xnor U3576 (N_3576,In_1512,N_1410);
xnor U3577 (N_3577,N_1974,In_1852);
nand U3578 (N_3578,N_575,N_740);
nor U3579 (N_3579,N_414,N_1121);
and U3580 (N_3580,In_3094,In_3589);
or U3581 (N_3581,In_4256,N_957);
and U3582 (N_3582,In_2233,N_462);
nor U3583 (N_3583,N_1810,N_377);
or U3584 (N_3584,N_1476,N_1578);
nand U3585 (N_3585,In_4135,N_797);
nand U3586 (N_3586,In_1341,In_4629);
and U3587 (N_3587,N_1839,In_2101);
nand U3588 (N_3588,N_1435,N_696);
nand U3589 (N_3589,N_205,N_266);
nor U3590 (N_3590,N_1687,N_1840);
nand U3591 (N_3591,N_1505,In_3531);
and U3592 (N_3592,N_693,N_1926);
or U3593 (N_3593,N_1722,In_281);
and U3594 (N_3594,N_446,N_450);
xnor U3595 (N_3595,N_102,N_1392);
nor U3596 (N_3596,In_1839,N_1235);
and U3597 (N_3597,N_1390,N_1528);
and U3598 (N_3598,In_1567,N_388);
or U3599 (N_3599,In_693,N_1976);
or U3600 (N_3600,In_1465,N_1631);
or U3601 (N_3601,N_350,N_927);
nor U3602 (N_3602,N_1089,In_2967);
nor U3603 (N_3603,N_1914,N_583);
or U3604 (N_3604,N_87,N_580);
nor U3605 (N_3605,N_210,N_1326);
or U3606 (N_3606,In_167,In_4926);
and U3607 (N_3607,N_1912,In_3647);
nand U3608 (N_3608,N_552,In_3351);
or U3609 (N_3609,N_1395,In_1270);
nor U3610 (N_3610,In_1636,N_317);
nand U3611 (N_3611,N_1638,In_2316);
or U3612 (N_3612,N_1375,In_2990);
or U3613 (N_3613,N_202,N_765);
nand U3614 (N_3614,N_1472,N_596);
nor U3615 (N_3615,N_308,N_1618);
xor U3616 (N_3616,N_883,In_3272);
nand U3617 (N_3617,In_3346,In_3960);
nand U3618 (N_3618,N_413,In_3016);
nor U3619 (N_3619,N_185,N_1678);
and U3620 (N_3620,N_805,In_1462);
and U3621 (N_3621,N_382,N_1463);
xor U3622 (N_3622,N_978,In_1517);
nor U3623 (N_3623,In_1747,N_1520);
nor U3624 (N_3624,N_1097,N_1474);
nand U3625 (N_3625,N_291,N_93);
nor U3626 (N_3626,In_2288,N_1143);
xor U3627 (N_3627,N_261,N_1075);
or U3628 (N_3628,N_1914,N_890);
or U3629 (N_3629,N_1932,In_2108);
nor U3630 (N_3630,N_86,N_367);
nor U3631 (N_3631,N_873,In_661);
or U3632 (N_3632,N_1905,In_758);
or U3633 (N_3633,N_1435,In_4248);
nor U3634 (N_3634,N_1577,N_400);
nand U3635 (N_3635,N_884,In_913);
or U3636 (N_3636,N_1846,N_1690);
nor U3637 (N_3637,N_1735,N_819);
or U3638 (N_3638,N_1484,In_920);
nor U3639 (N_3639,In_1400,N_1710);
or U3640 (N_3640,N_1360,In_4651);
or U3641 (N_3641,N_1420,In_3922);
nand U3642 (N_3642,N_1296,In_4162);
or U3643 (N_3643,N_542,N_1542);
xnor U3644 (N_3644,In_2817,N_511);
xor U3645 (N_3645,N_1372,N_1735);
nor U3646 (N_3646,N_1504,In_1);
nor U3647 (N_3647,In_2775,N_332);
nand U3648 (N_3648,N_1767,In_4358);
or U3649 (N_3649,N_1627,N_1219);
nor U3650 (N_3650,N_469,N_1738);
nor U3651 (N_3651,In_820,In_334);
xnor U3652 (N_3652,N_938,N_62);
and U3653 (N_3653,N_1946,N_1849);
and U3654 (N_3654,In_4160,N_1840);
and U3655 (N_3655,In_4036,In_4157);
nand U3656 (N_3656,N_1087,N_1315);
and U3657 (N_3657,N_518,N_1807);
nand U3658 (N_3658,N_41,In_2376);
and U3659 (N_3659,N_1316,N_194);
or U3660 (N_3660,N_1167,N_1649);
or U3661 (N_3661,N_1045,N_627);
nand U3662 (N_3662,N_178,N_36);
xnor U3663 (N_3663,N_1339,N_1047);
or U3664 (N_3664,In_3077,N_13);
nor U3665 (N_3665,N_1782,N_377);
nand U3666 (N_3666,In_3609,N_23);
xor U3667 (N_3667,N_1685,In_436);
xor U3668 (N_3668,N_1419,In_1998);
and U3669 (N_3669,N_1354,In_478);
and U3670 (N_3670,N_857,N_1063);
nor U3671 (N_3671,N_896,In_1842);
nand U3672 (N_3672,N_1050,In_3511);
nand U3673 (N_3673,In_2825,N_1799);
xor U3674 (N_3674,N_1276,In_3828);
nor U3675 (N_3675,In_3213,In_3272);
nor U3676 (N_3676,N_1710,N_218);
and U3677 (N_3677,N_214,N_549);
xnor U3678 (N_3678,N_1397,N_1720);
xnor U3679 (N_3679,N_1968,N_459);
nor U3680 (N_3680,In_1989,N_1812);
and U3681 (N_3681,In_4851,In_237);
or U3682 (N_3682,N_1767,N_38);
nand U3683 (N_3683,N_1435,N_158);
nand U3684 (N_3684,In_4726,In_52);
and U3685 (N_3685,In_3312,N_1741);
or U3686 (N_3686,In_4752,N_887);
or U3687 (N_3687,N_1391,N_72);
and U3688 (N_3688,In_4756,N_83);
and U3689 (N_3689,N_1091,In_588);
nor U3690 (N_3690,N_628,N_293);
or U3691 (N_3691,N_914,In_1980);
nor U3692 (N_3692,N_1527,In_4447);
nor U3693 (N_3693,In_269,N_842);
nor U3694 (N_3694,N_1722,In_2593);
xnor U3695 (N_3695,N_1008,In_4694);
and U3696 (N_3696,N_652,N_305);
or U3697 (N_3697,In_3242,N_207);
and U3698 (N_3698,N_1267,N_1911);
xor U3699 (N_3699,N_1829,In_3143);
and U3700 (N_3700,In_4012,In_2364);
or U3701 (N_3701,N_838,N_1471);
and U3702 (N_3702,N_1323,N_746);
nor U3703 (N_3703,In_3092,In_1439);
and U3704 (N_3704,In_3242,N_192);
nand U3705 (N_3705,N_1334,In_3815);
and U3706 (N_3706,N_1679,N_822);
nand U3707 (N_3707,N_1276,N_1105);
nand U3708 (N_3708,N_32,In_1998);
nor U3709 (N_3709,N_1210,N_1756);
or U3710 (N_3710,N_10,N_1552);
nor U3711 (N_3711,N_675,N_859);
and U3712 (N_3712,N_1722,N_483);
nand U3713 (N_3713,N_1491,N_1730);
or U3714 (N_3714,N_813,N_222);
nor U3715 (N_3715,N_1927,In_1492);
xnor U3716 (N_3716,N_1560,N_925);
and U3717 (N_3717,In_4058,In_1680);
nand U3718 (N_3718,N_1548,N_740);
or U3719 (N_3719,N_1575,N_675);
or U3720 (N_3720,N_1492,In_4433);
xnor U3721 (N_3721,In_306,N_497);
xor U3722 (N_3722,N_1693,N_1935);
xor U3723 (N_3723,N_703,In_3749);
nand U3724 (N_3724,N_592,In_4151);
and U3725 (N_3725,N_833,In_4392);
xnor U3726 (N_3726,In_4720,N_1645);
xnor U3727 (N_3727,N_1381,N_1738);
and U3728 (N_3728,N_856,N_1767);
nor U3729 (N_3729,In_3298,In_800);
xor U3730 (N_3730,N_579,N_93);
nor U3731 (N_3731,N_748,N_914);
nor U3732 (N_3732,N_1829,N_306);
xor U3733 (N_3733,N_721,In_1434);
nor U3734 (N_3734,N_1030,N_1505);
or U3735 (N_3735,N_1487,In_4926);
and U3736 (N_3736,N_1998,N_1975);
nor U3737 (N_3737,In_4689,N_592);
or U3738 (N_3738,In_1853,N_1220);
or U3739 (N_3739,In_2824,In_1078);
xnor U3740 (N_3740,N_259,In_2672);
and U3741 (N_3741,N_888,N_717);
and U3742 (N_3742,In_3010,In_4697);
xor U3743 (N_3743,In_2846,In_3701);
nand U3744 (N_3744,N_48,N_1858);
or U3745 (N_3745,N_1870,N_3);
xnor U3746 (N_3746,N_494,In_820);
xor U3747 (N_3747,In_3106,N_1487);
nor U3748 (N_3748,N_243,N_1862);
xnor U3749 (N_3749,N_151,In_848);
xor U3750 (N_3750,N_989,In_3041);
nor U3751 (N_3751,In_292,N_1944);
or U3752 (N_3752,N_1707,N_153);
nand U3753 (N_3753,N_1539,N_1736);
nand U3754 (N_3754,N_476,N_1414);
or U3755 (N_3755,In_2352,In_535);
xor U3756 (N_3756,N_1550,N_1378);
or U3757 (N_3757,N_1079,In_1434);
nand U3758 (N_3758,N_77,In_4476);
xnor U3759 (N_3759,In_3062,N_1);
and U3760 (N_3760,N_190,In_3092);
and U3761 (N_3761,In_4587,N_581);
and U3762 (N_3762,In_3877,N_1887);
nor U3763 (N_3763,In_653,In_4689);
nor U3764 (N_3764,N_971,In_3495);
or U3765 (N_3765,N_584,In_1972);
xnor U3766 (N_3766,N_734,N_1989);
or U3767 (N_3767,In_2875,N_195);
nor U3768 (N_3768,In_4317,N_287);
or U3769 (N_3769,N_1143,N_266);
xor U3770 (N_3770,N_1110,N_211);
nand U3771 (N_3771,In_2159,N_1034);
and U3772 (N_3772,In_3425,N_1695);
and U3773 (N_3773,N_252,N_1486);
or U3774 (N_3774,In_748,N_1371);
nor U3775 (N_3775,N_167,In_1624);
xor U3776 (N_3776,N_307,N_1352);
nor U3777 (N_3777,In_3799,N_900);
xor U3778 (N_3778,N_172,N_1464);
nand U3779 (N_3779,In_1462,N_90);
nor U3780 (N_3780,N_1353,N_115);
nand U3781 (N_3781,In_2710,N_206);
nor U3782 (N_3782,In_478,N_435);
xor U3783 (N_3783,N_1098,N_338);
xnor U3784 (N_3784,N_798,N_256);
and U3785 (N_3785,N_1043,In_3130);
and U3786 (N_3786,In_4181,In_2165);
xor U3787 (N_3787,In_4154,N_1897);
nor U3788 (N_3788,N_297,In_1909);
xor U3789 (N_3789,N_1418,In_2004);
and U3790 (N_3790,N_726,N_943);
and U3791 (N_3791,In_432,N_729);
and U3792 (N_3792,N_208,N_867);
or U3793 (N_3793,N_1571,In_3952);
or U3794 (N_3794,N_1222,N_1482);
and U3795 (N_3795,N_152,N_468);
xnor U3796 (N_3796,N_1485,In_4215);
nand U3797 (N_3797,In_2377,In_440);
nor U3798 (N_3798,N_875,In_1322);
or U3799 (N_3799,N_577,In_492);
nor U3800 (N_3800,N_1030,In_2505);
nand U3801 (N_3801,N_454,N_685);
xor U3802 (N_3802,N_1452,N_608);
nand U3803 (N_3803,N_1189,N_144);
and U3804 (N_3804,N_1552,N_1213);
nor U3805 (N_3805,In_2650,N_135);
nor U3806 (N_3806,N_1315,N_5);
xnor U3807 (N_3807,N_1793,N_162);
and U3808 (N_3808,N_1584,In_591);
or U3809 (N_3809,In_3137,N_1037);
and U3810 (N_3810,N_1023,N_580);
nor U3811 (N_3811,In_2455,N_1436);
and U3812 (N_3812,N_218,N_1622);
xnor U3813 (N_3813,In_1142,In_4724);
nor U3814 (N_3814,N_51,N_1392);
xnor U3815 (N_3815,N_601,N_1514);
or U3816 (N_3816,N_231,In_3328);
and U3817 (N_3817,N_678,In_556);
xnor U3818 (N_3818,N_1072,N_688);
nor U3819 (N_3819,N_1446,In_3086);
nand U3820 (N_3820,In_1103,In_1415);
and U3821 (N_3821,N_1500,N_1417);
xnor U3822 (N_3822,N_1269,N_1334);
and U3823 (N_3823,N_1940,N_1208);
xnor U3824 (N_3824,N_1181,N_1505);
and U3825 (N_3825,In_3921,N_1928);
and U3826 (N_3826,In_2216,N_1396);
xnor U3827 (N_3827,N_809,N_555);
or U3828 (N_3828,N_58,N_1282);
and U3829 (N_3829,N_693,N_303);
xnor U3830 (N_3830,N_988,N_442);
nor U3831 (N_3831,N_991,N_1625);
nand U3832 (N_3832,N_683,In_824);
xnor U3833 (N_3833,In_1649,N_1880);
nand U3834 (N_3834,N_894,N_1388);
nor U3835 (N_3835,N_1413,N_1705);
and U3836 (N_3836,In_1096,N_1207);
nand U3837 (N_3837,N_1214,N_636);
and U3838 (N_3838,N_499,N_185);
and U3839 (N_3839,N_1430,N_844);
or U3840 (N_3840,N_1993,In_4612);
or U3841 (N_3841,N_1743,N_1587);
or U3842 (N_3842,In_2250,In_869);
nand U3843 (N_3843,In_1267,In_2430);
nand U3844 (N_3844,N_1294,In_3346);
or U3845 (N_3845,N_299,N_524);
and U3846 (N_3846,N_449,In_2737);
nor U3847 (N_3847,N_63,N_1960);
xnor U3848 (N_3848,In_4225,In_4756);
nand U3849 (N_3849,N_992,N_1814);
nand U3850 (N_3850,In_1079,N_119);
and U3851 (N_3851,In_3841,N_1067);
or U3852 (N_3852,In_127,In_2786);
nand U3853 (N_3853,In_3060,In_4643);
nor U3854 (N_3854,N_1546,N_271);
and U3855 (N_3855,In_4327,N_1276);
xor U3856 (N_3856,N_929,N_603);
and U3857 (N_3857,N_1871,N_629);
nand U3858 (N_3858,N_43,N_472);
and U3859 (N_3859,N_145,In_3991);
nand U3860 (N_3860,N_371,N_844);
and U3861 (N_3861,In_647,N_1761);
and U3862 (N_3862,In_885,N_1384);
nor U3863 (N_3863,In_4227,In_941);
nor U3864 (N_3864,In_3952,In_3213);
nand U3865 (N_3865,In_2945,N_1159);
xnor U3866 (N_3866,In_1569,In_2178);
xor U3867 (N_3867,N_957,N_236);
nor U3868 (N_3868,N_276,N_1429);
and U3869 (N_3869,In_4088,N_1444);
or U3870 (N_3870,N_1804,N_1239);
or U3871 (N_3871,N_1677,N_341);
xor U3872 (N_3872,N_1758,N_1017);
and U3873 (N_3873,N_1239,N_1884);
nand U3874 (N_3874,N_83,N_1326);
or U3875 (N_3875,N_106,N_34);
and U3876 (N_3876,N_1080,In_1660);
nor U3877 (N_3877,In_2291,N_1087);
and U3878 (N_3878,N_1728,N_373);
and U3879 (N_3879,In_2851,N_883);
xor U3880 (N_3880,N_1573,N_1648);
xor U3881 (N_3881,N_1689,N_73);
or U3882 (N_3882,N_1642,N_905);
xor U3883 (N_3883,N_1314,In_4697);
or U3884 (N_3884,N_1819,In_3045);
and U3885 (N_3885,N_1365,N_99);
nand U3886 (N_3886,In_3457,N_652);
and U3887 (N_3887,N_270,N_1692);
nand U3888 (N_3888,N_1468,N_1004);
xnor U3889 (N_3889,N_1054,In_791);
and U3890 (N_3890,N_513,In_1030);
nor U3891 (N_3891,N_1451,N_1780);
and U3892 (N_3892,N_1927,N_709);
or U3893 (N_3893,In_584,In_1836);
or U3894 (N_3894,N_969,N_1512);
nand U3895 (N_3895,N_797,In_2686);
or U3896 (N_3896,N_147,In_425);
nand U3897 (N_3897,N_968,In_709);
nor U3898 (N_3898,In_760,N_1679);
or U3899 (N_3899,N_1254,N_871);
nor U3900 (N_3900,N_358,N_627);
or U3901 (N_3901,N_345,N_337);
nand U3902 (N_3902,N_1323,N_1424);
xor U3903 (N_3903,N_894,In_3641);
xnor U3904 (N_3904,N_1575,N_12);
and U3905 (N_3905,In_4851,N_856);
and U3906 (N_3906,In_2238,N_683);
and U3907 (N_3907,N_499,In_867);
nand U3908 (N_3908,N_658,In_1852);
or U3909 (N_3909,In_3272,N_95);
xor U3910 (N_3910,N_263,In_3805);
xor U3911 (N_3911,N_739,N_1076);
and U3912 (N_3912,N_1247,In_1747);
xor U3913 (N_3913,In_2113,In_584);
xor U3914 (N_3914,N_358,In_736);
and U3915 (N_3915,N_625,N_1108);
and U3916 (N_3916,In_728,N_1944);
or U3917 (N_3917,N_76,N_490);
or U3918 (N_3918,N_551,In_4414);
xnor U3919 (N_3919,N_36,In_4160);
or U3920 (N_3920,In_4527,In_1045);
xor U3921 (N_3921,N_1386,N_1266);
xor U3922 (N_3922,In_2710,In_3936);
or U3923 (N_3923,N_1501,In_2593);
nor U3924 (N_3924,In_804,In_2120);
nand U3925 (N_3925,In_1481,N_679);
xnor U3926 (N_3926,N_809,N_830);
xnor U3927 (N_3927,In_1593,In_3502);
or U3928 (N_3928,In_3457,In_2498);
xnor U3929 (N_3929,In_2374,N_1258);
nand U3930 (N_3930,In_2305,In_3566);
nand U3931 (N_3931,In_3879,N_133);
xnor U3932 (N_3932,In_3039,N_575);
xor U3933 (N_3933,N_240,In_824);
and U3934 (N_3934,N_1951,In_3873);
xor U3935 (N_3935,N_1770,In_3214);
nor U3936 (N_3936,N_518,N_182);
xor U3937 (N_3937,In_4716,N_1187);
nand U3938 (N_3938,N_1781,N_263);
xor U3939 (N_3939,N_970,In_3357);
nor U3940 (N_3940,N_32,N_1134);
xor U3941 (N_3941,N_680,In_201);
and U3942 (N_3942,N_1990,In_4739);
nand U3943 (N_3943,N_33,In_4604);
or U3944 (N_3944,N_1526,In_4367);
nand U3945 (N_3945,In_3651,N_1127);
or U3946 (N_3946,N_305,N_798);
nand U3947 (N_3947,N_984,N_519);
xnor U3948 (N_3948,N_553,In_805);
or U3949 (N_3949,N_1090,N_595);
xor U3950 (N_3950,N_777,In_1838);
or U3951 (N_3951,In_3700,N_1830);
or U3952 (N_3952,N_802,N_1279);
nand U3953 (N_3953,N_744,N_411);
and U3954 (N_3954,N_842,N_834);
or U3955 (N_3955,N_479,N_1991);
xnor U3956 (N_3956,N_1219,In_1874);
nand U3957 (N_3957,N_1304,N_665);
xnor U3958 (N_3958,In_3589,In_388);
and U3959 (N_3959,N_1852,In_4198);
nor U3960 (N_3960,N_739,N_1545);
or U3961 (N_3961,N_586,In_2062);
or U3962 (N_3962,In_1330,In_2874);
or U3963 (N_3963,N_812,N_1971);
or U3964 (N_3964,N_1006,N_1479);
xor U3965 (N_3965,N_386,In_3952);
nor U3966 (N_3966,N_277,N_1379);
or U3967 (N_3967,N_1103,In_3502);
nand U3968 (N_3968,In_1988,In_882);
nand U3969 (N_3969,N_1328,N_1791);
or U3970 (N_3970,N_1423,In_2442);
and U3971 (N_3971,In_4591,In_3133);
xor U3972 (N_3972,N_250,In_4162);
xnor U3973 (N_3973,N_1113,N_1168);
nor U3974 (N_3974,N_788,N_1669);
nor U3975 (N_3975,N_295,In_402);
or U3976 (N_3976,In_3647,In_92);
xnor U3977 (N_3977,N_580,In_98);
or U3978 (N_3978,N_1771,N_588);
and U3979 (N_3979,N_1644,N_293);
or U3980 (N_3980,In_3330,N_1858);
nand U3981 (N_3981,N_964,N_1880);
or U3982 (N_3982,In_269,N_759);
and U3983 (N_3983,N_452,In_3084);
nand U3984 (N_3984,In_1390,N_1806);
or U3985 (N_3985,In_807,In_1943);
nand U3986 (N_3986,N_21,N_1323);
nor U3987 (N_3987,In_4048,N_1901);
xnor U3988 (N_3988,In_2305,N_1156);
nor U3989 (N_3989,N_1584,N_831);
xnor U3990 (N_3990,In_1593,N_187);
nor U3991 (N_3991,In_4623,In_3921);
and U3992 (N_3992,In_3094,N_383);
nand U3993 (N_3993,N_690,N_258);
or U3994 (N_3994,In_1622,In_4616);
nand U3995 (N_3995,In_1481,N_1653);
and U3996 (N_3996,N_1933,N_1536);
nand U3997 (N_3997,N_1181,N_1093);
or U3998 (N_3998,In_1837,In_4696);
and U3999 (N_3999,N_878,N_281);
xor U4000 (N_4000,N_3981,N_3127);
xnor U4001 (N_4001,N_3335,N_2811);
and U4002 (N_4002,N_2075,N_3016);
or U4003 (N_4003,N_3831,N_3217);
and U4004 (N_4004,N_2521,N_3697);
or U4005 (N_4005,N_3369,N_2434);
nor U4006 (N_4006,N_3634,N_2770);
and U4007 (N_4007,N_2640,N_2916);
and U4008 (N_4008,N_2619,N_2166);
and U4009 (N_4009,N_2278,N_3391);
or U4010 (N_4010,N_3511,N_2012);
xor U4011 (N_4011,N_3479,N_3885);
nand U4012 (N_4012,N_2847,N_2441);
xor U4013 (N_4013,N_3595,N_2169);
and U4014 (N_4014,N_2763,N_2622);
nor U4015 (N_4015,N_2766,N_3617);
nor U4016 (N_4016,N_3242,N_3917);
nand U4017 (N_4017,N_2021,N_2950);
or U4018 (N_4018,N_2605,N_3184);
nand U4019 (N_4019,N_3941,N_2782);
and U4020 (N_4020,N_2334,N_2436);
nand U4021 (N_4021,N_3019,N_2964);
nand U4022 (N_4022,N_2875,N_2479);
nand U4023 (N_4023,N_3290,N_2374);
xor U4024 (N_4024,N_3573,N_2616);
nor U4025 (N_4025,N_3091,N_2096);
nand U4026 (N_4026,N_2353,N_3112);
and U4027 (N_4027,N_3446,N_2234);
and U4028 (N_4028,N_2229,N_3560);
nand U4029 (N_4029,N_2803,N_2363);
nand U4030 (N_4030,N_2726,N_2073);
or U4031 (N_4031,N_2139,N_2011);
xor U4032 (N_4032,N_3599,N_2732);
and U4033 (N_4033,N_3604,N_2016);
or U4034 (N_4034,N_3864,N_3212);
xnor U4035 (N_4035,N_2462,N_2313);
or U4036 (N_4036,N_2404,N_3356);
or U4037 (N_4037,N_2131,N_2344);
or U4038 (N_4038,N_3418,N_2989);
xor U4039 (N_4039,N_3771,N_3909);
xor U4040 (N_4040,N_2596,N_2801);
or U4041 (N_4041,N_2394,N_3168);
and U4042 (N_4042,N_2113,N_3466);
nor U4043 (N_4043,N_2986,N_2284);
and U4044 (N_4044,N_3274,N_2635);
and U4045 (N_4045,N_3603,N_2905);
or U4046 (N_4046,N_3285,N_3877);
xnor U4047 (N_4047,N_2509,N_3336);
or U4048 (N_4048,N_3904,N_3304);
or U4049 (N_4049,N_3045,N_3481);
xnor U4050 (N_4050,N_3211,N_2062);
xnor U4051 (N_4051,N_2641,N_2032);
xor U4052 (N_4052,N_2220,N_3995);
nor U4053 (N_4053,N_3773,N_3913);
xnor U4054 (N_4054,N_3240,N_2427);
nand U4055 (N_4055,N_2528,N_3377);
nor U4056 (N_4056,N_3722,N_3987);
nor U4057 (N_4057,N_2807,N_3600);
and U4058 (N_4058,N_2380,N_3038);
nand U4059 (N_4059,N_2867,N_3145);
and U4060 (N_4060,N_3098,N_3507);
nor U4061 (N_4061,N_3120,N_2280);
nand U4062 (N_4062,N_3652,N_2292);
xnor U4063 (N_4063,N_3280,N_2729);
nand U4064 (N_4064,N_2754,N_2846);
xnor U4065 (N_4065,N_3401,N_2673);
xor U4066 (N_4066,N_2405,N_3751);
nand U4067 (N_4067,N_2718,N_2920);
or U4068 (N_4068,N_2655,N_2854);
and U4069 (N_4069,N_2649,N_3908);
nor U4070 (N_4070,N_2272,N_2094);
xnor U4071 (N_4071,N_2712,N_2667);
nor U4072 (N_4072,N_3496,N_3247);
and U4073 (N_4073,N_3064,N_3782);
nor U4074 (N_4074,N_3366,N_2213);
or U4075 (N_4075,N_3153,N_2158);
and U4076 (N_4076,N_3482,N_3135);
nand U4077 (N_4077,N_2736,N_2561);
nor U4078 (N_4078,N_2737,N_2076);
xnor U4079 (N_4079,N_2647,N_2201);
xnor U4080 (N_4080,N_3137,N_3934);
xnor U4081 (N_4081,N_3358,N_3616);
nor U4082 (N_4082,N_2473,N_2051);
nand U4083 (N_4083,N_3218,N_2396);
nand U4084 (N_4084,N_2670,N_3498);
or U4085 (N_4085,N_3974,N_3798);
or U4086 (N_4086,N_2908,N_2773);
and U4087 (N_4087,N_3583,N_2735);
or U4088 (N_4088,N_2199,N_2791);
xor U4089 (N_4089,N_3737,N_3655);
nand U4090 (N_4090,N_2568,N_3753);
nand U4091 (N_4091,N_2960,N_3223);
or U4092 (N_4092,N_2800,N_3291);
nand U4093 (N_4093,N_3769,N_3269);
nand U4094 (N_4094,N_2663,N_2402);
xor U4095 (N_4095,N_2290,N_3157);
or U4096 (N_4096,N_2042,N_3074);
nor U4097 (N_4097,N_3796,N_3793);
and U4098 (N_4098,N_3578,N_3822);
nor U4099 (N_4099,N_2820,N_2844);
nand U4100 (N_4100,N_2702,N_3533);
nor U4101 (N_4101,N_3850,N_3331);
nand U4102 (N_4102,N_2123,N_3107);
nor U4103 (N_4103,N_3976,N_3868);
xor U4104 (N_4104,N_3213,N_3204);
or U4105 (N_4105,N_2167,N_3491);
and U4106 (N_4106,N_3455,N_3740);
and U4107 (N_4107,N_2983,N_2634);
nor U4108 (N_4108,N_3100,N_3855);
or U4109 (N_4109,N_3897,N_3163);
and U4110 (N_4110,N_3915,N_2897);
nor U4111 (N_4111,N_3676,N_2625);
nor U4112 (N_4112,N_2410,N_2785);
or U4113 (N_4113,N_2236,N_3415);
nand U4114 (N_4114,N_2328,N_3489);
nand U4115 (N_4115,N_2739,N_2185);
xnor U4116 (N_4116,N_3182,N_2865);
xnor U4117 (N_4117,N_3375,N_3251);
or U4118 (N_4118,N_2343,N_2298);
or U4119 (N_4119,N_2164,N_2851);
nand U4120 (N_4120,N_3005,N_3633);
nand U4121 (N_4121,N_3924,N_3024);
or U4122 (N_4122,N_3436,N_2923);
nand U4123 (N_4123,N_3619,N_2102);
or U4124 (N_4124,N_2239,N_2698);
or U4125 (N_4125,N_2332,N_3084);
nand U4126 (N_4126,N_2238,N_3283);
and U4127 (N_4127,N_3774,N_3273);
or U4128 (N_4128,N_3330,N_3004);
xor U4129 (N_4129,N_3015,N_2013);
nand U4130 (N_4130,N_2931,N_2703);
and U4131 (N_4131,N_2881,N_2928);
xnor U4132 (N_4132,N_3313,N_3900);
xnor U4133 (N_4133,N_3985,N_3714);
xnor U4134 (N_4134,N_2015,N_2771);
xnor U4135 (N_4135,N_3276,N_2799);
nor U4136 (N_4136,N_2997,N_3757);
xnor U4137 (N_4137,N_3720,N_2098);
nor U4138 (N_4138,N_3195,N_2850);
and U4139 (N_4139,N_3928,N_3539);
or U4140 (N_4140,N_3413,N_3986);
nor U4141 (N_4141,N_2688,N_3011);
nand U4142 (N_4142,N_2361,N_3231);
nor U4143 (N_4143,N_3427,N_2961);
and U4144 (N_4144,N_2002,N_2432);
and U4145 (N_4145,N_2318,N_3143);
and U4146 (N_4146,N_2864,N_3989);
or U4147 (N_4147,N_2795,N_3667);
nor U4148 (N_4148,N_3215,N_2775);
nand U4149 (N_4149,N_3054,N_3140);
or U4150 (N_4150,N_3660,N_3661);
and U4151 (N_4151,N_3233,N_3859);
nor U4152 (N_4152,N_2504,N_3390);
xor U4153 (N_4153,N_2564,N_3160);
nor U4154 (N_4154,N_3947,N_2492);
xnor U4155 (N_4155,N_3741,N_2079);
and U4156 (N_4156,N_2535,N_2705);
nor U4157 (N_4157,N_2887,N_3359);
nor U4158 (N_4158,N_3226,N_3065);
or U4159 (N_4159,N_2682,N_3543);
nor U4160 (N_4160,N_2288,N_2637);
and U4161 (N_4161,N_2194,N_2884);
or U4162 (N_4162,N_2812,N_2805);
nand U4163 (N_4163,N_3621,N_2553);
nand U4164 (N_4164,N_3259,N_2781);
xnor U4165 (N_4165,N_3002,N_2268);
xor U4166 (N_4166,N_2306,N_2891);
nor U4167 (N_4167,N_3063,N_2942);
and U4168 (N_4168,N_3853,N_2206);
xnor U4169 (N_4169,N_2172,N_3190);
xor U4170 (N_4170,N_2685,N_2233);
nor U4171 (N_4171,N_3136,N_2074);
or U4172 (N_4172,N_3288,N_2868);
nor U4173 (N_4173,N_3310,N_2943);
or U4174 (N_4174,N_3736,N_2838);
nand U4175 (N_4175,N_2582,N_2996);
and U4176 (N_4176,N_3587,N_3969);
nor U4177 (N_4177,N_2317,N_2182);
and U4178 (N_4178,N_3705,N_3665);
nor U4179 (N_4179,N_3955,N_3944);
and U4180 (N_4180,N_3344,N_2728);
xor U4181 (N_4181,N_2995,N_3349);
xor U4182 (N_4182,N_3445,N_2010);
or U4183 (N_4183,N_2889,N_3875);
nand U4184 (N_4184,N_2150,N_2751);
nand U4185 (N_4185,N_3684,N_3938);
nand U4186 (N_4186,N_2835,N_2497);
nand U4187 (N_4187,N_2362,N_2692);
xor U4188 (N_4188,N_3264,N_2629);
or U4189 (N_4189,N_3836,N_2722);
or U4190 (N_4190,N_3382,N_2612);
nand U4191 (N_4191,N_3116,N_3800);
and U4192 (N_4192,N_2817,N_2953);
or U4193 (N_4193,N_2885,N_2690);
and U4194 (N_4194,N_3109,N_2547);
xor U4195 (N_4195,N_2904,N_3959);
nor U4196 (N_4196,N_3918,N_2484);
and U4197 (N_4197,N_3151,N_2072);
xor U4198 (N_4198,N_2639,N_2910);
nor U4199 (N_4199,N_3365,N_2638);
nor U4200 (N_4200,N_3039,N_2365);
and U4201 (N_4201,N_3253,N_2901);
nand U4202 (N_4202,N_3817,N_2871);
nand U4203 (N_4203,N_3526,N_2527);
nand U4204 (N_4204,N_3698,N_3544);
and U4205 (N_4205,N_2176,N_3034);
or U4206 (N_4206,N_2709,N_2376);
or U4207 (N_4207,N_2412,N_2157);
xnor U4208 (N_4208,N_2575,N_2495);
or U4209 (N_4209,N_2257,N_3085);
and U4210 (N_4210,N_3721,N_2463);
nand U4211 (N_4211,N_3819,N_3452);
nand U4212 (N_4212,N_2069,N_3531);
nand U4213 (N_4213,N_2768,N_3815);
nor U4214 (N_4214,N_3248,N_2962);
xnor U4215 (N_4215,N_2939,N_3271);
nand U4216 (N_4216,N_2117,N_3397);
xnor U4217 (N_4217,N_2159,N_2843);
and U4218 (N_4218,N_3060,N_3144);
xor U4219 (N_4219,N_2447,N_3936);
nor U4220 (N_4220,N_3582,N_2711);
xnor U4221 (N_4221,N_2546,N_2385);
and U4222 (N_4222,N_3429,N_2531);
and U4223 (N_4223,N_3139,N_2584);
nand U4224 (N_4224,N_2777,N_2727);
xnor U4225 (N_4225,N_2337,N_3338);
and U4226 (N_4226,N_2876,N_3300);
xor U4227 (N_4227,N_2422,N_2033);
xor U4228 (N_4228,N_3830,N_2295);
and U4229 (N_4229,N_2745,N_2302);
nand U4230 (N_4230,N_2697,N_2603);
or U4231 (N_4231,N_3219,N_3188);
nor U4232 (N_4232,N_2813,N_2112);
xnor U4233 (N_4233,N_3732,N_2026);
or U4234 (N_4234,N_2118,N_3871);
and U4235 (N_4235,N_2987,N_3393);
or U4236 (N_4236,N_2578,N_3095);
xnor U4237 (N_4237,N_3685,N_2360);
and U4238 (N_4238,N_2248,N_3653);
xor U4239 (N_4239,N_2235,N_3572);
or U4240 (N_4240,N_3933,N_3072);
nand U4241 (N_4241,N_3922,N_2966);
xnor U4242 (N_4242,N_2925,N_2401);
or U4243 (N_4243,N_2107,N_2959);
or U4244 (N_4244,N_3912,N_2853);
nor U4245 (N_4245,N_2128,N_3444);
and U4246 (N_4246,N_3983,N_3891);
nor U4247 (N_4247,N_2384,N_3733);
xor U4248 (N_4248,N_3605,N_2429);
nand U4249 (N_4249,N_3268,N_3225);
nor U4250 (N_4250,N_2308,N_2273);
xor U4251 (N_4251,N_2140,N_3053);
xnor U4252 (N_4252,N_3516,N_3606);
nor U4253 (N_4253,N_2888,N_3687);
nor U4254 (N_4254,N_2188,N_3241);
nor U4255 (N_4255,N_2103,N_2517);
nand U4256 (N_4256,N_2091,N_3164);
nor U4257 (N_4257,N_2963,N_2440);
and U4258 (N_4258,N_3132,N_2862);
nand U4259 (N_4259,N_2717,N_3235);
nor U4260 (N_4260,N_3088,N_2264);
xor U4261 (N_4261,N_3786,N_2842);
and U4262 (N_4262,N_2678,N_3416);
nand U4263 (N_4263,N_3159,N_2304);
nor U4264 (N_4264,N_3592,N_3022);
and U4265 (N_4265,N_2758,N_2573);
and U4266 (N_4266,N_2615,N_3238);
or U4267 (N_4267,N_3860,N_2592);
nand U4268 (N_4268,N_2689,N_3766);
nand U4269 (N_4269,N_3325,N_2408);
or U4270 (N_4270,N_3282,N_2913);
xor U4271 (N_4271,N_3048,N_2058);
nor U4272 (N_4272,N_3387,N_2407);
nor U4273 (N_4273,N_3298,N_2071);
nor U4274 (N_4274,N_2255,N_2000);
and U4275 (N_4275,N_2765,N_3585);
nor U4276 (N_4276,N_3333,N_3301);
nand U4277 (N_4277,N_3772,N_2217);
nor U4278 (N_4278,N_2311,N_2154);
nor U4279 (N_4279,N_2787,N_3399);
nor U4280 (N_4280,N_2794,N_2597);
or U4281 (N_4281,N_2796,N_3326);
nand U4282 (N_4282,N_2469,N_3406);
and U4283 (N_4283,N_3747,N_2121);
and U4284 (N_4284,N_2645,N_3492);
or U4285 (N_4285,N_3236,N_3297);
and U4286 (N_4286,N_3978,N_2183);
and U4287 (N_4287,N_2924,N_2769);
nor U4288 (N_4288,N_2415,N_3169);
nor U4289 (N_4289,N_2945,N_2968);
xor U4290 (N_4290,N_2970,N_3594);
or U4291 (N_4291,N_2554,N_3111);
or U4292 (N_4292,N_2675,N_2626);
nand U4293 (N_4293,N_2565,N_3635);
or U4294 (N_4294,N_2253,N_2927);
or U4295 (N_4295,N_3467,N_3318);
xor U4296 (N_4296,N_3475,N_3322);
xnor U4297 (N_4297,N_2330,N_3404);
nor U4298 (N_4298,N_2082,N_2496);
nand U4299 (N_4299,N_2661,N_3662);
nand U4300 (N_4300,N_3823,N_2522);
and U4301 (N_4301,N_2674,N_2216);
nand U4302 (N_4302,N_2355,N_2814);
xor U4303 (N_4303,N_3453,N_2877);
nor U4304 (N_4304,N_3106,N_2100);
nor U4305 (N_4305,N_2538,N_3825);
or U4306 (N_4306,N_3051,N_3530);
nor U4307 (N_4307,N_3443,N_3672);
and U4308 (N_4308,N_2453,N_3659);
nor U4309 (N_4309,N_2633,N_2226);
and U4310 (N_4310,N_3468,N_3804);
nor U4311 (N_4311,N_3795,N_3442);
or U4312 (N_4312,N_2822,N_3636);
and U4313 (N_4313,N_3348,N_3465);
or U4314 (N_4314,N_2764,N_2613);
xor U4315 (N_4315,N_2602,N_2006);
nand U4316 (N_4316,N_2507,N_3726);
and U4317 (N_4317,N_3861,N_3688);
xnor U4318 (N_4318,N_2030,N_3787);
nor U4319 (N_4319,N_3538,N_3729);
and U4320 (N_4320,N_3451,N_3477);
nand U4321 (N_4321,N_2065,N_3104);
and U4322 (N_4322,N_2145,N_2136);
xnor U4323 (N_4323,N_3612,N_2018);
and U4324 (N_4324,N_3767,N_2577);
and U4325 (N_4325,N_2286,N_2654);
xnor U4326 (N_4326,N_3888,N_2896);
xnor U4327 (N_4327,N_3829,N_2237);
and U4328 (N_4328,N_2798,N_3889);
nand U4329 (N_4329,N_2300,N_3327);
nor U4330 (N_4330,N_2211,N_2543);
nor U4331 (N_4331,N_2915,N_3546);
and U4332 (N_4332,N_3898,N_3345);
and U4333 (N_4333,N_3258,N_2526);
nor U4334 (N_4334,N_3833,N_2687);
or U4335 (N_4335,N_2994,N_3047);
nand U4336 (N_4336,N_2364,N_2515);
xor U4337 (N_4337,N_2333,N_3716);
nand U4338 (N_4338,N_2919,N_2656);
xor U4339 (N_4339,N_3096,N_2246);
xor U4340 (N_4340,N_3666,N_3478);
or U4341 (N_4341,N_3781,N_2124);
xnor U4342 (N_4342,N_3613,N_2144);
nor U4343 (N_4343,N_2342,N_2872);
nor U4344 (N_4344,N_2624,N_3435);
nand U4345 (N_4345,N_2341,N_3176);
or U4346 (N_4346,N_3487,N_2165);
nand U4347 (N_4347,N_3008,N_2917);
and U4348 (N_4348,N_3960,N_2829);
and U4349 (N_4349,N_2585,N_3816);
or U4350 (N_4350,N_3837,N_2886);
or U4351 (N_4351,N_2816,N_2057);
nand U4352 (N_4352,N_2390,N_3824);
nand U4353 (N_4353,N_2086,N_3841);
and U4354 (N_4354,N_2031,N_3615);
nand U4355 (N_4355,N_2975,N_3321);
and U4356 (N_4356,N_3675,N_2828);
or U4357 (N_4357,N_3073,N_2265);
xor U4358 (N_4358,N_3308,N_3673);
and U4359 (N_4359,N_3049,N_2413);
nor U4360 (N_4360,N_3984,N_3407);
nand U4361 (N_4361,N_2276,N_3523);
nor U4362 (N_4362,N_3440,N_3430);
nor U4363 (N_4363,N_2529,N_2153);
nor U4364 (N_4364,N_2379,N_2214);
xnor U4365 (N_4365,N_3654,N_3059);
nor U4366 (N_4366,N_3244,N_2358);
nand U4367 (N_4367,N_3602,N_3062);
and U4368 (N_4368,N_3328,N_2599);
and U4369 (N_4369,N_3809,N_3857);
and U4370 (N_4370,N_2967,N_2783);
or U4371 (N_4371,N_2433,N_2357);
xnor U4372 (N_4372,N_2556,N_3149);
xnor U4373 (N_4373,N_3532,N_2090);
nand U4374 (N_4374,N_3239,N_2600);
and U4375 (N_4375,N_2303,N_3770);
nand U4376 (N_4376,N_2438,N_3294);
and U4377 (N_4377,N_2632,N_2007);
nor U4378 (N_4378,N_3628,N_3171);
nand U4379 (N_4379,N_2693,N_2400);
nand U4380 (N_4380,N_2126,N_2178);
or U4381 (N_4381,N_3521,N_3993);
xor U4382 (N_4382,N_2448,N_3856);
nand U4383 (N_4383,N_2569,N_3843);
nand U4384 (N_4384,N_2259,N_3563);
or U4385 (N_4385,N_2204,N_3964);
xnor U4386 (N_4386,N_2747,N_3760);
or U4387 (N_4387,N_3880,N_2558);
xor U4388 (N_4388,N_3117,N_2369);
and U4389 (N_4389,N_3930,N_2137);
nor U4390 (N_4390,N_3363,N_3035);
xor U4391 (N_4391,N_3923,N_2659);
xor U4392 (N_4392,N_2081,N_2147);
xor U4393 (N_4393,N_3971,N_3314);
xnor U4394 (N_4394,N_2499,N_3033);
nand U4395 (N_4395,N_2371,N_2969);
nor U4396 (N_4396,N_2426,N_2988);
or U4397 (N_4397,N_2261,N_3082);
nor U4398 (N_4398,N_2808,N_2156);
nor U4399 (N_4399,N_3500,N_2325);
nor U4400 (N_4400,N_2269,N_2116);
nand U4401 (N_4401,N_2707,N_2594);
and U4402 (N_4402,N_3303,N_2845);
and U4403 (N_4403,N_3166,N_3812);
and U4404 (N_4404,N_3907,N_2314);
xor U4405 (N_4405,N_3081,N_2038);
nor U4406 (N_4406,N_3126,N_3512);
nand U4407 (N_4407,N_3609,N_3932);
xor U4408 (N_4408,N_2373,N_3014);
xnor U4409 (N_4409,N_2759,N_3682);
nand U4410 (N_4410,N_3307,N_2824);
nor U4411 (N_4411,N_2834,N_3863);
or U4412 (N_4412,N_2485,N_3805);
xnor U4413 (N_4413,N_2549,N_2351);
nand U4414 (N_4414,N_2425,N_3341);
or U4415 (N_4415,N_3138,N_3006);
or U4416 (N_4416,N_2723,N_2019);
and U4417 (N_4417,N_3370,N_2498);
nor U4418 (N_4418,N_2819,N_3246);
nor U4419 (N_4419,N_2283,N_3958);
nor U4420 (N_4420,N_3542,N_2162);
and U4421 (N_4421,N_2841,N_3170);
or U4422 (N_4422,N_2097,N_3565);
xor U4423 (N_4423,N_2833,N_2532);
nand U4424 (N_4424,N_2731,N_3133);
or U4425 (N_4425,N_3638,N_3179);
nand U4426 (N_4426,N_3663,N_3518);
and U4427 (N_4427,N_2669,N_2772);
or U4428 (N_4428,N_3101,N_2104);
nand U4429 (N_4429,N_2457,N_3631);
nor U4430 (N_4430,N_2648,N_2451);
and U4431 (N_4431,N_2101,N_2974);
xor U4432 (N_4432,N_3398,N_2541);
nor U4433 (N_4433,N_2366,N_2720);
nand U4434 (N_4434,N_2738,N_2022);
or U4435 (N_4435,N_3141,N_3568);
xor U4436 (N_4436,N_3210,N_2428);
or U4437 (N_4437,N_3742,N_3146);
or U4438 (N_4438,N_2858,N_2548);
or U4439 (N_4439,N_3319,N_3540);
nor U4440 (N_4440,N_2471,N_2870);
nor U4441 (N_4441,N_3206,N_3895);
xnor U4442 (N_4442,N_3952,N_2588);
xnor U4443 (N_4443,N_2001,N_3691);
and U4444 (N_4444,N_2976,N_3010);
xor U4445 (N_4445,N_2068,N_3224);
nor U4446 (N_4446,N_2430,N_3265);
nand U4447 (N_4447,N_3130,N_2508);
and U4448 (N_4448,N_2034,N_2119);
or U4449 (N_4449,N_3625,N_2598);
and U4450 (N_4450,N_2570,N_3237);
and U4451 (N_4451,N_2207,N_3337);
and U4452 (N_4452,N_3846,N_3873);
or U4453 (N_4453,N_2721,N_3693);
and U4454 (N_4454,N_3092,N_2143);
nand U4455 (N_4455,N_3678,N_2906);
and U4456 (N_4456,N_3755,N_3570);
nor U4457 (N_4457,N_3394,N_3966);
nand U4458 (N_4458,N_2181,N_3746);
xnor U4459 (N_4459,N_3524,N_3998);
nor U4460 (N_4460,N_2866,N_2024);
or U4461 (N_4461,N_2452,N_3789);
and U4462 (N_4462,N_2608,N_3980);
nand U4463 (N_4463,N_2830,N_3180);
xnor U4464 (N_4464,N_2345,N_2513);
nor U4465 (N_4465,N_2417,N_3514);
and U4466 (N_4466,N_2391,N_3175);
xnor U4467 (N_4467,N_2198,N_2696);
xor U4468 (N_4468,N_3354,N_3994);
and U4469 (N_4469,N_2761,N_2270);
and U4470 (N_4470,N_3041,N_3447);
or U4471 (N_4471,N_2409,N_2083);
and U4472 (N_4472,N_3469,N_3400);
or U4473 (N_4473,N_3576,N_3368);
nor U4474 (N_4474,N_2395,N_3968);
and U4475 (N_4475,N_2540,N_3097);
nand U4476 (N_4476,N_3845,N_2134);
or U4477 (N_4477,N_2932,N_2378);
or U4478 (N_4478,N_2827,N_3937);
or U4479 (N_4479,N_3277,N_3528);
and U4480 (N_4480,N_3174,N_2551);
or U4481 (N_4481,N_2232,N_2981);
xnor U4482 (N_4482,N_2978,N_3456);
nand U4483 (N_4483,N_3943,N_2744);
xor U4484 (N_4484,N_3738,N_2852);
or U4485 (N_4485,N_3128,N_3910);
and U4486 (N_4486,N_2574,N_2523);
nand U4487 (N_4487,N_3234,N_3428);
xnor U4488 (N_4488,N_2444,N_2601);
xnor U4489 (N_4489,N_2704,N_2701);
and U4490 (N_4490,N_3536,N_3173);
and U4491 (N_4491,N_2490,N_2055);
and U4492 (N_4492,N_3087,N_3758);
nand U4493 (N_4493,N_3385,N_2338);
nand U4494 (N_4494,N_3586,N_3186);
nand U4495 (N_4495,N_2859,N_3199);
nand U4496 (N_4496,N_2831,N_2218);
nor U4497 (N_4497,N_3916,N_3718);
xor U4498 (N_4498,N_3222,N_2948);
nand U4499 (N_4499,N_2628,N_2790);
nand U4500 (N_4500,N_3461,N_2386);
or U4501 (N_4501,N_3706,N_2133);
xnor U4502 (N_4502,N_2152,N_3708);
xor U4503 (N_4503,N_2804,N_2135);
nor U4504 (N_4504,N_3797,N_3821);
and U4505 (N_4505,N_2809,N_3508);
xor U4506 (N_4506,N_2109,N_2356);
xnor U4507 (N_4507,N_3367,N_2487);
nor U4508 (N_4508,N_3957,N_3501);
nand U4509 (N_4509,N_2971,N_3656);
nand U4510 (N_4510,N_3921,N_2329);
or U4511 (N_4511,N_2676,N_2050);
xnor U4512 (N_4512,N_3036,N_2653);
nor U4513 (N_4513,N_3901,N_3162);
and U4514 (N_4514,N_2475,N_2179);
and U4515 (N_4515,N_3086,N_3715);
nor U4516 (N_4516,N_3649,N_3003);
nor U4517 (N_4517,N_3581,N_2175);
or U4518 (N_4518,N_3920,N_3438);
nor U4519 (N_4519,N_3079,N_3431);
or U4520 (N_4520,N_2651,N_2187);
and U4521 (N_4521,N_3973,N_3748);
or U4522 (N_4522,N_2423,N_3948);
nand U4523 (N_4523,N_3858,N_2168);
and U4524 (N_4524,N_3323,N_3967);
nand U4525 (N_4525,N_2346,N_3623);
or U4526 (N_4526,N_3739,N_3346);
nand U4527 (N_4527,N_2014,N_3262);
or U4528 (N_4528,N_2719,N_3472);
xnor U4529 (N_4529,N_2231,N_3881);
or U4530 (N_4530,N_2581,N_2972);
or U4531 (N_4531,N_2446,N_3590);
and U4532 (N_4532,N_2005,N_3839);
nor U4533 (N_4533,N_2715,N_3250);
nor U4534 (N_4534,N_3078,N_2335);
and U4535 (N_4535,N_3571,N_2713);
nand U4536 (N_4536,N_3263,N_2559);
xor U4537 (N_4537,N_3409,N_3124);
or U4538 (N_4538,N_2579,N_2512);
xnor U4539 (N_4539,N_2895,N_3735);
xnor U4540 (N_4540,N_3694,N_2614);
nor U4541 (N_4541,N_2909,N_2310);
xor U4542 (N_4542,N_2110,N_3306);
or U4543 (N_4543,N_2586,N_3458);
nand U4544 (N_4544,N_3148,N_2802);
xnor U4545 (N_4545,N_3712,N_2710);
or U4546 (N_4546,N_2312,N_3704);
or U4547 (N_4547,N_3360,N_2511);
nor U4548 (N_4548,N_3417,N_2571);
nor U4549 (N_4549,N_2027,N_3488);
nor U4550 (N_4550,N_2580,N_3305);
xor U4551 (N_4551,N_2668,N_3644);
nand U4552 (N_4552,N_3266,N_3061);
nor U4553 (N_4553,N_2029,N_2940);
or U4554 (N_4554,N_2750,N_3037);
xnor U4555 (N_4555,N_3953,N_2472);
or U4556 (N_4556,N_3187,N_3181);
nor U4557 (N_4557,N_3125,N_3353);
xnor U4558 (N_4558,N_2476,N_3775);
xnor U4559 (N_4559,N_3069,N_2869);
or U4560 (N_4560,N_3515,N_3316);
or U4561 (N_4561,N_2860,N_2367);
nand U4562 (N_4562,N_2437,N_2227);
xor U4563 (N_4563,N_3977,N_3744);
xnor U4564 (N_4564,N_2926,N_2424);
and U4565 (N_4565,N_3867,N_2557);
or U4566 (N_4566,N_3588,N_3031);
and U4567 (N_4567,N_2562,N_3992);
nand U4568 (N_4568,N_3420,N_2224);
nor U4569 (N_4569,N_2903,N_2724);
or U4570 (N_4570,N_2085,N_2730);
or U4571 (N_4571,N_3598,N_3249);
and U4572 (N_4572,N_3110,N_3765);
xnor U4573 (N_4573,N_3245,N_3641);
xor U4574 (N_4574,N_2780,N_3068);
or U4575 (N_4575,N_2241,N_2258);
or U4576 (N_4576,N_3876,N_3962);
or U4577 (N_4577,N_3449,N_2044);
nand U4578 (N_4578,N_3851,N_2826);
and U4579 (N_4579,N_3848,N_2810);
xor U4580 (N_4580,N_3332,N_3878);
and U4581 (N_4581,N_2786,N_3339);
nand U4582 (N_4582,N_2171,N_2757);
nand U4583 (N_4583,N_3752,N_2461);
or U4584 (N_4584,N_2525,N_2954);
xnor U4585 (N_4585,N_2478,N_3554);
nor U4586 (N_4586,N_2849,N_2228);
or U4587 (N_4587,N_3474,N_3899);
or U4588 (N_4588,N_2008,N_2679);
nand U4589 (N_4589,N_2125,N_3221);
xor U4590 (N_4590,N_3485,N_3030);
and U4591 (N_4591,N_3701,N_3459);
or U4592 (N_4592,N_3949,N_2208);
and U4593 (N_4593,N_3392,N_2080);
xor U4594 (N_4594,N_3852,N_2662);
nand U4595 (N_4595,N_2322,N_2274);
xnor U4596 (N_4596,N_3711,N_3228);
nor U4597 (N_4597,N_3378,N_3302);
xnor U4598 (N_4598,N_3870,N_2706);
nand U4599 (N_4599,N_2219,N_2481);
or U4600 (N_4600,N_2911,N_3778);
or U4601 (N_4601,N_2297,N_3754);
and U4602 (N_4602,N_2944,N_3674);
xnor U4603 (N_4603,N_3820,N_2454);
xor U4604 (N_4604,N_2174,N_3396);
or U4605 (N_4605,N_2200,N_2623);
nand U4606 (N_4606,N_2900,N_3593);
xnor U4607 (N_4607,N_3988,N_3847);
nand U4608 (N_4608,N_3556,N_3768);
nand U4609 (N_4609,N_2650,N_2946);
nand U4610 (N_4610,N_3890,N_2323);
nand U4611 (N_4611,N_2054,N_3874);
nor U4612 (N_4612,N_2488,N_3896);
nor U4613 (N_4613,N_2046,N_3503);
or U4614 (N_4614,N_2445,N_2936);
nand U4615 (N_4615,N_2331,N_2319);
xor U4616 (N_4616,N_2340,N_3272);
xor U4617 (N_4617,N_2749,N_2088);
nor U4618 (N_4618,N_2714,N_3645);
nor U4619 (N_4619,N_3454,N_2035);
and U4620 (N_4620,N_2316,N_2460);
xnor U4621 (N_4621,N_2129,N_3077);
xor U4622 (N_4622,N_3105,N_3651);
nand U4623 (N_4623,N_3637,N_3929);
nor U4624 (N_4624,N_3679,N_2242);
and U4625 (N_4625,N_2421,N_2105);
or U4626 (N_4626,N_3886,N_2991);
nand U4627 (N_4627,N_3050,N_3364);
nand U4628 (N_4628,N_3750,N_2933);
and U4629 (N_4629,N_3642,N_2177);
xor U4630 (N_4630,N_3414,N_3702);
or U4631 (N_4631,N_2245,N_3381);
xor U4632 (N_4632,N_3183,N_3083);
or U4633 (N_4633,N_2658,N_3725);
xnor U4634 (N_4634,N_3055,N_3788);
xor U4635 (N_4635,N_2193,N_3121);
and U4636 (N_4636,N_3486,N_3552);
nand U4637 (N_4637,N_3564,N_3887);
or U4638 (N_4638,N_2510,N_3471);
xor U4639 (N_4639,N_2474,N_2247);
or U4640 (N_4640,N_2230,N_2477);
and U4641 (N_4641,N_3562,N_3408);
xnor U4642 (N_4642,N_2583,N_2740);
and U4643 (N_4643,N_3906,N_3457);
or U4644 (N_4644,N_2952,N_3286);
or U4645 (N_4645,N_2630,N_3558);
nor U4646 (N_4646,N_2665,N_3347);
or U4647 (N_4647,N_2493,N_2064);
nor U4648 (N_4648,N_2542,N_3925);
nand U4649 (N_4649,N_2003,N_2307);
and U4650 (N_4650,N_2122,N_3557);
xnor U4651 (N_4651,N_2040,N_3703);
nand U4652 (N_4652,N_2349,N_3351);
nor U4653 (N_4653,N_2725,N_3762);
nand U4654 (N_4654,N_3630,N_2130);
xor U4655 (N_4655,N_3189,N_2036);
nand U4656 (N_4656,N_2756,N_2631);
xor U4657 (N_4657,N_2192,N_2215);
xnor U4658 (N_4658,N_3161,N_3713);
or U4659 (N_4659,N_2671,N_2611);
nor U4660 (N_4660,N_3260,N_2443);
xor U4661 (N_4661,N_2590,N_2977);
xnor U4662 (N_4662,N_2832,N_2818);
xnor U4663 (N_4663,N_3089,N_3032);
and U4664 (N_4664,N_2294,N_3803);
nor U4665 (N_4665,N_2127,N_3278);
nand U4666 (N_4666,N_3559,N_3042);
nand U4667 (N_4667,N_2203,N_2053);
nand U4668 (N_4668,N_3209,N_2466);
and U4669 (N_4669,N_3692,N_2550);
nand U4670 (N_4670,N_3892,N_3777);
nand U4671 (N_4671,N_2092,N_3029);
xor U4672 (N_4672,N_2752,N_3312);
xnor U4673 (N_4673,N_3317,N_3448);
or U4674 (N_4674,N_3473,N_3057);
and U4675 (N_4675,N_2142,N_3267);
nand U4676 (N_4676,N_3950,N_3596);
and U4677 (N_4677,N_3256,N_3517);
nand U4678 (N_4678,N_3759,N_2778);
or U4679 (N_4679,N_2695,N_3320);
xnor U4680 (N_4680,N_2106,N_3646);
xnor U4681 (N_4681,N_3919,N_2762);
nand U4682 (N_4682,N_2882,N_3167);
xor U4683 (N_4683,N_3842,N_2985);
and U4684 (N_4684,N_3940,N_2716);
or U4685 (N_4685,N_3480,N_2938);
and U4686 (N_4686,N_2839,N_3840);
nor U4687 (N_4687,N_3080,N_3802);
and U4688 (N_4688,N_2643,N_3389);
nand U4689 (N_4689,N_3441,N_2642);
nand U4690 (N_4690,N_2617,N_2099);
and U4691 (N_4691,N_3261,N_3216);
nand U4692 (N_4692,N_3380,N_3727);
or U4693 (N_4693,N_2591,N_3529);
and U4694 (N_4694,N_3996,N_3671);
xnor U4695 (N_4695,N_2209,N_2025);
and U4696 (N_4696,N_3411,N_2043);
xnor U4697 (N_4697,N_3935,N_2252);
and U4698 (N_4698,N_2392,N_3178);
and U4699 (N_4699,N_2982,N_3142);
nor U4700 (N_4700,N_3790,N_3119);
nor U4701 (N_4701,N_2486,N_3311);
or U4702 (N_4702,N_2327,N_3811);
and U4703 (N_4703,N_2533,N_3058);
and U4704 (N_4704,N_3502,N_2530);
xor U4705 (N_4705,N_3835,N_2857);
and U4706 (N_4706,N_2646,N_3419);
and U4707 (N_4707,N_3490,N_3611);
xor U4708 (N_4708,N_2059,N_3695);
nand U4709 (N_4709,N_2470,N_2815);
nand U4710 (N_4710,N_2482,N_2873);
nor U4711 (N_4711,N_2368,N_3395);
or U4712 (N_4712,N_2694,N_3201);
or U4713 (N_4713,N_2604,N_3574);
or U4714 (N_4714,N_2792,N_2262);
nand U4715 (N_4715,N_3731,N_3108);
nand U4716 (N_4716,N_2060,N_3567);
nor U4717 (N_4717,N_2899,N_3723);
and U4718 (N_4718,N_3643,N_3470);
xnor U4719 (N_4719,N_2383,N_2161);
xor U4720 (N_4720,N_2930,N_3961);
or U4721 (N_4721,N_2277,N_2045);
nand U4722 (N_4722,N_2941,N_2387);
and U4723 (N_4723,N_3743,N_3090);
xnor U4724 (N_4724,N_2260,N_2291);
xor U4725 (N_4725,N_2595,N_2743);
and U4726 (N_4726,N_3991,N_2500);
xor U4727 (N_4727,N_3854,N_2406);
or U4728 (N_4728,N_2382,N_3818);
xnor U4729 (N_4729,N_3550,N_3028);
and U4730 (N_4730,N_2459,N_3513);
or U4731 (N_4731,N_2880,N_3070);
nand U4732 (N_4732,N_2893,N_3893);
xor U4733 (N_4733,N_3527,N_3763);
and U4734 (N_4734,N_3295,N_3102);
nor U4735 (N_4735,N_2660,N_3826);
and U4736 (N_4736,N_2618,N_2282);
or U4737 (N_4737,N_3927,N_3009);
and U4738 (N_4738,N_2593,N_2992);
or U4739 (N_4739,N_2115,N_3914);
nand U4740 (N_4740,N_2821,N_2958);
or U4741 (N_4741,N_3203,N_3293);
nand U4742 (N_4742,N_2879,N_3926);
or U4743 (N_4743,N_3882,N_2502);
or U4744 (N_4744,N_2912,N_2666);
nand U4745 (N_4745,N_2160,N_2352);
nand U4746 (N_4746,N_2244,N_2285);
nand U4747 (N_4747,N_2004,N_2491);
xor U4748 (N_4748,N_2146,N_2979);
or U4749 (N_4749,N_2132,N_2375);
xor U4750 (N_4750,N_3350,N_2170);
and U4751 (N_4751,N_3202,N_3580);
xnor U4752 (N_4752,N_3808,N_3191);
and U4753 (N_4753,N_2271,N_2684);
xor U4754 (N_4754,N_2700,N_3801);
nand U4755 (N_4755,N_2095,N_2483);
and U4756 (N_4756,N_3872,N_3340);
nor U4757 (N_4757,N_2063,N_3954);
nor U4758 (N_4758,N_2196,N_3677);
and U4759 (N_4759,N_3099,N_3147);
and U4760 (N_4760,N_3198,N_2305);
and U4761 (N_4761,N_2420,N_2464);
or U4762 (N_4762,N_2644,N_2878);
nor U4763 (N_4763,N_3056,N_2902);
and U4764 (N_4764,N_3043,N_2348);
xor U4765 (N_4765,N_3997,N_3525);
nand U4766 (N_4766,N_2537,N_3052);
nor U4767 (N_4767,N_2456,N_3730);
or U4768 (N_4768,N_3421,N_3690);
nand U4769 (N_4769,N_3021,N_2397);
nor U4770 (N_4770,N_3255,N_2544);
nand U4771 (N_4771,N_3879,N_2120);
or U4772 (N_4772,N_3807,N_3114);
and U4773 (N_4773,N_3547,N_2949);
nor U4774 (N_4774,N_2516,N_3664);
or U4775 (N_4775,N_2336,N_3292);
nor U4776 (N_4776,N_3123,N_3749);
or U4777 (N_4777,N_3208,N_3869);
nor U4778 (N_4778,N_2505,N_3956);
or U4779 (N_4779,N_2465,N_2173);
and U4780 (N_4780,N_3905,N_3728);
or U4781 (N_4781,N_2250,N_3134);
and U4782 (N_4782,N_2503,N_2567);
nor U4783 (N_4783,N_3680,N_3724);
nand U4784 (N_4784,N_3717,N_3129);
xor U4785 (N_4785,N_3970,N_2856);
nand U4786 (N_4786,N_3023,N_3902);
and U4787 (N_4787,N_2836,N_2066);
xnor U4788 (N_4788,N_2691,N_3650);
xnor U4789 (N_4789,N_3001,N_2414);
nand U4790 (N_4790,N_2047,N_3230);
nor U4791 (N_4791,N_3719,N_2753);
and U4792 (N_4792,N_2148,N_3371);
nor U4793 (N_4793,N_3155,N_2403);
xnor U4794 (N_4794,N_2251,N_3284);
or U4795 (N_4795,N_2070,N_2301);
or U4796 (N_4796,N_3668,N_3152);
or U4797 (N_4797,N_3426,N_2190);
or U4798 (N_4798,N_3115,N_2973);
and U4799 (N_4799,N_3172,N_3462);
or U4800 (N_4800,N_2195,N_2221);
nand U4801 (N_4801,N_3780,N_3424);
and U4802 (N_4802,N_3700,N_2956);
nand U4803 (N_4803,N_3939,N_2999);
or U4804 (N_4804,N_2254,N_3463);
or U4805 (N_4805,N_2797,N_3535);
xnor U4806 (N_4806,N_2017,N_3497);
nor U4807 (N_4807,N_2184,N_3555);
xnor U4808 (N_4808,N_3946,N_3632);
or U4809 (N_4809,N_3504,N_2089);
or U4810 (N_4810,N_2672,N_3624);
or U4811 (N_4811,N_2914,N_3761);
nor U4812 (N_4812,N_2514,N_3270);
nand U4813 (N_4813,N_3066,N_2326);
xor U4814 (N_4814,N_2411,N_2494);
nand U4815 (N_4815,N_2520,N_3834);
nand U4816 (N_4816,N_3566,N_3756);
xnor U4817 (N_4817,N_3150,N_2606);
nor U4818 (N_4818,N_2049,N_2212);
or U4819 (N_4819,N_3509,N_2957);
or U4820 (N_4820,N_3931,N_3018);
and U4821 (N_4821,N_3194,N_3776);
nor U4822 (N_4822,N_3537,N_2052);
xor U4823 (N_4823,N_2784,N_3046);
nor U4824 (N_4824,N_3158,N_2324);
and U4825 (N_4825,N_3483,N_2566);
or U4826 (N_4826,N_3044,N_3520);
and U4827 (N_4827,N_3289,N_3352);
or U4828 (N_4828,N_2418,N_3207);
and U4829 (N_4829,N_3785,N_3227);
nand U4830 (N_4830,N_3197,N_3118);
nor U4831 (N_4831,N_2518,N_2398);
nor U4832 (N_4832,N_2610,N_2296);
or U4833 (N_4833,N_2287,N_3275);
xor U4834 (N_4834,N_2222,N_2138);
and U4835 (N_4835,N_3707,N_3553);
nand U4836 (N_4836,N_2377,N_3865);
and U4837 (N_4837,N_3017,N_2084);
xor U4838 (N_4838,N_2686,N_2205);
nor U4839 (N_4839,N_3591,N_3607);
nand U4840 (N_4840,N_2965,N_3000);
or U4841 (N_4841,N_2289,N_2890);
and U4842 (N_4842,N_3437,N_3627);
xor U4843 (N_4843,N_2621,N_2793);
or U4844 (N_4844,N_2848,N_2937);
nor U4845 (N_4845,N_2048,N_2534);
nor U4846 (N_4846,N_2267,N_2898);
nand U4847 (N_4847,N_3494,N_3476);
nor U4848 (N_4848,N_2056,N_3579);
nor U4849 (N_4849,N_3999,N_2468);
xor U4850 (N_4850,N_2393,N_2951);
xor U4851 (N_4851,N_3067,N_3548);
nand U4852 (N_4852,N_2627,N_3026);
nor U4853 (N_4853,N_2572,N_3884);
nand U4854 (N_4854,N_3639,N_2748);
or U4855 (N_4855,N_3614,N_2155);
nor U4856 (N_4856,N_3534,N_3200);
nor U4857 (N_4857,N_2388,N_2746);
and U4858 (N_4858,N_2734,N_2149);
nand U4859 (N_4859,N_2993,N_3779);
xnor U4860 (N_4860,N_2435,N_2921);
xor U4861 (N_4861,N_2087,N_3629);
nand U4862 (N_4862,N_3257,N_3681);
nand U4863 (N_4863,N_2563,N_2359);
nor U4864 (N_4864,N_3622,N_2299);
nor U4865 (N_4865,N_3357,N_3122);
nand U4866 (N_4866,N_3362,N_3220);
or U4867 (N_4867,N_3287,N_2041);
nand U4868 (N_4868,N_2419,N_3252);
and U4869 (N_4869,N_3784,N_2874);
or U4870 (N_4870,N_3683,N_2293);
and U4871 (N_4871,N_2114,N_3386);
xor U4872 (N_4872,N_3696,N_2489);
and U4873 (N_4873,N_3040,N_2225);
and U4874 (N_4874,N_3894,N_3343);
xor U4875 (N_4875,N_2028,N_3154);
nand U4876 (N_4876,N_2955,N_3185);
nand U4877 (N_4877,N_2840,N_3945);
xor U4878 (N_4878,N_3071,N_2760);
and U4879 (N_4879,N_2664,N_3296);
nor U4880 (N_4880,N_3669,N_3281);
or U4881 (N_4881,N_3329,N_3423);
and U4882 (N_4882,N_2249,N_3794);
nand U4883 (N_4883,N_2863,N_2243);
nor U4884 (N_4884,N_3156,N_3832);
nor U4885 (N_4885,N_2990,N_2067);
nor U4886 (N_4886,N_3626,N_2281);
or U4887 (N_4887,N_2699,N_2163);
and U4888 (N_4888,N_3814,N_2883);
nand U4889 (N_4889,N_3388,N_3965);
nand U4890 (N_4890,N_2825,N_2539);
xor U4891 (N_4891,N_3214,N_2907);
nor U4892 (N_4892,N_3361,N_2077);
and U4893 (N_4893,N_3601,N_3094);
nor U4894 (N_4894,N_3972,N_2370);
xnor U4895 (N_4895,N_2210,N_2151);
nand U4896 (N_4896,N_2309,N_3510);
or U4897 (N_4897,N_2449,N_3193);
nor U4898 (N_4898,N_2350,N_3686);
nand U4899 (N_4899,N_3710,N_3658);
and U4900 (N_4900,N_2381,N_3577);
and U4901 (N_4901,N_2755,N_3484);
or U4902 (N_4902,N_2536,N_3493);
nand U4903 (N_4903,N_2039,N_2180);
and U4904 (N_4904,N_3020,N_3229);
nor U4905 (N_4905,N_3433,N_3131);
xnor U4906 (N_4906,N_3575,N_2023);
and U4907 (N_4907,N_3334,N_3076);
nand U4908 (N_4908,N_2321,N_3838);
nand U4909 (N_4909,N_3384,N_2372);
nand U4910 (N_4910,N_3495,N_2922);
or U4911 (N_4911,N_2620,N_3075);
xor U4912 (N_4912,N_2892,N_3551);
or U4913 (N_4913,N_2609,N_3990);
and U4914 (N_4914,N_3103,N_2256);
and U4915 (N_4915,N_2683,N_2501);
or U4916 (N_4916,N_2186,N_2266);
nand U4917 (N_4917,N_2788,N_3745);
nand U4918 (N_4918,N_3519,N_3608);
xnor U4919 (N_4919,N_2389,N_2708);
nor U4920 (N_4920,N_3324,N_2837);
nor U4921 (N_4921,N_3439,N_3866);
or U4922 (N_4922,N_2354,N_3844);
nor U4923 (N_4923,N_2680,N_3093);
xnor U4924 (N_4924,N_2020,N_3410);
and U4925 (N_4925,N_3791,N_3975);
or U4926 (N_4926,N_2458,N_2202);
xor U4927 (N_4927,N_2767,N_3810);
xor U4928 (N_4928,N_2855,N_3734);
or U4929 (N_4929,N_2657,N_2191);
nor U4930 (N_4930,N_3432,N_3549);
or U4931 (N_4931,N_2552,N_3903);
and U4932 (N_4932,N_3618,N_2947);
xor U4933 (N_4933,N_3309,N_3464);
xnor U4934 (N_4934,N_2519,N_3806);
nand U4935 (N_4935,N_3709,N_3849);
or U4936 (N_4936,N_2589,N_3610);
xnor U4937 (N_4937,N_3764,N_3620);
xor U4938 (N_4938,N_2197,N_2587);
and U4939 (N_4939,N_3951,N_3113);
or U4940 (N_4940,N_2442,N_3499);
nand U4941 (N_4941,N_2431,N_3597);
nand U4942 (N_4942,N_2275,N_3799);
nand U4943 (N_4943,N_3545,N_3355);
nand U4944 (N_4944,N_2480,N_2189);
xnor U4945 (N_4945,N_2506,N_2576);
nor U4946 (N_4946,N_3402,N_3648);
nor U4947 (N_4947,N_3657,N_3376);
nor U4948 (N_4948,N_3232,N_2108);
and U4949 (N_4949,N_3383,N_2861);
and U4950 (N_4950,N_3783,N_2823);
nand U4951 (N_4951,N_2560,N_2223);
or U4952 (N_4952,N_2416,N_2037);
and U4953 (N_4953,N_3165,N_2141);
xor U4954 (N_4954,N_2347,N_3911);
or U4955 (N_4955,N_3569,N_3027);
or U4956 (N_4956,N_3373,N_3374);
xor U4957 (N_4957,N_2545,N_3192);
nor U4958 (N_4958,N_2935,N_2555);
nand U4959 (N_4959,N_2320,N_3670);
nand U4960 (N_4960,N_3196,N_3025);
nor U4961 (N_4961,N_2998,N_3982);
and U4962 (N_4962,N_3425,N_3205);
and U4963 (N_4963,N_3541,N_2806);
and U4964 (N_4964,N_3979,N_3522);
or U4965 (N_4965,N_3450,N_3883);
or U4966 (N_4966,N_3689,N_2078);
and U4967 (N_4967,N_2741,N_3177);
nand U4968 (N_4968,N_2677,N_3342);
nand U4969 (N_4969,N_2774,N_3372);
nand U4970 (N_4970,N_2279,N_3561);
and U4971 (N_4971,N_2524,N_2009);
or U4972 (N_4972,N_2636,N_2929);
nor U4973 (N_4973,N_2061,N_3403);
or U4974 (N_4974,N_3699,N_2240);
or U4975 (N_4975,N_2399,N_3405);
or U4976 (N_4976,N_3963,N_3460);
nand U4977 (N_4977,N_2742,N_3412);
and U4978 (N_4978,N_2450,N_2455);
or U4979 (N_4979,N_2263,N_2980);
nor U4980 (N_4980,N_3827,N_3792);
nor U4981 (N_4981,N_2652,N_3254);
nor U4982 (N_4982,N_2918,N_2111);
nor U4983 (N_4983,N_2681,N_3647);
xor U4984 (N_4984,N_3506,N_2607);
or U4985 (N_4985,N_2467,N_2093);
nand U4986 (N_4986,N_3379,N_3434);
nor U4987 (N_4987,N_2439,N_3012);
xnor U4988 (N_4988,N_2984,N_2934);
and U4989 (N_4989,N_3505,N_3640);
or U4990 (N_4990,N_2894,N_3942);
nand U4991 (N_4991,N_2733,N_3007);
or U4992 (N_4992,N_3315,N_3243);
nand U4993 (N_4993,N_2776,N_3862);
nor U4994 (N_4994,N_2779,N_3813);
nand U4995 (N_4995,N_2339,N_2789);
nor U4996 (N_4996,N_3013,N_3299);
nor U4997 (N_4997,N_3279,N_3584);
and U4998 (N_4998,N_3589,N_3422);
nor U4999 (N_4999,N_2315,N_3828);
nand U5000 (N_5000,N_2834,N_2334);
nand U5001 (N_5001,N_2599,N_3589);
or U5002 (N_5002,N_2605,N_2825);
nand U5003 (N_5003,N_2583,N_2161);
xor U5004 (N_5004,N_2421,N_2661);
nand U5005 (N_5005,N_3242,N_3311);
or U5006 (N_5006,N_2748,N_3455);
or U5007 (N_5007,N_3169,N_3184);
nand U5008 (N_5008,N_2270,N_2194);
or U5009 (N_5009,N_2479,N_2365);
and U5010 (N_5010,N_2944,N_2924);
xor U5011 (N_5011,N_2429,N_2301);
nor U5012 (N_5012,N_3258,N_2252);
nand U5013 (N_5013,N_3886,N_2645);
xor U5014 (N_5014,N_2331,N_2459);
nand U5015 (N_5015,N_2394,N_3754);
or U5016 (N_5016,N_3721,N_2368);
nand U5017 (N_5017,N_3258,N_3357);
xor U5018 (N_5018,N_3809,N_3437);
nor U5019 (N_5019,N_2922,N_3060);
nand U5020 (N_5020,N_3486,N_2589);
and U5021 (N_5021,N_3833,N_3703);
and U5022 (N_5022,N_3214,N_2006);
nand U5023 (N_5023,N_3374,N_3487);
or U5024 (N_5024,N_2554,N_2752);
or U5025 (N_5025,N_3187,N_2650);
xor U5026 (N_5026,N_3488,N_3364);
nor U5027 (N_5027,N_3619,N_3214);
or U5028 (N_5028,N_3316,N_3335);
nor U5029 (N_5029,N_2217,N_3469);
or U5030 (N_5030,N_2340,N_2798);
nand U5031 (N_5031,N_3446,N_3328);
and U5032 (N_5032,N_3788,N_2973);
xor U5033 (N_5033,N_3333,N_2917);
nand U5034 (N_5034,N_2221,N_2926);
xnor U5035 (N_5035,N_3126,N_2538);
nand U5036 (N_5036,N_3530,N_3738);
nor U5037 (N_5037,N_3667,N_3482);
and U5038 (N_5038,N_3689,N_3917);
nand U5039 (N_5039,N_2526,N_3594);
or U5040 (N_5040,N_2518,N_3139);
nand U5041 (N_5041,N_2322,N_3702);
nor U5042 (N_5042,N_3406,N_2159);
and U5043 (N_5043,N_2371,N_2261);
nand U5044 (N_5044,N_2053,N_2192);
and U5045 (N_5045,N_2178,N_2252);
and U5046 (N_5046,N_3438,N_3159);
xnor U5047 (N_5047,N_3008,N_2045);
xnor U5048 (N_5048,N_2366,N_2562);
nor U5049 (N_5049,N_3075,N_3174);
nand U5050 (N_5050,N_2406,N_3964);
or U5051 (N_5051,N_2375,N_2247);
and U5052 (N_5052,N_3725,N_3527);
and U5053 (N_5053,N_3596,N_2980);
xnor U5054 (N_5054,N_3471,N_3428);
nand U5055 (N_5055,N_2263,N_2637);
and U5056 (N_5056,N_3326,N_2047);
xnor U5057 (N_5057,N_2225,N_3446);
nor U5058 (N_5058,N_2203,N_2504);
nand U5059 (N_5059,N_2713,N_3970);
nand U5060 (N_5060,N_2863,N_2803);
nor U5061 (N_5061,N_3239,N_3834);
nand U5062 (N_5062,N_2891,N_2706);
and U5063 (N_5063,N_2647,N_3738);
or U5064 (N_5064,N_2319,N_2158);
and U5065 (N_5065,N_2143,N_3221);
nor U5066 (N_5066,N_2050,N_3719);
nand U5067 (N_5067,N_3248,N_3679);
or U5068 (N_5068,N_3023,N_3226);
xnor U5069 (N_5069,N_2916,N_2069);
and U5070 (N_5070,N_2166,N_2186);
and U5071 (N_5071,N_3176,N_2551);
or U5072 (N_5072,N_2505,N_2904);
nor U5073 (N_5073,N_3581,N_3436);
or U5074 (N_5074,N_3099,N_2145);
nor U5075 (N_5075,N_2888,N_3988);
and U5076 (N_5076,N_2315,N_3425);
nand U5077 (N_5077,N_2418,N_2928);
nand U5078 (N_5078,N_2257,N_3862);
or U5079 (N_5079,N_3017,N_3202);
nand U5080 (N_5080,N_2303,N_3923);
or U5081 (N_5081,N_3250,N_2729);
or U5082 (N_5082,N_2015,N_3433);
xnor U5083 (N_5083,N_3169,N_3276);
nor U5084 (N_5084,N_2449,N_2787);
and U5085 (N_5085,N_2529,N_3926);
and U5086 (N_5086,N_3615,N_3244);
or U5087 (N_5087,N_2117,N_3416);
nor U5088 (N_5088,N_3189,N_2209);
or U5089 (N_5089,N_2138,N_3303);
nand U5090 (N_5090,N_3196,N_3356);
and U5091 (N_5091,N_3407,N_2139);
and U5092 (N_5092,N_3826,N_3638);
nand U5093 (N_5093,N_2390,N_2465);
nor U5094 (N_5094,N_3042,N_3563);
xnor U5095 (N_5095,N_3050,N_3268);
nor U5096 (N_5096,N_3885,N_2233);
nand U5097 (N_5097,N_2779,N_3505);
xnor U5098 (N_5098,N_2043,N_2778);
nor U5099 (N_5099,N_3259,N_3994);
or U5100 (N_5100,N_3112,N_3421);
nor U5101 (N_5101,N_3825,N_3167);
xnor U5102 (N_5102,N_2954,N_2178);
xnor U5103 (N_5103,N_3634,N_2988);
and U5104 (N_5104,N_2175,N_3348);
and U5105 (N_5105,N_2346,N_2235);
nand U5106 (N_5106,N_3098,N_2830);
or U5107 (N_5107,N_2053,N_3555);
or U5108 (N_5108,N_2332,N_3598);
nand U5109 (N_5109,N_2689,N_3420);
nand U5110 (N_5110,N_2098,N_2314);
nand U5111 (N_5111,N_2371,N_3683);
or U5112 (N_5112,N_2141,N_3022);
nor U5113 (N_5113,N_3914,N_2951);
nand U5114 (N_5114,N_2195,N_2836);
xor U5115 (N_5115,N_2472,N_2119);
nor U5116 (N_5116,N_3661,N_3976);
nor U5117 (N_5117,N_2478,N_3596);
xor U5118 (N_5118,N_2974,N_3289);
xor U5119 (N_5119,N_3531,N_3550);
nand U5120 (N_5120,N_2665,N_2859);
or U5121 (N_5121,N_3748,N_2249);
xor U5122 (N_5122,N_3222,N_3909);
and U5123 (N_5123,N_2095,N_2306);
and U5124 (N_5124,N_2085,N_3430);
or U5125 (N_5125,N_2648,N_2782);
and U5126 (N_5126,N_2454,N_3560);
or U5127 (N_5127,N_3028,N_2458);
nor U5128 (N_5128,N_3598,N_3242);
nand U5129 (N_5129,N_2669,N_3191);
or U5130 (N_5130,N_3594,N_2413);
xnor U5131 (N_5131,N_2296,N_2329);
nor U5132 (N_5132,N_3645,N_3545);
and U5133 (N_5133,N_3570,N_3890);
xor U5134 (N_5134,N_3639,N_3070);
and U5135 (N_5135,N_2520,N_3125);
nor U5136 (N_5136,N_3175,N_3448);
and U5137 (N_5137,N_3821,N_2440);
nor U5138 (N_5138,N_3405,N_2518);
and U5139 (N_5139,N_3402,N_2799);
nand U5140 (N_5140,N_3547,N_2348);
and U5141 (N_5141,N_2367,N_2286);
nor U5142 (N_5142,N_2599,N_3829);
nor U5143 (N_5143,N_3303,N_3083);
nor U5144 (N_5144,N_3957,N_3970);
and U5145 (N_5145,N_3152,N_2831);
nand U5146 (N_5146,N_3069,N_2249);
and U5147 (N_5147,N_2207,N_3191);
and U5148 (N_5148,N_3864,N_3062);
and U5149 (N_5149,N_2972,N_3573);
or U5150 (N_5150,N_2454,N_2726);
xnor U5151 (N_5151,N_3290,N_2644);
and U5152 (N_5152,N_2657,N_3026);
or U5153 (N_5153,N_2835,N_2209);
nand U5154 (N_5154,N_2608,N_2120);
nand U5155 (N_5155,N_3060,N_3337);
xor U5156 (N_5156,N_2438,N_3195);
nor U5157 (N_5157,N_2283,N_3960);
or U5158 (N_5158,N_3776,N_2709);
or U5159 (N_5159,N_2652,N_2379);
or U5160 (N_5160,N_3103,N_2094);
nand U5161 (N_5161,N_2360,N_3185);
and U5162 (N_5162,N_2096,N_2810);
or U5163 (N_5163,N_2537,N_3325);
and U5164 (N_5164,N_3186,N_2384);
nand U5165 (N_5165,N_3308,N_3509);
nor U5166 (N_5166,N_2073,N_3868);
nand U5167 (N_5167,N_3639,N_2961);
nand U5168 (N_5168,N_2714,N_2801);
nand U5169 (N_5169,N_2051,N_3788);
nor U5170 (N_5170,N_2598,N_2253);
and U5171 (N_5171,N_3210,N_3387);
and U5172 (N_5172,N_2369,N_2478);
or U5173 (N_5173,N_3503,N_2594);
nand U5174 (N_5174,N_3053,N_2932);
nor U5175 (N_5175,N_3481,N_2281);
and U5176 (N_5176,N_3992,N_3675);
nand U5177 (N_5177,N_2929,N_2208);
xnor U5178 (N_5178,N_2956,N_3550);
nand U5179 (N_5179,N_2062,N_2918);
or U5180 (N_5180,N_3635,N_3057);
and U5181 (N_5181,N_3249,N_2578);
nor U5182 (N_5182,N_3574,N_3488);
nor U5183 (N_5183,N_2072,N_3995);
and U5184 (N_5184,N_3182,N_2385);
xor U5185 (N_5185,N_3419,N_3590);
nand U5186 (N_5186,N_2758,N_3496);
nor U5187 (N_5187,N_2429,N_3384);
and U5188 (N_5188,N_3462,N_2534);
and U5189 (N_5189,N_3952,N_2701);
xnor U5190 (N_5190,N_2480,N_2664);
and U5191 (N_5191,N_2094,N_2910);
xnor U5192 (N_5192,N_2668,N_2994);
nor U5193 (N_5193,N_2652,N_2829);
or U5194 (N_5194,N_2044,N_3927);
nor U5195 (N_5195,N_2562,N_3515);
and U5196 (N_5196,N_2714,N_3277);
nand U5197 (N_5197,N_2418,N_3120);
nand U5198 (N_5198,N_2688,N_3122);
nor U5199 (N_5199,N_2526,N_2613);
xor U5200 (N_5200,N_3252,N_2647);
or U5201 (N_5201,N_3643,N_3971);
and U5202 (N_5202,N_3402,N_3217);
and U5203 (N_5203,N_2322,N_2992);
or U5204 (N_5204,N_2928,N_2338);
xnor U5205 (N_5205,N_3000,N_2709);
or U5206 (N_5206,N_3861,N_2583);
xnor U5207 (N_5207,N_3318,N_2790);
nor U5208 (N_5208,N_3140,N_2909);
and U5209 (N_5209,N_3277,N_3228);
xor U5210 (N_5210,N_3290,N_3563);
or U5211 (N_5211,N_2755,N_2859);
xnor U5212 (N_5212,N_3445,N_2437);
xnor U5213 (N_5213,N_3577,N_2351);
nor U5214 (N_5214,N_2223,N_3802);
nand U5215 (N_5215,N_2111,N_2063);
nand U5216 (N_5216,N_3482,N_2962);
xnor U5217 (N_5217,N_3648,N_3124);
nand U5218 (N_5218,N_3636,N_2917);
nor U5219 (N_5219,N_2093,N_3408);
nand U5220 (N_5220,N_2815,N_3454);
or U5221 (N_5221,N_3920,N_3756);
and U5222 (N_5222,N_2427,N_3964);
nand U5223 (N_5223,N_2039,N_3354);
xnor U5224 (N_5224,N_2843,N_2128);
or U5225 (N_5225,N_2192,N_3177);
nor U5226 (N_5226,N_3414,N_2275);
nand U5227 (N_5227,N_3559,N_3333);
and U5228 (N_5228,N_3186,N_2007);
nand U5229 (N_5229,N_3388,N_3328);
nand U5230 (N_5230,N_2804,N_2166);
nor U5231 (N_5231,N_2290,N_3413);
nor U5232 (N_5232,N_2794,N_2323);
xnor U5233 (N_5233,N_2961,N_2206);
and U5234 (N_5234,N_2511,N_3079);
and U5235 (N_5235,N_2389,N_2907);
xnor U5236 (N_5236,N_3269,N_2644);
nand U5237 (N_5237,N_3557,N_2769);
nand U5238 (N_5238,N_3835,N_3439);
xnor U5239 (N_5239,N_2571,N_3211);
nand U5240 (N_5240,N_3949,N_2306);
nor U5241 (N_5241,N_3540,N_3524);
nor U5242 (N_5242,N_3082,N_2820);
nor U5243 (N_5243,N_2097,N_2669);
nor U5244 (N_5244,N_2949,N_3208);
nor U5245 (N_5245,N_2389,N_2541);
or U5246 (N_5246,N_2380,N_3077);
nand U5247 (N_5247,N_2514,N_3172);
nand U5248 (N_5248,N_3396,N_3694);
nor U5249 (N_5249,N_2621,N_2178);
or U5250 (N_5250,N_2759,N_2738);
nand U5251 (N_5251,N_3787,N_2210);
nor U5252 (N_5252,N_3991,N_2174);
xnor U5253 (N_5253,N_2946,N_2233);
or U5254 (N_5254,N_3667,N_2258);
nand U5255 (N_5255,N_2104,N_2370);
xnor U5256 (N_5256,N_3519,N_3726);
or U5257 (N_5257,N_3530,N_3950);
nor U5258 (N_5258,N_2867,N_2838);
nor U5259 (N_5259,N_2476,N_2377);
nand U5260 (N_5260,N_3973,N_2873);
or U5261 (N_5261,N_3355,N_3319);
xor U5262 (N_5262,N_3639,N_3814);
nand U5263 (N_5263,N_2941,N_2287);
and U5264 (N_5264,N_3926,N_2914);
xnor U5265 (N_5265,N_2879,N_3955);
nand U5266 (N_5266,N_3443,N_3319);
nand U5267 (N_5267,N_2910,N_3927);
or U5268 (N_5268,N_2438,N_3058);
nor U5269 (N_5269,N_2196,N_3230);
and U5270 (N_5270,N_3910,N_3657);
nor U5271 (N_5271,N_2964,N_3871);
nand U5272 (N_5272,N_3767,N_2694);
nor U5273 (N_5273,N_3952,N_3558);
or U5274 (N_5274,N_2292,N_3953);
nand U5275 (N_5275,N_3903,N_3773);
or U5276 (N_5276,N_3872,N_3353);
nor U5277 (N_5277,N_2323,N_3520);
xnor U5278 (N_5278,N_2763,N_2007);
nor U5279 (N_5279,N_3144,N_2348);
xor U5280 (N_5280,N_3536,N_2026);
or U5281 (N_5281,N_2421,N_2937);
or U5282 (N_5282,N_3410,N_2838);
nor U5283 (N_5283,N_2363,N_2648);
nor U5284 (N_5284,N_3982,N_3208);
nand U5285 (N_5285,N_3280,N_3959);
xnor U5286 (N_5286,N_3266,N_2087);
xor U5287 (N_5287,N_2473,N_3554);
xor U5288 (N_5288,N_3777,N_2810);
nand U5289 (N_5289,N_3827,N_3540);
nand U5290 (N_5290,N_3957,N_3592);
xor U5291 (N_5291,N_3456,N_2797);
nor U5292 (N_5292,N_3010,N_3711);
and U5293 (N_5293,N_3632,N_3565);
xor U5294 (N_5294,N_3787,N_3651);
nand U5295 (N_5295,N_3015,N_2584);
nand U5296 (N_5296,N_2233,N_3553);
or U5297 (N_5297,N_2239,N_3647);
nand U5298 (N_5298,N_2452,N_2540);
nor U5299 (N_5299,N_3777,N_2656);
xnor U5300 (N_5300,N_2144,N_3598);
and U5301 (N_5301,N_2936,N_2908);
or U5302 (N_5302,N_2174,N_2265);
xnor U5303 (N_5303,N_3492,N_3941);
xor U5304 (N_5304,N_2710,N_2928);
nor U5305 (N_5305,N_2262,N_3097);
xnor U5306 (N_5306,N_3056,N_2919);
xnor U5307 (N_5307,N_3529,N_3510);
or U5308 (N_5308,N_2981,N_2703);
and U5309 (N_5309,N_3988,N_3784);
nor U5310 (N_5310,N_2849,N_3170);
nor U5311 (N_5311,N_2871,N_3251);
or U5312 (N_5312,N_3654,N_2996);
or U5313 (N_5313,N_3424,N_2828);
xnor U5314 (N_5314,N_3497,N_3855);
or U5315 (N_5315,N_2992,N_2924);
and U5316 (N_5316,N_2977,N_2580);
nor U5317 (N_5317,N_2003,N_2533);
xor U5318 (N_5318,N_2583,N_3057);
xnor U5319 (N_5319,N_2163,N_3766);
or U5320 (N_5320,N_3178,N_2564);
nand U5321 (N_5321,N_2916,N_2146);
or U5322 (N_5322,N_3491,N_2803);
nand U5323 (N_5323,N_2870,N_2130);
and U5324 (N_5324,N_3094,N_2509);
and U5325 (N_5325,N_2439,N_2261);
nand U5326 (N_5326,N_3981,N_3857);
xnor U5327 (N_5327,N_2241,N_3466);
nor U5328 (N_5328,N_2303,N_2051);
nor U5329 (N_5329,N_3356,N_3800);
or U5330 (N_5330,N_2334,N_3852);
or U5331 (N_5331,N_2023,N_2824);
and U5332 (N_5332,N_2213,N_2893);
nand U5333 (N_5333,N_2414,N_3270);
and U5334 (N_5334,N_3427,N_2162);
nor U5335 (N_5335,N_3613,N_3837);
or U5336 (N_5336,N_2111,N_2186);
or U5337 (N_5337,N_2886,N_2786);
xor U5338 (N_5338,N_2529,N_3022);
or U5339 (N_5339,N_3273,N_3461);
xnor U5340 (N_5340,N_3401,N_3992);
xnor U5341 (N_5341,N_2750,N_3166);
and U5342 (N_5342,N_3459,N_2656);
and U5343 (N_5343,N_3991,N_2949);
nor U5344 (N_5344,N_3314,N_2016);
nor U5345 (N_5345,N_3202,N_3868);
xnor U5346 (N_5346,N_2122,N_3017);
or U5347 (N_5347,N_3394,N_2863);
xor U5348 (N_5348,N_3544,N_2642);
xnor U5349 (N_5349,N_2391,N_3399);
and U5350 (N_5350,N_2016,N_2524);
and U5351 (N_5351,N_3859,N_2534);
nand U5352 (N_5352,N_3662,N_2012);
nand U5353 (N_5353,N_3765,N_3142);
nor U5354 (N_5354,N_2730,N_3030);
xnor U5355 (N_5355,N_2620,N_3874);
nand U5356 (N_5356,N_3083,N_2765);
nor U5357 (N_5357,N_2711,N_2488);
and U5358 (N_5358,N_3917,N_2822);
nand U5359 (N_5359,N_2261,N_2877);
or U5360 (N_5360,N_2483,N_3289);
nor U5361 (N_5361,N_3361,N_2063);
and U5362 (N_5362,N_2002,N_2894);
nor U5363 (N_5363,N_2369,N_2413);
nor U5364 (N_5364,N_3135,N_3890);
and U5365 (N_5365,N_3258,N_3983);
nor U5366 (N_5366,N_2276,N_3980);
and U5367 (N_5367,N_3009,N_2900);
nor U5368 (N_5368,N_3349,N_2915);
xnor U5369 (N_5369,N_3153,N_3374);
nor U5370 (N_5370,N_3524,N_3624);
xor U5371 (N_5371,N_3079,N_3597);
xor U5372 (N_5372,N_2002,N_2859);
nor U5373 (N_5373,N_3373,N_3110);
xnor U5374 (N_5374,N_2093,N_2820);
or U5375 (N_5375,N_2242,N_2899);
xnor U5376 (N_5376,N_2803,N_2230);
xnor U5377 (N_5377,N_2689,N_2356);
or U5378 (N_5378,N_3875,N_3653);
or U5379 (N_5379,N_3891,N_3164);
and U5380 (N_5380,N_2779,N_3226);
nor U5381 (N_5381,N_3743,N_3987);
or U5382 (N_5382,N_3867,N_2258);
nand U5383 (N_5383,N_2185,N_3121);
and U5384 (N_5384,N_3990,N_3068);
xnor U5385 (N_5385,N_3913,N_2876);
nor U5386 (N_5386,N_2727,N_3129);
nand U5387 (N_5387,N_3918,N_2382);
nor U5388 (N_5388,N_3902,N_3943);
xnor U5389 (N_5389,N_2387,N_2561);
and U5390 (N_5390,N_3187,N_2819);
xor U5391 (N_5391,N_2841,N_3736);
nand U5392 (N_5392,N_3525,N_2615);
nor U5393 (N_5393,N_3214,N_3705);
or U5394 (N_5394,N_2605,N_3202);
nand U5395 (N_5395,N_2633,N_2041);
xnor U5396 (N_5396,N_3792,N_2398);
nor U5397 (N_5397,N_2621,N_3108);
nand U5398 (N_5398,N_2236,N_2201);
nand U5399 (N_5399,N_2469,N_3013);
xnor U5400 (N_5400,N_2292,N_2195);
xnor U5401 (N_5401,N_2839,N_2108);
or U5402 (N_5402,N_3820,N_2330);
or U5403 (N_5403,N_3550,N_3843);
xnor U5404 (N_5404,N_2684,N_2417);
nand U5405 (N_5405,N_3256,N_3254);
xor U5406 (N_5406,N_3216,N_3016);
or U5407 (N_5407,N_3337,N_2144);
nor U5408 (N_5408,N_3216,N_3036);
nor U5409 (N_5409,N_2927,N_3469);
and U5410 (N_5410,N_3907,N_2543);
and U5411 (N_5411,N_3251,N_2512);
or U5412 (N_5412,N_3303,N_2449);
and U5413 (N_5413,N_2919,N_2789);
xnor U5414 (N_5414,N_2450,N_2608);
xnor U5415 (N_5415,N_2961,N_2221);
nand U5416 (N_5416,N_2607,N_2008);
and U5417 (N_5417,N_2722,N_3706);
and U5418 (N_5418,N_2692,N_2261);
and U5419 (N_5419,N_2002,N_2855);
nor U5420 (N_5420,N_2219,N_2445);
nand U5421 (N_5421,N_2076,N_2711);
xnor U5422 (N_5422,N_3952,N_2921);
xnor U5423 (N_5423,N_2863,N_2763);
xor U5424 (N_5424,N_2041,N_3494);
xor U5425 (N_5425,N_2240,N_2248);
nor U5426 (N_5426,N_2574,N_2930);
or U5427 (N_5427,N_3462,N_3525);
nor U5428 (N_5428,N_2325,N_2679);
xnor U5429 (N_5429,N_3846,N_3975);
or U5430 (N_5430,N_2738,N_2135);
nor U5431 (N_5431,N_3958,N_3001);
nor U5432 (N_5432,N_3944,N_3744);
nor U5433 (N_5433,N_2257,N_3737);
xnor U5434 (N_5434,N_2055,N_3173);
nand U5435 (N_5435,N_3748,N_3175);
or U5436 (N_5436,N_2469,N_2813);
or U5437 (N_5437,N_2870,N_3764);
and U5438 (N_5438,N_2539,N_3762);
and U5439 (N_5439,N_3322,N_3702);
nand U5440 (N_5440,N_2199,N_2894);
and U5441 (N_5441,N_2397,N_3777);
and U5442 (N_5442,N_2512,N_2872);
nand U5443 (N_5443,N_2883,N_3823);
xnor U5444 (N_5444,N_2760,N_3749);
xor U5445 (N_5445,N_3207,N_2624);
or U5446 (N_5446,N_2993,N_3161);
and U5447 (N_5447,N_3013,N_3327);
nor U5448 (N_5448,N_2295,N_3179);
nand U5449 (N_5449,N_3023,N_3985);
or U5450 (N_5450,N_3593,N_2649);
nor U5451 (N_5451,N_3782,N_3598);
nand U5452 (N_5452,N_2310,N_3351);
or U5453 (N_5453,N_3593,N_3019);
nand U5454 (N_5454,N_3564,N_2398);
xnor U5455 (N_5455,N_2753,N_2254);
nor U5456 (N_5456,N_2608,N_2504);
nand U5457 (N_5457,N_2451,N_3608);
nand U5458 (N_5458,N_3636,N_2667);
nand U5459 (N_5459,N_3341,N_2867);
nand U5460 (N_5460,N_3671,N_3216);
nand U5461 (N_5461,N_3744,N_3807);
nor U5462 (N_5462,N_3356,N_2011);
nand U5463 (N_5463,N_2595,N_3609);
and U5464 (N_5464,N_3280,N_3821);
nand U5465 (N_5465,N_3946,N_3853);
nor U5466 (N_5466,N_3672,N_3764);
and U5467 (N_5467,N_2351,N_3710);
xnor U5468 (N_5468,N_2613,N_2376);
nand U5469 (N_5469,N_2289,N_3149);
nand U5470 (N_5470,N_3394,N_2963);
nand U5471 (N_5471,N_3922,N_2687);
xnor U5472 (N_5472,N_2537,N_2574);
nor U5473 (N_5473,N_3683,N_3859);
nand U5474 (N_5474,N_3158,N_2479);
xnor U5475 (N_5475,N_3053,N_2885);
nand U5476 (N_5476,N_2015,N_2652);
nor U5477 (N_5477,N_2010,N_3832);
or U5478 (N_5478,N_2929,N_3949);
nand U5479 (N_5479,N_3679,N_3767);
nand U5480 (N_5480,N_3863,N_3626);
nor U5481 (N_5481,N_2374,N_2129);
nand U5482 (N_5482,N_2883,N_2260);
nor U5483 (N_5483,N_2014,N_3994);
or U5484 (N_5484,N_3520,N_3684);
or U5485 (N_5485,N_2029,N_2378);
nand U5486 (N_5486,N_3655,N_3786);
nor U5487 (N_5487,N_3884,N_2994);
xnor U5488 (N_5488,N_3653,N_2194);
nor U5489 (N_5489,N_2038,N_2250);
nor U5490 (N_5490,N_2162,N_2345);
and U5491 (N_5491,N_3564,N_3206);
nor U5492 (N_5492,N_2501,N_2668);
or U5493 (N_5493,N_3175,N_2272);
or U5494 (N_5494,N_2518,N_2691);
nor U5495 (N_5495,N_2005,N_2278);
xnor U5496 (N_5496,N_3172,N_3538);
or U5497 (N_5497,N_2337,N_3744);
nor U5498 (N_5498,N_3606,N_3865);
nor U5499 (N_5499,N_3939,N_3203);
nor U5500 (N_5500,N_2653,N_3195);
and U5501 (N_5501,N_2435,N_2968);
nor U5502 (N_5502,N_3384,N_2251);
nor U5503 (N_5503,N_3714,N_2816);
nand U5504 (N_5504,N_2657,N_2973);
or U5505 (N_5505,N_2167,N_3445);
nor U5506 (N_5506,N_2006,N_3691);
nand U5507 (N_5507,N_2993,N_3418);
or U5508 (N_5508,N_2497,N_2978);
nand U5509 (N_5509,N_2037,N_3746);
and U5510 (N_5510,N_2467,N_2618);
and U5511 (N_5511,N_3937,N_2700);
nand U5512 (N_5512,N_3971,N_2409);
xor U5513 (N_5513,N_2770,N_2708);
nand U5514 (N_5514,N_3466,N_2597);
and U5515 (N_5515,N_3442,N_3710);
nand U5516 (N_5516,N_3947,N_3917);
nand U5517 (N_5517,N_3491,N_3197);
nand U5518 (N_5518,N_2432,N_2132);
xor U5519 (N_5519,N_2723,N_3515);
or U5520 (N_5520,N_2679,N_3156);
or U5521 (N_5521,N_3132,N_2018);
and U5522 (N_5522,N_2729,N_3145);
nand U5523 (N_5523,N_3324,N_3478);
or U5524 (N_5524,N_2923,N_3680);
nand U5525 (N_5525,N_3497,N_2842);
nand U5526 (N_5526,N_2180,N_2815);
and U5527 (N_5527,N_2158,N_2920);
xor U5528 (N_5528,N_3302,N_2632);
nand U5529 (N_5529,N_3586,N_2081);
xnor U5530 (N_5530,N_3545,N_3959);
or U5531 (N_5531,N_3917,N_2888);
xnor U5532 (N_5532,N_2894,N_3656);
and U5533 (N_5533,N_3447,N_2666);
and U5534 (N_5534,N_3051,N_2295);
xor U5535 (N_5535,N_2033,N_3342);
xnor U5536 (N_5536,N_2452,N_3552);
nand U5537 (N_5537,N_3659,N_2988);
nor U5538 (N_5538,N_2682,N_2140);
and U5539 (N_5539,N_3693,N_3749);
xor U5540 (N_5540,N_3177,N_3134);
nor U5541 (N_5541,N_2741,N_3759);
and U5542 (N_5542,N_3560,N_3928);
or U5543 (N_5543,N_2774,N_2072);
nand U5544 (N_5544,N_3147,N_3284);
xnor U5545 (N_5545,N_2833,N_3320);
nand U5546 (N_5546,N_2908,N_3113);
xor U5547 (N_5547,N_3671,N_2091);
or U5548 (N_5548,N_3148,N_2836);
nor U5549 (N_5549,N_3490,N_3581);
xnor U5550 (N_5550,N_3386,N_2222);
and U5551 (N_5551,N_3874,N_2572);
or U5552 (N_5552,N_2902,N_2538);
xor U5553 (N_5553,N_3940,N_3850);
or U5554 (N_5554,N_2911,N_3747);
or U5555 (N_5555,N_3208,N_3688);
nor U5556 (N_5556,N_2227,N_3646);
xnor U5557 (N_5557,N_2447,N_3933);
and U5558 (N_5558,N_2375,N_3143);
nand U5559 (N_5559,N_3986,N_2560);
nor U5560 (N_5560,N_3897,N_2824);
or U5561 (N_5561,N_2436,N_3928);
nand U5562 (N_5562,N_2153,N_3768);
nor U5563 (N_5563,N_3218,N_2390);
or U5564 (N_5564,N_2868,N_3515);
or U5565 (N_5565,N_2472,N_3742);
nand U5566 (N_5566,N_3412,N_2629);
xor U5567 (N_5567,N_2635,N_3679);
or U5568 (N_5568,N_3382,N_2856);
and U5569 (N_5569,N_3874,N_2025);
and U5570 (N_5570,N_2467,N_3102);
nor U5571 (N_5571,N_2552,N_2302);
nand U5572 (N_5572,N_3484,N_2305);
nand U5573 (N_5573,N_3492,N_3212);
xor U5574 (N_5574,N_3999,N_3686);
and U5575 (N_5575,N_3869,N_2547);
or U5576 (N_5576,N_3834,N_3483);
nor U5577 (N_5577,N_3230,N_2610);
nand U5578 (N_5578,N_2905,N_2041);
nor U5579 (N_5579,N_3737,N_2730);
and U5580 (N_5580,N_3022,N_3117);
or U5581 (N_5581,N_2146,N_2007);
xnor U5582 (N_5582,N_2571,N_3065);
and U5583 (N_5583,N_3035,N_3702);
nor U5584 (N_5584,N_3494,N_3839);
xor U5585 (N_5585,N_3822,N_2905);
or U5586 (N_5586,N_2880,N_3722);
xnor U5587 (N_5587,N_3949,N_2373);
nor U5588 (N_5588,N_2383,N_3853);
nor U5589 (N_5589,N_2204,N_3871);
xor U5590 (N_5590,N_3116,N_2652);
or U5591 (N_5591,N_2209,N_3970);
nand U5592 (N_5592,N_3044,N_2345);
nand U5593 (N_5593,N_2280,N_3703);
nor U5594 (N_5594,N_3562,N_2091);
nor U5595 (N_5595,N_2037,N_2905);
nand U5596 (N_5596,N_2296,N_2218);
and U5597 (N_5597,N_3376,N_3206);
nand U5598 (N_5598,N_3275,N_2104);
and U5599 (N_5599,N_2131,N_2180);
xor U5600 (N_5600,N_2863,N_2297);
or U5601 (N_5601,N_2522,N_3751);
nand U5602 (N_5602,N_2351,N_3935);
nand U5603 (N_5603,N_2266,N_2069);
or U5604 (N_5604,N_3930,N_2044);
nor U5605 (N_5605,N_2078,N_2506);
or U5606 (N_5606,N_2432,N_2848);
nor U5607 (N_5607,N_3781,N_2711);
xor U5608 (N_5608,N_3149,N_2953);
xnor U5609 (N_5609,N_2138,N_2327);
or U5610 (N_5610,N_3776,N_2938);
and U5611 (N_5611,N_2302,N_3538);
xnor U5612 (N_5612,N_2108,N_2870);
nand U5613 (N_5613,N_2933,N_3990);
nor U5614 (N_5614,N_2942,N_2681);
xor U5615 (N_5615,N_2288,N_2715);
nor U5616 (N_5616,N_2261,N_2342);
nand U5617 (N_5617,N_2607,N_2881);
and U5618 (N_5618,N_2179,N_3123);
or U5619 (N_5619,N_3807,N_2117);
nor U5620 (N_5620,N_3055,N_2888);
nand U5621 (N_5621,N_2400,N_3963);
nor U5622 (N_5622,N_3409,N_3611);
xnor U5623 (N_5623,N_3215,N_2376);
nor U5624 (N_5624,N_2799,N_3806);
xnor U5625 (N_5625,N_2182,N_2256);
or U5626 (N_5626,N_3393,N_3676);
nor U5627 (N_5627,N_2546,N_3974);
nand U5628 (N_5628,N_2682,N_3776);
nor U5629 (N_5629,N_2379,N_2012);
and U5630 (N_5630,N_3878,N_3061);
nor U5631 (N_5631,N_2001,N_2154);
and U5632 (N_5632,N_3402,N_3364);
and U5633 (N_5633,N_2708,N_3646);
nand U5634 (N_5634,N_2676,N_2260);
nand U5635 (N_5635,N_2841,N_2111);
or U5636 (N_5636,N_3487,N_3019);
nand U5637 (N_5637,N_3983,N_2982);
and U5638 (N_5638,N_3772,N_2108);
and U5639 (N_5639,N_3160,N_3214);
or U5640 (N_5640,N_2985,N_2961);
xor U5641 (N_5641,N_2882,N_2748);
and U5642 (N_5642,N_3637,N_3669);
nand U5643 (N_5643,N_3993,N_2238);
nor U5644 (N_5644,N_2653,N_3816);
xnor U5645 (N_5645,N_2130,N_3868);
and U5646 (N_5646,N_3260,N_3332);
nor U5647 (N_5647,N_2603,N_3450);
xor U5648 (N_5648,N_3605,N_2576);
or U5649 (N_5649,N_3878,N_2741);
or U5650 (N_5650,N_3780,N_3804);
and U5651 (N_5651,N_3540,N_2380);
nand U5652 (N_5652,N_3035,N_2023);
or U5653 (N_5653,N_2590,N_2518);
nor U5654 (N_5654,N_2626,N_3060);
or U5655 (N_5655,N_3238,N_3203);
xnor U5656 (N_5656,N_2927,N_3676);
or U5657 (N_5657,N_2144,N_3307);
nor U5658 (N_5658,N_2639,N_2190);
nand U5659 (N_5659,N_3588,N_3209);
xor U5660 (N_5660,N_2120,N_3766);
and U5661 (N_5661,N_3458,N_3270);
nor U5662 (N_5662,N_3288,N_2924);
or U5663 (N_5663,N_3535,N_3285);
xor U5664 (N_5664,N_2594,N_2705);
and U5665 (N_5665,N_2219,N_2148);
nand U5666 (N_5666,N_2999,N_2567);
xor U5667 (N_5667,N_2039,N_2372);
and U5668 (N_5668,N_3573,N_3113);
xor U5669 (N_5669,N_3226,N_2688);
nand U5670 (N_5670,N_2970,N_3942);
or U5671 (N_5671,N_2279,N_3278);
nor U5672 (N_5672,N_2472,N_3607);
and U5673 (N_5673,N_2451,N_2365);
nor U5674 (N_5674,N_3253,N_2691);
xor U5675 (N_5675,N_2731,N_3152);
and U5676 (N_5676,N_2709,N_3958);
and U5677 (N_5677,N_2299,N_3117);
nor U5678 (N_5678,N_2657,N_3980);
nor U5679 (N_5679,N_2769,N_3304);
and U5680 (N_5680,N_3408,N_2632);
nand U5681 (N_5681,N_3446,N_2339);
or U5682 (N_5682,N_2332,N_3811);
or U5683 (N_5683,N_2245,N_2673);
or U5684 (N_5684,N_2559,N_3501);
and U5685 (N_5685,N_3539,N_3128);
nand U5686 (N_5686,N_2003,N_3861);
or U5687 (N_5687,N_2468,N_3085);
nand U5688 (N_5688,N_3981,N_3563);
nand U5689 (N_5689,N_2933,N_3526);
or U5690 (N_5690,N_3778,N_3979);
and U5691 (N_5691,N_3735,N_3688);
nor U5692 (N_5692,N_2269,N_2165);
nor U5693 (N_5693,N_3960,N_2272);
xor U5694 (N_5694,N_3949,N_2981);
xor U5695 (N_5695,N_3530,N_3519);
xor U5696 (N_5696,N_3879,N_3430);
nand U5697 (N_5697,N_3973,N_2709);
nand U5698 (N_5698,N_3674,N_2338);
xnor U5699 (N_5699,N_2025,N_2824);
or U5700 (N_5700,N_3559,N_3571);
or U5701 (N_5701,N_2469,N_3578);
xor U5702 (N_5702,N_2361,N_2006);
or U5703 (N_5703,N_3458,N_3943);
nor U5704 (N_5704,N_3041,N_3818);
xor U5705 (N_5705,N_3198,N_2675);
xnor U5706 (N_5706,N_2967,N_2768);
or U5707 (N_5707,N_3840,N_3138);
and U5708 (N_5708,N_3934,N_2807);
nor U5709 (N_5709,N_3567,N_3698);
and U5710 (N_5710,N_3343,N_3915);
nand U5711 (N_5711,N_3737,N_3766);
and U5712 (N_5712,N_3435,N_3805);
nand U5713 (N_5713,N_2812,N_2493);
nand U5714 (N_5714,N_3027,N_2045);
nor U5715 (N_5715,N_2252,N_3475);
or U5716 (N_5716,N_2569,N_2022);
or U5717 (N_5717,N_3058,N_2712);
or U5718 (N_5718,N_3984,N_2933);
xnor U5719 (N_5719,N_2561,N_3134);
nor U5720 (N_5720,N_2193,N_2342);
nand U5721 (N_5721,N_2199,N_3713);
nand U5722 (N_5722,N_3224,N_3601);
or U5723 (N_5723,N_2137,N_2987);
and U5724 (N_5724,N_2903,N_2829);
xnor U5725 (N_5725,N_2894,N_3971);
nor U5726 (N_5726,N_2409,N_3020);
or U5727 (N_5727,N_2940,N_2348);
nor U5728 (N_5728,N_2459,N_2296);
and U5729 (N_5729,N_2410,N_3498);
or U5730 (N_5730,N_2019,N_3713);
nor U5731 (N_5731,N_2612,N_2793);
and U5732 (N_5732,N_3799,N_3786);
and U5733 (N_5733,N_2472,N_3513);
nand U5734 (N_5734,N_2407,N_3508);
xnor U5735 (N_5735,N_3599,N_2899);
and U5736 (N_5736,N_3824,N_2618);
xor U5737 (N_5737,N_3026,N_2170);
nor U5738 (N_5738,N_2430,N_3669);
nor U5739 (N_5739,N_3327,N_3681);
or U5740 (N_5740,N_3308,N_3505);
nor U5741 (N_5741,N_2863,N_2146);
nand U5742 (N_5742,N_2034,N_3288);
or U5743 (N_5743,N_3881,N_3401);
xnor U5744 (N_5744,N_2092,N_3073);
or U5745 (N_5745,N_3490,N_3485);
and U5746 (N_5746,N_2002,N_2987);
and U5747 (N_5747,N_3599,N_3836);
and U5748 (N_5748,N_2378,N_3923);
or U5749 (N_5749,N_2308,N_3709);
and U5750 (N_5750,N_2626,N_2571);
or U5751 (N_5751,N_3659,N_2144);
nand U5752 (N_5752,N_3002,N_2239);
or U5753 (N_5753,N_2402,N_2139);
or U5754 (N_5754,N_3756,N_2961);
xnor U5755 (N_5755,N_3161,N_2469);
or U5756 (N_5756,N_2194,N_3254);
xnor U5757 (N_5757,N_3338,N_3817);
xor U5758 (N_5758,N_3559,N_3636);
or U5759 (N_5759,N_2401,N_3760);
nor U5760 (N_5760,N_2264,N_3524);
nand U5761 (N_5761,N_3168,N_2983);
xor U5762 (N_5762,N_3616,N_2916);
xor U5763 (N_5763,N_2115,N_2736);
and U5764 (N_5764,N_2968,N_3349);
xnor U5765 (N_5765,N_3373,N_3462);
or U5766 (N_5766,N_3951,N_2672);
and U5767 (N_5767,N_2099,N_3759);
xnor U5768 (N_5768,N_3460,N_3178);
or U5769 (N_5769,N_3718,N_2831);
nor U5770 (N_5770,N_3152,N_2778);
xor U5771 (N_5771,N_3947,N_2613);
or U5772 (N_5772,N_3385,N_2139);
xnor U5773 (N_5773,N_2865,N_2402);
and U5774 (N_5774,N_2943,N_2511);
nor U5775 (N_5775,N_2097,N_3661);
nand U5776 (N_5776,N_3204,N_2262);
nand U5777 (N_5777,N_2903,N_2544);
nor U5778 (N_5778,N_2387,N_3410);
nand U5779 (N_5779,N_3589,N_3276);
nor U5780 (N_5780,N_2710,N_2110);
nand U5781 (N_5781,N_3270,N_3730);
nor U5782 (N_5782,N_3392,N_3779);
nand U5783 (N_5783,N_3981,N_2030);
nor U5784 (N_5784,N_2787,N_3669);
nor U5785 (N_5785,N_2626,N_2087);
or U5786 (N_5786,N_2074,N_2579);
xor U5787 (N_5787,N_3622,N_3235);
nor U5788 (N_5788,N_3237,N_2559);
and U5789 (N_5789,N_3214,N_2110);
xor U5790 (N_5790,N_2017,N_2520);
or U5791 (N_5791,N_3258,N_2824);
and U5792 (N_5792,N_2077,N_2229);
xor U5793 (N_5793,N_3027,N_2574);
or U5794 (N_5794,N_2287,N_2073);
nand U5795 (N_5795,N_2612,N_3243);
xor U5796 (N_5796,N_3837,N_2665);
and U5797 (N_5797,N_3123,N_2722);
and U5798 (N_5798,N_2705,N_3331);
xnor U5799 (N_5799,N_3532,N_2255);
and U5800 (N_5800,N_3153,N_2053);
and U5801 (N_5801,N_2260,N_3806);
nand U5802 (N_5802,N_3394,N_2710);
xnor U5803 (N_5803,N_2030,N_3337);
and U5804 (N_5804,N_2013,N_2649);
and U5805 (N_5805,N_2989,N_2116);
nand U5806 (N_5806,N_3280,N_3029);
nand U5807 (N_5807,N_3130,N_3595);
nor U5808 (N_5808,N_3160,N_3543);
nor U5809 (N_5809,N_2362,N_2497);
or U5810 (N_5810,N_3653,N_2756);
and U5811 (N_5811,N_3794,N_2259);
or U5812 (N_5812,N_2953,N_2972);
and U5813 (N_5813,N_2424,N_2761);
and U5814 (N_5814,N_3013,N_3684);
nand U5815 (N_5815,N_2392,N_2553);
nor U5816 (N_5816,N_3945,N_3749);
or U5817 (N_5817,N_2446,N_2740);
and U5818 (N_5818,N_2575,N_2842);
or U5819 (N_5819,N_2240,N_2814);
and U5820 (N_5820,N_2161,N_3564);
nor U5821 (N_5821,N_2688,N_3340);
nor U5822 (N_5822,N_2308,N_3484);
nor U5823 (N_5823,N_3045,N_2424);
nor U5824 (N_5824,N_3161,N_2394);
or U5825 (N_5825,N_2755,N_3134);
xor U5826 (N_5826,N_3035,N_2253);
and U5827 (N_5827,N_2609,N_3495);
or U5828 (N_5828,N_2709,N_2266);
or U5829 (N_5829,N_3011,N_2509);
nand U5830 (N_5830,N_2500,N_3484);
xnor U5831 (N_5831,N_2302,N_3711);
nand U5832 (N_5832,N_2982,N_3606);
nor U5833 (N_5833,N_2496,N_3588);
xnor U5834 (N_5834,N_3083,N_2595);
xor U5835 (N_5835,N_3653,N_3447);
nor U5836 (N_5836,N_2811,N_3990);
or U5837 (N_5837,N_2415,N_3981);
nand U5838 (N_5838,N_2714,N_3232);
xnor U5839 (N_5839,N_3412,N_3396);
or U5840 (N_5840,N_3167,N_3845);
xor U5841 (N_5841,N_2381,N_3302);
or U5842 (N_5842,N_2431,N_3593);
or U5843 (N_5843,N_2581,N_3946);
xnor U5844 (N_5844,N_3506,N_3233);
or U5845 (N_5845,N_3899,N_2687);
nand U5846 (N_5846,N_2379,N_3393);
or U5847 (N_5847,N_3711,N_3691);
or U5848 (N_5848,N_2687,N_3065);
nand U5849 (N_5849,N_2652,N_2590);
nor U5850 (N_5850,N_2129,N_2839);
or U5851 (N_5851,N_2864,N_3554);
xor U5852 (N_5852,N_2139,N_3867);
or U5853 (N_5853,N_3120,N_3332);
nand U5854 (N_5854,N_3720,N_3311);
and U5855 (N_5855,N_3711,N_3919);
nor U5856 (N_5856,N_2195,N_3232);
nor U5857 (N_5857,N_2959,N_2252);
or U5858 (N_5858,N_2705,N_3547);
or U5859 (N_5859,N_2923,N_2234);
nand U5860 (N_5860,N_2479,N_3794);
or U5861 (N_5861,N_3588,N_2408);
xnor U5862 (N_5862,N_3155,N_2737);
xor U5863 (N_5863,N_3203,N_2099);
nand U5864 (N_5864,N_2467,N_2940);
xor U5865 (N_5865,N_2157,N_3494);
xnor U5866 (N_5866,N_2614,N_2968);
or U5867 (N_5867,N_2379,N_2680);
or U5868 (N_5868,N_3291,N_3238);
nor U5869 (N_5869,N_2881,N_3145);
or U5870 (N_5870,N_3582,N_2756);
xor U5871 (N_5871,N_3978,N_3928);
xor U5872 (N_5872,N_3962,N_3008);
or U5873 (N_5873,N_3156,N_2711);
nand U5874 (N_5874,N_3083,N_2513);
xor U5875 (N_5875,N_3999,N_2435);
nand U5876 (N_5876,N_3353,N_2095);
or U5877 (N_5877,N_3611,N_3788);
or U5878 (N_5878,N_2982,N_3508);
nor U5879 (N_5879,N_3915,N_2423);
nor U5880 (N_5880,N_3917,N_2046);
or U5881 (N_5881,N_3674,N_2615);
or U5882 (N_5882,N_2873,N_2264);
nor U5883 (N_5883,N_3593,N_3793);
nand U5884 (N_5884,N_2842,N_2836);
nand U5885 (N_5885,N_2021,N_3528);
nor U5886 (N_5886,N_2440,N_2090);
nor U5887 (N_5887,N_2085,N_3669);
nor U5888 (N_5888,N_3219,N_2819);
or U5889 (N_5889,N_3617,N_2865);
nor U5890 (N_5890,N_2602,N_3561);
and U5891 (N_5891,N_2669,N_3502);
and U5892 (N_5892,N_2388,N_3042);
nand U5893 (N_5893,N_3185,N_2110);
and U5894 (N_5894,N_3698,N_2238);
nor U5895 (N_5895,N_3967,N_2113);
nor U5896 (N_5896,N_3945,N_2846);
or U5897 (N_5897,N_3614,N_2407);
nor U5898 (N_5898,N_2576,N_2280);
nand U5899 (N_5899,N_2005,N_3097);
xor U5900 (N_5900,N_3849,N_3051);
or U5901 (N_5901,N_3472,N_3578);
nand U5902 (N_5902,N_2128,N_2263);
and U5903 (N_5903,N_3163,N_2378);
xnor U5904 (N_5904,N_3701,N_2122);
xnor U5905 (N_5905,N_2546,N_3877);
nor U5906 (N_5906,N_2314,N_3175);
nand U5907 (N_5907,N_3008,N_3194);
nor U5908 (N_5908,N_2205,N_3904);
nor U5909 (N_5909,N_2166,N_2016);
nor U5910 (N_5910,N_2173,N_3490);
and U5911 (N_5911,N_2459,N_3824);
xnor U5912 (N_5912,N_2411,N_3221);
and U5913 (N_5913,N_2220,N_3044);
and U5914 (N_5914,N_3414,N_3711);
xnor U5915 (N_5915,N_3790,N_2185);
nand U5916 (N_5916,N_2652,N_2425);
nor U5917 (N_5917,N_3820,N_2877);
nor U5918 (N_5918,N_2283,N_3654);
nor U5919 (N_5919,N_2607,N_3422);
xor U5920 (N_5920,N_3509,N_2579);
xnor U5921 (N_5921,N_2880,N_2365);
xnor U5922 (N_5922,N_3728,N_3459);
nor U5923 (N_5923,N_3341,N_3478);
nor U5924 (N_5924,N_2905,N_2514);
xor U5925 (N_5925,N_2528,N_3091);
and U5926 (N_5926,N_3943,N_2436);
xor U5927 (N_5927,N_3999,N_3711);
and U5928 (N_5928,N_3344,N_3292);
and U5929 (N_5929,N_2830,N_2468);
nor U5930 (N_5930,N_3391,N_3221);
nand U5931 (N_5931,N_3811,N_2101);
and U5932 (N_5932,N_3612,N_2578);
nor U5933 (N_5933,N_2142,N_2918);
xor U5934 (N_5934,N_3679,N_3007);
nand U5935 (N_5935,N_3049,N_3208);
xor U5936 (N_5936,N_3792,N_3489);
nand U5937 (N_5937,N_3343,N_2034);
and U5938 (N_5938,N_2586,N_3339);
and U5939 (N_5939,N_2922,N_3478);
nor U5940 (N_5940,N_2395,N_2864);
nand U5941 (N_5941,N_3323,N_2795);
and U5942 (N_5942,N_3207,N_3684);
nor U5943 (N_5943,N_3846,N_3296);
xor U5944 (N_5944,N_3681,N_3960);
or U5945 (N_5945,N_2248,N_2127);
nor U5946 (N_5946,N_2379,N_3629);
nor U5947 (N_5947,N_3645,N_3349);
and U5948 (N_5948,N_2911,N_3943);
nor U5949 (N_5949,N_2782,N_3314);
and U5950 (N_5950,N_3869,N_2272);
xnor U5951 (N_5951,N_2161,N_3977);
nand U5952 (N_5952,N_3298,N_3213);
or U5953 (N_5953,N_3210,N_3487);
nand U5954 (N_5954,N_2503,N_3732);
nand U5955 (N_5955,N_2153,N_3114);
nor U5956 (N_5956,N_3545,N_3990);
and U5957 (N_5957,N_3602,N_2631);
xnor U5958 (N_5958,N_2047,N_2461);
and U5959 (N_5959,N_2705,N_2458);
nand U5960 (N_5960,N_2001,N_2138);
and U5961 (N_5961,N_2917,N_2233);
nand U5962 (N_5962,N_3662,N_2820);
and U5963 (N_5963,N_2602,N_3299);
or U5964 (N_5964,N_2862,N_2280);
nand U5965 (N_5965,N_2924,N_3513);
nor U5966 (N_5966,N_2943,N_2628);
nor U5967 (N_5967,N_2163,N_3675);
and U5968 (N_5968,N_2420,N_2463);
nor U5969 (N_5969,N_2197,N_2595);
xor U5970 (N_5970,N_2611,N_3293);
nand U5971 (N_5971,N_2266,N_3562);
and U5972 (N_5972,N_2112,N_3303);
xnor U5973 (N_5973,N_3627,N_2041);
nor U5974 (N_5974,N_3415,N_3872);
and U5975 (N_5975,N_2554,N_3363);
nor U5976 (N_5976,N_3764,N_3237);
xor U5977 (N_5977,N_3518,N_3558);
nand U5978 (N_5978,N_2678,N_3968);
nand U5979 (N_5979,N_3815,N_3187);
xor U5980 (N_5980,N_3480,N_2402);
nand U5981 (N_5981,N_3067,N_3572);
xor U5982 (N_5982,N_3365,N_2307);
or U5983 (N_5983,N_3012,N_3656);
or U5984 (N_5984,N_3547,N_2139);
and U5985 (N_5985,N_2226,N_2158);
or U5986 (N_5986,N_2832,N_3549);
nand U5987 (N_5987,N_2425,N_2290);
xor U5988 (N_5988,N_2832,N_2669);
or U5989 (N_5989,N_2507,N_2068);
nor U5990 (N_5990,N_2616,N_2028);
xnor U5991 (N_5991,N_3443,N_2139);
or U5992 (N_5992,N_3686,N_3978);
nand U5993 (N_5993,N_2218,N_2622);
nand U5994 (N_5994,N_2994,N_2460);
nor U5995 (N_5995,N_3474,N_2889);
xor U5996 (N_5996,N_3921,N_3944);
nor U5997 (N_5997,N_2725,N_3032);
nand U5998 (N_5998,N_2651,N_2987);
and U5999 (N_5999,N_2266,N_3871);
and U6000 (N_6000,N_4502,N_4790);
nor U6001 (N_6001,N_4134,N_5426);
nor U6002 (N_6002,N_5369,N_4160);
nand U6003 (N_6003,N_4114,N_4563);
nor U6004 (N_6004,N_4353,N_4212);
or U6005 (N_6005,N_4735,N_4571);
and U6006 (N_6006,N_4412,N_5852);
and U6007 (N_6007,N_4254,N_5061);
or U6008 (N_6008,N_4466,N_5218);
or U6009 (N_6009,N_4984,N_5608);
xnor U6010 (N_6010,N_5554,N_5766);
and U6011 (N_6011,N_4697,N_4183);
xnor U6012 (N_6012,N_5094,N_4847);
nand U6013 (N_6013,N_4054,N_5434);
and U6014 (N_6014,N_5036,N_4390);
nand U6015 (N_6015,N_5082,N_5022);
xor U6016 (N_6016,N_4728,N_4998);
and U6017 (N_6017,N_4995,N_4845);
nor U6018 (N_6018,N_5731,N_5655);
and U6019 (N_6019,N_5124,N_5170);
or U6020 (N_6020,N_4100,N_4976);
or U6021 (N_6021,N_4932,N_5443);
nand U6022 (N_6022,N_5619,N_5786);
nor U6023 (N_6023,N_4622,N_4078);
nand U6024 (N_6024,N_5853,N_5588);
nand U6025 (N_6025,N_4742,N_5138);
and U6026 (N_6026,N_4848,N_4020);
or U6027 (N_6027,N_4526,N_4717);
or U6028 (N_6028,N_4626,N_4323);
and U6029 (N_6029,N_4970,N_5215);
and U6030 (N_6030,N_5859,N_4248);
and U6031 (N_6031,N_5530,N_5103);
and U6032 (N_6032,N_4364,N_4438);
xnor U6033 (N_6033,N_5308,N_5778);
nand U6034 (N_6034,N_4744,N_5359);
or U6035 (N_6035,N_5845,N_4555);
nand U6036 (N_6036,N_4266,N_4301);
nand U6037 (N_6037,N_5381,N_5558);
or U6038 (N_6038,N_5519,N_5352);
or U6039 (N_6039,N_5505,N_5898);
or U6040 (N_6040,N_5687,N_4543);
and U6041 (N_6041,N_5172,N_5970);
nor U6042 (N_6042,N_4376,N_5884);
nor U6043 (N_6043,N_4320,N_5221);
xnor U6044 (N_6044,N_4570,N_4608);
and U6045 (N_6045,N_5544,N_5160);
or U6046 (N_6046,N_4494,N_5962);
and U6047 (N_6047,N_4792,N_5823);
xnor U6048 (N_6048,N_5900,N_4077);
or U6049 (N_6049,N_5803,N_5870);
xor U6050 (N_6050,N_5326,N_4913);
nor U6051 (N_6051,N_4377,N_5329);
or U6052 (N_6052,N_5165,N_5211);
and U6053 (N_6053,N_4396,N_4544);
nor U6054 (N_6054,N_4972,N_4861);
and U6055 (N_6055,N_4647,N_4954);
nor U6056 (N_6056,N_5273,N_5034);
and U6057 (N_6057,N_4684,N_5942);
or U6058 (N_6058,N_5562,N_5837);
and U6059 (N_6059,N_5468,N_4476);
and U6060 (N_6060,N_4680,N_4380);
or U6061 (N_6061,N_4854,N_4302);
nor U6062 (N_6062,N_4127,N_5903);
nor U6063 (N_6063,N_5427,N_4569);
and U6064 (N_6064,N_5716,N_4794);
xnor U6065 (N_6065,N_4188,N_4362);
xor U6066 (N_6066,N_5939,N_4517);
and U6067 (N_6067,N_4057,N_4853);
or U6068 (N_6068,N_5781,N_5760);
xor U6069 (N_6069,N_4395,N_4391);
nor U6070 (N_6070,N_4927,N_5254);
or U6071 (N_6071,N_4619,N_4048);
xnor U6072 (N_6072,N_4843,N_5700);
nor U6073 (N_6073,N_5998,N_5624);
or U6074 (N_6074,N_4340,N_4582);
and U6075 (N_6075,N_5964,N_4941);
or U6076 (N_6076,N_5343,N_5388);
nand U6077 (N_6077,N_5508,N_5446);
nor U6078 (N_6078,N_5983,N_4169);
nand U6079 (N_6079,N_5593,N_5166);
or U6080 (N_6080,N_5088,N_4785);
or U6081 (N_6081,N_4558,N_4331);
nand U6082 (N_6082,N_4102,N_4673);
xor U6083 (N_6083,N_5051,N_5956);
or U6084 (N_6084,N_5444,N_5918);
or U6085 (N_6085,N_4978,N_5754);
xor U6086 (N_6086,N_4479,N_4112);
xnor U6087 (N_6087,N_5228,N_4999);
xor U6088 (N_6088,N_5191,N_4501);
nand U6089 (N_6089,N_5590,N_4117);
nand U6090 (N_6090,N_5285,N_5794);
nand U6091 (N_6091,N_4222,N_4789);
xor U6092 (N_6092,N_4240,N_5889);
and U6093 (N_6093,N_4430,N_4791);
nand U6094 (N_6094,N_5693,N_5431);
and U6095 (N_6095,N_4458,N_4909);
nor U6096 (N_6096,N_4170,N_5628);
nor U6097 (N_6097,N_5332,N_4341);
xnor U6098 (N_6098,N_5576,N_5076);
and U6099 (N_6099,N_5950,N_4454);
or U6100 (N_6100,N_5489,N_4547);
nor U6101 (N_6101,N_4229,N_5216);
xnor U6102 (N_6102,N_5722,N_5994);
xnor U6103 (N_6103,N_5389,N_4284);
or U6104 (N_6104,N_5230,N_5579);
nor U6105 (N_6105,N_5682,N_5187);
or U6106 (N_6106,N_4421,N_5915);
nand U6107 (N_6107,N_5630,N_5605);
xor U6108 (N_6108,N_4311,N_4016);
nor U6109 (N_6109,N_4403,N_5050);
xor U6110 (N_6110,N_5398,N_5313);
nand U6111 (N_6111,N_4085,N_5250);
xnor U6112 (N_6112,N_4486,N_4452);
xor U6113 (N_6113,N_5328,N_4948);
nand U6114 (N_6114,N_5458,N_5163);
nor U6115 (N_6115,N_5146,N_4910);
and U6116 (N_6116,N_4669,N_4326);
or U6117 (N_6117,N_4951,N_5551);
nand U6118 (N_6118,N_5395,N_5346);
nor U6119 (N_6119,N_5137,N_4295);
xnor U6120 (N_6120,N_5143,N_4262);
and U6121 (N_6121,N_5635,N_4782);
nand U6122 (N_6122,N_5568,N_5141);
xor U6123 (N_6123,N_4268,N_4131);
nor U6124 (N_6124,N_4217,N_5932);
xnor U6125 (N_6125,N_4345,N_5473);
xnor U6126 (N_6126,N_5467,N_4404);
nor U6127 (N_6127,N_4679,N_5820);
nor U6128 (N_6128,N_5817,N_4318);
nor U6129 (N_6129,N_5023,N_5487);
nor U6130 (N_6130,N_5106,N_4500);
xor U6131 (N_6131,N_4309,N_5673);
xor U6132 (N_6132,N_5614,N_5459);
nand U6133 (N_6133,N_4576,N_5641);
xnor U6134 (N_6134,N_4330,N_5456);
and U6135 (N_6135,N_4294,N_4914);
or U6136 (N_6136,N_4524,N_4889);
and U6137 (N_6137,N_5861,N_5149);
or U6138 (N_6138,N_4444,N_4825);
or U6139 (N_6139,N_5776,N_4161);
or U6140 (N_6140,N_5771,N_4716);
and U6141 (N_6141,N_5144,N_4880);
nand U6142 (N_6142,N_4327,N_4413);
nand U6143 (N_6143,N_5710,N_4319);
nand U6144 (N_6144,N_4689,N_5816);
nand U6145 (N_6145,N_5765,N_4397);
nand U6146 (N_6146,N_4930,N_4042);
xnor U6147 (N_6147,N_5309,N_4233);
or U6148 (N_6148,N_4139,N_4906);
nand U6149 (N_6149,N_4965,N_5122);
nor U6150 (N_6150,N_5205,N_4540);
and U6151 (N_6151,N_4786,N_4975);
or U6152 (N_6152,N_4893,N_5252);
and U6153 (N_6153,N_5013,N_5663);
and U6154 (N_6154,N_4993,N_5793);
or U6155 (N_6155,N_5890,N_4314);
nor U6156 (N_6156,N_4801,N_4382);
xor U6157 (N_6157,N_5872,N_5694);
nand U6158 (N_6158,N_4687,N_5319);
xnor U6159 (N_6159,N_4067,N_5356);
nand U6160 (N_6160,N_5524,N_4819);
and U6161 (N_6161,N_4712,N_5780);
xnor U6162 (N_6162,N_4267,N_4565);
nor U6163 (N_6163,N_5463,N_4264);
and U6164 (N_6164,N_4151,N_4671);
xor U6165 (N_6165,N_4892,N_4710);
and U6166 (N_6166,N_4656,N_5967);
or U6167 (N_6167,N_5186,N_4305);
nor U6168 (N_6168,N_5249,N_5464);
and U6169 (N_6169,N_4211,N_4823);
nor U6170 (N_6170,N_5741,N_5941);
nand U6171 (N_6171,N_5110,N_4886);
nor U6172 (N_6172,N_5053,N_4554);
and U6173 (N_6173,N_4840,N_4245);
and U6174 (N_6174,N_4778,N_5449);
nor U6175 (N_6175,N_4659,N_5606);
or U6176 (N_6176,N_4291,N_5599);
nand U6177 (N_6177,N_5212,N_4002);
nand U6178 (N_6178,N_5441,N_5038);
xnor U6179 (N_6179,N_5404,N_5183);
xor U6180 (N_6180,N_5934,N_4488);
nor U6181 (N_6181,N_4401,N_4009);
nor U6182 (N_6182,N_4113,N_4159);
xnor U6183 (N_6183,N_4763,N_4257);
nor U6184 (N_6184,N_4428,N_4864);
and U6185 (N_6185,N_5098,N_5235);
nand U6186 (N_6186,N_4798,N_5337);
xnor U6187 (N_6187,N_4770,N_5016);
and U6188 (N_6188,N_4172,N_4130);
or U6189 (N_6189,N_4224,N_5792);
and U6190 (N_6190,N_4231,N_4899);
nor U6191 (N_6191,N_4882,N_5798);
or U6192 (N_6192,N_4468,N_5429);
xnor U6193 (N_6193,N_4624,N_5583);
xnor U6194 (N_6194,N_5288,N_5685);
nor U6195 (N_6195,N_5929,N_4695);
or U6196 (N_6196,N_4491,N_5435);
and U6197 (N_6197,N_4507,N_5946);
nand U6198 (N_6198,N_4214,N_5018);
nor U6199 (N_6199,N_5035,N_4908);
xor U6200 (N_6200,N_5638,N_4181);
and U6201 (N_6201,N_4709,N_4734);
and U6202 (N_6202,N_5156,N_4064);
and U6203 (N_6203,N_5512,N_5711);
xnor U6204 (N_6204,N_4981,N_4835);
nand U6205 (N_6205,N_5533,N_5277);
or U6206 (N_6206,N_4106,N_5737);
nor U6207 (N_6207,N_4903,N_5738);
nand U6208 (N_6208,N_5148,N_5931);
nor U6209 (N_6209,N_5827,N_4123);
and U6210 (N_6210,N_4164,N_5531);
and U6211 (N_6211,N_5145,N_5071);
nor U6212 (N_6212,N_4585,N_5151);
or U6213 (N_6213,N_4748,N_5897);
xnor U6214 (N_6214,N_5123,N_5797);
and U6215 (N_6215,N_5225,N_5510);
nand U6216 (N_6216,N_5140,N_4133);
and U6217 (N_6217,N_5095,N_5571);
or U6218 (N_6218,N_5750,N_5080);
nand U6219 (N_6219,N_5430,N_4347);
and U6220 (N_6220,N_5822,N_5069);
xnor U6221 (N_6221,N_5992,N_5589);
xor U6222 (N_6222,N_4101,N_4061);
and U6223 (N_6223,N_4460,N_4472);
xnor U6224 (N_6224,N_5350,N_4858);
or U6225 (N_6225,N_4645,N_5303);
nor U6226 (N_6226,N_4079,N_5732);
nand U6227 (N_6227,N_5011,N_5008);
or U6228 (N_6228,N_4887,N_5073);
nand U6229 (N_6229,N_5142,N_4283);
and U6230 (N_6230,N_4944,N_5159);
nor U6231 (N_6231,N_5925,N_4149);
nor U6232 (N_6232,N_4884,N_4752);
nor U6233 (N_6233,N_5860,N_4487);
nand U6234 (N_6234,N_5960,N_5854);
xnor U6235 (N_6235,N_4832,N_5670);
or U6236 (N_6236,N_5930,N_5234);
or U6237 (N_6237,N_5947,N_5938);
nor U6238 (N_6238,N_5301,N_4361);
and U6239 (N_6239,N_5111,N_5002);
and U6240 (N_6240,N_4611,N_5971);
or U6241 (N_6241,N_5155,N_4150);
nand U6242 (N_6242,N_5747,N_5789);
or U6243 (N_6243,N_4029,N_4722);
xnor U6244 (N_6244,N_4325,N_5119);
and U6245 (N_6245,N_5500,N_5916);
nand U6246 (N_6246,N_4553,N_5196);
or U6247 (N_6247,N_4003,N_4793);
nor U6248 (N_6248,N_4046,N_4186);
nor U6249 (N_6249,N_5813,N_4334);
and U6250 (N_6250,N_5661,N_5244);
xnor U6251 (N_6251,N_4031,N_5958);
and U6252 (N_6252,N_5263,N_5657);
nor U6253 (N_6253,N_5271,N_4510);
nor U6254 (N_6254,N_5819,N_4044);
or U6255 (N_6255,N_5746,N_5604);
and U6256 (N_6256,N_4751,N_4152);
xnor U6257 (N_6257,N_4306,N_4333);
or U6258 (N_6258,N_4166,N_5841);
xor U6259 (N_6259,N_5180,N_5314);
or U6260 (N_6260,N_5704,N_4766);
nand U6261 (N_6261,N_4588,N_5953);
and U6262 (N_6262,N_5865,N_4282);
and U6263 (N_6263,N_4414,N_5391);
or U6264 (N_6264,N_5949,N_5979);
or U6265 (N_6265,N_5969,N_5012);
nor U6266 (N_6266,N_5880,N_5296);
or U6267 (N_6267,N_5136,N_5534);
xnor U6268 (N_6268,N_4090,N_5806);
nand U6269 (N_6269,N_4157,N_4411);
xor U6270 (N_6270,N_5004,N_4234);
or U6271 (N_6271,N_5203,N_5447);
or U6272 (N_6272,N_5691,N_4530);
xor U6273 (N_6273,N_5718,N_5563);
and U6274 (N_6274,N_5227,N_5543);
and U6275 (N_6275,N_5681,N_4804);
xnor U6276 (N_6276,N_4097,N_4288);
and U6277 (N_6277,N_4053,N_4531);
nor U6278 (N_6278,N_5349,N_4655);
nand U6279 (N_6279,N_5466,N_5056);
xor U6280 (N_6280,N_5269,N_4691);
or U6281 (N_6281,N_4607,N_5762);
and U6282 (N_6282,N_5214,N_4860);
nand U6283 (N_6283,N_4200,N_4045);
and U6284 (N_6284,N_4099,N_5802);
and U6285 (N_6285,N_4521,N_5089);
nor U6286 (N_6286,N_5178,N_5096);
nand U6287 (N_6287,N_5192,N_4818);
or U6288 (N_6288,N_4508,N_4600);
nand U6289 (N_6289,N_5304,N_4776);
nor U6290 (N_6290,N_5413,N_4399);
nand U6291 (N_6291,N_5729,N_5863);
xor U6292 (N_6292,N_5424,N_5715);
xor U6293 (N_6293,N_4897,N_5363);
and U6294 (N_6294,N_4220,N_5127);
nand U6295 (N_6295,N_4637,N_5795);
xor U6296 (N_6296,N_5198,N_5945);
nand U6297 (N_6297,N_5659,N_5584);
and U6298 (N_6298,N_4762,N_5724);
nand U6299 (N_6299,N_4095,N_5092);
or U6300 (N_6300,N_4273,N_4179);
or U6301 (N_6301,N_4246,N_5321);
xnor U6302 (N_6302,N_4992,N_5952);
xnor U6303 (N_6303,N_5617,N_5209);
and U6304 (N_6304,N_4070,N_5514);
nor U6305 (N_6305,N_4829,N_4872);
xnor U6306 (N_6306,N_4155,N_5570);
xnor U6307 (N_6307,N_4303,N_4643);
and U6308 (N_6308,N_5298,N_5284);
or U6309 (N_6309,N_4378,N_4049);
or U6310 (N_6310,N_5636,N_4514);
nand U6311 (N_6311,N_4012,N_5882);
xor U6312 (N_6312,N_5922,N_4136);
xnor U6313 (N_6313,N_4055,N_4809);
nor U6314 (N_6314,N_4846,N_5849);
nand U6315 (N_6315,N_4481,N_4419);
nor U6316 (N_6316,N_4145,N_5936);
or U6317 (N_6317,N_4219,N_5014);
nor U6318 (N_6318,N_4560,N_5387);
nor U6319 (N_6319,N_5448,N_4589);
nor U6320 (N_6320,N_5428,N_4107);
nand U6321 (N_6321,N_5913,N_4703);
nand U6322 (N_6322,N_4496,N_4740);
nor U6323 (N_6323,N_5883,N_5370);
nor U6324 (N_6324,N_5257,N_5276);
or U6325 (N_6325,N_5567,N_5300);
nor U6326 (N_6326,N_4158,N_5208);
xnor U6327 (N_6327,N_4928,N_5695);
and U6328 (N_6328,N_5461,N_4803);
xnor U6329 (N_6329,N_5409,N_4387);
nand U6330 (N_6330,N_4852,N_4259);
nand U6331 (N_6331,N_4286,N_4416);
nand U6332 (N_6332,N_4435,N_5068);
xnor U6333 (N_6333,N_5414,N_4062);
and U6334 (N_6334,N_4453,N_5855);
and U6335 (N_6335,N_5161,N_4727);
nand U6336 (N_6336,N_5674,N_5364);
xor U6337 (N_6337,N_4739,N_5442);
and U6338 (N_6338,N_5272,N_4478);
xor U6339 (N_6339,N_5380,N_5907);
xor U6340 (N_6340,N_5000,N_5646);
and U6341 (N_6341,N_5041,N_5643);
nand U6342 (N_6342,N_4642,N_4651);
nor U6343 (N_6343,N_4346,N_5399);
xor U6344 (N_6344,N_4868,N_4105);
nor U6345 (N_6345,N_5618,N_4147);
nor U6346 (N_6346,N_4584,N_5767);
nand U6347 (N_6347,N_5537,N_5648);
or U6348 (N_6348,N_5675,N_4779);
or U6349 (N_6349,N_5220,N_4745);
and U6350 (N_6350,N_5996,N_4807);
or U6351 (N_6351,N_4678,N_5226);
xor U6352 (N_6352,N_5382,N_5749);
xnor U6353 (N_6353,N_5997,N_4081);
xnor U6354 (N_6354,N_5895,N_5239);
xor U6355 (N_6355,N_5465,N_5805);
nor U6356 (N_6356,N_5282,N_4681);
xnor U6357 (N_6357,N_4672,N_5680);
nor U6358 (N_6358,N_5185,N_5164);
nand U6359 (N_6359,N_4389,N_5631);
nor U6360 (N_6360,N_4512,N_5017);
or U6361 (N_6361,N_5190,N_4074);
xor U6362 (N_6362,N_5469,N_5727);
nand U6363 (N_6363,N_4879,N_4797);
and U6364 (N_6364,N_5482,N_4445);
nand U6365 (N_6365,N_5720,N_5154);
nor U6366 (N_6366,N_5879,N_5102);
xor U6367 (N_6367,N_5105,N_4010);
nand U6368 (N_6368,N_5042,N_4765);
nor U6369 (N_6369,N_4606,N_5553);
nor U6370 (N_6370,N_5494,N_5264);
nor U6371 (N_6371,N_5743,N_5305);
nand U6372 (N_6372,N_5392,N_4663);
nor U6373 (N_6373,N_4644,N_5848);
xor U6374 (N_6374,N_5977,N_5561);
or U6375 (N_6375,N_4237,N_5402);
nor U6376 (N_6376,N_4122,N_5133);
nand U6377 (N_6377,N_5756,N_4426);
or U6378 (N_6378,N_4603,N_5620);
xor U6379 (N_6379,N_4076,N_4800);
and U6380 (N_6380,N_4109,N_4406);
nor U6381 (N_6381,N_5677,N_5361);
nor U6382 (N_6382,N_5785,N_5603);
nand U6383 (N_6383,N_5063,N_4961);
xnor U6384 (N_6384,N_4506,N_4256);
and U6385 (N_6385,N_5341,N_4218);
nand U6386 (N_6386,N_4281,N_5782);
and U6387 (N_6387,N_5705,N_5703);
and U6388 (N_6388,N_5333,N_4519);
nor U6389 (N_6389,N_4648,N_5416);
and U6390 (N_6390,N_5697,N_4698);
nor U6391 (N_6391,N_5664,N_4427);
nand U6392 (N_6392,N_5957,N_4736);
xor U6393 (N_6393,N_4418,N_5299);
or U6394 (N_6394,N_4292,N_4128);
nand U6395 (N_6395,N_4400,N_5838);
xnor U6396 (N_6396,N_5773,N_5520);
or U6397 (N_6397,N_4636,N_5892);
xor U6398 (N_6398,N_5091,N_5005);
nand U6399 (N_6399,N_4541,N_5748);
nor U6400 (N_6400,N_4911,N_5373);
and U6401 (N_6401,N_4652,N_5078);
or U6402 (N_6402,N_5176,N_5219);
nand U6403 (N_6403,N_4821,N_4310);
nor U6404 (N_6404,N_5809,N_5826);
nand U6405 (N_6405,N_5824,N_4888);
and U6406 (N_6406,N_5107,N_4940);
or U6407 (N_6407,N_5052,N_4360);
nor U6408 (N_6408,N_5856,N_4338);
xor U6409 (N_6409,N_5592,N_4733);
xnor U6410 (N_6410,N_5498,N_4083);
and U6411 (N_6411,N_5323,N_5810);
nand U6412 (N_6412,N_5310,N_5851);
or U6413 (N_6413,N_5600,N_4705);
or U6414 (N_6414,N_5734,N_5517);
or U6415 (N_6415,N_4328,N_5258);
and U6416 (N_6416,N_4827,N_5601);
and U6417 (N_6417,N_4943,N_4828);
or U6418 (N_6418,N_5118,N_4119);
or U6419 (N_6419,N_5397,N_4878);
or U6420 (N_6420,N_4269,N_5815);
nand U6421 (N_6421,N_4690,N_5204);
nor U6422 (N_6422,N_4896,N_5480);
nand U6423 (N_6423,N_4881,N_4238);
nor U6424 (N_6424,N_4820,N_5832);
nand U6425 (N_6425,N_5656,N_5259);
nand U6426 (N_6426,N_5479,N_5575);
nand U6427 (N_6427,N_4545,N_5550);
nor U6428 (N_6428,N_4047,N_5294);
or U6429 (N_6429,N_5497,N_4750);
xnor U6430 (N_6430,N_5976,N_5385);
xnor U6431 (N_6431,N_5758,N_4959);
xnor U6432 (N_6432,N_4796,N_5322);
xor U6433 (N_6433,N_5831,N_5800);
nand U6434 (N_6434,N_5905,N_5116);
and U6435 (N_6435,N_4165,N_4720);
nand U6436 (N_6436,N_4590,N_5169);
and U6437 (N_6437,N_4277,N_5602);
or U6438 (N_6438,N_4202,N_4601);
nand U6439 (N_6439,N_5084,N_4731);
xor U6440 (N_6440,N_5496,N_5290);
or U6441 (N_6441,N_4808,N_5060);
and U6442 (N_6442,N_5281,N_4191);
nand U6443 (N_6443,N_4205,N_5981);
and U6444 (N_6444,N_5569,N_4358);
xor U6445 (N_6445,N_4904,N_5491);
or U6446 (N_6446,N_4308,N_5596);
xor U6447 (N_6447,N_4317,N_5024);
nor U6448 (N_6448,N_5317,N_4261);
xnor U6449 (N_6449,N_4103,N_5899);
or U6450 (N_6450,N_5814,N_5150);
and U6451 (N_6451,N_5026,N_5162);
xor U6452 (N_6452,N_4810,N_5763);
or U6453 (N_6453,N_5481,N_4026);
and U6454 (N_6454,N_5706,N_5108);
nand U6455 (N_6455,N_4824,N_5696);
and U6456 (N_6456,N_4520,N_4140);
and U6457 (N_6457,N_4321,N_5223);
xnor U6458 (N_6458,N_4104,N_4208);
xor U6459 (N_6459,N_5445,N_4356);
xor U6460 (N_6460,N_5966,N_4990);
xor U6461 (N_6461,N_5523,N_5739);
nor U6462 (N_6462,N_5477,N_4271);
xor U6463 (N_6463,N_4926,N_4339);
or U6464 (N_6464,N_5289,N_5113);
or U6465 (N_6465,N_5097,N_4863);
or U6466 (N_6466,N_4293,N_5504);
nand U6467 (N_6467,N_5779,N_4539);
xor U6468 (N_6468,N_5460,N_5280);
nand U6469 (N_6469,N_4329,N_5059);
nand U6470 (N_6470,N_4116,N_4875);
or U6471 (N_6471,N_5559,N_5632);
or U6472 (N_6472,N_5541,N_4957);
nand U6473 (N_6473,N_4125,N_4883);
xor U6474 (N_6474,N_5846,N_5440);
and U6475 (N_6475,N_4394,N_5316);
nor U6476 (N_6476,N_4477,N_5989);
nand U6477 (N_6477,N_4210,N_4255);
nand U6478 (N_6478,N_5256,N_4143);
nand U6479 (N_6479,N_5422,N_4425);
or U6480 (N_6480,N_4213,N_4244);
or U6481 (N_6481,N_5407,N_4753);
nor U6482 (N_6482,N_5513,N_4686);
and U6483 (N_6483,N_5896,N_4110);
xor U6484 (N_6484,N_4955,N_5044);
or U6485 (N_6485,N_4019,N_4971);
and U6486 (N_6486,N_5654,N_5240);
xnor U6487 (N_6487,N_4620,N_5406);
and U6488 (N_6488,N_4721,N_4027);
xnor U6489 (N_6489,N_4298,N_5525);
and U6490 (N_6490,N_5425,N_4304);
and U6491 (N_6491,N_5003,N_4204);
nand U6492 (N_6492,N_5833,N_5283);
nand U6493 (N_6493,N_4967,N_4788);
nor U6494 (N_6494,N_5134,N_4838);
nor U6495 (N_6495,N_5557,N_4694);
and U6496 (N_6496,N_5279,N_4028);
xor U6497 (N_6497,N_5708,N_5761);
nand U6498 (N_6498,N_5331,N_5790);
and U6499 (N_6499,N_4646,N_4597);
nor U6500 (N_6500,N_4035,N_4933);
or U6501 (N_6501,N_5135,N_4441);
and U6502 (N_6502,N_4473,N_4718);
xnor U6503 (N_6503,N_4977,N_5031);
nor U6504 (N_6504,N_5484,N_5902);
and U6505 (N_6505,N_4537,N_4443);
or U6506 (N_6506,N_5421,N_5408);
nor U6507 (N_6507,N_4371,N_5678);
nand U6508 (N_6508,N_4811,N_4552);
nor U6509 (N_6509,N_4579,N_4918);
nand U6510 (N_6510,N_5188,N_5307);
nor U6511 (N_6511,N_5158,N_5207);
and U6512 (N_6512,N_4274,N_4760);
nand U6513 (N_6513,N_4433,N_5470);
or U6514 (N_6514,N_5759,N_5045);
xnor U6515 (N_6515,N_5037,N_5951);
or U6516 (N_6516,N_4300,N_4724);
nand U6517 (N_6517,N_5079,N_5501);
xnor U6518 (N_6518,N_5125,N_5194);
or U6519 (N_6519,N_4594,N_4316);
or U6520 (N_6520,N_4704,N_5652);
nor U6521 (N_6521,N_5075,N_4994);
and U6522 (N_6522,N_5522,N_4439);
nand U6523 (N_6523,N_5535,N_5062);
or U6524 (N_6524,N_4442,N_5086);
nor U6525 (N_6525,N_4640,N_4124);
xnor U6526 (N_6526,N_4523,N_4974);
xor U6527 (N_6527,N_5432,N_5247);
xnor U6528 (N_6528,N_5577,N_5261);
nand U6529 (N_6529,N_4532,N_5622);
and U6530 (N_6530,N_5412,N_4163);
and U6531 (N_6531,N_4024,N_5348);
nand U6532 (N_6532,N_5390,N_4758);
nor U6533 (N_6533,N_5634,N_5384);
nand U6534 (N_6534,N_4153,N_4577);
nor U6535 (N_6535,N_5327,N_5336);
nor U6536 (N_6536,N_5410,N_4688);
nor U6537 (N_6537,N_5893,N_5286);
or U6538 (N_6538,N_5083,N_4243);
nand U6539 (N_6539,N_5842,N_4372);
xnor U6540 (N_6540,N_5365,N_5229);
or U6541 (N_6541,N_5450,N_4805);
xnor U6542 (N_6542,N_4253,N_5115);
nand U6543 (N_6543,N_4175,N_5923);
nor U6544 (N_6544,N_5112,N_5796);
or U6545 (N_6545,N_4297,N_4021);
and U6546 (N_6546,N_5030,N_5457);
nor U6547 (N_6547,N_5649,N_4859);
and U6548 (N_6548,N_4670,N_4870);
or U6549 (N_6549,N_4568,N_4743);
xnor U6550 (N_6550,N_4968,N_4461);
or U6551 (N_6551,N_5735,N_4167);
xor U6552 (N_6552,N_4815,N_4056);
and U6553 (N_6553,N_4635,N_4215);
nor U6554 (N_6554,N_5334,N_4041);
xor U6555 (N_6555,N_4176,N_4767);
and U6556 (N_6556,N_5818,N_5043);
or U6557 (N_6557,N_5131,N_4900);
nand U6558 (N_6558,N_4509,N_5572);
or U6559 (N_6559,N_4187,N_4385);
or U6560 (N_6560,N_4831,N_5713);
and U6561 (N_6561,N_5199,N_5338);
xor U6562 (N_6562,N_4676,N_5368);
nor U6563 (N_6563,N_5270,N_4907);
xor U6564 (N_6564,N_4296,N_5736);
nor U6565 (N_6565,N_4137,N_4459);
or U6566 (N_6566,N_4275,N_5650);
nor U6567 (N_6567,N_5521,N_5645);
and U6568 (N_6568,N_5857,N_5875);
xor U6569 (N_6569,N_5275,N_4596);
nor U6570 (N_6570,N_5132,N_4368);
xnor U6571 (N_6571,N_5728,N_4280);
nand U6572 (N_6572,N_5753,N_4355);
or U6573 (N_6573,N_4307,N_4917);
nand U6574 (N_6574,N_5087,N_4230);
or U6575 (N_6575,N_4276,N_5744);
nand U6576 (N_6576,N_4232,N_5536);
or U6577 (N_6577,N_4956,N_4402);
nor U6578 (N_6578,N_4641,N_5742);
xnor U6579 (N_6579,N_5943,N_5676);
xor U6580 (N_6580,N_5597,N_5835);
or U6581 (N_6581,N_4515,N_5615);
xnor U6582 (N_6582,N_4953,N_4732);
xnor U6583 (N_6583,N_5217,N_4484);
or U6584 (N_6584,N_5948,N_5339);
nor U6585 (N_6585,N_5940,N_4657);
and U6586 (N_6586,N_5978,N_4573);
xnor U6587 (N_6587,N_4032,N_4901);
nand U6588 (N_6588,N_4982,N_5699);
and U6589 (N_6589,N_5242,N_4923);
nor U6590 (N_6590,N_5120,N_4729);
nand U6591 (N_6591,N_4795,N_5419);
xor U6592 (N_6592,N_4759,N_4920);
or U6593 (N_6593,N_4609,N_4625);
or U6594 (N_6594,N_4142,N_4036);
and U6595 (N_6595,N_4772,N_4602);
or U6596 (N_6596,N_4455,N_4450);
and U6597 (N_6597,N_4658,N_4258);
xor U6598 (N_6598,N_5702,N_5182);
xnor U6599 (N_6599,N_4348,N_4916);
xor U6600 (N_6600,N_5552,N_4154);
nand U6601 (N_6601,N_5901,N_4518);
or U6602 (N_6602,N_5104,N_5688);
or U6603 (N_6603,N_4495,N_5921);
or U6604 (N_6604,N_4367,N_5325);
or U6605 (N_6605,N_5908,N_4986);
or U6606 (N_6606,N_4337,N_4365);
or U6607 (N_6607,N_4583,N_4764);
or U6608 (N_6608,N_5485,N_5121);
and U6609 (N_6609,N_5376,N_5213);
xnor U6610 (N_6610,N_4925,N_4236);
or U6611 (N_6611,N_5292,N_5057);
nand U6612 (N_6612,N_5020,N_4533);
nand U6613 (N_6613,N_4592,N_5394);
nand U6614 (N_6614,N_4008,N_5752);
nor U6615 (N_6615,N_4171,N_5709);
and U6616 (N_6616,N_5206,N_4905);
or U6617 (N_6617,N_5453,N_5358);
nor U6618 (N_6618,N_4873,N_4575);
xor U6619 (N_6619,N_4538,N_5028);
nor U6620 (N_6620,N_5251,N_4015);
nand U6621 (N_6621,N_5914,N_5667);
nor U6622 (N_6622,N_4120,N_5126);
xnor U6623 (N_6623,N_4420,N_5607);
nand U6624 (N_6624,N_5495,N_4783);
or U6625 (N_6625,N_4177,N_5184);
nor U6626 (N_6626,N_5302,N_4633);
nor U6627 (N_6627,N_4664,N_4885);
and U6628 (N_6628,N_4837,N_5926);
nor U6629 (N_6629,N_5917,N_4492);
nand U6630 (N_6630,N_4223,N_4771);
or U6631 (N_6631,N_4185,N_4949);
nand U6632 (N_6632,N_5974,N_4610);
nand U6633 (N_6633,N_5511,N_5690);
xnor U6634 (N_6634,N_5344,N_4639);
and U6635 (N_6635,N_5117,N_5887);
nand U6636 (N_6636,N_5725,N_5015);
nor U6637 (N_6637,N_4535,N_5375);
nor U6638 (N_6638,N_5529,N_5633);
and U6639 (N_6639,N_4946,N_4912);
and U6640 (N_6640,N_4525,N_4073);
or U6641 (N_6641,N_5651,N_5128);
or U6642 (N_6642,N_4960,N_5243);
nor U6643 (N_6643,N_4018,N_4239);
and U6644 (N_6644,N_5721,N_5010);
xnor U6645 (N_6645,N_5455,N_5764);
and U6646 (N_6646,N_4816,N_5237);
nor U6647 (N_6647,N_5787,N_5555);
nor U6648 (N_6648,N_5109,N_4263);
xnor U6649 (N_6649,N_5799,N_5345);
and U6650 (N_6650,N_5714,N_5973);
and U6651 (N_6651,N_4384,N_4964);
nand U6652 (N_6652,N_5807,N_5492);
and U6653 (N_6653,N_5420,N_4668);
nand U6654 (N_6654,N_5866,N_4058);
nor U6655 (N_6655,N_5871,N_5791);
nand U6656 (N_6656,N_5598,N_4937);
nand U6657 (N_6657,N_4516,N_5662);
or U6658 (N_6658,N_5665,N_5019);
nand U6659 (N_6659,N_4251,N_5245);
nand U6660 (N_6660,N_5545,N_4942);
and U6661 (N_6661,N_5171,N_5984);
and U6662 (N_6662,N_4621,N_4814);
nor U6663 (N_6663,N_5486,N_4604);
nor U6664 (N_6664,N_4522,N_4871);
xor U6665 (N_6665,N_4405,N_4919);
xor U6666 (N_6666,N_4551,N_4108);
and U6667 (N_6667,N_4534,N_4952);
and U6668 (N_6668,N_5878,N_4072);
and U6669 (N_6669,N_5374,N_4561);
xnor U6670 (N_6670,N_4634,N_5168);
xnor U6671 (N_6671,N_4674,N_5658);
or U6672 (N_6672,N_4931,N_4802);
nor U6673 (N_6673,N_5471,N_5623);
nor U6674 (N_6674,N_4004,N_4702);
nand U6675 (N_6675,N_5454,N_4040);
or U6676 (N_6676,N_4432,N_4312);
or U6677 (N_6677,N_5238,N_4826);
nor U6678 (N_6678,N_5587,N_4599);
nand U6679 (N_6679,N_5222,N_4060);
or U6680 (N_6680,N_4661,N_4249);
and U6681 (N_6681,N_4063,N_5712);
nand U6682 (N_6682,N_5642,N_5367);
nand U6683 (N_6683,N_4991,N_4207);
xnor U6684 (N_6684,N_4963,N_4746);
nand U6685 (N_6685,N_5153,N_5189);
or U6686 (N_6686,N_5644,N_4247);
nor U6687 (N_6687,N_5927,N_5995);
nand U6688 (N_6688,N_4683,N_5287);
nand U6689 (N_6689,N_5175,N_5812);
nor U6690 (N_6690,N_4780,N_4784);
xor U6691 (N_6691,N_4366,N_4902);
xor U6692 (N_6692,N_5772,N_4874);
and U6693 (N_6693,N_4556,N_4051);
xnor U6694 (N_6694,N_4000,N_4629);
or U6695 (N_6695,N_5181,N_4336);
xor U6696 (N_6696,N_5064,N_4546);
nand U6697 (N_6697,N_5232,N_5507);
xnor U6698 (N_6698,N_5542,N_4692);
nor U6699 (N_6699,N_5478,N_4138);
and U6700 (N_6700,N_4527,N_5847);
nor U6701 (N_6701,N_4528,N_4408);
nor U6702 (N_6702,N_5403,N_5527);
nand U6703 (N_6703,N_4605,N_4065);
and U6704 (N_6704,N_4052,N_4437);
or U6705 (N_6705,N_4851,N_5210);
nand U6706 (N_6706,N_5560,N_5912);
nand U6707 (N_6707,N_5894,N_5937);
and U6708 (N_6708,N_4011,N_4335);
nor U6709 (N_6709,N_4457,N_5268);
or U6710 (N_6710,N_5101,N_4034);
and U6711 (N_6711,N_4936,N_4638);
nor U6712 (N_6712,N_5532,N_5629);
nor U6713 (N_6713,N_5248,N_4322);
nand U6714 (N_6714,N_4386,N_4714);
and U6715 (N_6715,N_5985,N_4369);
or U6716 (N_6716,N_5566,N_4869);
nor U6717 (N_6717,N_4086,N_5072);
nand U6718 (N_6718,N_4446,N_4270);
nor U6719 (N_6719,N_5436,N_4983);
xnor U6720 (N_6720,N_4069,N_5692);
nand U6721 (N_6721,N_5548,N_4162);
or U6722 (N_6722,N_5415,N_5029);
or U6723 (N_6723,N_5689,N_4618);
nand U6724 (N_6724,N_5609,N_5476);
and U6725 (N_6725,N_4505,N_4662);
xnor U6726 (N_6726,N_4374,N_5701);
nand U6727 (N_6727,N_4969,N_4980);
and U6728 (N_6728,N_4915,N_4014);
xor U6729 (N_6729,N_4498,N_4195);
xor U6730 (N_6730,N_5362,N_4451);
or U6731 (N_6731,N_4193,N_5393);
and U6732 (N_6732,N_5293,N_4562);
and U6733 (N_6733,N_5881,N_4354);
or U6734 (N_6734,N_4192,N_5528);
nand U6735 (N_6735,N_4504,N_4039);
nor U6736 (N_6736,N_5811,N_5935);
nand U6737 (N_6737,N_5372,N_5065);
or U6738 (N_6738,N_4370,N_5626);
xor U6739 (N_6739,N_4180,N_4856);
nand U6740 (N_6740,N_5357,N_4289);
nand U6741 (N_6741,N_4707,N_4375);
or U6742 (N_6742,N_5850,N_5265);
xor U6743 (N_6743,N_4615,N_4482);
nand U6744 (N_6744,N_5821,N_4649);
or U6745 (N_6745,N_4895,N_4862);
nand U6746 (N_6746,N_4037,N_5048);
nor U6747 (N_6747,N_4489,N_5564);
and U6748 (N_6748,N_5438,N_4146);
or U6749 (N_6749,N_5986,N_4726);
or U6750 (N_6750,N_4945,N_4757);
nand U6751 (N_6751,N_4866,N_4092);
or U6752 (N_6752,N_5745,N_5174);
nor U6753 (N_6753,N_5862,N_4549);
and U6754 (N_6754,N_4754,N_4388);
nor U6755 (N_6755,N_4806,N_4747);
nor U6756 (N_6756,N_4315,N_4352);
or U6757 (N_6757,N_4761,N_5769);
xor U6758 (N_6758,N_4350,N_5200);
and U6759 (N_6759,N_4587,N_5193);
xor U6760 (N_6760,N_5843,N_4774);
nor U6761 (N_6761,N_5093,N_4775);
nor U6762 (N_6762,N_5173,N_5556);
nor U6763 (N_6763,N_4417,N_5757);
nor U6764 (N_6764,N_5707,N_4693);
nor U6765 (N_6765,N_4429,N_5506);
nand U6766 (N_6766,N_4632,N_4227);
nand U6767 (N_6767,N_5581,N_5231);
xnor U6768 (N_6768,N_4799,N_4436);
or U6769 (N_6769,N_5864,N_4513);
nor U6770 (N_6770,N_4080,N_5867);
and U6771 (N_6771,N_5582,N_4890);
nor U6772 (N_6772,N_4196,N_4001);
or U6773 (N_6773,N_4935,N_5233);
or U6774 (N_6774,N_5474,N_4542);
or U6775 (N_6775,N_4398,N_5462);
xnor U6776 (N_6776,N_5129,N_4675);
xnor U6777 (N_6777,N_4115,N_4557);
nor U6778 (N_6778,N_5518,N_4030);
or U6779 (N_6779,N_5928,N_4756);
or U6780 (N_6780,N_5335,N_4059);
and U6781 (N_6781,N_5669,N_4836);
nand U6782 (N_6782,N_5640,N_4973);
nor U6783 (N_6783,N_5411,N_4250);
nor U6784 (N_6784,N_4817,N_4088);
xnor U6785 (N_6785,N_4068,N_4265);
xor U6786 (N_6786,N_5904,N_4593);
nor U6787 (N_6787,N_4129,N_4839);
xor U6788 (N_6788,N_5924,N_4464);
nand U6789 (N_6789,N_5074,N_5058);
nand U6790 (N_6790,N_5910,N_5100);
xnor U6791 (N_6791,N_5295,N_5090);
and U6792 (N_6792,N_5980,N_5236);
xnor U6793 (N_6793,N_4025,N_4448);
xnor U6794 (N_6794,N_4650,N_5291);
or U6795 (N_6795,N_5627,N_4174);
nand U6796 (N_6796,N_5266,N_4084);
and U6797 (N_6797,N_5401,N_4548);
nor U6798 (N_6798,N_4410,N_5330);
nand U6799 (N_6799,N_5297,N_5580);
nand U6800 (N_6800,N_4121,N_4228);
nand U6801 (N_6801,N_4595,N_5647);
or U6802 (N_6802,N_5538,N_4700);
or U6803 (N_6803,N_5671,N_5726);
nand U6804 (N_6804,N_4381,N_4066);
and U6805 (N_6805,N_5099,N_5920);
or U6806 (N_6806,N_5972,N_4290);
xor U6807 (N_6807,N_4682,N_4203);
nand U6808 (N_6808,N_5312,N_5911);
xnor U6809 (N_6809,N_5698,N_5770);
and U6810 (N_6810,N_5377,N_4921);
nor U6811 (N_6811,N_4867,N_4344);
or U6812 (N_6812,N_4924,N_5130);
nor U6813 (N_6813,N_5255,N_5625);
and U6814 (N_6814,N_4781,N_4156);
nand U6815 (N_6815,N_5547,N_5526);
nor U6816 (N_6816,N_4434,N_4841);
nand U6817 (N_6817,N_5047,N_4225);
xnor U6818 (N_6818,N_4456,N_5515);
xor U6819 (N_6819,N_5613,N_4424);
nand U6820 (N_6820,N_5906,N_5888);
or U6821 (N_6821,N_4715,N_5828);
nor U6822 (N_6822,N_4469,N_5653);
xnor U6823 (N_6823,N_5502,N_5488);
nand U6824 (N_6824,N_4812,N_4988);
xor U6825 (N_6825,N_4987,N_5610);
and U6826 (N_6826,N_5774,N_5565);
nor U6827 (N_6827,N_4332,N_4007);
nor U6828 (N_6828,N_5717,N_4979);
nand U6829 (N_6829,N_4235,N_5383);
nor U6830 (N_6830,N_4934,N_5877);
nor U6831 (N_6831,N_5311,N_4833);
and U6832 (N_6832,N_5686,N_4876);
and U6833 (N_6833,N_5267,N_5039);
nand U6834 (N_6834,N_4929,N_4730);
and U6835 (N_6835,N_5021,N_4877);
nand U6836 (N_6836,N_4194,N_4939);
or U6837 (N_6837,N_4503,N_5433);
nand U6838 (N_6838,N_5539,N_5891);
xnor U6839 (N_6839,N_5733,N_5452);
or U6840 (N_6840,N_4363,N_4490);
nor U6841 (N_6841,N_5355,N_5152);
nor U6842 (N_6842,N_5483,N_5873);
or U6843 (N_6843,N_5177,N_5801);
and U6844 (N_6844,N_5157,N_5876);
or U6845 (N_6845,N_5027,N_4666);
nor U6846 (N_6846,N_4474,N_4699);
and U6847 (N_6847,N_5993,N_4598);
and U6848 (N_6848,N_5007,N_4178);
or U6849 (N_6849,N_4324,N_5740);
or U6850 (N_6850,N_5081,N_4493);
or U6851 (N_6851,N_4198,N_5197);
xor U6852 (N_6852,N_4091,N_5585);
and U6853 (N_6853,N_4738,N_4665);
or U6854 (N_6854,N_4849,N_4850);
nand U6855 (N_6855,N_4777,N_5869);
nand U6856 (N_6856,N_4449,N_5342);
and U6857 (N_6857,N_5001,N_4550);
nand U6858 (N_6858,N_5595,N_5179);
nor U6859 (N_6859,N_4685,N_5278);
nand U6860 (N_6860,N_4075,N_4422);
and U6861 (N_6861,N_4630,N_4950);
or U6862 (N_6862,N_4813,N_5591);
and U6863 (N_6863,N_5668,N_5253);
xnor U6864 (N_6864,N_5775,N_5241);
and U6865 (N_6865,N_4415,N_4612);
nor U6866 (N_6866,N_4141,N_5224);
and U6867 (N_6867,N_5988,N_4996);
nor U6868 (N_6868,N_4201,N_5516);
or U6869 (N_6869,N_4483,N_4572);
xnor U6870 (N_6870,N_4467,N_4586);
or U6871 (N_6871,N_4252,N_5683);
xnor U6872 (N_6872,N_4343,N_5933);
xor U6873 (N_6873,N_4299,N_5808);
or U6874 (N_6874,N_5147,N_4567);
nor U6875 (N_6875,N_4578,N_5006);
nor U6876 (N_6876,N_5660,N_4132);
and U6877 (N_6877,N_5195,N_4216);
or U6878 (N_6878,N_4842,N_5360);
nand U6879 (N_6879,N_5755,N_5954);
nand U6880 (N_6880,N_4272,N_4098);
and U6881 (N_6881,N_4725,N_4708);
nor U6882 (N_6882,N_5959,N_5546);
or U6883 (N_6883,N_5858,N_4087);
or U6884 (N_6884,N_5054,N_5066);
and U6885 (N_6885,N_4947,N_5637);
xnor U6886 (N_6886,N_5991,N_4287);
nor U6887 (N_6887,N_4043,N_4865);
or U6888 (N_6888,N_5379,N_5616);
xnor U6889 (N_6889,N_4653,N_4023);
xor U6890 (N_6890,N_5201,N_4844);
nand U6891 (N_6891,N_5353,N_5751);
and U6892 (N_6892,N_5417,N_5503);
xor U6893 (N_6893,N_5788,N_5423);
nand U6894 (N_6894,N_4898,N_4342);
nor U6895 (N_6895,N_4190,N_4769);
nand U6896 (N_6896,N_5840,N_4144);
and U6897 (N_6897,N_4966,N_5371);
xor U6898 (N_6898,N_4357,N_5509);
nor U6899 (N_6899,N_4536,N_5684);
nor U6900 (N_6900,N_5070,N_4148);
nor U6901 (N_6901,N_5999,N_4564);
nand U6902 (N_6902,N_5836,N_5033);
nor U6903 (N_6903,N_4094,N_4830);
nor U6904 (N_6904,N_4089,N_4677);
or U6905 (N_6905,N_5274,N_4184);
xnor U6906 (N_6906,N_5306,N_5077);
or U6907 (N_6907,N_4475,N_4580);
xnor U6908 (N_6908,N_4529,N_5405);
nand U6909 (N_6909,N_4465,N_5784);
or U6910 (N_6910,N_4711,N_4962);
and U6911 (N_6911,N_5202,N_5965);
xnor U6912 (N_6912,N_5386,N_4997);
nor U6913 (N_6913,N_4447,N_4511);
nor U6914 (N_6914,N_5621,N_4226);
or U6915 (N_6915,N_5067,N_4857);
nand U6916 (N_6916,N_4701,N_5493);
or U6917 (N_6917,N_4199,N_4440);
or U6918 (N_6918,N_5354,N_4082);
and U6919 (N_6919,N_4480,N_5825);
and U6920 (N_6920,N_4566,N_4135);
nor U6921 (N_6921,N_5315,N_4922);
or U6922 (N_6922,N_5723,N_4197);
xnor U6923 (N_6923,N_5549,N_5612);
nand U6924 (N_6924,N_4737,N_4260);
or U6925 (N_6925,N_4423,N_5987);
xor U6926 (N_6926,N_5777,N_4696);
nor U6927 (N_6927,N_4894,N_5540);
nor U6928 (N_6928,N_5085,N_5574);
or U6929 (N_6929,N_4938,N_4168);
nand U6930 (N_6930,N_4470,N_5968);
xor U6931 (N_6931,N_4471,N_5829);
nor U6932 (N_6932,N_4279,N_5366);
nand U6933 (N_6933,N_4613,N_4559);
or U6934 (N_6934,N_5961,N_5167);
nand U6935 (N_6935,N_5578,N_4581);
nor U6936 (N_6936,N_4741,N_4242);
xnor U6937 (N_6937,N_5783,N_5594);
and U6938 (N_6938,N_5032,N_5025);
or U6939 (N_6939,N_5730,N_4383);
or U6940 (N_6940,N_5262,N_5639);
and U6941 (N_6941,N_4462,N_4017);
or U6942 (N_6942,N_4118,N_4379);
xor U6943 (N_6943,N_4038,N_5885);
or U6944 (N_6944,N_5418,N_4660);
nand U6945 (N_6945,N_5246,N_5451);
nand U6946 (N_6946,N_4126,N_4768);
xnor U6947 (N_6947,N_4005,N_5874);
nand U6948 (N_6948,N_4713,N_5834);
nand U6949 (N_6949,N_4706,N_4392);
and U6950 (N_6950,N_5114,N_4431);
nor U6951 (N_6951,N_5586,N_4359);
or U6952 (N_6952,N_4499,N_5990);
nand U6953 (N_6953,N_4313,N_4182);
and U6954 (N_6954,N_5844,N_4096);
nand U6955 (N_6955,N_4463,N_4013);
and U6956 (N_6956,N_5886,N_4787);
or U6957 (N_6957,N_5666,N_4497);
and U6958 (N_6958,N_4616,N_4349);
or U6959 (N_6959,N_4093,N_5040);
nand U6960 (N_6960,N_4855,N_4050);
xor U6961 (N_6961,N_4209,N_5768);
nor U6962 (N_6962,N_4989,N_5573);
and U6963 (N_6963,N_4409,N_4591);
nand U6964 (N_6964,N_5955,N_5318);
xor U6965 (N_6965,N_4628,N_4206);
nand U6966 (N_6966,N_4958,N_5351);
or U6967 (N_6967,N_4773,N_5378);
or U6968 (N_6968,N_4755,N_4749);
xnor U6969 (N_6969,N_5679,N_4173);
nand U6970 (N_6970,N_4407,N_5046);
and U6971 (N_6971,N_4189,N_5982);
nor U6972 (N_6972,N_5347,N_5400);
nand U6973 (N_6973,N_4614,N_5396);
nand U6974 (N_6974,N_5868,N_5944);
or U6975 (N_6975,N_4631,N_4723);
or U6976 (N_6976,N_4485,N_5055);
nand U6977 (N_6977,N_5919,N_4834);
nor U6978 (N_6978,N_4627,N_5472);
xor U6979 (N_6979,N_5049,N_4373);
nand U6980 (N_6980,N_5139,N_5475);
and U6981 (N_6981,N_4022,N_5672);
xor U6982 (N_6982,N_4278,N_5804);
nand U6983 (N_6983,N_4285,N_5830);
xor U6984 (N_6984,N_4719,N_5324);
or U6985 (N_6985,N_5009,N_4985);
nand U6986 (N_6986,N_5320,N_5719);
xnor U6987 (N_6987,N_5439,N_4574);
and U6988 (N_6988,N_5975,N_4667);
xnor U6989 (N_6989,N_4623,N_4822);
or U6990 (N_6990,N_4221,N_4351);
or U6991 (N_6991,N_5963,N_4071);
nand U6992 (N_6992,N_5909,N_4891);
nor U6993 (N_6993,N_5611,N_4241);
and U6994 (N_6994,N_5839,N_5437);
xnor U6995 (N_6995,N_4006,N_4617);
or U6996 (N_6996,N_4393,N_5260);
nor U6997 (N_6997,N_5499,N_4111);
nand U6998 (N_6998,N_5340,N_5490);
xnor U6999 (N_6999,N_4033,N_4654);
nor U7000 (N_7000,N_5701,N_4543);
nand U7001 (N_7001,N_5934,N_5955);
or U7002 (N_7002,N_4390,N_4290);
nor U7003 (N_7003,N_5972,N_5984);
nand U7004 (N_7004,N_5791,N_5054);
nand U7005 (N_7005,N_5762,N_5038);
nand U7006 (N_7006,N_4081,N_4591);
nor U7007 (N_7007,N_5231,N_5761);
xor U7008 (N_7008,N_5394,N_5674);
or U7009 (N_7009,N_4057,N_4003);
or U7010 (N_7010,N_4144,N_4376);
nand U7011 (N_7011,N_5376,N_4513);
and U7012 (N_7012,N_5418,N_5341);
nand U7013 (N_7013,N_4142,N_4198);
or U7014 (N_7014,N_5659,N_4094);
nor U7015 (N_7015,N_4142,N_4529);
nor U7016 (N_7016,N_4180,N_5113);
or U7017 (N_7017,N_4742,N_5192);
nor U7018 (N_7018,N_4133,N_4498);
and U7019 (N_7019,N_5541,N_5810);
and U7020 (N_7020,N_4080,N_5975);
and U7021 (N_7021,N_4922,N_4406);
nand U7022 (N_7022,N_4105,N_5172);
xor U7023 (N_7023,N_5505,N_4913);
and U7024 (N_7024,N_4301,N_5420);
and U7025 (N_7025,N_4665,N_4245);
xor U7026 (N_7026,N_4428,N_5226);
xor U7027 (N_7027,N_5305,N_4404);
nor U7028 (N_7028,N_4840,N_5629);
xnor U7029 (N_7029,N_5778,N_4683);
xnor U7030 (N_7030,N_5575,N_5508);
xnor U7031 (N_7031,N_4148,N_5988);
nor U7032 (N_7032,N_4798,N_4021);
nor U7033 (N_7033,N_4654,N_4264);
or U7034 (N_7034,N_4587,N_5901);
or U7035 (N_7035,N_5602,N_4599);
nor U7036 (N_7036,N_4309,N_4439);
nand U7037 (N_7037,N_4001,N_4297);
nand U7038 (N_7038,N_4417,N_4859);
or U7039 (N_7039,N_5592,N_5794);
or U7040 (N_7040,N_5239,N_5383);
and U7041 (N_7041,N_5847,N_4368);
or U7042 (N_7042,N_5112,N_5336);
or U7043 (N_7043,N_4936,N_5089);
nand U7044 (N_7044,N_4752,N_5862);
nor U7045 (N_7045,N_4674,N_4814);
nand U7046 (N_7046,N_5398,N_5043);
or U7047 (N_7047,N_5365,N_5371);
or U7048 (N_7048,N_4528,N_4620);
xor U7049 (N_7049,N_4272,N_5827);
and U7050 (N_7050,N_5004,N_4123);
nand U7051 (N_7051,N_5997,N_4840);
and U7052 (N_7052,N_5410,N_4531);
or U7053 (N_7053,N_4690,N_4883);
nand U7054 (N_7054,N_5466,N_5481);
nand U7055 (N_7055,N_4068,N_5236);
nor U7056 (N_7056,N_4007,N_4733);
nor U7057 (N_7057,N_5630,N_5133);
or U7058 (N_7058,N_4067,N_5080);
nor U7059 (N_7059,N_5931,N_5745);
xnor U7060 (N_7060,N_5070,N_4692);
nand U7061 (N_7061,N_4491,N_5386);
and U7062 (N_7062,N_5051,N_5950);
nor U7063 (N_7063,N_4793,N_4292);
nand U7064 (N_7064,N_5467,N_5863);
or U7065 (N_7065,N_5859,N_5630);
xnor U7066 (N_7066,N_5479,N_4885);
xor U7067 (N_7067,N_5310,N_4794);
nor U7068 (N_7068,N_5844,N_5656);
xnor U7069 (N_7069,N_4098,N_5633);
nand U7070 (N_7070,N_4089,N_5097);
or U7071 (N_7071,N_5357,N_4599);
or U7072 (N_7072,N_5511,N_4305);
or U7073 (N_7073,N_4828,N_4928);
xnor U7074 (N_7074,N_4499,N_5123);
xor U7075 (N_7075,N_5472,N_5589);
and U7076 (N_7076,N_5623,N_4541);
and U7077 (N_7077,N_5896,N_5351);
and U7078 (N_7078,N_5637,N_5262);
or U7079 (N_7079,N_5193,N_4423);
and U7080 (N_7080,N_4941,N_5647);
xor U7081 (N_7081,N_5414,N_5900);
nor U7082 (N_7082,N_4150,N_5046);
nand U7083 (N_7083,N_4836,N_4994);
or U7084 (N_7084,N_5109,N_5174);
and U7085 (N_7085,N_4959,N_4789);
nor U7086 (N_7086,N_5293,N_4393);
xor U7087 (N_7087,N_4318,N_4836);
nand U7088 (N_7088,N_5497,N_5441);
and U7089 (N_7089,N_5380,N_5583);
xor U7090 (N_7090,N_5922,N_5208);
xnor U7091 (N_7091,N_4628,N_5326);
nor U7092 (N_7092,N_5072,N_4926);
nand U7093 (N_7093,N_4613,N_4414);
nor U7094 (N_7094,N_4737,N_4682);
xnor U7095 (N_7095,N_4237,N_5202);
nor U7096 (N_7096,N_4540,N_5034);
nor U7097 (N_7097,N_5024,N_5740);
nor U7098 (N_7098,N_5202,N_5838);
nand U7099 (N_7099,N_5306,N_5727);
or U7100 (N_7100,N_4654,N_5726);
nand U7101 (N_7101,N_5380,N_4154);
xor U7102 (N_7102,N_4368,N_4190);
and U7103 (N_7103,N_5201,N_4002);
nor U7104 (N_7104,N_4756,N_5101);
nor U7105 (N_7105,N_4872,N_4081);
nand U7106 (N_7106,N_5087,N_4984);
nor U7107 (N_7107,N_5667,N_5535);
nor U7108 (N_7108,N_5330,N_5970);
nand U7109 (N_7109,N_5561,N_5455);
and U7110 (N_7110,N_4990,N_5377);
nor U7111 (N_7111,N_5933,N_5902);
and U7112 (N_7112,N_4801,N_4109);
and U7113 (N_7113,N_5219,N_5856);
or U7114 (N_7114,N_5778,N_4500);
xor U7115 (N_7115,N_4699,N_5193);
nand U7116 (N_7116,N_5088,N_4104);
or U7117 (N_7117,N_5405,N_5481);
nor U7118 (N_7118,N_5314,N_5485);
or U7119 (N_7119,N_4091,N_5788);
nand U7120 (N_7120,N_4319,N_4656);
and U7121 (N_7121,N_5886,N_5591);
nand U7122 (N_7122,N_4042,N_4095);
or U7123 (N_7123,N_5589,N_5940);
and U7124 (N_7124,N_5980,N_4982);
or U7125 (N_7125,N_5134,N_4233);
nor U7126 (N_7126,N_5444,N_5082);
or U7127 (N_7127,N_5056,N_4708);
nand U7128 (N_7128,N_4672,N_5455);
nor U7129 (N_7129,N_4099,N_4454);
or U7130 (N_7130,N_4735,N_5461);
nand U7131 (N_7131,N_4811,N_4034);
or U7132 (N_7132,N_5754,N_5874);
or U7133 (N_7133,N_5986,N_4756);
nand U7134 (N_7134,N_4723,N_4790);
nor U7135 (N_7135,N_4876,N_5722);
or U7136 (N_7136,N_4487,N_5590);
nor U7137 (N_7137,N_4313,N_4388);
xor U7138 (N_7138,N_5396,N_4200);
nor U7139 (N_7139,N_4231,N_4429);
xnor U7140 (N_7140,N_4636,N_4442);
and U7141 (N_7141,N_5391,N_4872);
or U7142 (N_7142,N_4950,N_5381);
or U7143 (N_7143,N_4885,N_4139);
and U7144 (N_7144,N_5766,N_5128);
and U7145 (N_7145,N_4142,N_4589);
and U7146 (N_7146,N_4327,N_4751);
nor U7147 (N_7147,N_4239,N_4815);
or U7148 (N_7148,N_4738,N_4504);
nor U7149 (N_7149,N_5760,N_5641);
nand U7150 (N_7150,N_4512,N_4314);
or U7151 (N_7151,N_5863,N_4535);
and U7152 (N_7152,N_4900,N_5297);
and U7153 (N_7153,N_5019,N_4297);
and U7154 (N_7154,N_5179,N_5357);
or U7155 (N_7155,N_5511,N_5169);
nand U7156 (N_7156,N_5670,N_4621);
or U7157 (N_7157,N_4117,N_4053);
nor U7158 (N_7158,N_4787,N_4975);
and U7159 (N_7159,N_5767,N_5992);
xor U7160 (N_7160,N_4571,N_5020);
or U7161 (N_7161,N_5249,N_5530);
and U7162 (N_7162,N_4846,N_5944);
nand U7163 (N_7163,N_4305,N_5999);
or U7164 (N_7164,N_5936,N_4935);
or U7165 (N_7165,N_4553,N_5687);
nand U7166 (N_7166,N_4953,N_4420);
nand U7167 (N_7167,N_4672,N_4552);
or U7168 (N_7168,N_5308,N_5552);
and U7169 (N_7169,N_4871,N_5933);
nor U7170 (N_7170,N_5953,N_5496);
and U7171 (N_7171,N_5461,N_5224);
xnor U7172 (N_7172,N_5437,N_4806);
xor U7173 (N_7173,N_4919,N_4525);
xor U7174 (N_7174,N_5169,N_5165);
or U7175 (N_7175,N_4914,N_4666);
xor U7176 (N_7176,N_5493,N_4982);
xor U7177 (N_7177,N_5794,N_4150);
nand U7178 (N_7178,N_4417,N_4933);
and U7179 (N_7179,N_5752,N_5448);
xor U7180 (N_7180,N_4965,N_5949);
nand U7181 (N_7181,N_5212,N_4144);
or U7182 (N_7182,N_5486,N_5034);
or U7183 (N_7183,N_4908,N_5856);
and U7184 (N_7184,N_4078,N_4415);
nand U7185 (N_7185,N_4508,N_4947);
nand U7186 (N_7186,N_5514,N_4143);
or U7187 (N_7187,N_5403,N_4895);
and U7188 (N_7188,N_4375,N_5963);
or U7189 (N_7189,N_5496,N_5923);
xor U7190 (N_7190,N_4981,N_5308);
xor U7191 (N_7191,N_5082,N_4357);
xnor U7192 (N_7192,N_5850,N_5910);
xor U7193 (N_7193,N_4875,N_4922);
nor U7194 (N_7194,N_5003,N_4189);
xnor U7195 (N_7195,N_4983,N_4450);
nor U7196 (N_7196,N_5071,N_4048);
nor U7197 (N_7197,N_4361,N_4438);
xor U7198 (N_7198,N_4185,N_4508);
xnor U7199 (N_7199,N_5917,N_4959);
or U7200 (N_7200,N_5677,N_5782);
nand U7201 (N_7201,N_4298,N_4687);
nand U7202 (N_7202,N_4902,N_5613);
xor U7203 (N_7203,N_5046,N_5353);
nand U7204 (N_7204,N_5674,N_5206);
xnor U7205 (N_7205,N_5490,N_4557);
and U7206 (N_7206,N_4881,N_4235);
and U7207 (N_7207,N_5256,N_4292);
xnor U7208 (N_7208,N_5738,N_5187);
xor U7209 (N_7209,N_5721,N_5912);
xnor U7210 (N_7210,N_5432,N_5736);
and U7211 (N_7211,N_4553,N_5726);
nand U7212 (N_7212,N_5981,N_4008);
xnor U7213 (N_7213,N_5949,N_5206);
nand U7214 (N_7214,N_4088,N_4719);
nand U7215 (N_7215,N_4699,N_4492);
xnor U7216 (N_7216,N_5284,N_5481);
or U7217 (N_7217,N_4879,N_5859);
nand U7218 (N_7218,N_4653,N_4088);
nand U7219 (N_7219,N_5391,N_5353);
or U7220 (N_7220,N_5531,N_4720);
nand U7221 (N_7221,N_5390,N_4291);
nor U7222 (N_7222,N_4999,N_5545);
nor U7223 (N_7223,N_5423,N_5362);
nor U7224 (N_7224,N_5733,N_4375);
and U7225 (N_7225,N_4790,N_4750);
nand U7226 (N_7226,N_4847,N_5319);
and U7227 (N_7227,N_5385,N_5094);
nand U7228 (N_7228,N_4485,N_4250);
nor U7229 (N_7229,N_4176,N_5416);
nor U7230 (N_7230,N_4169,N_4738);
xnor U7231 (N_7231,N_4016,N_4832);
or U7232 (N_7232,N_5416,N_5523);
or U7233 (N_7233,N_5124,N_5516);
nor U7234 (N_7234,N_5760,N_5501);
xor U7235 (N_7235,N_5458,N_4170);
xnor U7236 (N_7236,N_5027,N_4117);
nand U7237 (N_7237,N_5660,N_4451);
and U7238 (N_7238,N_5701,N_5454);
nor U7239 (N_7239,N_5544,N_5169);
or U7240 (N_7240,N_5332,N_5004);
and U7241 (N_7241,N_5806,N_5539);
nand U7242 (N_7242,N_4434,N_5793);
xor U7243 (N_7243,N_5107,N_4645);
xor U7244 (N_7244,N_4748,N_5659);
nand U7245 (N_7245,N_4200,N_4823);
and U7246 (N_7246,N_5576,N_5903);
or U7247 (N_7247,N_5761,N_4509);
and U7248 (N_7248,N_5799,N_4841);
and U7249 (N_7249,N_4147,N_5877);
xnor U7250 (N_7250,N_5399,N_5848);
xor U7251 (N_7251,N_5921,N_4633);
and U7252 (N_7252,N_4292,N_4481);
nand U7253 (N_7253,N_5081,N_5717);
nor U7254 (N_7254,N_5014,N_5583);
nand U7255 (N_7255,N_4829,N_5440);
nand U7256 (N_7256,N_4819,N_5123);
and U7257 (N_7257,N_5172,N_5090);
and U7258 (N_7258,N_4869,N_5105);
and U7259 (N_7259,N_5506,N_4456);
or U7260 (N_7260,N_5695,N_4113);
and U7261 (N_7261,N_5338,N_4311);
and U7262 (N_7262,N_4987,N_4823);
nand U7263 (N_7263,N_5458,N_4812);
xor U7264 (N_7264,N_5505,N_5504);
nand U7265 (N_7265,N_4621,N_4911);
xnor U7266 (N_7266,N_5442,N_4416);
or U7267 (N_7267,N_4468,N_4783);
nor U7268 (N_7268,N_5363,N_5208);
nor U7269 (N_7269,N_5535,N_4465);
or U7270 (N_7270,N_5860,N_4865);
or U7271 (N_7271,N_4814,N_5590);
xnor U7272 (N_7272,N_4342,N_5602);
nor U7273 (N_7273,N_5618,N_4212);
or U7274 (N_7274,N_4063,N_5486);
nor U7275 (N_7275,N_4038,N_4355);
xor U7276 (N_7276,N_5582,N_4735);
or U7277 (N_7277,N_5627,N_5125);
and U7278 (N_7278,N_5963,N_5688);
nor U7279 (N_7279,N_5574,N_4422);
or U7280 (N_7280,N_4276,N_5916);
xnor U7281 (N_7281,N_4120,N_5739);
nor U7282 (N_7282,N_5493,N_4955);
and U7283 (N_7283,N_4729,N_5551);
nor U7284 (N_7284,N_5710,N_5745);
nor U7285 (N_7285,N_5027,N_4332);
xor U7286 (N_7286,N_5612,N_4394);
nor U7287 (N_7287,N_5512,N_4664);
nand U7288 (N_7288,N_4632,N_5001);
nand U7289 (N_7289,N_4406,N_5036);
xor U7290 (N_7290,N_5381,N_5348);
xnor U7291 (N_7291,N_5385,N_4294);
nor U7292 (N_7292,N_4369,N_4495);
nor U7293 (N_7293,N_5493,N_5206);
nor U7294 (N_7294,N_4514,N_4208);
and U7295 (N_7295,N_5366,N_5727);
nor U7296 (N_7296,N_5672,N_4941);
nor U7297 (N_7297,N_5983,N_5519);
xnor U7298 (N_7298,N_4859,N_4075);
nand U7299 (N_7299,N_5771,N_4060);
nor U7300 (N_7300,N_5875,N_5871);
xor U7301 (N_7301,N_5238,N_5551);
and U7302 (N_7302,N_5462,N_5468);
and U7303 (N_7303,N_5380,N_5837);
and U7304 (N_7304,N_4885,N_5934);
nor U7305 (N_7305,N_5905,N_4067);
xnor U7306 (N_7306,N_5551,N_5695);
nor U7307 (N_7307,N_5665,N_4675);
and U7308 (N_7308,N_5804,N_5480);
nand U7309 (N_7309,N_5005,N_4525);
and U7310 (N_7310,N_4228,N_5766);
nor U7311 (N_7311,N_4020,N_4022);
xnor U7312 (N_7312,N_4448,N_5556);
and U7313 (N_7313,N_5418,N_5519);
or U7314 (N_7314,N_5378,N_4753);
or U7315 (N_7315,N_5890,N_4827);
or U7316 (N_7316,N_4226,N_4006);
nand U7317 (N_7317,N_5687,N_4994);
nor U7318 (N_7318,N_4258,N_5914);
xnor U7319 (N_7319,N_5574,N_4387);
and U7320 (N_7320,N_4652,N_4385);
xnor U7321 (N_7321,N_4014,N_5878);
xor U7322 (N_7322,N_5678,N_5896);
or U7323 (N_7323,N_5486,N_4803);
or U7324 (N_7324,N_4555,N_4023);
or U7325 (N_7325,N_4507,N_5566);
nor U7326 (N_7326,N_4073,N_5674);
nor U7327 (N_7327,N_5905,N_4497);
nor U7328 (N_7328,N_4724,N_5261);
nand U7329 (N_7329,N_4868,N_5760);
xor U7330 (N_7330,N_4094,N_5691);
nand U7331 (N_7331,N_4947,N_5535);
nor U7332 (N_7332,N_4096,N_4684);
and U7333 (N_7333,N_5152,N_5981);
xnor U7334 (N_7334,N_4999,N_4091);
nand U7335 (N_7335,N_5020,N_5366);
nor U7336 (N_7336,N_4187,N_4113);
nand U7337 (N_7337,N_5085,N_5867);
nor U7338 (N_7338,N_4386,N_5094);
nor U7339 (N_7339,N_5855,N_5919);
xnor U7340 (N_7340,N_5347,N_5043);
or U7341 (N_7341,N_4840,N_4892);
and U7342 (N_7342,N_5671,N_4638);
nor U7343 (N_7343,N_4321,N_4802);
xnor U7344 (N_7344,N_5061,N_4251);
nand U7345 (N_7345,N_4858,N_5426);
nand U7346 (N_7346,N_5647,N_5729);
nand U7347 (N_7347,N_4666,N_5267);
or U7348 (N_7348,N_5901,N_4463);
nand U7349 (N_7349,N_5337,N_4564);
and U7350 (N_7350,N_4751,N_4643);
xnor U7351 (N_7351,N_4724,N_4619);
nand U7352 (N_7352,N_4597,N_4661);
or U7353 (N_7353,N_5428,N_5578);
xnor U7354 (N_7354,N_5532,N_4491);
or U7355 (N_7355,N_4152,N_4322);
xor U7356 (N_7356,N_5827,N_5830);
nor U7357 (N_7357,N_4553,N_4531);
and U7358 (N_7358,N_5796,N_5776);
xor U7359 (N_7359,N_5563,N_4149);
and U7360 (N_7360,N_5087,N_4549);
xor U7361 (N_7361,N_4732,N_5108);
nor U7362 (N_7362,N_5948,N_5285);
or U7363 (N_7363,N_4452,N_4265);
xnor U7364 (N_7364,N_5674,N_5993);
xnor U7365 (N_7365,N_5200,N_5042);
or U7366 (N_7366,N_5666,N_5641);
or U7367 (N_7367,N_5329,N_4052);
or U7368 (N_7368,N_4799,N_5041);
and U7369 (N_7369,N_5825,N_4647);
nand U7370 (N_7370,N_5135,N_5105);
or U7371 (N_7371,N_4802,N_4866);
nand U7372 (N_7372,N_4005,N_5827);
nand U7373 (N_7373,N_4918,N_4984);
xor U7374 (N_7374,N_5066,N_4376);
nand U7375 (N_7375,N_4730,N_4432);
xnor U7376 (N_7376,N_5299,N_4679);
or U7377 (N_7377,N_5268,N_5629);
or U7378 (N_7378,N_5338,N_4600);
nand U7379 (N_7379,N_5176,N_5525);
or U7380 (N_7380,N_5601,N_5701);
nor U7381 (N_7381,N_5654,N_5328);
or U7382 (N_7382,N_5540,N_5884);
and U7383 (N_7383,N_5002,N_5098);
nor U7384 (N_7384,N_5027,N_4100);
xor U7385 (N_7385,N_4722,N_4600);
or U7386 (N_7386,N_5570,N_5460);
and U7387 (N_7387,N_4147,N_4607);
or U7388 (N_7388,N_4110,N_4742);
xnor U7389 (N_7389,N_5724,N_4256);
or U7390 (N_7390,N_5028,N_5121);
or U7391 (N_7391,N_4017,N_4635);
or U7392 (N_7392,N_5241,N_5875);
and U7393 (N_7393,N_5458,N_5656);
xor U7394 (N_7394,N_5583,N_4695);
nand U7395 (N_7395,N_5157,N_5364);
xor U7396 (N_7396,N_4075,N_5567);
nand U7397 (N_7397,N_5203,N_4530);
or U7398 (N_7398,N_5698,N_4631);
and U7399 (N_7399,N_4948,N_4778);
and U7400 (N_7400,N_5075,N_4229);
or U7401 (N_7401,N_5524,N_4451);
nor U7402 (N_7402,N_4212,N_5364);
nand U7403 (N_7403,N_4536,N_4258);
nor U7404 (N_7404,N_4240,N_4223);
nand U7405 (N_7405,N_5674,N_5983);
nor U7406 (N_7406,N_4607,N_5008);
nor U7407 (N_7407,N_5533,N_5758);
or U7408 (N_7408,N_5812,N_4178);
and U7409 (N_7409,N_5922,N_5016);
xnor U7410 (N_7410,N_4011,N_4945);
nand U7411 (N_7411,N_4688,N_5348);
nand U7412 (N_7412,N_5861,N_5622);
xor U7413 (N_7413,N_5251,N_5802);
nand U7414 (N_7414,N_4943,N_4017);
nor U7415 (N_7415,N_4772,N_5925);
and U7416 (N_7416,N_4275,N_4896);
nor U7417 (N_7417,N_4636,N_5928);
and U7418 (N_7418,N_4263,N_5184);
nor U7419 (N_7419,N_5993,N_5728);
or U7420 (N_7420,N_5170,N_4568);
nor U7421 (N_7421,N_5718,N_4423);
or U7422 (N_7422,N_4904,N_5897);
xnor U7423 (N_7423,N_4510,N_5863);
nor U7424 (N_7424,N_5817,N_4226);
or U7425 (N_7425,N_5826,N_5315);
nand U7426 (N_7426,N_5825,N_5855);
nand U7427 (N_7427,N_4413,N_5026);
or U7428 (N_7428,N_4319,N_5783);
and U7429 (N_7429,N_4041,N_4963);
and U7430 (N_7430,N_5561,N_4878);
and U7431 (N_7431,N_5463,N_5893);
xnor U7432 (N_7432,N_4328,N_4482);
or U7433 (N_7433,N_4216,N_5198);
or U7434 (N_7434,N_5391,N_5654);
and U7435 (N_7435,N_5211,N_5844);
nor U7436 (N_7436,N_5838,N_5327);
nor U7437 (N_7437,N_4582,N_5818);
and U7438 (N_7438,N_4432,N_4761);
nand U7439 (N_7439,N_4241,N_5128);
or U7440 (N_7440,N_5765,N_4631);
and U7441 (N_7441,N_5112,N_5643);
nor U7442 (N_7442,N_5297,N_5560);
nor U7443 (N_7443,N_4108,N_4411);
xnor U7444 (N_7444,N_5781,N_4307);
xnor U7445 (N_7445,N_4754,N_5989);
and U7446 (N_7446,N_4369,N_4036);
xor U7447 (N_7447,N_4581,N_5159);
xnor U7448 (N_7448,N_5063,N_5299);
or U7449 (N_7449,N_5231,N_5431);
and U7450 (N_7450,N_5538,N_4229);
nor U7451 (N_7451,N_4305,N_4925);
nor U7452 (N_7452,N_4566,N_5942);
xor U7453 (N_7453,N_5415,N_4527);
nand U7454 (N_7454,N_4872,N_4539);
and U7455 (N_7455,N_5064,N_5491);
and U7456 (N_7456,N_4650,N_5403);
or U7457 (N_7457,N_4781,N_4782);
and U7458 (N_7458,N_5149,N_5296);
xnor U7459 (N_7459,N_5390,N_5521);
nand U7460 (N_7460,N_5683,N_4004);
xnor U7461 (N_7461,N_4835,N_5144);
xor U7462 (N_7462,N_5121,N_5727);
xor U7463 (N_7463,N_5180,N_4443);
or U7464 (N_7464,N_4457,N_4992);
nor U7465 (N_7465,N_5147,N_5381);
xnor U7466 (N_7466,N_4466,N_4015);
and U7467 (N_7467,N_5966,N_4619);
and U7468 (N_7468,N_5485,N_5756);
nand U7469 (N_7469,N_4320,N_4802);
and U7470 (N_7470,N_4100,N_5920);
or U7471 (N_7471,N_4083,N_5007);
or U7472 (N_7472,N_4878,N_4155);
xnor U7473 (N_7473,N_4531,N_4834);
and U7474 (N_7474,N_4476,N_5532);
or U7475 (N_7475,N_5656,N_4890);
nand U7476 (N_7476,N_4129,N_5909);
or U7477 (N_7477,N_4253,N_5070);
xnor U7478 (N_7478,N_5836,N_5510);
nand U7479 (N_7479,N_5427,N_4872);
xnor U7480 (N_7480,N_4958,N_4211);
or U7481 (N_7481,N_4971,N_5358);
xor U7482 (N_7482,N_5245,N_5845);
xor U7483 (N_7483,N_5754,N_4687);
nor U7484 (N_7484,N_4172,N_4878);
and U7485 (N_7485,N_5097,N_5016);
or U7486 (N_7486,N_4235,N_5860);
xor U7487 (N_7487,N_5342,N_4383);
nand U7488 (N_7488,N_5287,N_4034);
and U7489 (N_7489,N_4274,N_4330);
and U7490 (N_7490,N_4915,N_5441);
or U7491 (N_7491,N_5674,N_4495);
or U7492 (N_7492,N_4626,N_5349);
nor U7493 (N_7493,N_4113,N_5281);
xnor U7494 (N_7494,N_5828,N_4312);
or U7495 (N_7495,N_4202,N_4444);
nor U7496 (N_7496,N_5014,N_4838);
and U7497 (N_7497,N_4494,N_4933);
nor U7498 (N_7498,N_4004,N_5629);
nor U7499 (N_7499,N_4699,N_4922);
xnor U7500 (N_7500,N_4921,N_5366);
or U7501 (N_7501,N_4228,N_5590);
or U7502 (N_7502,N_5178,N_4787);
xnor U7503 (N_7503,N_4097,N_4811);
and U7504 (N_7504,N_4256,N_5188);
xor U7505 (N_7505,N_5361,N_5307);
and U7506 (N_7506,N_4392,N_5949);
and U7507 (N_7507,N_5097,N_5893);
and U7508 (N_7508,N_4681,N_4060);
and U7509 (N_7509,N_4712,N_4219);
and U7510 (N_7510,N_4430,N_5592);
nor U7511 (N_7511,N_4069,N_5172);
xnor U7512 (N_7512,N_4882,N_4560);
or U7513 (N_7513,N_5280,N_4777);
and U7514 (N_7514,N_4689,N_5239);
xor U7515 (N_7515,N_5445,N_4662);
nor U7516 (N_7516,N_4553,N_5979);
nand U7517 (N_7517,N_4266,N_5465);
and U7518 (N_7518,N_4024,N_5375);
xnor U7519 (N_7519,N_5982,N_5785);
or U7520 (N_7520,N_4448,N_4371);
nand U7521 (N_7521,N_4185,N_4769);
and U7522 (N_7522,N_4952,N_5546);
nor U7523 (N_7523,N_5626,N_4991);
nand U7524 (N_7524,N_5184,N_4508);
or U7525 (N_7525,N_4449,N_4878);
nand U7526 (N_7526,N_5294,N_4637);
xor U7527 (N_7527,N_4300,N_4338);
nor U7528 (N_7528,N_4179,N_5199);
or U7529 (N_7529,N_4397,N_5796);
nand U7530 (N_7530,N_4992,N_4183);
and U7531 (N_7531,N_5227,N_5420);
or U7532 (N_7532,N_5396,N_5500);
nor U7533 (N_7533,N_5373,N_5194);
nand U7534 (N_7534,N_5704,N_5258);
nor U7535 (N_7535,N_4253,N_5555);
xor U7536 (N_7536,N_5066,N_4343);
nand U7537 (N_7537,N_4514,N_5851);
nor U7538 (N_7538,N_5759,N_5283);
and U7539 (N_7539,N_5101,N_4337);
and U7540 (N_7540,N_4823,N_4380);
or U7541 (N_7541,N_5651,N_5767);
and U7542 (N_7542,N_5435,N_5690);
or U7543 (N_7543,N_4258,N_5708);
and U7544 (N_7544,N_4501,N_4130);
and U7545 (N_7545,N_5600,N_5159);
or U7546 (N_7546,N_4973,N_4473);
xor U7547 (N_7547,N_4920,N_4929);
nand U7548 (N_7548,N_5859,N_4601);
nand U7549 (N_7549,N_4900,N_4661);
or U7550 (N_7550,N_4032,N_5055);
and U7551 (N_7551,N_4873,N_4319);
and U7552 (N_7552,N_4229,N_5242);
xor U7553 (N_7553,N_4447,N_4387);
nor U7554 (N_7554,N_4852,N_5233);
and U7555 (N_7555,N_5997,N_4896);
nor U7556 (N_7556,N_4008,N_4997);
and U7557 (N_7557,N_4177,N_5196);
nand U7558 (N_7558,N_4955,N_5132);
or U7559 (N_7559,N_5281,N_4156);
nor U7560 (N_7560,N_4851,N_5921);
and U7561 (N_7561,N_5739,N_5890);
xor U7562 (N_7562,N_4280,N_5692);
xor U7563 (N_7563,N_4379,N_4971);
nand U7564 (N_7564,N_5218,N_5631);
nand U7565 (N_7565,N_4065,N_5734);
nand U7566 (N_7566,N_5585,N_4603);
xor U7567 (N_7567,N_5631,N_4746);
nand U7568 (N_7568,N_5612,N_4688);
nor U7569 (N_7569,N_5408,N_4072);
or U7570 (N_7570,N_5842,N_4540);
nor U7571 (N_7571,N_5030,N_4130);
or U7572 (N_7572,N_5031,N_4824);
and U7573 (N_7573,N_5055,N_5753);
nand U7574 (N_7574,N_5788,N_4075);
or U7575 (N_7575,N_5062,N_5859);
xnor U7576 (N_7576,N_4177,N_5209);
nand U7577 (N_7577,N_4726,N_5110);
or U7578 (N_7578,N_5366,N_4473);
xor U7579 (N_7579,N_4079,N_4698);
nor U7580 (N_7580,N_5940,N_4883);
and U7581 (N_7581,N_4748,N_4790);
nor U7582 (N_7582,N_4605,N_5293);
xor U7583 (N_7583,N_4023,N_4974);
nand U7584 (N_7584,N_4309,N_4463);
xor U7585 (N_7585,N_5569,N_4042);
or U7586 (N_7586,N_4241,N_5402);
nand U7587 (N_7587,N_5488,N_5250);
or U7588 (N_7588,N_5435,N_5382);
or U7589 (N_7589,N_5645,N_4636);
nor U7590 (N_7590,N_5448,N_4525);
xor U7591 (N_7591,N_5489,N_5028);
or U7592 (N_7592,N_5422,N_5425);
and U7593 (N_7593,N_4085,N_5421);
nor U7594 (N_7594,N_5640,N_4676);
or U7595 (N_7595,N_5289,N_5627);
xor U7596 (N_7596,N_5040,N_5441);
xnor U7597 (N_7597,N_4759,N_4267);
xnor U7598 (N_7598,N_5938,N_4778);
xnor U7599 (N_7599,N_5397,N_5321);
xnor U7600 (N_7600,N_5946,N_4950);
or U7601 (N_7601,N_5097,N_4648);
or U7602 (N_7602,N_4476,N_4613);
or U7603 (N_7603,N_5440,N_5347);
xor U7604 (N_7604,N_5695,N_4949);
and U7605 (N_7605,N_5908,N_5491);
or U7606 (N_7606,N_5210,N_4160);
nand U7607 (N_7607,N_4236,N_5852);
nand U7608 (N_7608,N_4671,N_5701);
xnor U7609 (N_7609,N_4828,N_5322);
or U7610 (N_7610,N_5088,N_4114);
or U7611 (N_7611,N_5389,N_4685);
xor U7612 (N_7612,N_4028,N_5265);
nand U7613 (N_7613,N_4349,N_5312);
or U7614 (N_7614,N_5207,N_4731);
nor U7615 (N_7615,N_4311,N_4056);
or U7616 (N_7616,N_4858,N_5502);
nand U7617 (N_7617,N_5086,N_4141);
nand U7618 (N_7618,N_5164,N_5439);
and U7619 (N_7619,N_4960,N_5541);
or U7620 (N_7620,N_4712,N_4897);
nor U7621 (N_7621,N_4469,N_5047);
nor U7622 (N_7622,N_4110,N_5359);
and U7623 (N_7623,N_4280,N_5129);
and U7624 (N_7624,N_5892,N_4954);
and U7625 (N_7625,N_5455,N_4464);
and U7626 (N_7626,N_5339,N_5738);
and U7627 (N_7627,N_4608,N_5345);
nand U7628 (N_7628,N_5845,N_5067);
nor U7629 (N_7629,N_5690,N_5024);
or U7630 (N_7630,N_4064,N_4565);
or U7631 (N_7631,N_4263,N_4012);
nor U7632 (N_7632,N_5300,N_4079);
nand U7633 (N_7633,N_5606,N_4683);
nand U7634 (N_7634,N_5337,N_5603);
xnor U7635 (N_7635,N_5765,N_5804);
xnor U7636 (N_7636,N_4735,N_5388);
and U7637 (N_7637,N_5708,N_4498);
nor U7638 (N_7638,N_5428,N_4476);
nand U7639 (N_7639,N_5501,N_5487);
xnor U7640 (N_7640,N_4637,N_5235);
xor U7641 (N_7641,N_4635,N_5704);
and U7642 (N_7642,N_4763,N_5484);
or U7643 (N_7643,N_4030,N_4801);
or U7644 (N_7644,N_5080,N_4758);
or U7645 (N_7645,N_5050,N_4462);
nor U7646 (N_7646,N_4235,N_4610);
nand U7647 (N_7647,N_5026,N_5470);
xnor U7648 (N_7648,N_4552,N_5067);
xnor U7649 (N_7649,N_5429,N_4131);
and U7650 (N_7650,N_4516,N_5014);
xor U7651 (N_7651,N_4854,N_5557);
and U7652 (N_7652,N_4946,N_4954);
xor U7653 (N_7653,N_5218,N_5920);
or U7654 (N_7654,N_4369,N_4795);
and U7655 (N_7655,N_4151,N_5634);
or U7656 (N_7656,N_4639,N_5863);
or U7657 (N_7657,N_4683,N_4924);
and U7658 (N_7658,N_4339,N_5831);
nor U7659 (N_7659,N_5232,N_5137);
or U7660 (N_7660,N_4903,N_4575);
or U7661 (N_7661,N_4976,N_5010);
nand U7662 (N_7662,N_4176,N_5504);
xnor U7663 (N_7663,N_4688,N_5630);
nand U7664 (N_7664,N_5826,N_4605);
nor U7665 (N_7665,N_5787,N_5298);
or U7666 (N_7666,N_4110,N_5046);
and U7667 (N_7667,N_5121,N_5297);
or U7668 (N_7668,N_4318,N_5379);
nand U7669 (N_7669,N_5110,N_5312);
nor U7670 (N_7670,N_5834,N_4576);
nand U7671 (N_7671,N_5751,N_4243);
xnor U7672 (N_7672,N_5163,N_5502);
and U7673 (N_7673,N_5460,N_4596);
xor U7674 (N_7674,N_4278,N_4451);
nand U7675 (N_7675,N_5256,N_4346);
nor U7676 (N_7676,N_5974,N_4164);
nand U7677 (N_7677,N_5854,N_4331);
or U7678 (N_7678,N_4757,N_4168);
and U7679 (N_7679,N_4728,N_4604);
nor U7680 (N_7680,N_5067,N_4669);
xnor U7681 (N_7681,N_5838,N_4136);
nand U7682 (N_7682,N_4819,N_4825);
nand U7683 (N_7683,N_5946,N_5620);
and U7684 (N_7684,N_4953,N_4274);
or U7685 (N_7685,N_4886,N_5883);
nand U7686 (N_7686,N_5433,N_5217);
nor U7687 (N_7687,N_4223,N_4555);
nand U7688 (N_7688,N_4960,N_5462);
nand U7689 (N_7689,N_4129,N_5984);
nand U7690 (N_7690,N_4267,N_4378);
and U7691 (N_7691,N_4238,N_5314);
nand U7692 (N_7692,N_4838,N_5607);
xor U7693 (N_7693,N_4481,N_5499);
nor U7694 (N_7694,N_4040,N_4959);
and U7695 (N_7695,N_4881,N_5496);
and U7696 (N_7696,N_4191,N_5417);
nor U7697 (N_7697,N_5302,N_4509);
and U7698 (N_7698,N_5575,N_5080);
nand U7699 (N_7699,N_5425,N_4519);
and U7700 (N_7700,N_5945,N_5103);
or U7701 (N_7701,N_4801,N_5210);
nor U7702 (N_7702,N_5830,N_4218);
and U7703 (N_7703,N_4218,N_5514);
nand U7704 (N_7704,N_5850,N_5544);
xnor U7705 (N_7705,N_4066,N_4855);
and U7706 (N_7706,N_4112,N_4809);
xnor U7707 (N_7707,N_4627,N_5778);
xor U7708 (N_7708,N_5155,N_4999);
xor U7709 (N_7709,N_5239,N_4080);
or U7710 (N_7710,N_4400,N_4888);
xor U7711 (N_7711,N_5293,N_5871);
xnor U7712 (N_7712,N_5370,N_5262);
and U7713 (N_7713,N_4878,N_5866);
and U7714 (N_7714,N_4064,N_4224);
or U7715 (N_7715,N_5414,N_4966);
nor U7716 (N_7716,N_5496,N_5267);
nor U7717 (N_7717,N_4147,N_4785);
nand U7718 (N_7718,N_4591,N_4800);
or U7719 (N_7719,N_4956,N_4726);
nor U7720 (N_7720,N_5576,N_4326);
xnor U7721 (N_7721,N_5338,N_4933);
xnor U7722 (N_7722,N_5961,N_5884);
nand U7723 (N_7723,N_5247,N_4333);
or U7724 (N_7724,N_5370,N_5082);
and U7725 (N_7725,N_4448,N_4115);
and U7726 (N_7726,N_4258,N_5096);
nand U7727 (N_7727,N_5677,N_4313);
nor U7728 (N_7728,N_5044,N_5381);
xor U7729 (N_7729,N_5273,N_4001);
or U7730 (N_7730,N_4570,N_5696);
and U7731 (N_7731,N_4795,N_5910);
nand U7732 (N_7732,N_5778,N_5606);
xor U7733 (N_7733,N_5259,N_4110);
or U7734 (N_7734,N_5679,N_5734);
nor U7735 (N_7735,N_5371,N_5020);
and U7736 (N_7736,N_4229,N_5672);
and U7737 (N_7737,N_5791,N_4155);
nor U7738 (N_7738,N_5578,N_4866);
and U7739 (N_7739,N_5739,N_4953);
and U7740 (N_7740,N_5994,N_4620);
or U7741 (N_7741,N_5094,N_5182);
nand U7742 (N_7742,N_5365,N_5271);
or U7743 (N_7743,N_4732,N_5034);
nor U7744 (N_7744,N_5062,N_5471);
xor U7745 (N_7745,N_4228,N_5265);
or U7746 (N_7746,N_4167,N_4212);
nor U7747 (N_7747,N_5423,N_4208);
and U7748 (N_7748,N_5350,N_5094);
xor U7749 (N_7749,N_4617,N_4675);
or U7750 (N_7750,N_5180,N_4247);
nor U7751 (N_7751,N_5529,N_5055);
xnor U7752 (N_7752,N_5244,N_4965);
nor U7753 (N_7753,N_4251,N_4451);
nand U7754 (N_7754,N_4447,N_5215);
nor U7755 (N_7755,N_5894,N_5441);
nand U7756 (N_7756,N_4682,N_4330);
xnor U7757 (N_7757,N_5974,N_4335);
nor U7758 (N_7758,N_5762,N_5084);
nand U7759 (N_7759,N_4500,N_5637);
and U7760 (N_7760,N_4809,N_5071);
nand U7761 (N_7761,N_4733,N_5340);
xnor U7762 (N_7762,N_5232,N_5939);
nand U7763 (N_7763,N_4622,N_5609);
and U7764 (N_7764,N_5712,N_4142);
xnor U7765 (N_7765,N_5817,N_5339);
nor U7766 (N_7766,N_5681,N_4623);
xnor U7767 (N_7767,N_5009,N_5076);
and U7768 (N_7768,N_5244,N_4073);
nor U7769 (N_7769,N_5680,N_5843);
xor U7770 (N_7770,N_5050,N_4169);
or U7771 (N_7771,N_4046,N_5937);
xor U7772 (N_7772,N_5301,N_4883);
or U7773 (N_7773,N_5828,N_5104);
and U7774 (N_7774,N_5145,N_4678);
or U7775 (N_7775,N_5117,N_4136);
and U7776 (N_7776,N_4441,N_4140);
nor U7777 (N_7777,N_5495,N_4057);
or U7778 (N_7778,N_4154,N_4528);
nor U7779 (N_7779,N_5465,N_5342);
and U7780 (N_7780,N_5161,N_4103);
nand U7781 (N_7781,N_5088,N_4877);
nor U7782 (N_7782,N_5172,N_4081);
nand U7783 (N_7783,N_4869,N_4323);
nor U7784 (N_7784,N_4268,N_5371);
or U7785 (N_7785,N_4289,N_4709);
or U7786 (N_7786,N_4353,N_5913);
nor U7787 (N_7787,N_5111,N_4525);
xor U7788 (N_7788,N_4409,N_4386);
xnor U7789 (N_7789,N_4225,N_5692);
or U7790 (N_7790,N_4517,N_4411);
nor U7791 (N_7791,N_5227,N_4157);
xor U7792 (N_7792,N_5190,N_4952);
nand U7793 (N_7793,N_4649,N_4236);
nand U7794 (N_7794,N_4151,N_4651);
or U7795 (N_7795,N_4355,N_4692);
nor U7796 (N_7796,N_4141,N_4195);
or U7797 (N_7797,N_5197,N_4373);
nand U7798 (N_7798,N_4907,N_4793);
nand U7799 (N_7799,N_5002,N_4773);
nand U7800 (N_7800,N_4552,N_5229);
and U7801 (N_7801,N_5867,N_5200);
and U7802 (N_7802,N_5786,N_5126);
or U7803 (N_7803,N_4136,N_5979);
nor U7804 (N_7804,N_5451,N_5190);
nor U7805 (N_7805,N_5026,N_4372);
nor U7806 (N_7806,N_4039,N_5903);
nand U7807 (N_7807,N_4427,N_5871);
nor U7808 (N_7808,N_5732,N_5668);
or U7809 (N_7809,N_4606,N_5962);
nor U7810 (N_7810,N_5455,N_4839);
xor U7811 (N_7811,N_4392,N_5073);
and U7812 (N_7812,N_4733,N_4797);
nand U7813 (N_7813,N_5200,N_4721);
and U7814 (N_7814,N_5491,N_5804);
and U7815 (N_7815,N_5814,N_5455);
and U7816 (N_7816,N_4133,N_5950);
and U7817 (N_7817,N_4898,N_5632);
nand U7818 (N_7818,N_5265,N_4181);
xnor U7819 (N_7819,N_4717,N_4701);
xor U7820 (N_7820,N_4999,N_5942);
nand U7821 (N_7821,N_5879,N_4169);
nor U7822 (N_7822,N_4142,N_5783);
nor U7823 (N_7823,N_4394,N_5435);
xor U7824 (N_7824,N_5168,N_4351);
nor U7825 (N_7825,N_4748,N_4319);
or U7826 (N_7826,N_4522,N_5559);
xor U7827 (N_7827,N_5245,N_4844);
nand U7828 (N_7828,N_4277,N_5933);
nand U7829 (N_7829,N_4590,N_5541);
nor U7830 (N_7830,N_4179,N_5326);
and U7831 (N_7831,N_5504,N_5981);
nor U7832 (N_7832,N_4445,N_5634);
xnor U7833 (N_7833,N_5700,N_5740);
and U7834 (N_7834,N_5430,N_5288);
and U7835 (N_7835,N_5041,N_5726);
or U7836 (N_7836,N_4772,N_5595);
or U7837 (N_7837,N_4417,N_4982);
and U7838 (N_7838,N_4846,N_5740);
or U7839 (N_7839,N_5981,N_5589);
nand U7840 (N_7840,N_5629,N_5520);
nand U7841 (N_7841,N_4981,N_5642);
or U7842 (N_7842,N_4571,N_5875);
nand U7843 (N_7843,N_5801,N_4929);
nand U7844 (N_7844,N_5399,N_4265);
and U7845 (N_7845,N_5427,N_5514);
and U7846 (N_7846,N_5047,N_5064);
nand U7847 (N_7847,N_4763,N_5044);
nor U7848 (N_7848,N_5860,N_5423);
and U7849 (N_7849,N_4653,N_5442);
nor U7850 (N_7850,N_5575,N_5316);
and U7851 (N_7851,N_4585,N_5189);
or U7852 (N_7852,N_4659,N_5401);
nor U7853 (N_7853,N_5971,N_4990);
or U7854 (N_7854,N_4430,N_5608);
and U7855 (N_7855,N_5482,N_4921);
nor U7856 (N_7856,N_4652,N_4404);
or U7857 (N_7857,N_4700,N_4473);
or U7858 (N_7858,N_5942,N_4540);
xor U7859 (N_7859,N_4148,N_5167);
nand U7860 (N_7860,N_5090,N_4288);
or U7861 (N_7861,N_4099,N_4913);
or U7862 (N_7862,N_4285,N_4529);
nor U7863 (N_7863,N_5241,N_5267);
and U7864 (N_7864,N_4513,N_4976);
and U7865 (N_7865,N_5000,N_5090);
xnor U7866 (N_7866,N_4844,N_4454);
or U7867 (N_7867,N_5871,N_4948);
nor U7868 (N_7868,N_5379,N_5908);
and U7869 (N_7869,N_4630,N_5854);
xnor U7870 (N_7870,N_5983,N_4473);
or U7871 (N_7871,N_4589,N_4012);
nor U7872 (N_7872,N_4675,N_5128);
or U7873 (N_7873,N_4824,N_5048);
and U7874 (N_7874,N_4824,N_4057);
and U7875 (N_7875,N_4204,N_5302);
or U7876 (N_7876,N_4206,N_4895);
xor U7877 (N_7877,N_4097,N_5086);
nor U7878 (N_7878,N_5993,N_4607);
or U7879 (N_7879,N_4683,N_4443);
xor U7880 (N_7880,N_5986,N_4770);
nand U7881 (N_7881,N_4521,N_5827);
and U7882 (N_7882,N_5445,N_4483);
nand U7883 (N_7883,N_5173,N_5396);
and U7884 (N_7884,N_5982,N_5026);
nor U7885 (N_7885,N_5216,N_4663);
or U7886 (N_7886,N_4934,N_5740);
and U7887 (N_7887,N_4317,N_4912);
or U7888 (N_7888,N_5485,N_4092);
nand U7889 (N_7889,N_4151,N_5810);
or U7890 (N_7890,N_4014,N_5037);
nand U7891 (N_7891,N_4450,N_4736);
and U7892 (N_7892,N_4980,N_4644);
and U7893 (N_7893,N_5663,N_4580);
xnor U7894 (N_7894,N_5190,N_5600);
nand U7895 (N_7895,N_5142,N_5089);
xor U7896 (N_7896,N_5732,N_4240);
nand U7897 (N_7897,N_5108,N_4575);
nor U7898 (N_7898,N_4902,N_4499);
or U7899 (N_7899,N_4881,N_5270);
or U7900 (N_7900,N_5270,N_4805);
or U7901 (N_7901,N_5661,N_5241);
xor U7902 (N_7902,N_5635,N_4432);
nand U7903 (N_7903,N_4819,N_5241);
nand U7904 (N_7904,N_5145,N_4273);
nor U7905 (N_7905,N_4782,N_4245);
nor U7906 (N_7906,N_5163,N_5179);
nor U7907 (N_7907,N_5070,N_4647);
or U7908 (N_7908,N_5942,N_5910);
or U7909 (N_7909,N_5383,N_5217);
or U7910 (N_7910,N_4714,N_5202);
or U7911 (N_7911,N_4475,N_5874);
and U7912 (N_7912,N_4103,N_4547);
nand U7913 (N_7913,N_4910,N_5833);
nor U7914 (N_7914,N_4004,N_5743);
nor U7915 (N_7915,N_4576,N_5086);
nor U7916 (N_7916,N_5115,N_5228);
or U7917 (N_7917,N_5011,N_5012);
or U7918 (N_7918,N_4616,N_5160);
xnor U7919 (N_7919,N_4478,N_5047);
or U7920 (N_7920,N_5543,N_4112);
and U7921 (N_7921,N_5254,N_4982);
or U7922 (N_7922,N_5309,N_4776);
and U7923 (N_7923,N_4501,N_5772);
nor U7924 (N_7924,N_5205,N_4451);
and U7925 (N_7925,N_4191,N_4097);
and U7926 (N_7926,N_4871,N_4942);
or U7927 (N_7927,N_5307,N_5299);
xnor U7928 (N_7928,N_5744,N_4927);
or U7929 (N_7929,N_4614,N_5252);
nand U7930 (N_7930,N_5910,N_5008);
nand U7931 (N_7931,N_4125,N_5953);
nor U7932 (N_7932,N_4394,N_5288);
and U7933 (N_7933,N_5244,N_5086);
nor U7934 (N_7934,N_4060,N_5937);
and U7935 (N_7935,N_4819,N_4136);
nor U7936 (N_7936,N_4197,N_5941);
and U7937 (N_7937,N_5023,N_5327);
nand U7938 (N_7938,N_5286,N_4496);
xor U7939 (N_7939,N_5725,N_5918);
or U7940 (N_7940,N_5703,N_4515);
or U7941 (N_7941,N_5755,N_5355);
or U7942 (N_7942,N_5262,N_5981);
nor U7943 (N_7943,N_5832,N_5980);
or U7944 (N_7944,N_4518,N_5650);
nor U7945 (N_7945,N_5702,N_5260);
nor U7946 (N_7946,N_5240,N_5455);
nor U7947 (N_7947,N_5998,N_5140);
and U7948 (N_7948,N_5616,N_4564);
nor U7949 (N_7949,N_5570,N_5992);
nor U7950 (N_7950,N_5935,N_4642);
or U7951 (N_7951,N_4139,N_4350);
nor U7952 (N_7952,N_5154,N_4268);
or U7953 (N_7953,N_4913,N_4778);
and U7954 (N_7954,N_5807,N_4503);
nor U7955 (N_7955,N_4370,N_5947);
xor U7956 (N_7956,N_5410,N_5622);
or U7957 (N_7957,N_5438,N_4750);
and U7958 (N_7958,N_5306,N_5008);
and U7959 (N_7959,N_5706,N_4340);
nand U7960 (N_7960,N_5772,N_5618);
nand U7961 (N_7961,N_4368,N_5473);
nand U7962 (N_7962,N_5403,N_5828);
or U7963 (N_7963,N_5864,N_4000);
or U7964 (N_7964,N_4472,N_5939);
or U7965 (N_7965,N_4786,N_5157);
and U7966 (N_7966,N_5888,N_4021);
and U7967 (N_7967,N_5419,N_4099);
nand U7968 (N_7968,N_4462,N_4375);
nand U7969 (N_7969,N_4097,N_5717);
or U7970 (N_7970,N_5287,N_5324);
xnor U7971 (N_7971,N_4327,N_4998);
xnor U7972 (N_7972,N_4442,N_4046);
xor U7973 (N_7973,N_5762,N_5703);
xor U7974 (N_7974,N_5543,N_4810);
nor U7975 (N_7975,N_5454,N_4097);
nor U7976 (N_7976,N_4981,N_4972);
and U7977 (N_7977,N_4207,N_4597);
or U7978 (N_7978,N_4008,N_5775);
nor U7979 (N_7979,N_4919,N_5252);
or U7980 (N_7980,N_5522,N_4947);
xnor U7981 (N_7981,N_5811,N_4733);
and U7982 (N_7982,N_4869,N_4859);
nand U7983 (N_7983,N_4242,N_4018);
nor U7984 (N_7984,N_4161,N_5842);
nand U7985 (N_7985,N_4687,N_5322);
xor U7986 (N_7986,N_4033,N_5930);
nor U7987 (N_7987,N_5983,N_4316);
nor U7988 (N_7988,N_5071,N_5444);
xnor U7989 (N_7989,N_4119,N_5522);
nor U7990 (N_7990,N_4367,N_5856);
nor U7991 (N_7991,N_4449,N_5983);
nor U7992 (N_7992,N_4211,N_4662);
and U7993 (N_7993,N_4585,N_5010);
and U7994 (N_7994,N_5330,N_5176);
nand U7995 (N_7995,N_4725,N_4613);
nand U7996 (N_7996,N_4596,N_5220);
nor U7997 (N_7997,N_4487,N_5135);
nor U7998 (N_7998,N_5772,N_5003);
and U7999 (N_7999,N_4653,N_5976);
xnor U8000 (N_8000,N_6326,N_7706);
nor U8001 (N_8001,N_7637,N_6173);
and U8002 (N_8002,N_7369,N_6303);
and U8003 (N_8003,N_6993,N_7237);
and U8004 (N_8004,N_7378,N_6599);
or U8005 (N_8005,N_6987,N_6439);
nor U8006 (N_8006,N_6750,N_6094);
nor U8007 (N_8007,N_6804,N_6084);
or U8008 (N_8008,N_6645,N_6376);
or U8009 (N_8009,N_6584,N_7830);
nor U8010 (N_8010,N_6871,N_6478);
nand U8011 (N_8011,N_7261,N_6216);
nand U8012 (N_8012,N_7405,N_7433);
or U8013 (N_8013,N_6503,N_7112);
or U8014 (N_8014,N_6996,N_6110);
or U8015 (N_8015,N_6267,N_6149);
nand U8016 (N_8016,N_7781,N_6946);
nor U8017 (N_8017,N_6279,N_6921);
or U8018 (N_8018,N_6277,N_6894);
nor U8019 (N_8019,N_6081,N_6906);
and U8020 (N_8020,N_7589,N_7460);
xnor U8021 (N_8021,N_6964,N_7734);
nor U8022 (N_8022,N_7095,N_6095);
and U8023 (N_8023,N_6014,N_7495);
xnor U8024 (N_8024,N_6926,N_7654);
xnor U8025 (N_8025,N_6783,N_7332);
xor U8026 (N_8026,N_6065,N_6238);
or U8027 (N_8027,N_7659,N_7121);
and U8028 (N_8028,N_6268,N_6514);
and U8029 (N_8029,N_6815,N_6892);
nand U8030 (N_8030,N_7043,N_6357);
xnor U8031 (N_8031,N_7187,N_7923);
or U8032 (N_8032,N_7558,N_6969);
nor U8033 (N_8033,N_6465,N_6294);
or U8034 (N_8034,N_7240,N_7918);
nor U8035 (N_8035,N_6600,N_6394);
nand U8036 (N_8036,N_7407,N_6811);
and U8037 (N_8037,N_6832,N_7638);
and U8038 (N_8038,N_6312,N_6248);
nand U8039 (N_8039,N_7166,N_7126);
and U8040 (N_8040,N_6835,N_7562);
nand U8041 (N_8041,N_6104,N_7373);
or U8042 (N_8042,N_6087,N_7245);
nand U8043 (N_8043,N_7531,N_6624);
nor U8044 (N_8044,N_7530,N_7356);
and U8045 (N_8045,N_7278,N_6893);
nor U8046 (N_8046,N_7564,N_6126);
xnor U8047 (N_8047,N_6122,N_6611);
nor U8048 (N_8048,N_7211,N_7521);
and U8049 (N_8049,N_6269,N_6009);
nor U8050 (N_8050,N_6435,N_7117);
nand U8051 (N_8051,N_6642,N_6912);
xnor U8052 (N_8052,N_6175,N_6239);
xnor U8053 (N_8053,N_7809,N_7444);
or U8054 (N_8054,N_6879,N_7581);
nand U8055 (N_8055,N_6025,N_6449);
nor U8056 (N_8056,N_7525,N_7340);
nor U8057 (N_8057,N_7168,N_6531);
xnor U8058 (N_8058,N_6548,N_7817);
nor U8059 (N_8059,N_7475,N_6870);
and U8060 (N_8060,N_7945,N_7891);
or U8061 (N_8061,N_7616,N_6627);
and U8062 (N_8062,N_6516,N_6457);
nor U8063 (N_8063,N_6693,N_6618);
or U8064 (N_8064,N_7459,N_6299);
nor U8065 (N_8065,N_6050,N_7160);
or U8066 (N_8066,N_7671,N_7762);
and U8067 (N_8067,N_6905,N_7238);
nor U8068 (N_8068,N_7142,N_7758);
or U8069 (N_8069,N_7973,N_6709);
xor U8070 (N_8070,N_7551,N_7700);
xnor U8071 (N_8071,N_6231,N_6535);
nand U8072 (N_8072,N_7191,N_7688);
and U8073 (N_8073,N_6150,N_6307);
nand U8074 (N_8074,N_7596,N_6393);
nor U8075 (N_8075,N_7962,N_6994);
xnor U8076 (N_8076,N_7389,N_6582);
nor U8077 (N_8077,N_7143,N_6913);
nor U8078 (N_8078,N_7736,N_7929);
nand U8079 (N_8079,N_7946,N_7508);
and U8080 (N_8080,N_7928,N_6495);
nor U8081 (N_8081,N_7546,N_6569);
and U8082 (N_8082,N_7726,N_6375);
nor U8083 (N_8083,N_7588,N_7539);
nand U8084 (N_8084,N_6447,N_7036);
nand U8085 (N_8085,N_6286,N_7430);
or U8086 (N_8086,N_7978,N_6614);
nand U8087 (N_8087,N_6358,N_6740);
and U8088 (N_8088,N_7154,N_6550);
or U8089 (N_8089,N_6469,N_7339);
or U8090 (N_8090,N_6718,N_7425);
nor U8091 (N_8091,N_7372,N_6021);
and U8092 (N_8092,N_7090,N_7974);
xnor U8093 (N_8093,N_7631,N_7364);
nor U8094 (N_8094,N_7451,N_6814);
or U8095 (N_8095,N_7257,N_6933);
nor U8096 (N_8096,N_6170,N_7391);
xor U8097 (N_8097,N_7100,N_7896);
nand U8098 (N_8098,N_6383,N_6800);
nor U8099 (N_8099,N_6732,N_7084);
nand U8100 (N_8100,N_7570,N_6491);
and U8101 (N_8101,N_7766,N_6107);
or U8102 (N_8102,N_6643,N_7741);
nor U8103 (N_8103,N_7560,N_6117);
nor U8104 (N_8104,N_6264,N_6978);
and U8105 (N_8105,N_6766,N_7657);
or U8106 (N_8106,N_7432,N_7975);
and U8107 (N_8107,N_6324,N_6436);
xor U8108 (N_8108,N_6445,N_6572);
xor U8109 (N_8109,N_7383,N_6951);
or U8110 (N_8110,N_7109,N_6806);
or U8111 (N_8111,N_6733,N_6121);
xor U8112 (N_8112,N_7162,N_6197);
or U8113 (N_8113,N_7698,N_7574);
xnor U8114 (N_8114,N_7010,N_6039);
nor U8115 (N_8115,N_7880,N_6075);
xnor U8116 (N_8116,N_6045,N_7579);
xor U8117 (N_8117,N_7445,N_7336);
nor U8118 (N_8118,N_6590,N_7963);
xnor U8119 (N_8119,N_7704,N_6213);
nor U8120 (N_8120,N_6844,N_7927);
or U8121 (N_8121,N_6164,N_7256);
xor U8122 (N_8122,N_6467,N_7371);
and U8123 (N_8123,N_6658,N_7153);
and U8124 (N_8124,N_6347,N_7346);
or U8125 (N_8125,N_6650,N_6079);
nand U8126 (N_8126,N_6966,N_7384);
or U8127 (N_8127,N_6024,N_6880);
nor U8128 (N_8128,N_7501,N_7158);
and U8129 (N_8129,N_6678,N_6096);
nand U8130 (N_8130,N_7934,N_6974);
xnor U8131 (N_8131,N_7966,N_7634);
nand U8132 (N_8132,N_7865,N_6027);
or U8133 (N_8133,N_7878,N_7790);
and U8134 (N_8134,N_6369,N_7715);
xnor U8135 (N_8135,N_7752,N_6952);
xor U8136 (N_8136,N_7620,N_7832);
or U8137 (N_8137,N_6040,N_7777);
nor U8138 (N_8138,N_7116,N_6301);
nor U8139 (N_8139,N_6723,N_6308);
nor U8140 (N_8140,N_6348,N_6203);
and U8141 (N_8141,N_7795,N_6147);
and U8142 (N_8142,N_7494,N_7788);
nand U8143 (N_8143,N_6717,N_7628);
or U8144 (N_8144,N_7210,N_6266);
and U8145 (N_8145,N_6072,N_6300);
xnor U8146 (N_8146,N_7070,N_7682);
nand U8147 (N_8147,N_7047,N_7661);
and U8148 (N_8148,N_6230,N_6706);
or U8149 (N_8149,N_7718,N_6061);
and U8150 (N_8150,N_7823,N_7839);
nand U8151 (N_8151,N_6249,N_6132);
nand U8152 (N_8152,N_7677,N_7075);
and U8153 (N_8153,N_6604,N_7587);
nor U8154 (N_8154,N_7511,N_7106);
nor U8155 (N_8155,N_7155,N_6633);
xor U8156 (N_8156,N_6275,N_6411);
xor U8157 (N_8157,N_7484,N_6533);
xnor U8158 (N_8158,N_7398,N_7426);
and U8159 (N_8159,N_6346,N_6448);
xor U8160 (N_8160,N_6846,N_6172);
nand U8161 (N_8161,N_6975,N_7710);
nor U8162 (N_8162,N_6217,N_7349);
xnor U8163 (N_8163,N_7246,N_6959);
or U8164 (N_8164,N_6787,N_6354);
and U8165 (N_8165,N_6875,N_7198);
xor U8166 (N_8166,N_7608,N_6339);
and U8167 (N_8167,N_6296,N_6404);
nor U8168 (N_8168,N_6454,N_7916);
nor U8169 (N_8169,N_7201,N_7768);
or U8170 (N_8170,N_7548,N_6373);
nand U8171 (N_8171,N_7183,N_6059);
or U8172 (N_8172,N_6685,N_7129);
xnor U8173 (N_8173,N_7933,N_7497);
nand U8174 (N_8174,N_6505,N_7785);
nand U8175 (N_8175,N_6444,N_7092);
and U8176 (N_8176,N_6847,N_7130);
xor U8177 (N_8177,N_6125,N_7816);
nand U8178 (N_8178,N_7236,N_7749);
xor U8179 (N_8179,N_6158,N_7134);
xor U8180 (N_8180,N_6588,N_6360);
or U8181 (N_8181,N_7877,N_6561);
nor U8182 (N_8182,N_6335,N_6100);
or U8183 (N_8183,N_6939,N_7406);
xor U8184 (N_8184,N_7217,N_6000);
and U8185 (N_8185,N_7771,N_6032);
nor U8186 (N_8186,N_6749,N_7863);
or U8187 (N_8187,N_6223,N_6257);
and U8188 (N_8188,N_7561,N_7469);
xor U8189 (N_8189,N_7655,N_7012);
nand U8190 (N_8190,N_6981,N_6547);
or U8191 (N_8191,N_6226,N_7003);
and U8192 (N_8192,N_7317,N_6509);
nor U8193 (N_8193,N_6649,N_6963);
and U8194 (N_8194,N_6641,N_7723);
or U8195 (N_8195,N_6234,N_6953);
or U8196 (N_8196,N_7556,N_7533);
or U8197 (N_8197,N_6005,N_6728);
xnor U8198 (N_8198,N_7983,N_6976);
or U8199 (N_8199,N_7305,N_6161);
and U8200 (N_8200,N_6507,N_6625);
or U8201 (N_8201,N_7189,N_7408);
nor U8202 (N_8202,N_6169,N_7778);
xnor U8203 (N_8203,N_6992,N_6011);
xnor U8204 (N_8204,N_6432,N_6295);
nor U8205 (N_8205,N_7977,N_7837);
and U8206 (N_8206,N_6263,N_7997);
or U8207 (N_8207,N_6779,N_6070);
or U8208 (N_8208,N_6304,N_6035);
nand U8209 (N_8209,N_6013,N_7428);
xnor U8210 (N_8210,N_7157,N_6560);
nor U8211 (N_8211,N_6873,N_6754);
and U8212 (N_8212,N_6413,N_6674);
nor U8213 (N_8213,N_7541,N_6519);
and U8214 (N_8214,N_7363,N_6058);
xor U8215 (N_8215,N_7024,N_6669);
and U8216 (N_8216,N_7271,N_6431);
nor U8217 (N_8217,N_7798,N_6481);
or U8218 (N_8218,N_7602,N_6757);
and U8219 (N_8219,N_6017,N_6640);
nor U8220 (N_8220,N_6379,N_7585);
or U8221 (N_8221,N_6475,N_6057);
xor U8222 (N_8222,N_6251,N_7080);
nand U8223 (N_8223,N_6416,N_7442);
and U8224 (N_8224,N_7825,N_6468);
xor U8225 (N_8225,N_7820,N_7632);
and U8226 (N_8226,N_7215,N_6386);
or U8227 (N_8227,N_7779,N_7503);
or U8228 (N_8228,N_7903,N_6452);
nor U8229 (N_8229,N_6099,N_6644);
or U8230 (N_8230,N_6528,N_7286);
and U8231 (N_8231,N_7213,N_6512);
nor U8232 (N_8232,N_6314,N_6559);
or U8233 (N_8233,N_7491,N_6850);
or U8234 (N_8234,N_6524,N_7293);
xor U8235 (N_8235,N_6105,N_7870);
nand U8236 (N_8236,N_7591,N_6372);
or U8237 (N_8237,N_6967,N_6711);
xor U8238 (N_8238,N_6704,N_6868);
or U8239 (N_8239,N_7619,N_7493);
nor U8240 (N_8240,N_7132,N_7476);
xnor U8241 (N_8241,N_7642,N_7601);
or U8242 (N_8242,N_6623,N_7526);
and U8243 (N_8243,N_7550,N_7102);
or U8244 (N_8244,N_7474,N_7611);
or U8245 (N_8245,N_6920,N_6710);
nand U8246 (N_8246,N_7329,N_7834);
xor U8247 (N_8247,N_6763,N_7051);
nand U8248 (N_8248,N_7625,N_6282);
or U8249 (N_8249,N_7592,N_7641);
and U8250 (N_8250,N_6546,N_6602);
and U8251 (N_8251,N_6159,N_6558);
and U8252 (N_8252,N_6720,N_7269);
nor U8253 (N_8253,N_7976,N_6288);
nor U8254 (N_8254,N_6729,N_6043);
or U8255 (N_8255,N_7829,N_7985);
or U8256 (N_8256,N_7480,N_6830);
nand U8257 (N_8257,N_6490,N_7139);
xor U8258 (N_8258,N_7279,N_6679);
or U8259 (N_8259,N_7453,N_6731);
and U8260 (N_8260,N_6818,N_7717);
xor U8261 (N_8261,N_6581,N_6714);
nand U8262 (N_8262,N_7085,N_6302);
and U8263 (N_8263,N_6826,N_7855);
nand U8264 (N_8264,N_6440,N_7145);
nor U8265 (N_8265,N_6422,N_6198);
or U8266 (N_8266,N_6453,N_6362);
nor U8267 (N_8267,N_7686,N_6055);
and U8268 (N_8268,N_7652,N_7354);
nand U8269 (N_8269,N_7909,N_7913);
nor U8270 (N_8270,N_6318,N_7969);
xor U8271 (N_8271,N_6607,N_6908);
xor U8272 (N_8272,N_6423,N_6367);
xor U8273 (N_8273,N_6770,N_7604);
nand U8274 (N_8274,N_6427,N_7427);
and U8275 (N_8275,N_7422,N_6135);
or U8276 (N_8276,N_7454,N_6193);
xor U8277 (N_8277,N_7052,N_7643);
nor U8278 (N_8278,N_7614,N_6773);
xor U8279 (N_8279,N_6137,N_6333);
and U8280 (N_8280,N_7041,N_6552);
and U8281 (N_8281,N_6789,N_7538);
xnor U8282 (N_8282,N_7315,N_6020);
nor U8283 (N_8283,N_7335,N_7420);
nand U8284 (N_8284,N_7489,N_6986);
or U8285 (N_8285,N_7379,N_6486);
nor U8286 (N_8286,N_7535,N_7889);
or U8287 (N_8287,N_7603,N_6661);
nand U8288 (N_8288,N_7290,N_7818);
nand U8289 (N_8289,N_6355,N_7300);
nor U8290 (N_8290,N_6224,N_7712);
xor U8291 (N_8291,N_6580,N_7044);
xor U8292 (N_8292,N_6605,N_6716);
xor U8293 (N_8293,N_7529,N_6639);
nand U8294 (N_8294,N_6368,N_7801);
nor U8295 (N_8295,N_6612,N_6666);
and U8296 (N_8296,N_7847,N_6016);
and U8297 (N_8297,N_7284,N_7852);
nor U8298 (N_8298,N_7496,N_6562);
or U8299 (N_8299,N_7872,N_7038);
or U8300 (N_8300,N_6931,N_7831);
or U8301 (N_8301,N_6918,N_6810);
and U8302 (N_8302,N_6023,N_7568);
and U8303 (N_8303,N_7076,N_7610);
and U8304 (N_8304,N_7727,N_7720);
xor U8305 (N_8305,N_6450,N_7824);
xor U8306 (N_8306,N_6289,N_6211);
or U8307 (N_8307,N_6089,N_7639);
nor U8308 (N_8308,N_6219,N_6077);
and U8309 (N_8309,N_7517,N_7234);
and U8310 (N_8310,N_7308,N_6442);
xor U8311 (N_8311,N_7876,N_7273);
nor U8312 (N_8312,N_7707,N_7202);
nor U8313 (N_8313,N_7396,N_7296);
xnor U8314 (N_8314,N_6510,N_6881);
nand U8315 (N_8315,N_6885,N_6929);
xor U8316 (N_8316,N_6593,N_6796);
nor U8317 (N_8317,N_7840,N_7507);
or U8318 (N_8318,N_6460,N_7998);
nand U8319 (N_8319,N_7243,N_7512);
and U8320 (N_8320,N_6668,N_7288);
and U8321 (N_8321,N_6807,N_7902);
nand U8322 (N_8322,N_6954,N_6555);
or U8323 (N_8323,N_7421,N_6759);
and U8324 (N_8324,N_7252,N_6934);
or U8325 (N_8325,N_7066,N_7714);
xor U8326 (N_8326,N_6220,N_7506);
nand U8327 (N_8327,N_7074,N_7833);
and U8328 (N_8328,N_6406,N_7443);
xor U8329 (N_8329,N_6725,N_7310);
nor U8330 (N_8330,N_7282,N_6340);
nand U8331 (N_8331,N_7730,N_7846);
xor U8332 (N_8332,N_7287,N_6909);
or U8333 (N_8333,N_7452,N_6565);
and U8334 (N_8334,N_7808,N_6425);
and U8335 (N_8335,N_7472,N_7586);
or U8336 (N_8336,N_6973,N_6616);
nor U8337 (N_8337,N_7146,N_6012);
and U8338 (N_8338,N_7776,N_6665);
xor U8339 (N_8339,N_6492,N_7487);
nor U8340 (N_8340,N_7223,N_6938);
or U8341 (N_8341,N_6060,N_7393);
nor U8342 (N_8342,N_6708,N_6280);
nand U8343 (N_8343,N_6374,N_7285);
or U8344 (N_8344,N_7239,N_7578);
and U8345 (N_8345,N_7093,N_6594);
or U8346 (N_8346,N_6222,N_7448);
xor U8347 (N_8347,N_6200,N_7225);
xnor U8348 (N_8348,N_6752,N_6941);
or U8349 (N_8349,N_7761,N_7137);
xnor U8350 (N_8350,N_7268,N_7792);
or U8351 (N_8351,N_6511,N_6388);
nor U8352 (N_8352,N_6417,N_7705);
nand U8353 (N_8353,N_6071,N_7662);
and U8354 (N_8354,N_7400,N_6656);
xor U8355 (N_8355,N_7681,N_6194);
or U8356 (N_8356,N_7952,N_7697);
or U8357 (N_8357,N_6746,N_7437);
nor U8358 (N_8358,N_7226,N_7206);
and U8359 (N_8359,N_7322,N_7381);
nor U8360 (N_8360,N_7193,N_6738);
xnor U8361 (N_8361,N_7783,N_7458);
and U8362 (N_8362,N_7415,N_6136);
and U8363 (N_8363,N_6364,N_7649);
and U8364 (N_8364,N_7735,N_7324);
nor U8365 (N_8365,N_7149,N_7993);
or U8366 (N_8366,N_6430,N_6745);
and U8367 (N_8367,N_7250,N_7552);
and U8368 (N_8368,N_7251,N_7810);
nor U8369 (N_8369,N_7575,N_6142);
nand U8370 (N_8370,N_6860,N_7684);
or U8371 (N_8371,N_7862,N_6769);
and U8372 (N_8372,N_7382,N_7742);
and U8373 (N_8373,N_6699,N_7351);
or U8374 (N_8374,N_6936,N_7786);
nor U8375 (N_8375,N_6278,N_6391);
and U8376 (N_8376,N_7576,N_6813);
or U8377 (N_8377,N_7151,N_7377);
nand U8378 (N_8378,N_7937,N_7418);
or U8379 (N_8379,N_6925,N_6958);
and U8380 (N_8380,N_6112,N_7685);
nor U8381 (N_8381,N_6972,N_6483);
xor U8382 (N_8382,N_7848,N_7417);
nor U8383 (N_8383,N_7680,N_6859);
and U8384 (N_8384,N_7150,N_6659);
and U8385 (N_8385,N_7035,N_7164);
nand U8386 (N_8386,N_7230,N_6521);
nand U8387 (N_8387,N_7607,N_6701);
nand U8388 (N_8388,N_6428,N_7163);
or U8389 (N_8389,N_7949,N_6323);
or U8390 (N_8390,N_6525,N_7402);
nor U8391 (N_8391,N_6983,N_7873);
or U8392 (N_8392,N_6522,N_7253);
xnor U8393 (N_8393,N_7866,N_6284);
nand U8394 (N_8394,N_6188,N_7037);
and U8395 (N_8395,N_6420,N_6466);
nor U8396 (N_8396,N_6237,N_6534);
nand U8397 (N_8397,N_7013,N_6629);
nand U8398 (N_8398,N_7486,N_7544);
nor U8399 (N_8399,N_6210,N_7964);
nand U8400 (N_8400,N_6207,N_6088);
nand U8401 (N_8401,N_6638,N_7921);
nor U8402 (N_8402,N_7875,N_6177);
and U8403 (N_8403,N_6019,N_6233);
and U8404 (N_8404,N_7200,N_6456);
or U8405 (N_8405,N_7483,N_7110);
nand U8406 (N_8406,N_7366,N_6948);
nor U8407 (N_8407,N_7636,N_7724);
nand U8408 (N_8408,N_7212,N_6195);
or U8409 (N_8409,N_7623,N_7283);
nand U8410 (N_8410,N_7951,N_7789);
or U8411 (N_8411,N_7753,N_7327);
nor U8412 (N_8412,N_7303,N_6046);
xor U8413 (N_8413,N_6113,N_6006);
xnor U8414 (N_8414,N_7731,N_6031);
nor U8415 (N_8415,N_6116,N_6760);
xor U8416 (N_8416,N_7879,N_6493);
and U8417 (N_8417,N_6585,N_7728);
nand U8418 (N_8418,N_7537,N_6683);
nor U8419 (N_8419,N_7748,N_7466);
and U8420 (N_8420,N_7196,N_7708);
or U8421 (N_8421,N_6834,N_6349);
or U8422 (N_8422,N_6256,N_6128);
xor U8423 (N_8423,N_7729,N_6979);
xnor U8424 (N_8424,N_7693,N_7656);
nor U8425 (N_8425,N_6971,N_6345);
nor U8426 (N_8426,N_6473,N_6803);
or U8427 (N_8427,N_6310,N_6897);
nand U8428 (N_8428,N_6008,N_7254);
or U8429 (N_8429,N_7672,N_7849);
or U8430 (N_8430,N_6053,N_6227);
nor U8431 (N_8431,N_7970,N_6438);
or U8432 (N_8432,N_7111,N_7416);
nand U8433 (N_8433,N_7029,N_7185);
and U8434 (N_8434,N_6353,N_7065);
nor U8435 (N_8435,N_6655,N_7812);
or U8436 (N_8436,N_6022,N_6378);
nand U8437 (N_8437,N_6778,N_6464);
and U8438 (N_8438,N_6397,N_7881);
nand U8439 (N_8439,N_7021,N_6380);
or U8440 (N_8440,N_7940,N_6703);
xor U8441 (N_8441,N_7965,N_7169);
nand U8442 (N_8442,N_7375,N_6229);
or U8443 (N_8443,N_6287,N_6341);
xnor U8444 (N_8444,N_7314,N_6596);
xnor U8445 (N_8445,N_7005,N_6790);
or U8446 (N_8446,N_6543,N_7249);
xnor U8447 (N_8447,N_6532,N_7468);
or U8448 (N_8448,N_7397,N_6474);
nor U8449 (N_8449,N_7667,N_7802);
or U8450 (N_8450,N_6856,N_6033);
nand U8451 (N_8451,N_7606,N_6823);
nor U8452 (N_8452,N_7431,N_7301);
nand U8453 (N_8453,N_6777,N_7441);
nor U8454 (N_8454,N_7456,N_7058);
or U8455 (N_8455,N_6184,N_6316);
or U8456 (N_8456,N_7376,N_6108);
nor U8457 (N_8457,N_6123,N_7205);
or U8458 (N_8458,N_7784,N_7757);
xor U8459 (N_8459,N_7302,N_6141);
and U8460 (N_8460,N_7888,N_7194);
xor U8461 (N_8461,N_7695,N_6129);
xor U8462 (N_8462,N_6657,N_7323);
xor U8463 (N_8463,N_7887,N_6739);
xor U8464 (N_8464,N_6178,N_6900);
and U8465 (N_8465,N_7743,N_7097);
nor U8466 (N_8466,N_6462,N_6118);
and U8467 (N_8467,N_7853,N_6407);
or U8468 (N_8468,N_7241,N_7759);
and U8469 (N_8469,N_6103,N_6851);
nand U8470 (N_8470,N_6878,N_6148);
nor U8471 (N_8471,N_7915,N_6477);
or U8472 (N_8472,N_6250,N_6459);
xnor U8473 (N_8473,N_6101,N_7519);
xor U8474 (N_8474,N_6822,N_7115);
and U8475 (N_8475,N_7411,N_6245);
nor U8476 (N_8476,N_6898,N_7954);
xnor U8477 (N_8477,N_7813,N_7390);
and U8478 (N_8478,N_7644,N_6001);
xor U8479 (N_8479,N_7227,N_7401);
nand U8480 (N_8480,N_6564,N_6888);
xnor U8481 (N_8481,N_7509,N_6330);
nor U8482 (N_8482,N_6361,N_7072);
nand U8483 (N_8483,N_6338,N_6566);
nand U8484 (N_8484,N_7125,N_7214);
and U8485 (N_8485,N_6630,N_6887);
or U8486 (N_8486,N_6365,N_6410);
or U8487 (N_8487,N_7958,N_7858);
nand U8488 (N_8488,N_7819,N_6619);
nand U8489 (N_8489,N_6646,N_6608);
nand U8490 (N_8490,N_7515,N_6651);
nor U8491 (N_8491,N_6907,N_6412);
nor U8492 (N_8492,N_7077,N_7844);
nand U8493 (N_8493,N_7091,N_7127);
and U8494 (N_8494,N_6753,N_6409);
nor U8495 (N_8495,N_6156,N_7199);
nor U8496 (N_8496,N_6496,N_7144);
nand U8497 (N_8497,N_6556,N_6864);
xnor U8498 (N_8498,N_7796,N_7510);
and U8499 (N_8499,N_6575,N_7646);
or U8500 (N_8500,N_7733,N_7086);
and U8501 (N_8501,N_7008,N_6927);
nor U8502 (N_8502,N_7955,N_6311);
nor U8503 (N_8503,N_6852,N_6190);
nor U8504 (N_8504,N_7716,N_7195);
and U8505 (N_8505,N_6741,N_7939);
nand U8506 (N_8506,N_7457,N_6849);
nor U8507 (N_8507,N_7703,N_6389);
xnor U8508 (N_8508,N_6883,N_7593);
and U8509 (N_8509,N_7598,N_7104);
and U8510 (N_8510,N_7713,N_6697);
nand U8511 (N_8511,N_6691,N_6451);
and U8512 (N_8512,N_7087,N_6950);
nand U8513 (N_8513,N_6111,N_7083);
xnor U8514 (N_8514,N_7488,N_6861);
nand U8515 (N_8515,N_7756,N_6313);
and U8516 (N_8516,N_7886,N_7263);
or U8517 (N_8517,N_6426,N_6841);
xor U8518 (N_8518,N_7412,N_7176);
or U8519 (N_8519,N_6446,N_7281);
or U8520 (N_8520,N_6082,N_6209);
nand U8521 (N_8521,N_6098,N_7764);
xor U8522 (N_8522,N_7449,N_6695);
xor U8523 (N_8523,N_6742,N_6513);
nor U8524 (N_8524,N_6673,N_6429);
or U8525 (N_8525,N_7919,N_7299);
or U8526 (N_8526,N_7136,N_6337);
or U8527 (N_8527,N_6501,N_6315);
and U8528 (N_8528,N_7774,N_7922);
and U8529 (N_8529,N_7666,N_6085);
or U8530 (N_8530,N_7871,N_7828);
nor U8531 (N_8531,N_7676,N_6387);
or U8532 (N_8532,N_7499,N_6677);
or U8533 (N_8533,N_6688,N_6797);
nor U8534 (N_8534,N_6327,N_6336);
xnor U8535 (N_8535,N_7306,N_6727);
and U8536 (N_8536,N_6003,N_6309);
nand U8537 (N_8537,N_6545,N_7920);
and U8538 (N_8538,N_6480,N_7479);
nand U8539 (N_8539,N_6636,N_6956);
or U8540 (N_8540,N_7309,N_7181);
or U8541 (N_8541,N_6418,N_6942);
nand U8542 (N_8542,N_7229,N_7118);
xor U8543 (N_8543,N_6597,N_7197);
xor U8544 (N_8544,N_7350,N_7590);
or U8545 (N_8545,N_6332,N_6181);
and U8546 (N_8546,N_7258,N_6798);
nor U8547 (N_8547,N_7333,N_6370);
nand U8548 (N_8548,N_7900,N_6405);
or U8549 (N_8549,N_7244,N_6403);
and U8550 (N_8550,N_7640,N_7259);
or U8551 (N_8551,N_7014,N_6603);
or U8552 (N_8552,N_7843,N_7532);
or U8553 (N_8553,N_7167,N_6499);
nand U8554 (N_8554,N_6080,N_6498);
nor U8555 (N_8555,N_6592,N_6102);
and U8556 (N_8556,N_6083,N_7152);
nand U8557 (N_8557,N_6615,N_7270);
xor U8558 (N_8558,N_6421,N_7057);
or U8559 (N_8559,N_7056,N_6890);
xor U8560 (N_8560,N_7359,N_7780);
nor U8561 (N_8561,N_6097,N_6036);
and U8562 (N_8562,N_7424,N_6788);
and U8563 (N_8563,N_7557,N_7721);
xnor U8564 (N_8564,N_6682,N_6034);
nand U8565 (N_8565,N_7122,N_6781);
and U8566 (N_8566,N_7663,N_6153);
nand U8567 (N_8567,N_7814,N_7912);
nand U8568 (N_8568,N_6281,N_6274);
nor U8569 (N_8569,N_6488,N_7019);
and U8570 (N_8570,N_6221,N_7826);
xnor U8571 (N_8571,N_6342,N_6702);
nor U8572 (N_8572,N_7318,N_7787);
xnor U8573 (N_8573,N_6772,N_6689);
nand U8574 (N_8574,N_6915,N_7648);
and U8575 (N_8575,N_6943,N_6204);
and U8576 (N_8576,N_7140,N_7320);
nor U8577 (N_8577,N_6601,N_7725);
nand U8578 (N_8578,N_7337,N_7203);
and U8579 (N_8579,N_6744,N_6479);
or U8580 (N_8580,N_6254,N_6960);
and U8581 (N_8581,N_6127,N_6845);
xor U8582 (N_8582,N_6007,N_7615);
nor U8583 (N_8583,N_6041,N_7280);
or U8584 (N_8584,N_6049,N_7536);
and U8585 (N_8585,N_7547,N_6829);
nor U8586 (N_8586,N_6352,N_7836);
nand U8587 (N_8587,N_6586,N_6433);
nor U8588 (N_8588,N_7683,N_7274);
and U8589 (N_8589,N_7992,N_7159);
xnor U8590 (N_8590,N_6395,N_7999);
or U8591 (N_8591,N_6494,N_7719);
nor U8592 (N_8592,N_6577,N_6359);
nand U8593 (N_8593,N_6351,N_6696);
xnor U8594 (N_8594,N_7932,N_7018);
or U8595 (N_8595,N_7367,N_6520);
xnor U8596 (N_8596,N_7180,N_7298);
xor U8597 (N_8597,N_6652,N_7775);
nand U8598 (N_8598,N_6808,N_7867);
or U8599 (N_8599,N_6817,N_7885);
nor U8600 (N_8600,N_6537,N_6476);
nand U8601 (N_8601,N_6205,N_6109);
nand U8602 (N_8602,N_7027,N_7219);
nand U8603 (N_8603,N_7312,N_6761);
nor U8604 (N_8604,N_6306,N_6131);
nor U8605 (N_8605,N_6206,N_6133);
nand U8606 (N_8606,N_7062,N_6648);
nand U8607 (N_8607,N_7000,N_7352);
nand U8608 (N_8608,N_7803,N_6401);
and U8609 (N_8609,N_6399,N_7368);
nor U8610 (N_8610,N_7358,N_7645);
or U8611 (N_8611,N_7291,N_6276);
nor U8612 (N_8612,N_6854,N_6518);
and U8613 (N_8613,N_6795,N_6026);
xnor U8614 (N_8614,N_7711,N_6877);
and U8615 (N_8615,N_7388,N_6270);
or U8616 (N_8616,N_6707,N_7904);
nand U8617 (N_8617,N_6232,N_7242);
and U8618 (N_8618,N_6824,N_7103);
nand U8619 (N_8619,N_6208,N_6199);
xnor U8620 (N_8620,N_7004,N_7738);
and U8621 (N_8621,N_7692,N_7069);
nor U8622 (N_8622,N_6086,N_6134);
nor U8623 (N_8623,N_6144,N_7914);
or U8624 (N_8624,N_7569,N_6356);
and U8625 (N_8625,N_7988,N_6736);
nor U8626 (N_8626,N_6246,N_6068);
nand U8627 (N_8627,N_7326,N_7319);
xor U8628 (N_8628,N_7386,N_6064);
nand U8629 (N_8629,N_6325,N_6628);
nand U8630 (N_8630,N_7811,N_6320);
or U8631 (N_8631,N_7022,N_7248);
xnor U8632 (N_8632,N_6485,N_6917);
or U8633 (N_8633,N_7138,N_6140);
nand U8634 (N_8634,N_7334,N_6821);
and U8635 (N_8635,N_6635,N_7861);
nor U8636 (N_8636,N_6980,N_6255);
or U8637 (N_8637,N_6637,N_6840);
nor U8638 (N_8638,N_7357,N_6955);
xor U8639 (N_8639,N_6843,N_7582);
nor U8640 (N_8640,N_7330,N_7821);
nand U8641 (N_8641,N_7073,N_6730);
and U8642 (N_8642,N_6998,N_7567);
nor U8643 (N_8643,N_7980,N_7907);
and U8644 (N_8644,N_6671,N_7015);
or U8645 (N_8645,N_6321,N_7668);
nand U8646 (N_8646,N_6319,N_7629);
and U8647 (N_8647,N_7114,N_7679);
nor U8648 (N_8648,N_6236,N_7895);
nand U8649 (N_8649,N_6201,N_6434);
and U8650 (N_8650,N_7842,N_6037);
and U8651 (N_8651,N_6765,N_6526);
and U8652 (N_8652,N_7020,N_7622);
nor U8653 (N_8653,N_6889,N_7765);
nor U8654 (N_8654,N_7996,N_7857);
or U8655 (N_8655,N_7805,N_7128);
xnor U8656 (N_8656,N_7972,N_7751);
nand U8657 (N_8657,N_7950,N_7986);
xor U8658 (N_8658,N_7647,N_7722);
nor U8659 (N_8659,N_6273,N_7032);
and U8660 (N_8660,N_7135,N_7942);
nand U8661 (N_8661,N_6831,N_6051);
and U8662 (N_8662,N_6692,N_7423);
xor U8663 (N_8663,N_7017,N_6816);
nor U8664 (N_8664,N_7247,N_6298);
nand U8665 (N_8665,N_6911,N_7696);
xor U8666 (N_8666,N_7635,N_7665);
and U8667 (N_8667,N_6945,N_6271);
and U8668 (N_8668,N_7583,N_6940);
nor U8669 (N_8669,N_6441,N_6331);
or U8670 (N_8670,N_6872,N_7209);
xnor U8671 (N_8671,N_6775,N_7874);
and U8672 (N_8672,N_7040,N_6502);
xor U8673 (N_8673,N_7770,N_7053);
nor U8674 (N_8674,N_6544,N_7864);
or U8675 (N_8675,N_6241,N_7860);
and U8676 (N_8676,N_7462,N_6780);
xnor U8677 (N_8677,N_7026,N_7991);
or U8678 (N_8678,N_7216,N_6672);
or U8679 (N_8679,N_7794,N_7182);
nor U8680 (N_8680,N_7113,N_6853);
xnor U8681 (N_8681,N_6554,N_7222);
nor U8682 (N_8682,N_7316,N_7011);
or U8683 (N_8683,N_7098,N_6764);
or U8684 (N_8684,N_6151,N_7470);
or U8685 (N_8685,N_6583,N_7935);
nand U8686 (N_8686,N_6317,N_6139);
and U8687 (N_8687,N_6857,N_6253);
or U8688 (N_8688,N_6768,N_7289);
xor U8689 (N_8689,N_7571,N_6214);
nand U8690 (N_8690,N_7908,N_7094);
nand U8691 (N_8691,N_6799,N_7906);
nand U8692 (N_8692,N_7627,N_7901);
xnor U8693 (N_8693,N_6377,N_7260);
nand U8694 (N_8694,N_7835,N_6793);
and U8695 (N_8695,N_6812,N_6961);
nor U8696 (N_8696,N_7573,N_7440);
and U8697 (N_8697,N_7502,N_7370);
or U8698 (N_8698,N_7362,N_6977);
nor U8699 (N_8699,N_6028,N_6919);
or U8700 (N_8700,N_6858,N_6063);
nand U8701 (N_8701,N_6984,N_7699);
nor U8702 (N_8702,N_6568,N_7409);
xor U8703 (N_8703,N_6621,N_7119);
and U8704 (N_8704,N_7687,N_7984);
nand U8705 (N_8705,N_6078,N_6291);
or U8706 (N_8706,N_7088,N_6508);
nor U8707 (N_8707,N_6902,N_6371);
and U8708 (N_8708,N_7353,N_6947);
and U8709 (N_8709,N_6837,N_7626);
nand U8710 (N_8710,N_7231,N_7485);
nor U8711 (N_8711,N_7171,N_6985);
nand U8712 (N_8712,N_7650,N_7653);
nand U8713 (N_8713,N_6228,N_6570);
xnor U8714 (N_8714,N_7767,N_6191);
nand U8715 (N_8715,N_7760,N_6785);
xor U8716 (N_8716,N_7989,N_6392);
xnor U8717 (N_8717,N_7208,N_7042);
or U8718 (N_8718,N_6748,N_7045);
or U8719 (N_8719,N_7514,N_7374);
and U8720 (N_8720,N_6054,N_6762);
nor U8721 (N_8721,N_6202,N_6914);
nor U8722 (N_8722,N_6712,N_6527);
nor U8723 (N_8723,N_6995,N_7554);
xor U8724 (N_8724,N_7577,N_6579);
nand U8725 (N_8725,N_6988,N_7089);
nand U8726 (N_8726,N_7931,N_7033);
xnor U8727 (N_8727,N_7549,N_7342);
nor U8728 (N_8728,N_6329,N_6989);
or U8729 (N_8729,N_7365,N_6350);
or U8730 (N_8730,N_7982,N_6472);
nand U8731 (N_8731,N_7264,N_7481);
nand U8732 (N_8732,N_7265,N_6461);
and U8733 (N_8733,N_6152,N_6662);
xor U8734 (N_8734,N_6155,N_7439);
nor U8735 (N_8735,N_7815,N_7967);
nor U8736 (N_8736,N_6622,N_7694);
and U8737 (N_8737,N_6747,N_6932);
and U8738 (N_8738,N_7763,N_7224);
nand U8739 (N_8739,N_7540,N_7905);
xnor U8740 (N_8740,N_7311,N_6455);
or U8741 (N_8741,N_7175,N_7419);
nand U8742 (N_8742,N_6171,N_7179);
or U8743 (N_8743,N_6827,N_6687);
nor U8744 (N_8744,N_6240,N_6782);
xnor U8745 (N_8745,N_7108,N_7123);
and U8746 (N_8746,N_7434,N_7255);
nand U8747 (N_8747,N_7791,N_6924);
nand U8748 (N_8748,N_6305,N_6999);
nor U8749 (N_8749,N_6261,N_6130);
nand U8750 (N_8750,N_7633,N_7321);
or U8751 (N_8751,N_7868,N_7232);
xnor U8752 (N_8752,N_6882,N_7691);
xor U8753 (N_8753,N_6167,N_7936);
nand U8754 (N_8754,N_6265,N_6567);
xor U8755 (N_8755,N_6923,N_6381);
and U8756 (N_8756,N_7061,N_6965);
nor U8757 (N_8757,N_6743,N_6573);
or U8758 (N_8758,N_7124,N_7341);
or U8759 (N_8759,N_6663,N_7170);
and U8760 (N_8760,N_6930,N_7294);
nor U8761 (N_8761,N_7624,N_7450);
and U8762 (N_8762,N_6866,N_7894);
nand U8763 (N_8763,N_7186,N_7740);
and U8764 (N_8764,N_7473,N_6015);
nor U8765 (N_8765,N_7559,N_7277);
nor U8766 (N_8766,N_7890,N_7690);
nor U8767 (N_8767,N_7678,N_7911);
nand U8768 (N_8768,N_6044,N_6018);
and U8769 (N_8769,N_7572,N_6517);
nand U8770 (N_8770,N_6163,N_6756);
and U8771 (N_8771,N_6384,N_7355);
xnor U8772 (N_8772,N_6004,N_7621);
xor U8773 (N_8773,N_6272,N_6062);
xor U8774 (N_8774,N_6398,N_7050);
xnor U8775 (N_8775,N_6244,N_7101);
or U8776 (N_8776,N_7347,N_6698);
nor U8777 (N_8777,N_7235,N_7147);
xor U8778 (N_8778,N_6292,N_7994);
xnor U8779 (N_8779,N_6504,N_6437);
or U8780 (N_8780,N_7161,N_6293);
or U8781 (N_8781,N_7267,N_7165);
or U8782 (N_8782,N_6523,N_6189);
nor U8783 (N_8783,N_6589,N_7295);
and U8784 (N_8784,N_6654,N_6713);
nand U8785 (N_8785,N_6540,N_7773);
nand U8786 (N_8786,N_7612,N_7800);
and U8787 (N_8787,N_6771,N_6157);
nor U8788 (N_8788,N_7141,N_7435);
or U8789 (N_8789,N_7542,N_7516);
nand U8790 (N_8790,N_6836,N_7944);
or U8791 (N_8791,N_6363,N_7500);
and U8792 (N_8792,N_7078,N_7599);
xnor U8793 (N_8793,N_6791,N_7553);
nor U8794 (N_8794,N_6595,N_6767);
or U8795 (N_8795,N_7505,N_6343);
and U8796 (N_8796,N_7584,N_7750);
xor U8797 (N_8797,N_6463,N_7067);
or U8798 (N_8798,N_6928,N_7838);
or U8799 (N_8799,N_6536,N_7461);
xor U8800 (N_8800,N_7995,N_6187);
xnor U8801 (N_8801,N_7049,N_7068);
nand U8802 (N_8802,N_6297,N_6408);
or U8803 (N_8803,N_6949,N_6506);
xor U8804 (N_8804,N_7987,N_6115);
nor U8805 (N_8805,N_7675,N_6076);
and U8806 (N_8806,N_6557,N_6613);
xor U8807 (N_8807,N_6848,N_7745);
nand U8808 (N_8808,N_7971,N_7048);
xnor U8809 (N_8809,N_6247,N_7899);
nor U8810 (N_8810,N_6676,N_6587);
and U8811 (N_8811,N_6591,N_7338);
and U8812 (N_8812,N_7297,N_6258);
and U8813 (N_8813,N_6322,N_6119);
nand U8814 (N_8814,N_7477,N_6610);
nor U8815 (N_8815,N_6146,N_6751);
nor U8816 (N_8816,N_7806,N_6092);
nor U8817 (N_8817,N_6471,N_6328);
nor U8818 (N_8818,N_7190,N_7859);
or U8819 (N_8819,N_7793,N_7006);
nor U8820 (N_8820,N_7410,N_7600);
nor U8821 (N_8821,N_7990,N_7465);
nor U8822 (N_8822,N_7737,N_6935);
nor U8823 (N_8823,N_6029,N_6755);
and U8824 (N_8824,N_7746,N_7580);
or U8825 (N_8825,N_6631,N_6576);
or U8826 (N_8826,N_7555,N_7563);
or U8827 (N_8827,N_7744,N_6869);
and U8828 (N_8828,N_7882,N_7099);
or U8829 (N_8829,N_6186,N_7025);
or U8830 (N_8830,N_6957,N_7002);
xor U8831 (N_8831,N_6876,N_6424);
and U8832 (N_8832,N_7063,N_7953);
and U8833 (N_8833,N_6606,N_7926);
xnor U8834 (N_8834,N_7845,N_7414);
nand U8835 (N_8835,N_7131,N_7081);
xor U8836 (N_8836,N_6833,N_6252);
or U8837 (N_8837,N_7272,N_6542);
and U8838 (N_8838,N_7046,N_7674);
nor U8839 (N_8839,N_7016,N_7148);
nand U8840 (N_8840,N_7220,N_6290);
or U8841 (N_8841,N_6114,N_6067);
and U8842 (N_8842,N_6563,N_6182);
or U8843 (N_8843,N_6090,N_7924);
or U8844 (N_8844,N_6443,N_6792);
or U8845 (N_8845,N_6842,N_6653);
nand U8846 (N_8846,N_7464,N_7394);
xor U8847 (N_8847,N_7897,N_7172);
nor U8848 (N_8848,N_7747,N_7804);
xnor U8849 (N_8849,N_6734,N_6982);
nand U8850 (N_8850,N_6530,N_6242);
nand U8851 (N_8851,N_7523,N_7941);
nand U8852 (N_8852,N_7522,N_7082);
or U8853 (N_8853,N_7807,N_7060);
or U8854 (N_8854,N_7266,N_7822);
nand U8855 (N_8855,N_6802,N_6056);
or U8856 (N_8856,N_6138,N_7968);
xnor U8857 (N_8857,N_6553,N_7446);
and U8858 (N_8858,N_6839,N_7609);
nor U8859 (N_8859,N_6904,N_6489);
nor U8860 (N_8860,N_6899,N_6180);
nor U8861 (N_8861,N_7133,N_6069);
nand U8862 (N_8862,N_7331,N_6819);
and U8863 (N_8863,N_7009,N_7981);
nand U8864 (N_8864,N_6154,N_6529);
xor U8865 (N_8865,N_7504,N_7769);
xnor U8866 (N_8866,N_7436,N_6002);
nor U8867 (N_8867,N_7947,N_7960);
and U8868 (N_8868,N_7701,N_6538);
or U8869 (N_8869,N_6776,N_7617);
nor U8870 (N_8870,N_7910,N_6042);
xor U8871 (N_8871,N_7023,N_6165);
nand U8872 (N_8872,N_7403,N_7304);
nand U8873 (N_8873,N_6215,N_7178);
nor U8874 (N_8874,N_6419,N_6482);
or U8875 (N_8875,N_6634,N_6174);
xor U8876 (N_8876,N_7651,N_7188);
or U8877 (N_8877,N_7438,N_7345);
and U8878 (N_8878,N_7177,N_6487);
xor U8879 (N_8879,N_6344,N_7797);
nor U8880 (N_8880,N_6758,N_6010);
xnor U8881 (N_8881,N_7385,N_6632);
xor U8882 (N_8882,N_6196,N_6617);
and U8883 (N_8883,N_6074,N_7455);
or U8884 (N_8884,N_7898,N_6598);
or U8885 (N_8885,N_6867,N_6183);
nor U8886 (N_8886,N_6366,N_7064);
or U8887 (N_8887,N_6539,N_7463);
nand U8888 (N_8888,N_7490,N_7772);
and U8889 (N_8889,N_7739,N_6091);
and U8890 (N_8890,N_6647,N_6901);
and U8891 (N_8891,N_7361,N_6400);
and U8892 (N_8892,N_6664,N_7001);
xor U8893 (N_8893,N_7597,N_6838);
or U8894 (N_8894,N_7658,N_6705);
or U8895 (N_8895,N_6855,N_7105);
nor U8896 (N_8896,N_7594,N_6578);
nor U8897 (N_8897,N_7513,N_6047);
nor U8898 (N_8898,N_6390,N_6212);
nor U8899 (N_8899,N_6414,N_6259);
nor U8900 (N_8900,N_6218,N_6551);
nor U8901 (N_8901,N_6145,N_7034);
nand U8902 (N_8902,N_7156,N_7492);
nor U8903 (N_8903,N_7884,N_7096);
xnor U8904 (N_8904,N_6402,N_6176);
nor U8905 (N_8905,N_7343,N_7079);
nor U8906 (N_8906,N_7669,N_6500);
nand U8907 (N_8907,N_7956,N_7754);
xnor U8908 (N_8908,N_6458,N_7233);
nand U8909 (N_8909,N_6895,N_6549);
or U8910 (N_8910,N_6944,N_7782);
or U8911 (N_8911,N_6382,N_7030);
and U8912 (N_8912,N_6675,N_7660);
nor U8913 (N_8913,N_7395,N_7228);
or U8914 (N_8914,N_7447,N_6660);
nand U8915 (N_8915,N_7527,N_7348);
and U8916 (N_8916,N_7387,N_7207);
nor U8917 (N_8917,N_7618,N_7276);
nand U8918 (N_8918,N_7689,N_7979);
or U8919 (N_8919,N_6066,N_6285);
or U8920 (N_8920,N_7702,N_6735);
nand U8921 (N_8921,N_6903,N_6724);
xnor U8922 (N_8922,N_6052,N_6185);
xnor U8923 (N_8923,N_7892,N_6262);
and U8924 (N_8924,N_6106,N_7850);
xor U8925 (N_8925,N_6916,N_7360);
nor U8926 (N_8926,N_7204,N_7925);
nor U8927 (N_8927,N_6283,N_6891);
and U8928 (N_8928,N_6626,N_7380);
or U8929 (N_8929,N_7732,N_6737);
nand U8930 (N_8930,N_7275,N_6726);
and U8931 (N_8931,N_7007,N_6192);
nor U8932 (N_8932,N_7221,N_6120);
xnor U8933 (N_8933,N_7392,N_6143);
nor U8934 (N_8934,N_6786,N_7528);
xor U8935 (N_8935,N_6825,N_6686);
and U8936 (N_8936,N_6166,N_6260);
nand U8937 (N_8937,N_7054,N_7192);
nor U8938 (N_8938,N_7482,N_7938);
nor U8939 (N_8939,N_6093,N_6609);
nand U8940 (N_8940,N_6124,N_7184);
xor U8941 (N_8941,N_7948,N_7961);
nand U8942 (N_8942,N_6620,N_7957);
nor U8943 (N_8943,N_7664,N_6162);
or U8944 (N_8944,N_6970,N_6396);
and U8945 (N_8945,N_7292,N_6680);
or U8946 (N_8946,N_6937,N_6801);
nor U8947 (N_8947,N_6073,N_7471);
or U8948 (N_8948,N_6991,N_7930);
nor U8949 (N_8949,N_7498,N_6497);
nor U8950 (N_8950,N_7518,N_7313);
or U8951 (N_8951,N_7325,N_6179);
or U8952 (N_8952,N_7107,N_7595);
nand U8953 (N_8953,N_6828,N_7827);
nand U8954 (N_8954,N_7670,N_7534);
or U8955 (N_8955,N_7893,N_6470);
and U8956 (N_8956,N_7709,N_6030);
nand U8957 (N_8957,N_6048,N_7071);
nand U8958 (N_8958,N_7613,N_7344);
xnor U8959 (N_8959,N_7524,N_6968);
and U8960 (N_8960,N_6910,N_6997);
xor U8961 (N_8961,N_6896,N_6667);
nand U8962 (N_8962,N_6809,N_6235);
nor U8963 (N_8963,N_7031,N_7545);
and U8964 (N_8964,N_6962,N_7478);
or U8965 (N_8965,N_7399,N_6820);
xnor U8966 (N_8966,N_7755,N_6715);
or U8967 (N_8967,N_6719,N_6684);
nor U8968 (N_8968,N_6484,N_6160);
and U8969 (N_8969,N_7413,N_7120);
or U8970 (N_8970,N_6694,N_7218);
nand U8971 (N_8971,N_7174,N_6515);
nor U8972 (N_8972,N_6243,N_6805);
or U8973 (N_8973,N_6385,N_7917);
nand U8974 (N_8974,N_7262,N_7307);
nand U8975 (N_8975,N_7429,N_6990);
xnor U8976 (N_8976,N_6225,N_7565);
xor U8977 (N_8977,N_7404,N_7959);
nand U8978 (N_8978,N_6784,N_7851);
xnor U8979 (N_8979,N_6415,N_6874);
or U8980 (N_8980,N_6700,N_6774);
xor U8981 (N_8981,N_7055,N_7799);
and U8982 (N_8982,N_7869,N_7566);
or U8983 (N_8983,N_6670,N_6571);
nor U8984 (N_8984,N_6681,N_7841);
nor U8985 (N_8985,N_7520,N_7467);
xor U8986 (N_8986,N_6863,N_6862);
nand U8987 (N_8987,N_7173,N_6541);
or U8988 (N_8988,N_7028,N_7605);
nor U8989 (N_8989,N_6884,N_6038);
or U8990 (N_8990,N_7854,N_7059);
nor U8991 (N_8991,N_6794,N_6922);
xor U8992 (N_8992,N_7856,N_6722);
nor U8993 (N_8993,N_6886,N_7328);
nor U8994 (N_8994,N_6721,N_7883);
or U8995 (N_8995,N_7943,N_6574);
and U8996 (N_8996,N_6690,N_7543);
and U8997 (N_8997,N_6865,N_7673);
and U8998 (N_8998,N_7039,N_6334);
and U8999 (N_8999,N_7630,N_6168);
nor U9000 (N_9000,N_6998,N_7921);
xnor U9001 (N_9001,N_6881,N_6657);
or U9002 (N_9002,N_7655,N_7942);
xor U9003 (N_9003,N_6062,N_7643);
xor U9004 (N_9004,N_6635,N_7349);
and U9005 (N_9005,N_6141,N_6386);
and U9006 (N_9006,N_7458,N_6519);
nor U9007 (N_9007,N_7902,N_6088);
nor U9008 (N_9008,N_6224,N_6168);
and U9009 (N_9009,N_6559,N_7069);
nor U9010 (N_9010,N_7245,N_7309);
xor U9011 (N_9011,N_7147,N_6248);
xor U9012 (N_9012,N_6345,N_6637);
or U9013 (N_9013,N_7759,N_7705);
nor U9014 (N_9014,N_6494,N_7354);
xor U9015 (N_9015,N_7700,N_7395);
nor U9016 (N_9016,N_7995,N_6780);
xor U9017 (N_9017,N_7116,N_6360);
nor U9018 (N_9018,N_6160,N_7498);
or U9019 (N_9019,N_6243,N_7064);
nor U9020 (N_9020,N_6962,N_7912);
or U9021 (N_9021,N_6731,N_6564);
nand U9022 (N_9022,N_6253,N_7834);
nand U9023 (N_9023,N_7717,N_6729);
xnor U9024 (N_9024,N_6405,N_7636);
nor U9025 (N_9025,N_7898,N_6618);
nor U9026 (N_9026,N_6491,N_6142);
and U9027 (N_9027,N_6937,N_6581);
nand U9028 (N_9028,N_6549,N_6824);
xor U9029 (N_9029,N_6483,N_6961);
nand U9030 (N_9030,N_6797,N_6513);
nand U9031 (N_9031,N_6517,N_6414);
and U9032 (N_9032,N_6277,N_7557);
xor U9033 (N_9033,N_7514,N_6435);
or U9034 (N_9034,N_6783,N_7977);
nor U9035 (N_9035,N_6580,N_6408);
nand U9036 (N_9036,N_6895,N_6962);
nor U9037 (N_9037,N_6630,N_7975);
and U9038 (N_9038,N_6400,N_6852);
nor U9039 (N_9039,N_6251,N_7968);
and U9040 (N_9040,N_6548,N_6552);
and U9041 (N_9041,N_7765,N_7979);
xnor U9042 (N_9042,N_7133,N_7223);
nand U9043 (N_9043,N_6649,N_7935);
xnor U9044 (N_9044,N_7120,N_6891);
nand U9045 (N_9045,N_7972,N_6649);
or U9046 (N_9046,N_6280,N_6112);
nor U9047 (N_9047,N_7608,N_6075);
and U9048 (N_9048,N_7896,N_7743);
xnor U9049 (N_9049,N_7888,N_6368);
nand U9050 (N_9050,N_6697,N_6157);
nor U9051 (N_9051,N_7139,N_6278);
or U9052 (N_9052,N_7192,N_7543);
nor U9053 (N_9053,N_6819,N_7677);
and U9054 (N_9054,N_6493,N_7455);
or U9055 (N_9055,N_7945,N_6338);
and U9056 (N_9056,N_6391,N_6687);
nor U9057 (N_9057,N_6536,N_6962);
nand U9058 (N_9058,N_7457,N_7909);
xnor U9059 (N_9059,N_6595,N_7601);
nand U9060 (N_9060,N_6205,N_7038);
nor U9061 (N_9061,N_7418,N_7074);
xor U9062 (N_9062,N_7579,N_7901);
nor U9063 (N_9063,N_7292,N_6482);
nand U9064 (N_9064,N_7742,N_7132);
or U9065 (N_9065,N_7808,N_6590);
and U9066 (N_9066,N_7577,N_7621);
nand U9067 (N_9067,N_7720,N_7782);
xnor U9068 (N_9068,N_7472,N_6085);
and U9069 (N_9069,N_7380,N_6995);
nor U9070 (N_9070,N_7268,N_6419);
nand U9071 (N_9071,N_7587,N_6994);
xor U9072 (N_9072,N_7271,N_7842);
nor U9073 (N_9073,N_7323,N_7268);
nor U9074 (N_9074,N_7053,N_6785);
nor U9075 (N_9075,N_6139,N_7248);
and U9076 (N_9076,N_6675,N_7273);
nand U9077 (N_9077,N_6103,N_6485);
or U9078 (N_9078,N_7565,N_7617);
nand U9079 (N_9079,N_6524,N_7935);
nor U9080 (N_9080,N_6021,N_7492);
or U9081 (N_9081,N_7445,N_7956);
nand U9082 (N_9082,N_6261,N_6599);
nand U9083 (N_9083,N_7109,N_6624);
or U9084 (N_9084,N_6366,N_6119);
nor U9085 (N_9085,N_6136,N_6654);
nor U9086 (N_9086,N_7726,N_7604);
nand U9087 (N_9087,N_6186,N_7896);
nand U9088 (N_9088,N_6613,N_7702);
nand U9089 (N_9089,N_7453,N_7468);
nor U9090 (N_9090,N_7680,N_6667);
nand U9091 (N_9091,N_6585,N_6320);
nand U9092 (N_9092,N_6765,N_7665);
xnor U9093 (N_9093,N_6250,N_6972);
nand U9094 (N_9094,N_7154,N_6856);
and U9095 (N_9095,N_7295,N_7920);
and U9096 (N_9096,N_7698,N_6899);
and U9097 (N_9097,N_7725,N_7710);
nor U9098 (N_9098,N_7152,N_7139);
xor U9099 (N_9099,N_7605,N_6326);
nand U9100 (N_9100,N_7066,N_7152);
nand U9101 (N_9101,N_7334,N_6110);
xor U9102 (N_9102,N_7020,N_7023);
and U9103 (N_9103,N_7626,N_7290);
nor U9104 (N_9104,N_7987,N_7206);
nand U9105 (N_9105,N_6897,N_7267);
xnor U9106 (N_9106,N_6875,N_6836);
nand U9107 (N_9107,N_6282,N_6664);
nand U9108 (N_9108,N_6389,N_7453);
and U9109 (N_9109,N_6116,N_7327);
nand U9110 (N_9110,N_6027,N_7308);
nand U9111 (N_9111,N_7752,N_7472);
xnor U9112 (N_9112,N_7527,N_7487);
nand U9113 (N_9113,N_7084,N_7759);
and U9114 (N_9114,N_6503,N_7981);
or U9115 (N_9115,N_7429,N_6301);
nor U9116 (N_9116,N_6364,N_7642);
or U9117 (N_9117,N_6505,N_6406);
and U9118 (N_9118,N_7831,N_6248);
nor U9119 (N_9119,N_6330,N_7855);
and U9120 (N_9120,N_7525,N_6643);
and U9121 (N_9121,N_7396,N_6665);
nand U9122 (N_9122,N_6603,N_6645);
and U9123 (N_9123,N_7036,N_7623);
xnor U9124 (N_9124,N_7810,N_7849);
xnor U9125 (N_9125,N_6201,N_6014);
and U9126 (N_9126,N_7274,N_7292);
or U9127 (N_9127,N_7054,N_6480);
nand U9128 (N_9128,N_6457,N_6352);
and U9129 (N_9129,N_6487,N_6258);
nand U9130 (N_9130,N_7608,N_7081);
and U9131 (N_9131,N_7369,N_6195);
nand U9132 (N_9132,N_7368,N_6561);
and U9133 (N_9133,N_6527,N_6877);
nand U9134 (N_9134,N_7886,N_6254);
and U9135 (N_9135,N_6536,N_7493);
nor U9136 (N_9136,N_6777,N_7032);
nand U9137 (N_9137,N_7763,N_7436);
or U9138 (N_9138,N_7251,N_7764);
nand U9139 (N_9139,N_6097,N_6132);
and U9140 (N_9140,N_7394,N_6424);
or U9141 (N_9141,N_6611,N_7252);
xnor U9142 (N_9142,N_6977,N_6631);
and U9143 (N_9143,N_7661,N_6708);
xnor U9144 (N_9144,N_7950,N_6381);
nand U9145 (N_9145,N_6761,N_6108);
and U9146 (N_9146,N_7683,N_7794);
or U9147 (N_9147,N_6539,N_6946);
nor U9148 (N_9148,N_6990,N_6849);
xnor U9149 (N_9149,N_7834,N_7245);
nand U9150 (N_9150,N_7280,N_6932);
or U9151 (N_9151,N_7077,N_6480);
nor U9152 (N_9152,N_6990,N_6300);
and U9153 (N_9153,N_6440,N_6253);
xnor U9154 (N_9154,N_6832,N_6551);
and U9155 (N_9155,N_6118,N_6804);
nor U9156 (N_9156,N_7804,N_7924);
nor U9157 (N_9157,N_6421,N_6727);
and U9158 (N_9158,N_6747,N_6714);
and U9159 (N_9159,N_6649,N_7783);
nor U9160 (N_9160,N_6284,N_7525);
and U9161 (N_9161,N_6699,N_6110);
and U9162 (N_9162,N_6305,N_6206);
or U9163 (N_9163,N_7207,N_7880);
xnor U9164 (N_9164,N_7775,N_7263);
and U9165 (N_9165,N_7924,N_6581);
or U9166 (N_9166,N_7336,N_7120);
nor U9167 (N_9167,N_7014,N_6265);
or U9168 (N_9168,N_6714,N_6477);
and U9169 (N_9169,N_6844,N_7367);
and U9170 (N_9170,N_7687,N_7847);
xor U9171 (N_9171,N_7871,N_7500);
nor U9172 (N_9172,N_7906,N_7083);
nand U9173 (N_9173,N_6457,N_7882);
nor U9174 (N_9174,N_7969,N_7375);
nand U9175 (N_9175,N_6154,N_6418);
and U9176 (N_9176,N_6081,N_7842);
xor U9177 (N_9177,N_6769,N_6657);
or U9178 (N_9178,N_7007,N_6763);
nand U9179 (N_9179,N_7340,N_6754);
xnor U9180 (N_9180,N_7320,N_7871);
or U9181 (N_9181,N_6927,N_7628);
nor U9182 (N_9182,N_6921,N_6622);
and U9183 (N_9183,N_6517,N_7861);
and U9184 (N_9184,N_7250,N_6617);
or U9185 (N_9185,N_6686,N_7927);
nand U9186 (N_9186,N_7915,N_7817);
or U9187 (N_9187,N_7375,N_7484);
and U9188 (N_9188,N_7775,N_6064);
xnor U9189 (N_9189,N_6951,N_6199);
xor U9190 (N_9190,N_6622,N_6302);
xnor U9191 (N_9191,N_7563,N_7451);
xnor U9192 (N_9192,N_7944,N_7874);
and U9193 (N_9193,N_6477,N_6058);
and U9194 (N_9194,N_6139,N_6364);
nor U9195 (N_9195,N_6918,N_7631);
nor U9196 (N_9196,N_6765,N_6626);
or U9197 (N_9197,N_7244,N_7994);
or U9198 (N_9198,N_6169,N_7376);
or U9199 (N_9199,N_6618,N_7019);
xnor U9200 (N_9200,N_7129,N_6353);
xnor U9201 (N_9201,N_6236,N_7082);
nor U9202 (N_9202,N_7385,N_6403);
xnor U9203 (N_9203,N_6129,N_7700);
nor U9204 (N_9204,N_7729,N_7861);
and U9205 (N_9205,N_7404,N_7070);
nand U9206 (N_9206,N_6230,N_7196);
and U9207 (N_9207,N_6078,N_7220);
xnor U9208 (N_9208,N_7908,N_6065);
or U9209 (N_9209,N_7902,N_6676);
or U9210 (N_9210,N_6650,N_6154);
and U9211 (N_9211,N_6541,N_7194);
and U9212 (N_9212,N_6474,N_7430);
or U9213 (N_9213,N_7075,N_7720);
nand U9214 (N_9214,N_6710,N_7087);
xnor U9215 (N_9215,N_6077,N_7975);
and U9216 (N_9216,N_7680,N_7895);
or U9217 (N_9217,N_6707,N_7442);
xor U9218 (N_9218,N_7830,N_6304);
nand U9219 (N_9219,N_7939,N_7204);
xnor U9220 (N_9220,N_6695,N_7938);
and U9221 (N_9221,N_6242,N_7861);
and U9222 (N_9222,N_7253,N_7337);
xor U9223 (N_9223,N_7019,N_6847);
nand U9224 (N_9224,N_7491,N_6181);
xnor U9225 (N_9225,N_6362,N_7300);
xor U9226 (N_9226,N_6294,N_6354);
or U9227 (N_9227,N_6142,N_7341);
and U9228 (N_9228,N_6811,N_6114);
xnor U9229 (N_9229,N_7887,N_6773);
or U9230 (N_9230,N_6994,N_6812);
and U9231 (N_9231,N_7987,N_6588);
or U9232 (N_9232,N_7438,N_6190);
nand U9233 (N_9233,N_6786,N_6604);
nor U9234 (N_9234,N_6661,N_7182);
or U9235 (N_9235,N_6543,N_7739);
nor U9236 (N_9236,N_7798,N_6622);
nor U9237 (N_9237,N_7565,N_6315);
nor U9238 (N_9238,N_6736,N_7278);
nor U9239 (N_9239,N_7180,N_6989);
and U9240 (N_9240,N_6480,N_6499);
xnor U9241 (N_9241,N_6881,N_6972);
nor U9242 (N_9242,N_7736,N_7833);
nor U9243 (N_9243,N_7494,N_7858);
or U9244 (N_9244,N_7093,N_7634);
or U9245 (N_9245,N_6518,N_7360);
nor U9246 (N_9246,N_7226,N_7915);
xor U9247 (N_9247,N_7179,N_7736);
nand U9248 (N_9248,N_6886,N_7594);
or U9249 (N_9249,N_7046,N_6390);
nor U9250 (N_9250,N_6850,N_6565);
xor U9251 (N_9251,N_6121,N_7436);
nand U9252 (N_9252,N_6840,N_7509);
or U9253 (N_9253,N_7130,N_7877);
xor U9254 (N_9254,N_7484,N_6395);
nand U9255 (N_9255,N_7262,N_6443);
nand U9256 (N_9256,N_6431,N_6028);
nor U9257 (N_9257,N_7140,N_7481);
and U9258 (N_9258,N_7526,N_6307);
nand U9259 (N_9259,N_6564,N_7283);
or U9260 (N_9260,N_6033,N_7055);
xnor U9261 (N_9261,N_6654,N_7457);
and U9262 (N_9262,N_6243,N_7216);
and U9263 (N_9263,N_6061,N_7653);
nand U9264 (N_9264,N_7018,N_7617);
and U9265 (N_9265,N_6504,N_6561);
nand U9266 (N_9266,N_7848,N_7913);
xor U9267 (N_9267,N_6347,N_7169);
or U9268 (N_9268,N_6833,N_7912);
nand U9269 (N_9269,N_7832,N_7489);
or U9270 (N_9270,N_6491,N_6002);
or U9271 (N_9271,N_7905,N_7570);
nor U9272 (N_9272,N_6758,N_7978);
and U9273 (N_9273,N_7315,N_7046);
xor U9274 (N_9274,N_7400,N_6400);
or U9275 (N_9275,N_6331,N_7684);
xnor U9276 (N_9276,N_6261,N_6133);
nor U9277 (N_9277,N_6497,N_6695);
xnor U9278 (N_9278,N_7323,N_7839);
xor U9279 (N_9279,N_6709,N_6946);
nor U9280 (N_9280,N_7993,N_6144);
nand U9281 (N_9281,N_6442,N_6265);
nor U9282 (N_9282,N_6040,N_6885);
nand U9283 (N_9283,N_6145,N_7610);
nor U9284 (N_9284,N_7714,N_6734);
xnor U9285 (N_9285,N_6454,N_6485);
nand U9286 (N_9286,N_6311,N_7529);
and U9287 (N_9287,N_6061,N_6686);
or U9288 (N_9288,N_7898,N_6429);
and U9289 (N_9289,N_6835,N_6815);
or U9290 (N_9290,N_7849,N_7710);
and U9291 (N_9291,N_7705,N_7037);
xnor U9292 (N_9292,N_7527,N_7875);
and U9293 (N_9293,N_7676,N_7853);
nand U9294 (N_9294,N_6586,N_7449);
xor U9295 (N_9295,N_7801,N_6225);
xor U9296 (N_9296,N_7378,N_6435);
xor U9297 (N_9297,N_7584,N_7404);
xnor U9298 (N_9298,N_6894,N_7881);
nand U9299 (N_9299,N_6315,N_6472);
and U9300 (N_9300,N_6618,N_7535);
xnor U9301 (N_9301,N_6697,N_6947);
or U9302 (N_9302,N_7294,N_6946);
and U9303 (N_9303,N_7106,N_7381);
and U9304 (N_9304,N_7352,N_6318);
or U9305 (N_9305,N_7999,N_6105);
nand U9306 (N_9306,N_7568,N_6716);
or U9307 (N_9307,N_7256,N_6255);
nor U9308 (N_9308,N_7181,N_6664);
nand U9309 (N_9309,N_6471,N_6634);
nor U9310 (N_9310,N_6262,N_6258);
or U9311 (N_9311,N_7652,N_6001);
or U9312 (N_9312,N_6768,N_7322);
nand U9313 (N_9313,N_6943,N_6667);
nand U9314 (N_9314,N_7173,N_6890);
nand U9315 (N_9315,N_7441,N_6664);
xor U9316 (N_9316,N_6519,N_6510);
and U9317 (N_9317,N_6551,N_7416);
xor U9318 (N_9318,N_7969,N_6197);
or U9319 (N_9319,N_6639,N_7707);
and U9320 (N_9320,N_7180,N_6739);
and U9321 (N_9321,N_7756,N_7912);
nor U9322 (N_9322,N_7074,N_7125);
nand U9323 (N_9323,N_7575,N_7914);
or U9324 (N_9324,N_7060,N_7221);
xor U9325 (N_9325,N_7638,N_6659);
nor U9326 (N_9326,N_7109,N_7607);
or U9327 (N_9327,N_7032,N_7565);
nand U9328 (N_9328,N_6007,N_7978);
or U9329 (N_9329,N_6876,N_6259);
nand U9330 (N_9330,N_6842,N_6164);
xnor U9331 (N_9331,N_6191,N_6066);
and U9332 (N_9332,N_6632,N_6565);
nor U9333 (N_9333,N_6675,N_7389);
and U9334 (N_9334,N_7682,N_7472);
or U9335 (N_9335,N_7459,N_6448);
and U9336 (N_9336,N_7498,N_7493);
or U9337 (N_9337,N_7617,N_6403);
and U9338 (N_9338,N_6037,N_6919);
nor U9339 (N_9339,N_7438,N_6890);
xnor U9340 (N_9340,N_6432,N_6322);
and U9341 (N_9341,N_6111,N_7055);
nand U9342 (N_9342,N_7670,N_6805);
xor U9343 (N_9343,N_7505,N_7711);
and U9344 (N_9344,N_6871,N_6924);
nand U9345 (N_9345,N_6987,N_7344);
and U9346 (N_9346,N_6973,N_6331);
or U9347 (N_9347,N_7998,N_7769);
nand U9348 (N_9348,N_6802,N_6299);
and U9349 (N_9349,N_7576,N_7453);
nand U9350 (N_9350,N_7524,N_6277);
nand U9351 (N_9351,N_7010,N_7196);
or U9352 (N_9352,N_6367,N_7488);
and U9353 (N_9353,N_7934,N_7473);
and U9354 (N_9354,N_7836,N_7581);
and U9355 (N_9355,N_6513,N_6877);
or U9356 (N_9356,N_7986,N_6275);
and U9357 (N_9357,N_7315,N_6980);
nand U9358 (N_9358,N_7301,N_6165);
xnor U9359 (N_9359,N_6946,N_6744);
nand U9360 (N_9360,N_6835,N_6581);
and U9361 (N_9361,N_6506,N_7574);
or U9362 (N_9362,N_7342,N_7737);
nor U9363 (N_9363,N_6538,N_7635);
nor U9364 (N_9364,N_7378,N_6423);
nand U9365 (N_9365,N_7235,N_6306);
nor U9366 (N_9366,N_7727,N_6432);
and U9367 (N_9367,N_7973,N_6465);
nor U9368 (N_9368,N_7293,N_7670);
nand U9369 (N_9369,N_6142,N_7162);
and U9370 (N_9370,N_7455,N_7545);
and U9371 (N_9371,N_6953,N_6850);
xnor U9372 (N_9372,N_7416,N_6063);
xor U9373 (N_9373,N_6624,N_7871);
or U9374 (N_9374,N_6087,N_6440);
xnor U9375 (N_9375,N_7723,N_7588);
and U9376 (N_9376,N_7837,N_7820);
nor U9377 (N_9377,N_6888,N_6194);
nand U9378 (N_9378,N_7624,N_7486);
xor U9379 (N_9379,N_6964,N_6874);
nand U9380 (N_9380,N_6064,N_7968);
xnor U9381 (N_9381,N_6858,N_7732);
and U9382 (N_9382,N_6713,N_6454);
xor U9383 (N_9383,N_6140,N_7354);
or U9384 (N_9384,N_7476,N_6006);
nand U9385 (N_9385,N_7976,N_7526);
nand U9386 (N_9386,N_6558,N_7289);
nand U9387 (N_9387,N_7727,N_7474);
nand U9388 (N_9388,N_7338,N_6563);
and U9389 (N_9389,N_7921,N_6675);
nand U9390 (N_9390,N_7359,N_6577);
and U9391 (N_9391,N_7832,N_7393);
or U9392 (N_9392,N_7999,N_7172);
and U9393 (N_9393,N_7404,N_6176);
or U9394 (N_9394,N_6138,N_6335);
nor U9395 (N_9395,N_6881,N_6621);
nand U9396 (N_9396,N_7837,N_7309);
nor U9397 (N_9397,N_6143,N_7512);
or U9398 (N_9398,N_7524,N_7995);
nand U9399 (N_9399,N_7632,N_6655);
or U9400 (N_9400,N_7175,N_6321);
nor U9401 (N_9401,N_6736,N_7135);
xnor U9402 (N_9402,N_7560,N_7536);
and U9403 (N_9403,N_7862,N_6337);
and U9404 (N_9404,N_6065,N_7501);
xor U9405 (N_9405,N_6548,N_7696);
xnor U9406 (N_9406,N_7805,N_6201);
xnor U9407 (N_9407,N_6712,N_7984);
or U9408 (N_9408,N_6074,N_6847);
nand U9409 (N_9409,N_7501,N_7541);
nand U9410 (N_9410,N_6182,N_7445);
and U9411 (N_9411,N_7464,N_7892);
xor U9412 (N_9412,N_6523,N_7778);
xnor U9413 (N_9413,N_6478,N_7581);
xor U9414 (N_9414,N_7853,N_7276);
or U9415 (N_9415,N_6361,N_6465);
nor U9416 (N_9416,N_7958,N_6462);
nand U9417 (N_9417,N_6759,N_7849);
nand U9418 (N_9418,N_6401,N_7694);
xnor U9419 (N_9419,N_6260,N_7096);
nor U9420 (N_9420,N_6348,N_6956);
and U9421 (N_9421,N_7975,N_6661);
xnor U9422 (N_9422,N_6784,N_7404);
or U9423 (N_9423,N_6421,N_6324);
or U9424 (N_9424,N_6750,N_7916);
nor U9425 (N_9425,N_7793,N_6316);
xor U9426 (N_9426,N_6461,N_7990);
and U9427 (N_9427,N_6467,N_7235);
nor U9428 (N_9428,N_6288,N_7123);
nor U9429 (N_9429,N_7653,N_7507);
and U9430 (N_9430,N_6653,N_7331);
or U9431 (N_9431,N_6623,N_7803);
xnor U9432 (N_9432,N_7428,N_6877);
and U9433 (N_9433,N_7482,N_6878);
nand U9434 (N_9434,N_7454,N_6563);
and U9435 (N_9435,N_6245,N_6861);
and U9436 (N_9436,N_7204,N_7003);
nor U9437 (N_9437,N_6651,N_6902);
xnor U9438 (N_9438,N_7075,N_7932);
or U9439 (N_9439,N_6337,N_7394);
nand U9440 (N_9440,N_6888,N_7895);
xnor U9441 (N_9441,N_7981,N_6502);
or U9442 (N_9442,N_7419,N_7301);
xnor U9443 (N_9443,N_6307,N_6855);
nor U9444 (N_9444,N_6746,N_7040);
xnor U9445 (N_9445,N_6614,N_6685);
nand U9446 (N_9446,N_7733,N_7667);
nand U9447 (N_9447,N_7957,N_6315);
and U9448 (N_9448,N_6309,N_7546);
or U9449 (N_9449,N_7969,N_6703);
nand U9450 (N_9450,N_6741,N_6482);
and U9451 (N_9451,N_6601,N_6013);
nand U9452 (N_9452,N_6154,N_6266);
xnor U9453 (N_9453,N_6549,N_6241);
and U9454 (N_9454,N_7789,N_6569);
or U9455 (N_9455,N_6793,N_7534);
xnor U9456 (N_9456,N_6114,N_6783);
and U9457 (N_9457,N_6470,N_7657);
xnor U9458 (N_9458,N_7557,N_7262);
nor U9459 (N_9459,N_6942,N_6382);
nand U9460 (N_9460,N_7588,N_7656);
nand U9461 (N_9461,N_7437,N_6166);
xnor U9462 (N_9462,N_7943,N_7666);
nor U9463 (N_9463,N_7973,N_6152);
nand U9464 (N_9464,N_6183,N_7934);
or U9465 (N_9465,N_6447,N_7370);
nand U9466 (N_9466,N_7176,N_7131);
xnor U9467 (N_9467,N_7256,N_7106);
xor U9468 (N_9468,N_7219,N_7892);
xor U9469 (N_9469,N_6862,N_7666);
nand U9470 (N_9470,N_6501,N_7288);
nand U9471 (N_9471,N_6658,N_7674);
or U9472 (N_9472,N_6420,N_7956);
nand U9473 (N_9473,N_6880,N_7518);
nor U9474 (N_9474,N_7125,N_7407);
and U9475 (N_9475,N_6517,N_6807);
and U9476 (N_9476,N_6826,N_6615);
xnor U9477 (N_9477,N_6891,N_7041);
nor U9478 (N_9478,N_6553,N_6099);
xor U9479 (N_9479,N_7332,N_7871);
nor U9480 (N_9480,N_6089,N_6922);
xnor U9481 (N_9481,N_6679,N_7999);
or U9482 (N_9482,N_6980,N_7769);
nand U9483 (N_9483,N_6140,N_7025);
or U9484 (N_9484,N_7899,N_6974);
xnor U9485 (N_9485,N_7332,N_7175);
or U9486 (N_9486,N_6635,N_7119);
or U9487 (N_9487,N_6098,N_6120);
or U9488 (N_9488,N_7682,N_6883);
nor U9489 (N_9489,N_6648,N_7570);
nor U9490 (N_9490,N_7422,N_7444);
and U9491 (N_9491,N_6136,N_7163);
xor U9492 (N_9492,N_7663,N_7594);
xor U9493 (N_9493,N_7514,N_6124);
and U9494 (N_9494,N_6285,N_7857);
or U9495 (N_9495,N_7897,N_7095);
nor U9496 (N_9496,N_7150,N_7666);
nor U9497 (N_9497,N_6173,N_7789);
nand U9498 (N_9498,N_6435,N_7687);
nor U9499 (N_9499,N_6457,N_7059);
and U9500 (N_9500,N_7855,N_6881);
xor U9501 (N_9501,N_7180,N_6163);
nand U9502 (N_9502,N_6169,N_6141);
and U9503 (N_9503,N_7930,N_6174);
or U9504 (N_9504,N_7469,N_6183);
xnor U9505 (N_9505,N_7088,N_6900);
or U9506 (N_9506,N_7066,N_6236);
nor U9507 (N_9507,N_6872,N_7594);
xnor U9508 (N_9508,N_6364,N_6286);
nand U9509 (N_9509,N_7333,N_7013);
nor U9510 (N_9510,N_7519,N_7029);
xor U9511 (N_9511,N_6706,N_6114);
or U9512 (N_9512,N_7352,N_7762);
nand U9513 (N_9513,N_6761,N_6751);
and U9514 (N_9514,N_6182,N_6300);
xor U9515 (N_9515,N_7451,N_6838);
xnor U9516 (N_9516,N_7022,N_6287);
nand U9517 (N_9517,N_6402,N_6595);
xnor U9518 (N_9518,N_6085,N_7928);
nand U9519 (N_9519,N_7870,N_7585);
nand U9520 (N_9520,N_6148,N_7879);
nor U9521 (N_9521,N_6547,N_6152);
nor U9522 (N_9522,N_7524,N_6237);
or U9523 (N_9523,N_6892,N_7542);
nand U9524 (N_9524,N_7684,N_7779);
xor U9525 (N_9525,N_7149,N_6604);
nand U9526 (N_9526,N_7163,N_6483);
and U9527 (N_9527,N_7125,N_6296);
nor U9528 (N_9528,N_7765,N_6798);
or U9529 (N_9529,N_6267,N_7428);
and U9530 (N_9530,N_6969,N_7337);
or U9531 (N_9531,N_6427,N_6748);
nor U9532 (N_9532,N_6840,N_7005);
or U9533 (N_9533,N_6689,N_6326);
or U9534 (N_9534,N_6023,N_7132);
and U9535 (N_9535,N_6844,N_6756);
xor U9536 (N_9536,N_6084,N_7415);
or U9537 (N_9537,N_7410,N_7186);
xor U9538 (N_9538,N_7026,N_7067);
xnor U9539 (N_9539,N_6333,N_6640);
nor U9540 (N_9540,N_7510,N_7899);
nor U9541 (N_9541,N_6584,N_7418);
xnor U9542 (N_9542,N_6794,N_7079);
nor U9543 (N_9543,N_7863,N_7154);
xnor U9544 (N_9544,N_7890,N_7218);
or U9545 (N_9545,N_6223,N_7185);
and U9546 (N_9546,N_7367,N_6453);
nand U9547 (N_9547,N_7001,N_6972);
xor U9548 (N_9548,N_7886,N_6506);
nand U9549 (N_9549,N_7412,N_7259);
nor U9550 (N_9550,N_6343,N_6674);
nor U9551 (N_9551,N_6320,N_6568);
nand U9552 (N_9552,N_7488,N_7154);
nor U9553 (N_9553,N_6156,N_7785);
or U9554 (N_9554,N_6735,N_7268);
and U9555 (N_9555,N_6443,N_6977);
and U9556 (N_9556,N_6139,N_6539);
nand U9557 (N_9557,N_7564,N_6142);
and U9558 (N_9558,N_7411,N_6233);
xor U9559 (N_9559,N_7350,N_7302);
nor U9560 (N_9560,N_7128,N_6424);
nand U9561 (N_9561,N_7044,N_6026);
and U9562 (N_9562,N_6617,N_7266);
nor U9563 (N_9563,N_6738,N_7944);
xnor U9564 (N_9564,N_6134,N_7885);
and U9565 (N_9565,N_7435,N_7078);
nor U9566 (N_9566,N_6311,N_7104);
and U9567 (N_9567,N_7919,N_7278);
and U9568 (N_9568,N_7804,N_6559);
nand U9569 (N_9569,N_6854,N_7834);
or U9570 (N_9570,N_7891,N_6040);
or U9571 (N_9571,N_6223,N_6556);
xor U9572 (N_9572,N_7833,N_6564);
nand U9573 (N_9573,N_6542,N_6926);
nor U9574 (N_9574,N_7460,N_6933);
or U9575 (N_9575,N_7194,N_6734);
xnor U9576 (N_9576,N_7998,N_6198);
xnor U9577 (N_9577,N_7338,N_6695);
or U9578 (N_9578,N_6710,N_7716);
and U9579 (N_9579,N_7111,N_7211);
and U9580 (N_9580,N_7569,N_6413);
and U9581 (N_9581,N_7280,N_7258);
nand U9582 (N_9582,N_7875,N_7759);
and U9583 (N_9583,N_6212,N_6714);
or U9584 (N_9584,N_6929,N_6342);
xnor U9585 (N_9585,N_6983,N_7948);
and U9586 (N_9586,N_7435,N_6551);
and U9587 (N_9587,N_7678,N_6249);
and U9588 (N_9588,N_6794,N_7448);
nor U9589 (N_9589,N_7168,N_7598);
and U9590 (N_9590,N_6950,N_6207);
or U9591 (N_9591,N_6600,N_6083);
nand U9592 (N_9592,N_6527,N_7147);
xnor U9593 (N_9593,N_7799,N_7925);
nand U9594 (N_9594,N_7380,N_6268);
nor U9595 (N_9595,N_7030,N_7831);
nand U9596 (N_9596,N_6926,N_6825);
or U9597 (N_9597,N_7465,N_7096);
xnor U9598 (N_9598,N_6851,N_6089);
and U9599 (N_9599,N_7921,N_7197);
xnor U9600 (N_9600,N_6761,N_6433);
nor U9601 (N_9601,N_7322,N_6380);
xnor U9602 (N_9602,N_7061,N_6528);
or U9603 (N_9603,N_6967,N_7810);
and U9604 (N_9604,N_7245,N_6120);
nor U9605 (N_9605,N_7649,N_7979);
nand U9606 (N_9606,N_7283,N_7724);
nor U9607 (N_9607,N_7987,N_6271);
and U9608 (N_9608,N_7806,N_7742);
xor U9609 (N_9609,N_6428,N_7487);
nand U9610 (N_9610,N_6670,N_6938);
and U9611 (N_9611,N_7420,N_7483);
xnor U9612 (N_9612,N_6156,N_7535);
and U9613 (N_9613,N_7557,N_7697);
or U9614 (N_9614,N_6599,N_7651);
or U9615 (N_9615,N_6800,N_6827);
and U9616 (N_9616,N_7382,N_6867);
or U9617 (N_9617,N_6697,N_7988);
nor U9618 (N_9618,N_7565,N_6214);
xor U9619 (N_9619,N_7177,N_6654);
xnor U9620 (N_9620,N_6278,N_6770);
and U9621 (N_9621,N_7170,N_7395);
nor U9622 (N_9622,N_6776,N_7110);
nor U9623 (N_9623,N_7896,N_6419);
and U9624 (N_9624,N_7933,N_7395);
or U9625 (N_9625,N_6074,N_6054);
and U9626 (N_9626,N_7664,N_7603);
nor U9627 (N_9627,N_6122,N_6138);
nor U9628 (N_9628,N_7471,N_7687);
xor U9629 (N_9629,N_6492,N_6515);
xnor U9630 (N_9630,N_6152,N_7906);
nand U9631 (N_9631,N_7424,N_7169);
or U9632 (N_9632,N_6627,N_7480);
and U9633 (N_9633,N_6535,N_7110);
and U9634 (N_9634,N_7826,N_6970);
and U9635 (N_9635,N_7294,N_6836);
nand U9636 (N_9636,N_6176,N_6968);
and U9637 (N_9637,N_7976,N_7532);
nor U9638 (N_9638,N_7563,N_7424);
and U9639 (N_9639,N_7354,N_6452);
and U9640 (N_9640,N_6741,N_7543);
and U9641 (N_9641,N_6536,N_6743);
nand U9642 (N_9642,N_7030,N_7062);
nand U9643 (N_9643,N_6592,N_6032);
xnor U9644 (N_9644,N_7010,N_6929);
xnor U9645 (N_9645,N_6145,N_7724);
nor U9646 (N_9646,N_7611,N_6841);
xor U9647 (N_9647,N_6160,N_6815);
and U9648 (N_9648,N_6439,N_7074);
and U9649 (N_9649,N_7683,N_6550);
nor U9650 (N_9650,N_6560,N_6255);
xnor U9651 (N_9651,N_7463,N_7818);
nand U9652 (N_9652,N_7087,N_7802);
or U9653 (N_9653,N_7406,N_7156);
or U9654 (N_9654,N_6071,N_6324);
or U9655 (N_9655,N_7821,N_6749);
nor U9656 (N_9656,N_7075,N_6525);
nand U9657 (N_9657,N_7122,N_6136);
nor U9658 (N_9658,N_7274,N_6846);
and U9659 (N_9659,N_7067,N_6310);
and U9660 (N_9660,N_7119,N_6290);
or U9661 (N_9661,N_7943,N_6342);
and U9662 (N_9662,N_7559,N_7755);
nand U9663 (N_9663,N_6283,N_6113);
nor U9664 (N_9664,N_6261,N_7928);
nand U9665 (N_9665,N_7895,N_7389);
nor U9666 (N_9666,N_7453,N_7572);
nand U9667 (N_9667,N_6447,N_6516);
nand U9668 (N_9668,N_6282,N_6310);
nand U9669 (N_9669,N_6111,N_6340);
and U9670 (N_9670,N_7653,N_7593);
and U9671 (N_9671,N_6644,N_6098);
xnor U9672 (N_9672,N_7594,N_7838);
nand U9673 (N_9673,N_6040,N_6315);
or U9674 (N_9674,N_6120,N_6028);
nor U9675 (N_9675,N_6358,N_7302);
nor U9676 (N_9676,N_7097,N_7749);
nand U9677 (N_9677,N_6105,N_7453);
xor U9678 (N_9678,N_7890,N_6692);
or U9679 (N_9679,N_7433,N_7115);
or U9680 (N_9680,N_6327,N_6016);
xnor U9681 (N_9681,N_7881,N_6588);
nor U9682 (N_9682,N_6830,N_6602);
nor U9683 (N_9683,N_7180,N_6437);
xor U9684 (N_9684,N_6455,N_7488);
nor U9685 (N_9685,N_7450,N_6069);
xor U9686 (N_9686,N_6276,N_6376);
and U9687 (N_9687,N_6783,N_7138);
and U9688 (N_9688,N_7176,N_6758);
xor U9689 (N_9689,N_6518,N_7426);
xnor U9690 (N_9690,N_6161,N_7464);
nand U9691 (N_9691,N_7789,N_7338);
nand U9692 (N_9692,N_7271,N_6293);
and U9693 (N_9693,N_7177,N_6028);
nand U9694 (N_9694,N_6196,N_7287);
xnor U9695 (N_9695,N_7232,N_6995);
or U9696 (N_9696,N_6802,N_6845);
or U9697 (N_9697,N_7155,N_7434);
nand U9698 (N_9698,N_7972,N_7802);
nand U9699 (N_9699,N_7724,N_7707);
or U9700 (N_9700,N_7921,N_6466);
nor U9701 (N_9701,N_7618,N_6175);
and U9702 (N_9702,N_6498,N_6981);
or U9703 (N_9703,N_6221,N_6154);
or U9704 (N_9704,N_7462,N_7418);
and U9705 (N_9705,N_6147,N_6837);
nor U9706 (N_9706,N_6668,N_7398);
xnor U9707 (N_9707,N_7563,N_6930);
xnor U9708 (N_9708,N_6369,N_6638);
or U9709 (N_9709,N_6482,N_6594);
nor U9710 (N_9710,N_7568,N_7620);
nor U9711 (N_9711,N_6981,N_7597);
and U9712 (N_9712,N_6355,N_7641);
xnor U9713 (N_9713,N_7923,N_6604);
nor U9714 (N_9714,N_7070,N_6681);
nand U9715 (N_9715,N_6716,N_6258);
and U9716 (N_9716,N_7005,N_7802);
and U9717 (N_9717,N_6856,N_7257);
nand U9718 (N_9718,N_6623,N_6905);
nand U9719 (N_9719,N_6653,N_6827);
or U9720 (N_9720,N_7455,N_6170);
and U9721 (N_9721,N_6316,N_6525);
nor U9722 (N_9722,N_6201,N_7430);
and U9723 (N_9723,N_6681,N_7172);
xor U9724 (N_9724,N_7060,N_6675);
nor U9725 (N_9725,N_6256,N_7217);
and U9726 (N_9726,N_7017,N_7780);
or U9727 (N_9727,N_6198,N_7574);
nor U9728 (N_9728,N_7137,N_6065);
nand U9729 (N_9729,N_7654,N_7436);
nor U9730 (N_9730,N_7840,N_7544);
nor U9731 (N_9731,N_6886,N_7819);
or U9732 (N_9732,N_7608,N_7863);
nor U9733 (N_9733,N_6734,N_6745);
xor U9734 (N_9734,N_6250,N_6993);
nand U9735 (N_9735,N_7081,N_7719);
and U9736 (N_9736,N_7371,N_7200);
or U9737 (N_9737,N_6153,N_7380);
and U9738 (N_9738,N_6585,N_6542);
xnor U9739 (N_9739,N_7000,N_6590);
or U9740 (N_9740,N_6384,N_6550);
or U9741 (N_9741,N_7128,N_7320);
and U9742 (N_9742,N_7361,N_7448);
xnor U9743 (N_9743,N_7948,N_6528);
nand U9744 (N_9744,N_6748,N_6134);
nand U9745 (N_9745,N_7520,N_7535);
xnor U9746 (N_9746,N_7487,N_7120);
and U9747 (N_9747,N_6362,N_7470);
or U9748 (N_9748,N_7359,N_6165);
xor U9749 (N_9749,N_6777,N_6248);
or U9750 (N_9750,N_7698,N_7585);
xor U9751 (N_9751,N_7658,N_7355);
nand U9752 (N_9752,N_6938,N_7055);
nor U9753 (N_9753,N_6062,N_7486);
xor U9754 (N_9754,N_7724,N_6545);
nand U9755 (N_9755,N_7542,N_7042);
nand U9756 (N_9756,N_6499,N_6309);
nor U9757 (N_9757,N_6270,N_7701);
and U9758 (N_9758,N_6420,N_6014);
nand U9759 (N_9759,N_7277,N_7011);
and U9760 (N_9760,N_6835,N_7443);
xor U9761 (N_9761,N_7728,N_6698);
xor U9762 (N_9762,N_7641,N_7190);
xnor U9763 (N_9763,N_6812,N_7824);
nand U9764 (N_9764,N_7316,N_6343);
nor U9765 (N_9765,N_7003,N_7391);
xor U9766 (N_9766,N_7723,N_7601);
and U9767 (N_9767,N_6008,N_7311);
or U9768 (N_9768,N_6409,N_7488);
or U9769 (N_9769,N_6923,N_7604);
nor U9770 (N_9770,N_6461,N_6396);
nor U9771 (N_9771,N_6845,N_7881);
nor U9772 (N_9772,N_6574,N_6299);
nor U9773 (N_9773,N_7947,N_7697);
or U9774 (N_9774,N_7215,N_7056);
and U9775 (N_9775,N_7551,N_7337);
and U9776 (N_9776,N_7038,N_7532);
xnor U9777 (N_9777,N_6025,N_7850);
or U9778 (N_9778,N_6028,N_6309);
or U9779 (N_9779,N_7155,N_7997);
xor U9780 (N_9780,N_7579,N_7397);
nor U9781 (N_9781,N_6155,N_7293);
and U9782 (N_9782,N_7512,N_6476);
nor U9783 (N_9783,N_7044,N_7130);
nor U9784 (N_9784,N_6447,N_7351);
and U9785 (N_9785,N_7348,N_7549);
xnor U9786 (N_9786,N_7071,N_6314);
and U9787 (N_9787,N_6581,N_6907);
xor U9788 (N_9788,N_6724,N_6629);
nand U9789 (N_9789,N_6445,N_7679);
xor U9790 (N_9790,N_7374,N_7255);
xnor U9791 (N_9791,N_7855,N_6073);
or U9792 (N_9792,N_6317,N_6717);
and U9793 (N_9793,N_7549,N_6559);
nor U9794 (N_9794,N_7962,N_7228);
or U9795 (N_9795,N_6319,N_7867);
nor U9796 (N_9796,N_7894,N_6566);
and U9797 (N_9797,N_7248,N_7512);
and U9798 (N_9798,N_6112,N_7275);
and U9799 (N_9799,N_7064,N_6156);
or U9800 (N_9800,N_7128,N_7558);
or U9801 (N_9801,N_7057,N_6314);
nor U9802 (N_9802,N_6530,N_7557);
nor U9803 (N_9803,N_7120,N_7216);
or U9804 (N_9804,N_7282,N_6790);
nor U9805 (N_9805,N_7065,N_7173);
nand U9806 (N_9806,N_7355,N_6198);
xnor U9807 (N_9807,N_6005,N_6684);
xor U9808 (N_9808,N_7956,N_6337);
or U9809 (N_9809,N_7655,N_7259);
xnor U9810 (N_9810,N_7171,N_6418);
or U9811 (N_9811,N_6581,N_7042);
nand U9812 (N_9812,N_6912,N_6539);
or U9813 (N_9813,N_6117,N_7948);
or U9814 (N_9814,N_7945,N_6956);
or U9815 (N_9815,N_7539,N_7323);
nor U9816 (N_9816,N_6912,N_6226);
xnor U9817 (N_9817,N_6341,N_6235);
and U9818 (N_9818,N_7953,N_7091);
nand U9819 (N_9819,N_6368,N_7226);
nand U9820 (N_9820,N_6179,N_7257);
xnor U9821 (N_9821,N_6958,N_7971);
or U9822 (N_9822,N_6313,N_7955);
and U9823 (N_9823,N_7569,N_6921);
or U9824 (N_9824,N_7884,N_7482);
nand U9825 (N_9825,N_7687,N_7435);
xnor U9826 (N_9826,N_6246,N_7791);
xor U9827 (N_9827,N_6270,N_7827);
nor U9828 (N_9828,N_6980,N_6401);
nand U9829 (N_9829,N_6131,N_7819);
nor U9830 (N_9830,N_7070,N_6073);
nor U9831 (N_9831,N_7416,N_6960);
nor U9832 (N_9832,N_7337,N_7432);
xor U9833 (N_9833,N_7604,N_6548);
and U9834 (N_9834,N_7348,N_7358);
or U9835 (N_9835,N_7734,N_6059);
and U9836 (N_9836,N_6027,N_6769);
nor U9837 (N_9837,N_7999,N_7586);
or U9838 (N_9838,N_6457,N_6298);
or U9839 (N_9839,N_7103,N_7306);
nor U9840 (N_9840,N_6443,N_6181);
xnor U9841 (N_9841,N_7952,N_6359);
xor U9842 (N_9842,N_6844,N_6373);
and U9843 (N_9843,N_6225,N_6533);
nor U9844 (N_9844,N_7816,N_7070);
or U9845 (N_9845,N_6824,N_6718);
and U9846 (N_9846,N_6416,N_7176);
or U9847 (N_9847,N_6613,N_7252);
xnor U9848 (N_9848,N_7720,N_7952);
or U9849 (N_9849,N_7744,N_7860);
and U9850 (N_9850,N_6208,N_7228);
nor U9851 (N_9851,N_6567,N_7180);
nand U9852 (N_9852,N_6749,N_6652);
and U9853 (N_9853,N_7089,N_7446);
xnor U9854 (N_9854,N_6916,N_6907);
or U9855 (N_9855,N_7155,N_7020);
nor U9856 (N_9856,N_7356,N_6145);
nor U9857 (N_9857,N_6808,N_6725);
nor U9858 (N_9858,N_6809,N_6617);
and U9859 (N_9859,N_7185,N_6407);
nand U9860 (N_9860,N_7208,N_7534);
and U9861 (N_9861,N_7819,N_6597);
or U9862 (N_9862,N_7248,N_6900);
xor U9863 (N_9863,N_7654,N_7573);
or U9864 (N_9864,N_7263,N_7553);
and U9865 (N_9865,N_7756,N_6506);
or U9866 (N_9866,N_6236,N_7965);
xnor U9867 (N_9867,N_7283,N_6735);
and U9868 (N_9868,N_6695,N_6875);
xor U9869 (N_9869,N_7860,N_7669);
or U9870 (N_9870,N_6915,N_7791);
nor U9871 (N_9871,N_6117,N_7839);
or U9872 (N_9872,N_6728,N_7056);
nand U9873 (N_9873,N_6049,N_7687);
nor U9874 (N_9874,N_6421,N_6273);
xor U9875 (N_9875,N_7480,N_7135);
xor U9876 (N_9876,N_6855,N_6387);
and U9877 (N_9877,N_6566,N_7615);
or U9878 (N_9878,N_6690,N_7009);
xnor U9879 (N_9879,N_7126,N_6135);
nor U9880 (N_9880,N_7032,N_6685);
xnor U9881 (N_9881,N_6138,N_6379);
or U9882 (N_9882,N_6873,N_7348);
or U9883 (N_9883,N_7912,N_7459);
xor U9884 (N_9884,N_6884,N_6701);
xor U9885 (N_9885,N_7516,N_6998);
and U9886 (N_9886,N_7016,N_6072);
nand U9887 (N_9887,N_7629,N_6418);
and U9888 (N_9888,N_7747,N_7410);
xnor U9889 (N_9889,N_6234,N_7397);
nand U9890 (N_9890,N_7590,N_7399);
nor U9891 (N_9891,N_6193,N_7250);
nor U9892 (N_9892,N_6529,N_6789);
and U9893 (N_9893,N_6011,N_6146);
and U9894 (N_9894,N_7451,N_6982);
xnor U9895 (N_9895,N_6788,N_6892);
xor U9896 (N_9896,N_7999,N_7783);
nor U9897 (N_9897,N_7420,N_6309);
nand U9898 (N_9898,N_7825,N_7614);
xor U9899 (N_9899,N_6094,N_7410);
or U9900 (N_9900,N_6045,N_6441);
xnor U9901 (N_9901,N_7392,N_7894);
nor U9902 (N_9902,N_7347,N_7602);
nand U9903 (N_9903,N_6340,N_6902);
and U9904 (N_9904,N_6263,N_6792);
nand U9905 (N_9905,N_6269,N_7412);
and U9906 (N_9906,N_7758,N_6728);
and U9907 (N_9907,N_6378,N_6355);
or U9908 (N_9908,N_6824,N_6055);
nor U9909 (N_9909,N_7083,N_7391);
nor U9910 (N_9910,N_6273,N_7728);
and U9911 (N_9911,N_7359,N_7516);
or U9912 (N_9912,N_7870,N_7705);
and U9913 (N_9913,N_6847,N_6999);
or U9914 (N_9914,N_7096,N_6014);
nor U9915 (N_9915,N_7084,N_6925);
xnor U9916 (N_9916,N_6463,N_6732);
nor U9917 (N_9917,N_6119,N_6576);
and U9918 (N_9918,N_7751,N_7634);
nand U9919 (N_9919,N_6693,N_6584);
nand U9920 (N_9920,N_6074,N_6771);
nor U9921 (N_9921,N_6293,N_7723);
nand U9922 (N_9922,N_7240,N_7364);
and U9923 (N_9923,N_7638,N_7696);
nand U9924 (N_9924,N_6485,N_7136);
and U9925 (N_9925,N_7479,N_7558);
or U9926 (N_9926,N_7501,N_7834);
nand U9927 (N_9927,N_7604,N_7776);
xor U9928 (N_9928,N_6734,N_7780);
xor U9929 (N_9929,N_6978,N_7292);
and U9930 (N_9930,N_6541,N_7220);
nand U9931 (N_9931,N_6143,N_7882);
or U9932 (N_9932,N_7636,N_7226);
and U9933 (N_9933,N_6621,N_7489);
xnor U9934 (N_9934,N_7734,N_6264);
and U9935 (N_9935,N_7583,N_6629);
or U9936 (N_9936,N_6005,N_6346);
xor U9937 (N_9937,N_6233,N_6443);
xor U9938 (N_9938,N_6146,N_7692);
nand U9939 (N_9939,N_6525,N_7948);
nor U9940 (N_9940,N_7160,N_7445);
nor U9941 (N_9941,N_7788,N_7371);
or U9942 (N_9942,N_6766,N_7156);
and U9943 (N_9943,N_6519,N_7034);
and U9944 (N_9944,N_6120,N_6566);
nor U9945 (N_9945,N_6355,N_6517);
and U9946 (N_9946,N_7453,N_7058);
nand U9947 (N_9947,N_6502,N_7411);
xnor U9948 (N_9948,N_6872,N_6563);
xor U9949 (N_9949,N_7142,N_6097);
nand U9950 (N_9950,N_6682,N_7494);
nor U9951 (N_9951,N_7335,N_7100);
or U9952 (N_9952,N_6970,N_7849);
or U9953 (N_9953,N_6002,N_6901);
nand U9954 (N_9954,N_6930,N_6196);
nor U9955 (N_9955,N_7923,N_6860);
and U9956 (N_9956,N_6611,N_6996);
nor U9957 (N_9957,N_7531,N_6788);
xnor U9958 (N_9958,N_6793,N_6919);
or U9959 (N_9959,N_6331,N_6886);
or U9960 (N_9960,N_7763,N_7556);
nor U9961 (N_9961,N_6835,N_7948);
nand U9962 (N_9962,N_7215,N_7247);
nor U9963 (N_9963,N_7205,N_7892);
or U9964 (N_9964,N_7396,N_6797);
or U9965 (N_9965,N_7912,N_7240);
xor U9966 (N_9966,N_6102,N_7187);
nand U9967 (N_9967,N_7159,N_7578);
nor U9968 (N_9968,N_7142,N_7839);
and U9969 (N_9969,N_6984,N_6230);
and U9970 (N_9970,N_7591,N_7149);
and U9971 (N_9971,N_6848,N_6061);
xnor U9972 (N_9972,N_6922,N_7912);
nor U9973 (N_9973,N_7173,N_7262);
xor U9974 (N_9974,N_7022,N_6911);
nor U9975 (N_9975,N_7555,N_6924);
nor U9976 (N_9976,N_6445,N_6579);
and U9977 (N_9977,N_7932,N_6752);
xnor U9978 (N_9978,N_7448,N_6363);
xnor U9979 (N_9979,N_7564,N_7906);
and U9980 (N_9980,N_7470,N_7673);
xnor U9981 (N_9981,N_6955,N_7910);
and U9982 (N_9982,N_7883,N_6676);
and U9983 (N_9983,N_7455,N_7091);
nand U9984 (N_9984,N_6119,N_6406);
and U9985 (N_9985,N_6430,N_7910);
nor U9986 (N_9986,N_6315,N_7337);
or U9987 (N_9987,N_6422,N_7252);
xnor U9988 (N_9988,N_7497,N_7463);
xor U9989 (N_9989,N_6395,N_6997);
nor U9990 (N_9990,N_6959,N_6083);
or U9991 (N_9991,N_6132,N_7417);
or U9992 (N_9992,N_6818,N_7576);
or U9993 (N_9993,N_6529,N_6913);
nand U9994 (N_9994,N_7045,N_6505);
nor U9995 (N_9995,N_7201,N_7444);
and U9996 (N_9996,N_6596,N_7534);
xnor U9997 (N_9997,N_6712,N_7772);
nand U9998 (N_9998,N_6977,N_7598);
nor U9999 (N_9999,N_6531,N_7158);
nor U10000 (N_10000,N_8268,N_9153);
or U10001 (N_10001,N_9352,N_8732);
and U10002 (N_10002,N_8960,N_8610);
and U10003 (N_10003,N_9090,N_9560);
and U10004 (N_10004,N_9821,N_9020);
xor U10005 (N_10005,N_9624,N_9377);
or U10006 (N_10006,N_9540,N_8481);
nor U10007 (N_10007,N_8194,N_9067);
nand U10008 (N_10008,N_9158,N_9634);
xnor U10009 (N_10009,N_8290,N_8835);
xnor U10010 (N_10010,N_9093,N_8172);
nor U10011 (N_10011,N_9263,N_9165);
or U10012 (N_10012,N_9446,N_8328);
or U10013 (N_10013,N_8095,N_8152);
nor U10014 (N_10014,N_9072,N_9187);
nand U10015 (N_10015,N_9959,N_9735);
and U10016 (N_10016,N_9648,N_8629);
nand U10017 (N_10017,N_8027,N_9291);
nand U10018 (N_10018,N_8797,N_9194);
or U10019 (N_10019,N_9611,N_9572);
or U10020 (N_10020,N_9069,N_8887);
or U10021 (N_10021,N_9864,N_9315);
or U10022 (N_10022,N_8740,N_9450);
nand U10023 (N_10023,N_9508,N_9924);
xor U10024 (N_10024,N_8421,N_8825);
nor U10025 (N_10025,N_9643,N_9167);
xnor U10026 (N_10026,N_8382,N_8641);
or U10027 (N_10027,N_9743,N_9030);
or U10028 (N_10028,N_8227,N_9038);
xnor U10029 (N_10029,N_9405,N_9454);
xor U10030 (N_10030,N_8489,N_8961);
nor U10031 (N_10031,N_8682,N_9596);
nor U10032 (N_10032,N_8075,N_8858);
and U10033 (N_10033,N_9637,N_8883);
and U10034 (N_10034,N_9497,N_8602);
and U10035 (N_10035,N_8153,N_9860);
or U10036 (N_10036,N_9827,N_8369);
and U10037 (N_10037,N_8265,N_8549);
xnor U10038 (N_10038,N_8403,N_9235);
xor U10039 (N_10039,N_9185,N_8730);
nand U10040 (N_10040,N_9073,N_9314);
and U10041 (N_10041,N_9669,N_8561);
nand U10042 (N_10042,N_9991,N_8218);
or U10043 (N_10043,N_9773,N_8266);
nor U10044 (N_10044,N_9685,N_8427);
xnor U10045 (N_10045,N_8673,N_9408);
or U10046 (N_10046,N_8762,N_8007);
nor U10047 (N_10047,N_8892,N_9488);
nor U10048 (N_10048,N_8243,N_9296);
nor U10049 (N_10049,N_9018,N_9653);
or U10050 (N_10050,N_9028,N_8263);
or U10051 (N_10051,N_9471,N_9892);
nor U10052 (N_10052,N_8923,N_9802);
nand U10053 (N_10053,N_9299,N_8217);
nand U10054 (N_10054,N_9032,N_8687);
and U10055 (N_10055,N_8970,N_9851);
xnor U10056 (N_10056,N_8969,N_9628);
or U10057 (N_10057,N_9337,N_9831);
xor U10058 (N_10058,N_8046,N_8792);
and U10059 (N_10059,N_8898,N_9681);
nor U10060 (N_10060,N_9520,N_9172);
nor U10061 (N_10061,N_8963,N_9576);
or U10062 (N_10062,N_8213,N_9799);
nand U10063 (N_10063,N_8800,N_8073);
nand U10064 (N_10064,N_8251,N_9253);
nor U10065 (N_10065,N_9380,N_9974);
xor U10066 (N_10066,N_8336,N_8259);
and U10067 (N_10067,N_9753,N_9651);
xor U10068 (N_10068,N_9922,N_9320);
nor U10069 (N_10069,N_9761,N_8175);
nand U10070 (N_10070,N_8933,N_8911);
nor U10071 (N_10071,N_8004,N_8181);
nand U10072 (N_10072,N_8434,N_9988);
or U10073 (N_10073,N_8138,N_8493);
xor U10074 (N_10074,N_8889,N_9638);
or U10075 (N_10075,N_8498,N_9074);
xor U10076 (N_10076,N_9688,N_9356);
and U10077 (N_10077,N_8768,N_9720);
and U10078 (N_10078,N_8927,N_8613);
nand U10079 (N_10079,N_8658,N_9837);
and U10080 (N_10080,N_9041,N_9117);
and U10081 (N_10081,N_8020,N_9661);
nand U10082 (N_10082,N_9191,N_9723);
nor U10083 (N_10083,N_9714,N_8793);
or U10084 (N_10084,N_8398,N_8503);
or U10085 (N_10085,N_9986,N_9911);
nor U10086 (N_10086,N_9566,N_8234);
nor U10087 (N_10087,N_8519,N_9905);
xor U10088 (N_10088,N_9290,N_8601);
nor U10089 (N_10089,N_9332,N_9123);
nand U10090 (N_10090,N_9822,N_8627);
nand U10091 (N_10091,N_8743,N_8529);
nor U10092 (N_10092,N_9607,N_9049);
nand U10093 (N_10093,N_8026,N_9774);
nor U10094 (N_10094,N_8537,N_8592);
and U10095 (N_10095,N_9573,N_8860);
nand U10096 (N_10096,N_8867,N_8907);
xor U10097 (N_10097,N_8338,N_9783);
nor U10098 (N_10098,N_9920,N_8484);
xnor U10099 (N_10099,N_8494,N_9690);
or U10100 (N_10100,N_9644,N_8813);
nor U10101 (N_10101,N_9978,N_9729);
or U10102 (N_10102,N_8558,N_9420);
nand U10103 (N_10103,N_9963,N_9391);
and U10104 (N_10104,N_8286,N_8754);
xnor U10105 (N_10105,N_8299,N_8291);
and U10106 (N_10106,N_9278,N_8106);
or U10107 (N_10107,N_9858,N_9138);
nor U10108 (N_10108,N_9015,N_9431);
nor U10109 (N_10109,N_9283,N_9602);
xnor U10110 (N_10110,N_8738,N_8876);
or U10111 (N_10111,N_8201,N_8991);
nor U10112 (N_10112,N_9843,N_8163);
xor U10113 (N_10113,N_8061,N_8639);
nand U10114 (N_10114,N_8567,N_8551);
and U10115 (N_10115,N_8716,N_9173);
and U10116 (N_10116,N_8147,N_9186);
or U10117 (N_10117,N_9812,N_9141);
and U10118 (N_10118,N_9294,N_8032);
and U10119 (N_10119,N_8984,N_8986);
or U10120 (N_10120,N_9594,N_9734);
xor U10121 (N_10121,N_9965,N_8118);
and U10122 (N_10122,N_8424,N_9244);
nor U10123 (N_10123,N_9946,N_8302);
xor U10124 (N_10124,N_8916,N_8304);
or U10125 (N_10125,N_8246,N_8553);
or U10126 (N_10126,N_8344,N_9042);
or U10127 (N_10127,N_9150,N_8736);
and U10128 (N_10128,N_8452,N_8620);
and U10129 (N_10129,N_8968,N_8456);
and U10130 (N_10130,N_9239,N_8919);
and U10131 (N_10131,N_8226,N_8733);
or U10132 (N_10132,N_8901,N_9108);
nor U10133 (N_10133,N_8411,N_9234);
nor U10134 (N_10134,N_9999,N_8895);
or U10135 (N_10135,N_9070,N_9895);
nand U10136 (N_10136,N_9993,N_9503);
xor U10137 (N_10137,N_9209,N_8185);
or U10138 (N_10138,N_8414,N_9045);
and U10139 (N_10139,N_8642,N_8113);
nor U10140 (N_10140,N_9262,N_9867);
and U10141 (N_10141,N_8440,N_8453);
and U10142 (N_10142,N_9137,N_8590);
xnor U10143 (N_10143,N_8647,N_8830);
xor U10144 (N_10144,N_9417,N_9749);
and U10145 (N_10145,N_8461,N_8231);
nor U10146 (N_10146,N_8050,N_8495);
xor U10147 (N_10147,N_8022,N_8996);
nor U10148 (N_10148,N_8978,N_9306);
or U10149 (N_10149,N_8011,N_9793);
xor U10150 (N_10150,N_9601,N_8047);
and U10151 (N_10151,N_9427,N_9094);
xnor U10152 (N_10152,N_9163,N_9495);
or U10153 (N_10153,N_8972,N_8446);
and U10154 (N_10154,N_9053,N_9449);
nand U10155 (N_10155,N_8973,N_8232);
nand U10156 (N_10156,N_9726,N_8509);
xor U10157 (N_10157,N_9679,N_9258);
nor U10158 (N_10158,N_8976,N_8038);
xnor U10159 (N_10159,N_9517,N_8086);
and U10160 (N_10160,N_9059,N_9511);
xnor U10161 (N_10161,N_8904,N_9272);
and U10162 (N_10162,N_8184,N_8831);
or U10163 (N_10163,N_9221,N_8807);
nor U10164 (N_10164,N_8315,N_8584);
xor U10165 (N_10165,N_8524,N_8873);
nand U10166 (N_10166,N_8173,N_8925);
or U10167 (N_10167,N_8532,N_9562);
nor U10168 (N_10168,N_8855,N_8404);
xor U10169 (N_10169,N_9586,N_8870);
or U10170 (N_10170,N_8186,N_9412);
or U10171 (N_10171,N_9918,N_9433);
and U10172 (N_10172,N_8838,N_9887);
or U10173 (N_10173,N_8205,N_9797);
xnor U10174 (N_10174,N_8099,N_8997);
and U10175 (N_10175,N_8428,N_9640);
and U10176 (N_10176,N_9788,N_9604);
or U10177 (N_10177,N_9512,N_8757);
or U10178 (N_10178,N_9621,N_8849);
xor U10179 (N_10179,N_9178,N_8745);
xnor U10180 (N_10180,N_9482,N_8527);
or U10181 (N_10181,N_8284,N_9614);
nor U10182 (N_10182,N_8300,N_8965);
xnor U10183 (N_10183,N_8264,N_8008);
and U10184 (N_10184,N_9410,N_9409);
or U10185 (N_10185,N_9204,N_9456);
xnor U10186 (N_10186,N_8024,N_8628);
or U10187 (N_10187,N_9225,N_9565);
and U10188 (N_10188,N_8706,N_9809);
and U10189 (N_10189,N_8985,N_9063);
nor U10190 (N_10190,N_8891,N_8164);
nor U10191 (N_10191,N_8822,N_9370);
nand U10192 (N_10192,N_9019,N_9981);
xnor U10193 (N_10193,N_9366,N_8115);
and U10194 (N_10194,N_8668,N_9666);
nor U10195 (N_10195,N_8517,N_9645);
nor U10196 (N_10196,N_9987,N_9099);
xor U10197 (N_10197,N_8789,N_9092);
xor U10198 (N_10198,N_8848,N_9131);
and U10199 (N_10199,N_9956,N_8770);
or U10200 (N_10200,N_8202,N_9457);
nor U10201 (N_10201,N_9564,N_8696);
xor U10202 (N_10202,N_9779,N_8671);
nor U10203 (N_10203,N_8018,N_8777);
and U10204 (N_10204,N_8079,N_8749);
nor U10205 (N_10205,N_9961,N_8123);
nand U10206 (N_10206,N_8223,N_9804);
and U10207 (N_10207,N_9780,N_8857);
xor U10208 (N_10208,N_9140,N_8649);
nor U10209 (N_10209,N_8017,N_9658);
or U10210 (N_10210,N_9071,N_8563);
nor U10211 (N_10211,N_8827,N_8943);
nor U10212 (N_10212,N_8541,N_8015);
nand U10213 (N_10213,N_9494,N_8323);
nand U10214 (N_10214,N_9750,N_8094);
or U10215 (N_10215,N_9989,N_8330);
or U10216 (N_10216,N_9732,N_8121);
xnor U10217 (N_10217,N_8168,N_9861);
nand U10218 (N_10218,N_9436,N_8272);
nand U10219 (N_10219,N_9309,N_8980);
nand U10220 (N_10220,N_9526,N_8611);
or U10221 (N_10221,N_9011,N_9311);
nor U10222 (N_10222,N_8297,N_8759);
nand U10223 (N_10223,N_8374,N_8235);
or U10224 (N_10224,N_8786,N_9098);
xnor U10225 (N_10225,N_8318,N_9208);
and U10226 (N_10226,N_9746,N_9817);
and U10227 (N_10227,N_9012,N_8699);
and U10228 (N_10228,N_8245,N_8307);
and U10229 (N_10229,N_9724,N_9663);
xor U10230 (N_10230,N_9033,N_9084);
xor U10231 (N_10231,N_9334,N_9075);
xnor U10232 (N_10232,N_9901,N_8847);
nand U10233 (N_10233,N_9752,N_9992);
and U10234 (N_10234,N_8132,N_8871);
nor U10235 (N_10235,N_9917,N_8994);
xnor U10236 (N_10236,N_9792,N_8693);
nor U10237 (N_10237,N_9659,N_8037);
nor U10238 (N_10238,N_9857,N_8387);
nand U10239 (N_10239,N_8937,N_9480);
nand U10240 (N_10240,N_9154,N_9673);
xor U10241 (N_10241,N_8347,N_8215);
nor U10242 (N_10242,N_8210,N_8229);
and U10243 (N_10243,N_8853,N_9313);
xor U10244 (N_10244,N_9678,N_8882);
nand U10245 (N_10245,N_9806,N_8005);
nor U10246 (N_10246,N_9671,N_9894);
nor U10247 (N_10247,N_9183,N_8310);
xor U10248 (N_10248,N_8479,N_8788);
nor U10249 (N_10249,N_8337,N_8364);
or U10250 (N_10250,N_9122,N_9630);
xnor U10251 (N_10251,N_9631,N_8169);
and U10252 (N_10252,N_9719,N_8400);
nor U10253 (N_10253,N_9425,N_9079);
and U10254 (N_10254,N_9318,N_8543);
or U10255 (N_10255,N_9738,N_8363);
and U10256 (N_10256,N_9979,N_8619);
nand U10257 (N_10257,N_9514,N_8460);
and U10258 (N_10258,N_8936,N_9504);
and U10259 (N_10259,N_9603,N_8220);
nand U10260 (N_10260,N_8995,N_8345);
nand U10261 (N_10261,N_9836,N_8091);
or U10262 (N_10262,N_9826,N_8145);
and U10263 (N_10263,N_8309,N_9364);
or U10264 (N_10264,N_8652,N_8396);
nor U10265 (N_10265,N_8864,N_8728);
xnor U10266 (N_10266,N_8033,N_9910);
and U10267 (N_10267,N_8683,N_9899);
xor U10268 (N_10268,N_9995,N_8760);
nor U10269 (N_10269,N_9051,N_8957);
or U10270 (N_10270,N_8114,N_9196);
and U10271 (N_10271,N_8540,N_8116);
nor U10272 (N_10272,N_9710,N_9013);
and U10273 (N_10273,N_9725,N_8029);
or U10274 (N_10274,N_9037,N_9932);
nor U10275 (N_10275,N_8816,N_8780);
nand U10276 (N_10276,N_9442,N_8081);
or U10277 (N_10277,N_8149,N_9257);
and U10278 (N_10278,N_8426,N_8093);
and U10279 (N_10279,N_9375,N_9636);
and U10280 (N_10280,N_8964,N_9950);
nor U10281 (N_10281,N_8470,N_8502);
or U10282 (N_10282,N_9229,N_9745);
nand U10283 (N_10283,N_9938,N_9810);
xnor U10284 (N_10284,N_9009,N_8052);
and U10285 (N_10285,N_8921,N_8270);
nand U10286 (N_10286,N_9324,N_9119);
xnor U10287 (N_10287,N_8763,N_9579);
or U10288 (N_10288,N_8260,N_9374);
xnor U10289 (N_10289,N_8276,N_9429);
nand U10290 (N_10290,N_9730,N_8370);
nand U10291 (N_10291,N_8097,N_8392);
nand U10292 (N_10292,N_8438,N_9023);
or U10293 (N_10293,N_8715,N_8962);
or U10294 (N_10294,N_8448,N_9365);
nand U10295 (N_10295,N_8562,N_8277);
xnor U10296 (N_10296,N_8311,N_8665);
xnor U10297 (N_10297,N_8166,N_8914);
and U10298 (N_10298,N_9944,N_8874);
nand U10299 (N_10299,N_9414,N_9468);
nor U10300 (N_10300,N_8319,N_9518);
or U10301 (N_10301,N_9884,N_8485);
or U10302 (N_10302,N_8579,N_9955);
nor U10303 (N_10303,N_9006,N_8817);
xor U10304 (N_10304,N_8274,N_8934);
xor U10305 (N_10305,N_9852,N_8836);
nor U10306 (N_10306,N_9578,N_9316);
nor U10307 (N_10307,N_8454,N_8912);
or U10308 (N_10308,N_8607,N_9966);
and U10309 (N_10309,N_9873,N_9325);
and U10310 (N_10310,N_8941,N_9040);
xor U10311 (N_10311,N_8525,N_8488);
and U10312 (N_10312,N_8950,N_9862);
nand U10313 (N_10313,N_9105,N_8557);
or U10314 (N_10314,N_9542,N_8308);
nand U10315 (N_10315,N_9559,N_8684);
and U10316 (N_10316,N_8059,N_9271);
nor U10317 (N_10317,N_8285,N_9904);
nand U10318 (N_10318,N_8935,N_9699);
xor U10319 (N_10319,N_9328,N_9189);
xor U10320 (N_10320,N_8672,N_8365);
nand U10321 (N_10321,N_8397,N_9242);
nor U10322 (N_10322,N_9491,N_9650);
nand U10323 (N_10323,N_8077,N_8784);
nor U10324 (N_10324,N_8151,N_8248);
or U10325 (N_10325,N_8704,N_8449);
or U10326 (N_10326,N_9385,N_8362);
nor U10327 (N_10327,N_9236,N_8262);
nand U10328 (N_10328,N_9487,N_8894);
nand U10329 (N_10329,N_8180,N_8124);
nor U10330 (N_10330,N_8069,N_9419);
nand U10331 (N_10331,N_8664,N_9421);
or U10332 (N_10332,N_8395,N_9129);
nand U10333 (N_10333,N_8866,N_8942);
and U10334 (N_10334,N_8595,N_8306);
or U10335 (N_10335,N_9548,N_9740);
or U10336 (N_10336,N_9536,N_9344);
xor U10337 (N_10337,N_9458,N_8320);
or U10338 (N_10338,N_9898,N_9200);
xor U10339 (N_10339,N_8134,N_9025);
and U10340 (N_10340,N_8071,N_9192);
or U10341 (N_10341,N_8289,N_8688);
nor U10342 (N_10342,N_9933,N_8522);
or U10343 (N_10343,N_9855,N_9358);
nor U10344 (N_10344,N_9849,N_9936);
and U10345 (N_10345,N_8242,N_9139);
nor U10346 (N_10346,N_9971,N_8966);
and U10347 (N_10347,N_9934,N_8615);
or U10348 (N_10348,N_8843,N_8303);
nor U10349 (N_10349,N_8513,N_9622);
nand U10350 (N_10350,N_8572,N_8820);
and U10351 (N_10351,N_8842,N_9581);
nor U10352 (N_10352,N_8025,N_8305);
or U10353 (N_10353,N_8998,N_9064);
or U10354 (N_10354,N_9289,N_8482);
nor U10355 (N_10355,N_9307,N_8516);
nor U10356 (N_10356,N_8500,N_8236);
or U10357 (N_10357,N_9055,N_9201);
and U10358 (N_10358,N_8694,N_8083);
nand U10359 (N_10359,N_9940,N_9465);
or U10360 (N_10360,N_8467,N_8954);
and U10361 (N_10361,N_9177,N_8491);
xor U10362 (N_10362,N_8811,N_8146);
and U10363 (N_10363,N_8352,N_9171);
or U10364 (N_10364,N_8556,N_9954);
xnor U10365 (N_10365,N_9452,N_8806);
and U10366 (N_10366,N_8252,N_9760);
nand U10367 (N_10367,N_8103,N_8361);
xnor U10368 (N_10368,N_8617,N_8293);
nor U10369 (N_10369,N_9169,N_9583);
nand U10370 (N_10370,N_9285,N_8885);
nor U10371 (N_10371,N_8512,N_8774);
and U10372 (N_10372,N_8486,N_8131);
and U10373 (N_10373,N_8711,N_8766);
and U10374 (N_10374,N_9001,N_9655);
nor U10375 (N_10375,N_8003,N_8437);
nor U10376 (N_10376,N_9460,N_8295);
and U10377 (N_10377,N_8926,N_9437);
xor U10378 (N_10378,N_9247,N_9813);
or U10379 (N_10379,N_8021,N_8707);
xnor U10380 (N_10380,N_9923,N_8433);
nand U10381 (N_10381,N_9880,N_9046);
xnor U10382 (N_10382,N_8141,N_8214);
xor U10383 (N_10383,N_9859,N_8267);
xnor U10384 (N_10384,N_9128,N_9692);
and U10385 (N_10385,N_8385,N_9403);
nor U10386 (N_10386,N_9909,N_9967);
and U10387 (N_10387,N_9453,N_9463);
nor U10388 (N_10388,N_9764,N_9915);
nor U10389 (N_10389,N_9372,N_9657);
or U10390 (N_10390,N_8193,N_9990);
nand U10391 (N_10391,N_9083,N_8769);
xor U10392 (N_10392,N_8288,N_9885);
and U10393 (N_10393,N_9287,N_8974);
nor U10394 (N_10394,N_9392,N_8700);
or U10395 (N_10395,N_8312,N_9284);
nand U10396 (N_10396,N_9275,N_8729);
xor U10397 (N_10397,N_9543,N_9769);
xor U10398 (N_10398,N_8862,N_8959);
nor U10399 (N_10399,N_9615,N_9903);
xnor U10400 (N_10400,N_8377,N_9230);
nor U10401 (N_10401,N_9619,N_9585);
or U10402 (N_10402,N_9396,N_8062);
and U10403 (N_10403,N_8501,N_9255);
xnor U10404 (N_10404,N_8313,N_9882);
nor U10405 (N_10405,N_8955,N_9478);
xnor U10406 (N_10406,N_8531,N_9026);
or U10407 (N_10407,N_8135,N_9082);
and U10408 (N_10408,N_9350,N_8971);
nor U10409 (N_10409,N_8329,N_8677);
xor U10410 (N_10410,N_8367,N_9606);
and U10411 (N_10411,N_9635,N_8987);
or U10412 (N_10412,N_9510,N_8508);
and U10413 (N_10413,N_8975,N_8321);
nand U10414 (N_10414,N_9097,N_8063);
nand U10415 (N_10415,N_8890,N_8042);
and U10416 (N_10416,N_9676,N_8076);
xor U10417 (N_10417,N_9820,N_8435);
nand U10418 (N_10418,N_8977,N_9238);
nand U10419 (N_10419,N_9202,N_9451);
or U10420 (N_10420,N_9913,N_8657);
nand U10421 (N_10421,N_8566,N_8040);
xor U10422 (N_10422,N_9840,N_8476);
nor U10423 (N_10423,N_8144,N_9223);
xor U10424 (N_10424,N_9387,N_9665);
xnor U10425 (N_10425,N_8165,N_8221);
xnor U10426 (N_10426,N_9144,N_8967);
nor U10427 (N_10427,N_8167,N_9116);
xor U10428 (N_10428,N_9700,N_8384);
and U10429 (N_10429,N_9664,N_9312);
or U10430 (N_10430,N_9524,N_8280);
or U10431 (N_10431,N_9516,N_9184);
and U10432 (N_10432,N_8691,N_9698);
and U10433 (N_10433,N_9142,N_9741);
nor U10434 (N_10434,N_8474,N_9632);
nand U10435 (N_10435,N_9672,N_9948);
nand U10436 (N_10436,N_8938,N_9689);
and U10437 (N_10437,N_9340,N_8350);
xor U10438 (N_10438,N_8717,N_9212);
xor U10439 (N_10439,N_8981,N_9853);
nand U10440 (N_10440,N_9462,N_8143);
nand U10441 (N_10441,N_8638,N_9343);
xnor U10442 (N_10442,N_8599,N_9633);
xnor U10443 (N_10443,N_8989,N_9771);
or U10444 (N_10444,N_8724,N_8709);
or U10445 (N_10445,N_9347,N_9589);
or U10446 (N_10446,N_8356,N_9975);
xnor U10447 (N_10447,N_9713,N_8102);
nor U10448 (N_10448,N_9742,N_9569);
xor U10449 (N_10449,N_8204,N_9521);
nor U10450 (N_10450,N_8982,N_8695);
or U10451 (N_10451,N_9856,N_8662);
nor U10452 (N_10452,N_8358,N_9757);
and U10453 (N_10453,N_9014,N_9155);
xor U10454 (N_10454,N_8399,N_8378);
nand U10455 (N_10455,N_9527,N_8101);
xor U10456 (N_10456,N_9850,N_9969);
and U10457 (N_10457,N_9121,N_8472);
and U10458 (N_10458,N_8908,N_9426);
nor U10459 (N_10459,N_9702,N_8910);
or U10460 (N_10460,N_9246,N_9345);
nand U10461 (N_10461,N_9393,N_8571);
nor U10462 (N_10462,N_9428,N_9149);
or U10463 (N_10463,N_8394,N_8580);
or U10464 (N_10464,N_9134,N_9088);
and U10465 (N_10465,N_9870,N_8576);
and U10466 (N_10466,N_8681,N_8692);
nor U10467 (N_10467,N_9866,N_9438);
nor U10468 (N_10468,N_8741,N_9228);
and U10469 (N_10469,N_9830,N_8869);
and U10470 (N_10470,N_9373,N_9383);
or U10471 (N_10471,N_8130,N_8030);
nand U10472 (N_10472,N_8407,N_8758);
and U10473 (N_10473,N_8000,N_9662);
or U10474 (N_10474,N_9519,N_8471);
nand U10475 (N_10475,N_8253,N_8366);
xor U10476 (N_10476,N_9835,N_9101);
or U10477 (N_10477,N_9381,N_9422);
and U10478 (N_10478,N_9709,N_8212);
xor U10479 (N_10479,N_9647,N_9441);
xnor U10480 (N_10480,N_8814,N_8155);
xnor U10481 (N_10481,N_8603,N_9361);
xor U10482 (N_10482,N_9027,N_8176);
and U10483 (N_10483,N_8057,N_8171);
or U10484 (N_10484,N_8316,N_9925);
xor U10485 (N_10485,N_9605,N_8339);
nor U10486 (N_10486,N_9513,N_8612);
or U10487 (N_10487,N_9962,N_9863);
xor U10488 (N_10488,N_9411,N_9776);
xor U10489 (N_10489,N_8355,N_8719);
nor U10490 (N_10490,N_8783,N_8346);
or U10491 (N_10491,N_8298,N_8012);
or U10492 (N_10492,N_9164,N_8159);
nand U10493 (N_10493,N_9609,N_8600);
xnor U10494 (N_10494,N_9264,N_8275);
nor U10495 (N_10495,N_9379,N_8920);
xnor U10496 (N_10496,N_9731,N_9890);
xnor U10497 (N_10497,N_8465,N_9168);
xor U10498 (N_10498,N_9106,N_9357);
nand U10499 (N_10499,N_8533,N_9277);
and U10500 (N_10500,N_8341,N_8209);
xnor U10501 (N_10501,N_9484,N_9219);
nor U10502 (N_10502,N_8958,N_8742);
nor U10503 (N_10503,N_8120,N_9362);
nor U10504 (N_10504,N_9031,N_9473);
xnor U10505 (N_10505,N_8080,N_8727);
xor U10506 (N_10506,N_8380,N_9386);
or U10507 (N_10507,N_9790,N_9811);
or U10508 (N_10508,N_9686,N_8430);
or U10509 (N_10509,N_8107,N_9485);
nor U10510 (N_10510,N_9044,N_9675);
and U10511 (N_10511,N_8405,N_8915);
nor U10512 (N_10512,N_9834,N_8604);
or U10513 (N_10513,N_8594,N_9353);
or U10514 (N_10514,N_8334,N_8585);
and U10515 (N_10515,N_9842,N_8009);
and U10516 (N_10516,N_9625,N_9390);
nand U10517 (N_10517,N_9878,N_9532);
and U10518 (N_10518,N_9509,N_9378);
nor U10519 (N_10519,N_8013,N_9216);
nand U10520 (N_10520,N_9841,N_8893);
nand U10521 (N_10521,N_9891,N_8840);
or U10522 (N_10522,N_8241,N_8279);
xnor U10523 (N_10523,N_9553,N_8475);
xnor U10524 (N_10524,N_8429,N_9507);
xor U10525 (N_10525,N_8633,N_9058);
nor U10526 (N_10526,N_8177,N_9010);
nor U10527 (N_10527,N_8478,N_9047);
nand U10528 (N_10528,N_9537,N_8863);
nand U10529 (N_10529,N_9443,N_8518);
and U10530 (N_10530,N_9958,N_8900);
nor U10531 (N_10531,N_8419,N_8578);
and U10532 (N_10532,N_8451,N_8596);
nand U10533 (N_10533,N_8422,N_9135);
and U10534 (N_10534,N_8413,N_9211);
or U10535 (N_10535,N_9224,N_8795);
or U10536 (N_10536,N_8483,N_9985);
nand U10537 (N_10537,N_9794,N_9558);
and U10538 (N_10538,N_9953,N_8206);
nor U10539 (N_10539,N_9754,N_9159);
nand U10540 (N_10540,N_8044,N_9571);
xor U10541 (N_10541,N_8539,N_8140);
or U10542 (N_10542,N_8538,N_8439);
and U10543 (N_10543,N_8028,N_9062);
xnor U10544 (N_10544,N_9775,N_9354);
nand U10545 (N_10545,N_9549,N_9941);
xor U10546 (N_10546,N_9879,N_9103);
or U10547 (N_10547,N_8877,N_9939);
xor U10548 (N_10548,N_8841,N_8778);
xor U10549 (N_10549,N_9706,N_9430);
and U10550 (N_10550,N_9801,N_8815);
or U10551 (N_10551,N_9095,N_8401);
nor U10552 (N_10552,N_9654,N_9825);
xnor U10553 (N_10553,N_9198,N_8856);
nand U10554 (N_10554,N_8983,N_8609);
or U10555 (N_10555,N_9937,N_9260);
nor U10556 (N_10556,N_8645,N_9534);
xor U10557 (N_10557,N_8497,N_9711);
nor U10558 (N_10558,N_8060,N_8331);
or U10559 (N_10559,N_8690,N_8386);
nand U10560 (N_10560,N_8678,N_9432);
xnor U10561 (N_10561,N_9308,N_9407);
nand U10562 (N_10562,N_8409,N_9680);
nand U10563 (N_10563,N_8105,N_8109);
xor U10564 (N_10564,N_9231,N_9496);
or U10565 (N_10565,N_8228,N_8765);
xor U10566 (N_10566,N_9175,N_9256);
xnor U10567 (N_10567,N_9973,N_8880);
nand U10568 (N_10568,N_8846,N_9156);
nand U10569 (N_10569,N_8203,N_8521);
nor U10570 (N_10570,N_8808,N_9319);
xnor U10571 (N_10571,N_8569,N_8156);
xor U10572 (N_10572,N_8773,N_8039);
nand U10573 (N_10573,N_9333,N_9002);
and U10574 (N_10574,N_8781,N_9300);
or U10575 (N_10575,N_8703,N_9715);
and U10576 (N_10576,N_8948,N_8906);
nor U10577 (N_10577,N_9886,N_8750);
xor U10578 (N_10578,N_8944,N_9004);
nor U10579 (N_10579,N_8746,N_8648);
nor U10580 (N_10580,N_8085,N_8679);
or U10581 (N_10581,N_8924,N_8661);
or U10582 (N_10582,N_9292,N_9912);
nand U10583 (N_10583,N_9434,N_8127);
and U10584 (N_10584,N_8634,N_8616);
and U10585 (N_10585,N_9592,N_8256);
nand U10586 (N_10586,N_9349,N_8542);
nand U10587 (N_10587,N_9035,N_9610);
xnor U10588 (N_10588,N_9217,N_8247);
or U10589 (N_10589,N_8111,N_8832);
nor U10590 (N_10590,N_8368,N_9376);
xor U10591 (N_10591,N_9591,N_8697);
nor U10592 (N_10592,N_8752,N_8930);
and U10593 (N_10593,N_8582,N_9404);
xor U10594 (N_10594,N_9523,N_9039);
xor U10595 (N_10595,N_8041,N_9444);
xnor U10596 (N_10596,N_8222,N_9384);
or U10597 (N_10597,N_8375,N_9214);
xor U10598 (N_10598,N_8499,N_8162);
nor U10599 (N_10599,N_9056,N_8126);
nand U10600 (N_10600,N_9218,N_8515);
or U10601 (N_10601,N_9399,N_8646);
nand U10602 (N_10602,N_8408,N_8575);
or U10603 (N_10603,N_8928,N_9445);
or U10604 (N_10604,N_8721,N_8187);
xnor U10605 (N_10605,N_8548,N_8294);
nand U10606 (N_10606,N_9947,N_9089);
xor U10607 (N_10607,N_9765,N_9266);
or U10608 (N_10608,N_9415,N_9931);
nor U10609 (N_10609,N_9907,N_9737);
or U10610 (N_10610,N_9252,N_9065);
nand U10611 (N_10611,N_9506,N_9896);
nor U10612 (N_10612,N_8070,N_8450);
nand U10613 (N_10613,N_8250,N_9424);
nor U10614 (N_10614,N_8506,N_9413);
nand U10615 (N_10615,N_8666,N_9701);
nor U10616 (N_10616,N_9888,N_9157);
xor U10617 (N_10617,N_9080,N_8618);
or U10618 (N_10618,N_8593,N_8631);
and U10619 (N_10619,N_8667,N_9416);
xnor U10620 (N_10620,N_8608,N_8473);
and U10621 (N_10621,N_8376,N_8545);
nand U10622 (N_10622,N_9943,N_9180);
xor U10623 (N_10623,N_9286,N_8104);
nor U10624 (N_10624,N_9336,N_8359);
and U10625 (N_10625,N_8314,N_8654);
and U10626 (N_10626,N_8335,N_9983);
or U10627 (N_10627,N_9977,N_9869);
and U10628 (N_10628,N_8296,N_9703);
nand U10629 (N_10629,N_9469,N_8096);
and U10630 (N_10630,N_9368,N_8865);
and U10631 (N_10631,N_9305,N_9828);
or U10632 (N_10632,N_8586,N_8992);
nor U10633 (N_10633,N_9575,N_8416);
nor U10634 (N_10634,N_9113,N_9626);
nor U10635 (N_10635,N_8755,N_9369);
or U10636 (N_10636,N_8918,N_9627);
and U10637 (N_10637,N_8142,N_8271);
nor U10638 (N_10638,N_8197,N_9908);
nor U10639 (N_10639,N_8343,N_9733);
nand U10640 (N_10640,N_9767,N_8993);
nand U10641 (N_10641,N_9829,N_8125);
and U10642 (N_10642,N_9736,N_9297);
or U10643 (N_10643,N_8244,N_8761);
or U10644 (N_10644,N_9132,N_9530);
nor U10645 (N_10645,N_9091,N_9115);
nor U10646 (N_10646,N_8614,N_8536);
or U10647 (N_10647,N_8273,N_9112);
and U10648 (N_10648,N_9997,N_9273);
or U10649 (N_10649,N_9772,N_9490);
nor U10650 (N_10650,N_8670,N_8014);
nor U10651 (N_10651,N_8023,N_9111);
nand U10652 (N_10652,N_9102,N_9248);
xnor U10653 (N_10653,N_9394,N_8787);
xor U10654 (N_10654,N_9016,N_8240);
xnor U10655 (N_10655,N_8884,N_9213);
nor U10656 (N_10656,N_9447,N_9854);
nor U10657 (N_10657,N_8861,N_8136);
xnor U10658 (N_10658,N_9876,N_9789);
and U10659 (N_10659,N_8066,N_8734);
nand U10660 (N_10660,N_9561,N_8821);
nand U10661 (N_10661,N_9599,N_9476);
nand U10662 (N_10662,N_9952,N_9751);
nor U10663 (N_10663,N_8951,N_9304);
nand U10664 (N_10664,N_8254,N_8238);
nand U10665 (N_10665,N_9024,N_9338);
xor U10666 (N_10666,N_9400,N_9203);
xnor U10667 (N_10667,N_8087,N_8161);
xor U10668 (N_10668,N_9261,N_8988);
and U10669 (N_10669,N_9188,N_9598);
nor U10670 (N_10670,N_8458,N_9170);
nand U10671 (N_10671,N_8301,N_8653);
and U10672 (N_10672,N_8802,N_9660);
xnor U10673 (N_10673,N_8705,N_9500);
or U10674 (N_10674,N_8036,N_8158);
and U10675 (N_10675,N_8148,N_8211);
and U10676 (N_10676,N_8845,N_8216);
xor U10677 (N_10677,N_9550,N_9241);
nor U10678 (N_10678,N_8282,N_9197);
and U10679 (N_10679,N_9919,N_9555);
xnor U10680 (N_10680,N_9048,N_9107);
nor U10681 (N_10681,N_9739,N_9942);
and U10682 (N_10682,N_8949,N_8388);
and U10683 (N_10683,N_9207,N_8431);
and U10684 (N_10684,N_8170,N_9744);
and U10685 (N_10685,N_8072,N_8534);
xnor U10686 (N_10686,N_8818,N_9846);
or U10687 (N_10687,N_9215,N_9382);
nor U10688 (N_10688,N_8735,N_9110);
nand U10689 (N_10689,N_8947,N_9652);
nand U10690 (N_10690,N_9464,N_8410);
nand U10691 (N_10691,N_9758,N_8568);
nor U10692 (N_10692,N_9718,N_8317);
or U10693 (N_10693,N_9781,N_8191);
nor U10694 (N_10694,N_8798,N_8581);
and U10695 (N_10695,N_8225,N_9727);
xnor U10696 (N_10696,N_9616,N_8953);
xnor U10697 (N_10697,N_8391,N_9670);
and U10698 (N_10698,N_9397,N_9557);
and U10699 (N_10699,N_8809,N_9597);
and U10700 (N_10700,N_8523,N_9815);
xnor U10701 (N_10701,N_8597,N_8468);
xnor U10702 (N_10702,N_9054,N_9448);
nor U10703 (N_10703,N_9022,N_8084);
nor U10704 (N_10704,N_8546,N_8663);
nor U10705 (N_10705,N_8725,N_8049);
nand U10706 (N_10706,N_8932,N_8656);
nor U10707 (N_10707,N_9282,N_8383);
or U10708 (N_10708,N_8574,N_8122);
xnor U10709 (N_10709,N_8196,N_8718);
and U10710 (N_10710,N_9249,N_9259);
xnor U10711 (N_10711,N_8999,N_9481);
and U10712 (N_10712,N_8931,N_8559);
and U10713 (N_10713,N_8514,N_8834);
or U10714 (N_10714,N_9818,N_9342);
and U10715 (N_10715,N_8708,N_8464);
nor U10716 (N_10716,N_9100,N_8731);
xor U10717 (N_10717,N_8200,N_9486);
nand U10718 (N_10718,N_9590,N_9639);
nor U10719 (N_10719,N_9819,N_9613);
xnor U10720 (N_10720,N_9533,N_8902);
and U10721 (N_10721,N_9649,N_9935);
or U10722 (N_10722,N_9323,N_8632);
and U10723 (N_10723,N_9329,N_8810);
or U10724 (N_10724,N_9077,N_9600);
or U10725 (N_10725,N_9756,N_9193);
nand U10726 (N_10726,N_9957,N_8852);
xor U10727 (N_10727,N_9483,N_8630);
and U10728 (N_10728,N_9960,N_8772);
xor U10729 (N_10729,N_9768,N_8098);
and U10730 (N_10730,N_8702,N_8710);
and U10731 (N_10731,N_9348,N_9435);
and U10732 (N_10732,N_9176,N_8393);
nand U10733 (N_10733,N_8824,N_9367);
xnor U10734 (N_10734,N_9161,N_9814);
nand U10735 (N_10735,N_9104,N_9220);
nor U10736 (N_10736,N_9976,N_9951);
nor U10737 (N_10737,N_9930,N_9868);
nand U10738 (N_10738,N_9574,N_8056);
or U10739 (N_10739,N_9848,N_8881);
and U10740 (N_10740,N_9568,N_8462);
nand U10741 (N_10741,N_9838,N_8373);
and U10742 (N_10742,N_8354,N_8292);
nor U10743 (N_10743,N_9021,N_9582);
nor U10744 (N_10744,N_9130,N_8447);
nand U10745 (N_10745,N_8249,N_9489);
or U10746 (N_10746,N_8160,N_8767);
and U10747 (N_10747,N_8389,N_9617);
nor U10748 (N_10748,N_8255,N_9674);
xor U10749 (N_10749,N_8764,N_8839);
or U10750 (N_10750,N_8010,N_8051);
and U10751 (N_10751,N_9470,N_8045);
xor U10752 (N_10752,N_9499,N_9222);
nor U10753 (N_10753,N_8833,N_8990);
and U10754 (N_10754,N_9406,N_9539);
or U10755 (N_10755,N_8756,N_8281);
nor U10756 (N_10756,N_8237,N_9008);
xor U10757 (N_10757,N_8199,N_8929);
nor U10758 (N_10758,N_9124,N_8939);
or U10759 (N_10759,N_9057,N_9972);
and U10760 (N_10760,N_8747,N_8190);
and U10761 (N_10761,N_8844,N_8896);
xnor U10762 (N_10762,N_8100,N_9874);
xnor U10763 (N_10763,N_8088,N_8360);
or U10764 (N_10764,N_9160,N_8390);
or U10765 (N_10765,N_8441,N_9538);
or U10766 (N_10766,N_9087,N_8660);
xnor U10767 (N_10767,N_9472,N_9327);
xor U10768 (N_10768,N_9233,N_9227);
xnor U10769 (N_10769,N_8698,N_8119);
nor U10770 (N_10770,N_8207,N_9151);
nor U10771 (N_10771,N_9078,N_8850);
xnor U10772 (N_10772,N_9147,N_8589);
and U10773 (N_10773,N_8117,N_8659);
nand U10774 (N_10774,N_9274,N_9317);
nand U10775 (N_10775,N_9467,N_9968);
and U10776 (N_10776,N_8195,N_9808);
nor U10777 (N_10777,N_9916,N_8685);
nor U10778 (N_10778,N_8805,N_9717);
or U10779 (N_10779,N_8325,N_8744);
and U10780 (N_10780,N_8208,N_9824);
nand U10781 (N_10781,N_9833,N_8644);
or U10782 (N_10782,N_8189,N_8128);
nor U10783 (N_10783,N_9541,N_9205);
nor U10784 (N_10784,N_8133,N_9784);
xnor U10785 (N_10785,N_8463,N_9563);
xor U10786 (N_10786,N_8192,N_8753);
nor U10787 (N_10787,N_8872,N_9683);
nand U10788 (N_10788,N_9298,N_9251);
nor U10789 (N_10789,N_9755,N_9206);
nor U10790 (N_10790,N_9455,N_8224);
nand U10791 (N_10791,N_8823,N_8090);
and U10792 (N_10792,N_9704,N_8726);
nor U10793 (N_10793,N_9330,N_9326);
and U10794 (N_10794,N_8689,N_9668);
xor U10795 (N_10795,N_9181,N_9096);
xor U10796 (N_10796,N_9402,N_8511);
and U10797 (N_10797,N_8560,N_9667);
and U10798 (N_10798,N_9145,N_9245);
xnor U10799 (N_10799,N_8353,N_8068);
nor U10800 (N_10800,N_8074,N_9694);
nor U10801 (N_10801,N_9525,N_9439);
nor U10802 (N_10802,N_9440,N_8065);
xnor U10803 (N_10803,N_8179,N_8794);
nor U10804 (N_10804,N_9707,N_9994);
and U10805 (N_10805,N_8477,N_8418);
or U10806 (N_10806,N_8888,N_9881);
nor U10807 (N_10807,N_9708,N_8859);
nor U10808 (N_10808,N_8804,N_8819);
nand U10809 (N_10809,N_8379,N_8676);
nor U10810 (N_10810,N_9697,N_8510);
or U10811 (N_10811,N_9136,N_9696);
or U10812 (N_10812,N_9778,N_8686);
nor U10813 (N_10813,N_8909,N_9545);
nand U10814 (N_10814,N_9865,N_8565);
nand U10815 (N_10815,N_9785,N_8879);
nor U10816 (N_10816,N_9477,N_9588);
nand U10817 (N_10817,N_8490,N_8505);
and U10818 (N_10818,N_9269,N_9267);
xnor U10819 (N_10819,N_8799,N_8415);
and U10820 (N_10820,N_9927,N_9893);
and U10821 (N_10821,N_9906,N_9900);
nor U10822 (N_10822,N_8054,N_9360);
and U10823 (N_10823,N_8019,N_8544);
and U10824 (N_10824,N_9528,N_9232);
or U10825 (N_10825,N_9547,N_9005);
or U10826 (N_10826,N_9928,N_9883);
and U10827 (N_10827,N_8129,N_9493);
xnor U10828 (N_10828,N_9515,N_8564);
nand U10829 (N_10829,N_8043,N_8913);
and U10830 (N_10830,N_9716,N_8828);
nand U10831 (N_10831,N_8530,N_8455);
nand U10832 (N_10832,N_8174,N_9301);
xnor U10833 (N_10833,N_9243,N_9921);
or U10834 (N_10834,N_8554,N_8552);
nand U10835 (N_10835,N_9322,N_9641);
or U10836 (N_10836,N_8089,N_8445);
nand U10837 (N_10837,N_8108,N_8459);
and U10838 (N_10838,N_9270,N_9174);
nor U10839 (N_10839,N_8157,N_8801);
or U10840 (N_10840,N_9580,N_9398);
nor U10841 (N_10841,N_8583,N_9086);
nor U10842 (N_10842,N_9293,N_8625);
or U10843 (N_10843,N_9182,N_9875);
or U10844 (N_10844,N_8064,N_9237);
xor U10845 (N_10845,N_9595,N_9061);
nor U10846 (N_10846,N_8342,N_8922);
or U10847 (N_10847,N_9798,N_9389);
xor U10848 (N_10848,N_8737,N_9302);
and U10849 (N_10849,N_9748,N_8001);
nor U10850 (N_10850,N_8640,N_8137);
or U10851 (N_10851,N_8526,N_9984);
xnor U10852 (N_10852,N_8348,N_8269);
nand U10853 (N_10853,N_8487,N_9423);
xor U10854 (N_10854,N_8680,N_9970);
or U10855 (N_10855,N_9341,N_8002);
and U10856 (N_10856,N_9577,N_9000);
xor U10857 (N_10857,N_9118,N_8550);
xnor U10858 (N_10858,N_9276,N_8945);
or U10859 (N_10859,N_9162,N_9029);
nand U10860 (N_10860,N_9268,N_8078);
and U10861 (N_10861,N_8406,N_9807);
xor U10862 (N_10862,N_9114,N_9152);
xor U10863 (N_10863,N_8714,N_9823);
nand U10864 (N_10864,N_8257,N_9498);
xnor U10865 (N_10865,N_9656,N_8425);
xnor U10866 (N_10866,N_9479,N_8598);
xnor U10867 (N_10867,N_8322,N_9982);
xnor U10868 (N_10868,N_9050,N_9677);
and U10869 (N_10869,N_9546,N_9133);
nor U10870 (N_10870,N_8333,N_9691);
and U10871 (N_10871,N_9612,N_8785);
xnor U10872 (N_10872,N_9786,N_9036);
nand U10873 (N_10873,N_8650,N_9593);
or U10874 (N_10874,N_8751,N_9567);
and U10875 (N_10875,N_9199,N_9371);
nand U10876 (N_10876,N_9335,N_8606);
nand U10877 (N_10877,N_9288,N_9210);
and U10878 (N_10878,N_8899,N_9926);
and U10879 (N_10879,N_9395,N_8092);
xnor U10880 (N_10880,N_8278,N_9017);
xor U10881 (N_10881,N_9847,N_9250);
xnor U10882 (N_10882,N_9544,N_9620);
xor U10883 (N_10883,N_9148,N_9766);
xor U10884 (N_10884,N_8803,N_8261);
nand U10885 (N_10885,N_8796,N_8878);
nor U10886 (N_10886,N_9265,N_8112);
or U10887 (N_10887,N_9179,N_9125);
and U10888 (N_10888,N_9280,N_9501);
nor U10889 (N_10889,N_8371,N_8332);
or U10890 (N_10890,N_9693,N_9805);
xor U10891 (N_10891,N_8055,N_9872);
xnor U10892 (N_10892,N_9721,N_8956);
or U10893 (N_10893,N_9007,N_9877);
or U10894 (N_10894,N_8031,N_8588);
nand U10895 (N_10895,N_9642,N_8837);
nand U10896 (N_10896,N_8504,N_9034);
xnor U10897 (N_10897,N_8791,N_9777);
nand U10898 (N_10898,N_9787,N_9845);
nand U10899 (N_10899,N_9623,N_9195);
nor U10900 (N_10900,N_9800,N_9303);
or U10901 (N_10901,N_8183,N_8016);
and U10902 (N_10902,N_9474,N_8258);
xor U10903 (N_10903,N_8712,N_9355);
or U10904 (N_10904,N_8720,N_8897);
xnor U10905 (N_10905,N_9902,N_8327);
or U10906 (N_10906,N_9712,N_9127);
xnor U10907 (N_10907,N_8875,N_9682);
nor U10908 (N_10908,N_9346,N_9832);
nor U10909 (N_10909,N_8457,N_8636);
or U10910 (N_10910,N_9551,N_8150);
xnor U10911 (N_10911,N_9339,N_9629);
nand U10912 (N_10912,N_8722,N_9401);
or U10913 (N_10913,N_8349,N_9949);
and U10914 (N_10914,N_8771,N_8420);
or U10915 (N_10915,N_8507,N_8035);
xor U10916 (N_10916,N_8623,N_9803);
nand U10917 (N_10917,N_8178,N_8605);
and U10918 (N_10918,N_9081,N_9043);
nand U10919 (N_10919,N_9695,N_8626);
nor U10920 (N_10920,N_8340,N_8198);
and U10921 (N_10921,N_9492,N_9120);
nand U10922 (N_10922,N_9747,N_8591);
or U10923 (N_10923,N_9254,N_9143);
xnor U10924 (N_10924,N_8674,N_9003);
and U10925 (N_10925,N_9466,N_9897);
and U10926 (N_10926,N_9554,N_8635);
or U10927 (N_10927,N_9687,N_9762);
nand U10928 (N_10928,N_9552,N_8952);
nor U10929 (N_10929,N_8006,N_8739);
and U10930 (N_10930,N_8573,N_8854);
nor U10931 (N_10931,N_8067,N_9359);
xnor U10932 (N_10932,N_8034,N_9240);
xor U10933 (N_10933,N_8469,N_8466);
nand U10934 (N_10934,N_8287,N_9770);
or U10935 (N_10935,N_8444,N_9759);
xnor U10936 (N_10936,N_9310,N_8324);
nor U10937 (N_10937,N_9166,N_8903);
and U10938 (N_10938,N_9068,N_8775);
and U10939 (N_10939,N_8417,N_8326);
xor U10940 (N_10940,N_8436,N_8812);
and U10941 (N_10941,N_9066,N_9475);
and U10942 (N_10942,N_8851,N_9998);
xnor U10943 (N_10943,N_8219,N_8675);
xor U10944 (N_10944,N_8082,N_9295);
xor U10945 (N_10945,N_8868,N_8230);
xor U10946 (N_10946,N_8239,N_9871);
nor U10947 (N_10947,N_9076,N_8535);
nand U10948 (N_10948,N_8979,N_8412);
nand U10949 (N_10949,N_9418,N_8905);
nor U10950 (N_10950,N_9126,N_9085);
xor U10951 (N_10951,N_8110,N_9796);
nor U10952 (N_10952,N_9646,N_8940);
nor U10953 (N_10953,N_8643,N_9535);
and U10954 (N_10954,N_9795,N_9705);
and U10955 (N_10955,N_9505,N_9929);
and U10956 (N_10956,N_9281,N_8053);
xor U10957 (N_10957,N_8351,N_8520);
and U10958 (N_10958,N_8829,N_8432);
or U10959 (N_10959,N_8790,N_8886);
xor U10960 (N_10960,N_8555,N_8779);
nor U10961 (N_10961,N_9502,N_8442);
or U10962 (N_10962,N_9584,N_8233);
xor U10963 (N_10963,N_9914,N_9618);
or U10964 (N_10964,N_8723,N_9522);
nand U10965 (N_10965,N_9531,N_9279);
xnor U10966 (N_10966,N_8577,N_8188);
and U10967 (N_10967,N_8480,N_9351);
nand U10968 (N_10968,N_9945,N_8621);
or U10969 (N_10969,N_8496,N_9782);
xor U10970 (N_10970,N_8776,N_8443);
or U10971 (N_10971,N_9109,N_8048);
xor U10972 (N_10972,N_8655,N_8547);
and U10973 (N_10973,N_9459,N_9608);
nand U10974 (N_10974,N_9964,N_9556);
xor U10975 (N_10975,N_8637,N_8381);
nor U10976 (N_10976,N_9146,N_9052);
nor U10977 (N_10977,N_8826,N_8917);
nand U10978 (N_10978,N_8154,N_9763);
nor U10979 (N_10979,N_9816,N_8402);
and U10980 (N_10980,N_8669,N_9321);
nand U10981 (N_10981,N_8946,N_8058);
nor U10982 (N_10982,N_8492,N_8423);
xor U10983 (N_10983,N_9587,N_9980);
and U10984 (N_10984,N_8283,N_9722);
xor U10985 (N_10985,N_9331,N_8782);
or U10986 (N_10986,N_9190,N_9570);
or U10987 (N_10987,N_9363,N_8570);
nand U10988 (N_10988,N_8651,N_8587);
xnor U10989 (N_10989,N_8622,N_8357);
xnor U10990 (N_10990,N_8528,N_8748);
nand U10991 (N_10991,N_9839,N_9388);
nand U10992 (N_10992,N_9728,N_9684);
or U10993 (N_10993,N_8182,N_9461);
and U10994 (N_10994,N_9529,N_9996);
or U10995 (N_10995,N_9060,N_8372);
nor U10996 (N_10996,N_9226,N_9791);
nor U10997 (N_10997,N_9889,N_8701);
nand U10998 (N_10998,N_9844,N_8624);
and U10999 (N_10999,N_8713,N_8139);
nand U11000 (N_11000,N_8354,N_9067);
or U11001 (N_11001,N_8627,N_9544);
and U11002 (N_11002,N_9880,N_9675);
xnor U11003 (N_11003,N_8867,N_9466);
nor U11004 (N_11004,N_9925,N_9864);
nor U11005 (N_11005,N_9055,N_8145);
nor U11006 (N_11006,N_8698,N_8382);
or U11007 (N_11007,N_8201,N_9943);
and U11008 (N_11008,N_8586,N_9083);
or U11009 (N_11009,N_8533,N_9941);
nand U11010 (N_11010,N_9571,N_9281);
nand U11011 (N_11011,N_9918,N_8305);
and U11012 (N_11012,N_9237,N_8801);
and U11013 (N_11013,N_8471,N_9399);
and U11014 (N_11014,N_9413,N_8780);
nor U11015 (N_11015,N_9192,N_9042);
nand U11016 (N_11016,N_8363,N_9144);
and U11017 (N_11017,N_8424,N_9191);
nand U11018 (N_11018,N_8906,N_8768);
and U11019 (N_11019,N_9992,N_8688);
and U11020 (N_11020,N_8936,N_9213);
xnor U11021 (N_11021,N_8232,N_8122);
nor U11022 (N_11022,N_8117,N_9737);
or U11023 (N_11023,N_9660,N_8530);
xnor U11024 (N_11024,N_8371,N_9187);
and U11025 (N_11025,N_8907,N_9457);
xnor U11026 (N_11026,N_9362,N_9468);
or U11027 (N_11027,N_9760,N_8901);
nand U11028 (N_11028,N_8292,N_8759);
or U11029 (N_11029,N_9764,N_8480);
xor U11030 (N_11030,N_8297,N_8663);
or U11031 (N_11031,N_8821,N_8961);
nand U11032 (N_11032,N_8443,N_8923);
or U11033 (N_11033,N_9329,N_9330);
nand U11034 (N_11034,N_9856,N_8610);
nand U11035 (N_11035,N_9157,N_8333);
nor U11036 (N_11036,N_8530,N_9417);
or U11037 (N_11037,N_8024,N_9739);
and U11038 (N_11038,N_8173,N_9320);
nand U11039 (N_11039,N_9080,N_8459);
nand U11040 (N_11040,N_9392,N_8509);
and U11041 (N_11041,N_8135,N_9724);
nand U11042 (N_11042,N_9240,N_9551);
nand U11043 (N_11043,N_8617,N_8010);
nand U11044 (N_11044,N_8847,N_9140);
nand U11045 (N_11045,N_8079,N_8483);
and U11046 (N_11046,N_9944,N_8902);
nand U11047 (N_11047,N_8870,N_9307);
and U11048 (N_11048,N_8484,N_8256);
or U11049 (N_11049,N_8528,N_8336);
nand U11050 (N_11050,N_9238,N_9784);
xor U11051 (N_11051,N_9270,N_9917);
nor U11052 (N_11052,N_9478,N_9449);
xnor U11053 (N_11053,N_9001,N_9754);
xor U11054 (N_11054,N_9397,N_9799);
nor U11055 (N_11055,N_9389,N_9916);
or U11056 (N_11056,N_8663,N_9175);
or U11057 (N_11057,N_9784,N_9761);
xnor U11058 (N_11058,N_8135,N_9377);
nor U11059 (N_11059,N_9743,N_9731);
and U11060 (N_11060,N_8993,N_9965);
or U11061 (N_11061,N_8897,N_8360);
nand U11062 (N_11062,N_9679,N_9933);
nand U11063 (N_11063,N_9991,N_9538);
nand U11064 (N_11064,N_8470,N_9101);
and U11065 (N_11065,N_8654,N_9755);
xor U11066 (N_11066,N_9342,N_9177);
or U11067 (N_11067,N_9961,N_9659);
or U11068 (N_11068,N_9643,N_8497);
nor U11069 (N_11069,N_8884,N_8030);
or U11070 (N_11070,N_9853,N_9071);
and U11071 (N_11071,N_9924,N_8132);
nor U11072 (N_11072,N_9236,N_8650);
nand U11073 (N_11073,N_9659,N_9223);
and U11074 (N_11074,N_8877,N_9873);
and U11075 (N_11075,N_8425,N_8114);
nor U11076 (N_11076,N_8571,N_9304);
nand U11077 (N_11077,N_9593,N_8178);
and U11078 (N_11078,N_9017,N_8101);
xor U11079 (N_11079,N_9435,N_9622);
and U11080 (N_11080,N_8895,N_9202);
nand U11081 (N_11081,N_9094,N_9448);
nand U11082 (N_11082,N_8219,N_8476);
or U11083 (N_11083,N_8015,N_9319);
nand U11084 (N_11084,N_8710,N_9222);
nor U11085 (N_11085,N_9746,N_9667);
xnor U11086 (N_11086,N_8673,N_8400);
xnor U11087 (N_11087,N_9724,N_8190);
and U11088 (N_11088,N_8663,N_9754);
and U11089 (N_11089,N_9012,N_8744);
or U11090 (N_11090,N_9160,N_9683);
nand U11091 (N_11091,N_8447,N_9174);
xnor U11092 (N_11092,N_9065,N_9338);
xor U11093 (N_11093,N_9070,N_8572);
nand U11094 (N_11094,N_8115,N_9482);
nor U11095 (N_11095,N_9078,N_9278);
nand U11096 (N_11096,N_8079,N_9657);
or U11097 (N_11097,N_9620,N_8779);
nand U11098 (N_11098,N_8986,N_8531);
xor U11099 (N_11099,N_8626,N_9378);
or U11100 (N_11100,N_9834,N_8522);
and U11101 (N_11101,N_9609,N_8660);
nor U11102 (N_11102,N_8328,N_9347);
xor U11103 (N_11103,N_8705,N_9153);
and U11104 (N_11104,N_8377,N_9304);
xor U11105 (N_11105,N_8111,N_8275);
nand U11106 (N_11106,N_8172,N_8209);
nand U11107 (N_11107,N_8578,N_8715);
or U11108 (N_11108,N_9257,N_9962);
nor U11109 (N_11109,N_8985,N_8621);
nor U11110 (N_11110,N_8113,N_9347);
and U11111 (N_11111,N_9553,N_9175);
and U11112 (N_11112,N_9998,N_8086);
xnor U11113 (N_11113,N_8657,N_9975);
xnor U11114 (N_11114,N_8744,N_8923);
and U11115 (N_11115,N_9200,N_8084);
nand U11116 (N_11116,N_8764,N_8725);
or U11117 (N_11117,N_8965,N_9310);
nor U11118 (N_11118,N_9264,N_9652);
nor U11119 (N_11119,N_8693,N_8195);
or U11120 (N_11120,N_9935,N_8043);
nor U11121 (N_11121,N_8321,N_9297);
or U11122 (N_11122,N_8848,N_8831);
xnor U11123 (N_11123,N_8145,N_9644);
xnor U11124 (N_11124,N_8453,N_8719);
and U11125 (N_11125,N_9367,N_8359);
or U11126 (N_11126,N_9854,N_8398);
nor U11127 (N_11127,N_8590,N_8977);
nand U11128 (N_11128,N_9247,N_8916);
or U11129 (N_11129,N_9900,N_9406);
nand U11130 (N_11130,N_8652,N_9913);
and U11131 (N_11131,N_9029,N_8140);
and U11132 (N_11132,N_8849,N_9541);
nand U11133 (N_11133,N_9468,N_9878);
xnor U11134 (N_11134,N_9094,N_8951);
and U11135 (N_11135,N_8461,N_8081);
nand U11136 (N_11136,N_8064,N_8713);
xnor U11137 (N_11137,N_9160,N_9857);
nand U11138 (N_11138,N_8991,N_9365);
or U11139 (N_11139,N_8476,N_9288);
and U11140 (N_11140,N_8344,N_9370);
xor U11141 (N_11141,N_9909,N_8976);
nor U11142 (N_11142,N_8406,N_9971);
nor U11143 (N_11143,N_9070,N_8686);
nor U11144 (N_11144,N_9939,N_8618);
nand U11145 (N_11145,N_9944,N_8771);
and U11146 (N_11146,N_9484,N_8285);
nor U11147 (N_11147,N_8392,N_8703);
xnor U11148 (N_11148,N_9672,N_8681);
xor U11149 (N_11149,N_9207,N_8887);
or U11150 (N_11150,N_9141,N_8890);
or U11151 (N_11151,N_9856,N_8846);
nand U11152 (N_11152,N_9138,N_9042);
nor U11153 (N_11153,N_8905,N_8844);
and U11154 (N_11154,N_9546,N_8951);
nand U11155 (N_11155,N_8795,N_9989);
xor U11156 (N_11156,N_9101,N_9769);
nand U11157 (N_11157,N_8277,N_8884);
or U11158 (N_11158,N_9818,N_8643);
nor U11159 (N_11159,N_9321,N_8055);
or U11160 (N_11160,N_9046,N_8749);
or U11161 (N_11161,N_8636,N_8295);
nand U11162 (N_11162,N_8926,N_9671);
and U11163 (N_11163,N_8936,N_9848);
xor U11164 (N_11164,N_8978,N_9299);
and U11165 (N_11165,N_8928,N_9184);
nand U11166 (N_11166,N_8613,N_8085);
xnor U11167 (N_11167,N_9155,N_9427);
and U11168 (N_11168,N_9509,N_8558);
or U11169 (N_11169,N_8220,N_9440);
xor U11170 (N_11170,N_8669,N_8097);
xor U11171 (N_11171,N_9970,N_8719);
nor U11172 (N_11172,N_9937,N_8511);
xor U11173 (N_11173,N_8189,N_8908);
and U11174 (N_11174,N_9800,N_9659);
xnor U11175 (N_11175,N_9865,N_9643);
nor U11176 (N_11176,N_8849,N_9990);
nor U11177 (N_11177,N_8936,N_8668);
xnor U11178 (N_11178,N_8381,N_9821);
and U11179 (N_11179,N_8980,N_9277);
xnor U11180 (N_11180,N_8266,N_8714);
xnor U11181 (N_11181,N_9327,N_8177);
and U11182 (N_11182,N_8750,N_9996);
nor U11183 (N_11183,N_8953,N_9490);
xor U11184 (N_11184,N_9655,N_9219);
xor U11185 (N_11185,N_8462,N_9131);
nand U11186 (N_11186,N_8611,N_8937);
xor U11187 (N_11187,N_9554,N_9044);
and U11188 (N_11188,N_8896,N_8573);
nor U11189 (N_11189,N_8249,N_8253);
nand U11190 (N_11190,N_9501,N_8096);
or U11191 (N_11191,N_8065,N_9808);
nor U11192 (N_11192,N_9960,N_8520);
or U11193 (N_11193,N_8568,N_9808);
and U11194 (N_11194,N_8079,N_8398);
and U11195 (N_11195,N_8747,N_8239);
nand U11196 (N_11196,N_9287,N_8451);
xor U11197 (N_11197,N_9631,N_8521);
nor U11198 (N_11198,N_8186,N_8746);
or U11199 (N_11199,N_8603,N_8243);
or U11200 (N_11200,N_8517,N_8129);
nor U11201 (N_11201,N_9264,N_9627);
nand U11202 (N_11202,N_9814,N_9199);
xor U11203 (N_11203,N_8209,N_8478);
xnor U11204 (N_11204,N_9374,N_8694);
and U11205 (N_11205,N_8546,N_8136);
nand U11206 (N_11206,N_9098,N_8296);
nand U11207 (N_11207,N_8516,N_8705);
xor U11208 (N_11208,N_9529,N_9049);
xnor U11209 (N_11209,N_8641,N_8743);
nor U11210 (N_11210,N_8134,N_9574);
nand U11211 (N_11211,N_8586,N_9793);
nand U11212 (N_11212,N_9975,N_9016);
nor U11213 (N_11213,N_8208,N_8611);
xor U11214 (N_11214,N_9645,N_9499);
or U11215 (N_11215,N_8805,N_9577);
or U11216 (N_11216,N_9456,N_9686);
nand U11217 (N_11217,N_9736,N_8293);
and U11218 (N_11218,N_8216,N_8588);
and U11219 (N_11219,N_8343,N_9008);
or U11220 (N_11220,N_9337,N_9207);
and U11221 (N_11221,N_9996,N_8167);
nor U11222 (N_11222,N_8403,N_9915);
nor U11223 (N_11223,N_8827,N_8573);
xnor U11224 (N_11224,N_9750,N_8104);
xor U11225 (N_11225,N_9500,N_9249);
and U11226 (N_11226,N_9932,N_9425);
or U11227 (N_11227,N_9179,N_8456);
nor U11228 (N_11228,N_9170,N_9606);
nor U11229 (N_11229,N_8566,N_9903);
xor U11230 (N_11230,N_8744,N_9300);
nor U11231 (N_11231,N_9468,N_8882);
nor U11232 (N_11232,N_9615,N_9571);
nor U11233 (N_11233,N_8854,N_9991);
and U11234 (N_11234,N_8261,N_9774);
xor U11235 (N_11235,N_8270,N_9275);
or U11236 (N_11236,N_8092,N_9481);
and U11237 (N_11237,N_8400,N_8541);
xnor U11238 (N_11238,N_8772,N_9052);
nor U11239 (N_11239,N_8460,N_8545);
or U11240 (N_11240,N_9883,N_9523);
nor U11241 (N_11241,N_9709,N_8022);
and U11242 (N_11242,N_8054,N_8351);
xnor U11243 (N_11243,N_8891,N_8085);
nor U11244 (N_11244,N_8234,N_9426);
or U11245 (N_11245,N_9704,N_8691);
or U11246 (N_11246,N_9530,N_8061);
nand U11247 (N_11247,N_8207,N_9132);
and U11248 (N_11248,N_9551,N_8226);
nor U11249 (N_11249,N_8447,N_9944);
nor U11250 (N_11250,N_9922,N_8248);
nand U11251 (N_11251,N_9659,N_8968);
nor U11252 (N_11252,N_9217,N_9137);
nor U11253 (N_11253,N_8192,N_8574);
or U11254 (N_11254,N_8047,N_9580);
or U11255 (N_11255,N_8339,N_9526);
nand U11256 (N_11256,N_9799,N_9646);
nor U11257 (N_11257,N_9601,N_9949);
and U11258 (N_11258,N_8112,N_8111);
nor U11259 (N_11259,N_8045,N_8895);
or U11260 (N_11260,N_8952,N_8782);
nand U11261 (N_11261,N_8212,N_8457);
nand U11262 (N_11262,N_9800,N_9053);
and U11263 (N_11263,N_9008,N_9235);
xor U11264 (N_11264,N_8043,N_9061);
xor U11265 (N_11265,N_9903,N_8042);
or U11266 (N_11266,N_8182,N_9656);
xnor U11267 (N_11267,N_9801,N_8101);
xnor U11268 (N_11268,N_9823,N_9018);
and U11269 (N_11269,N_8063,N_9849);
xnor U11270 (N_11270,N_8339,N_8127);
or U11271 (N_11271,N_9206,N_9407);
nand U11272 (N_11272,N_9876,N_9961);
and U11273 (N_11273,N_8746,N_9576);
and U11274 (N_11274,N_8584,N_8140);
xor U11275 (N_11275,N_8927,N_8413);
and U11276 (N_11276,N_8615,N_8053);
nand U11277 (N_11277,N_8453,N_9581);
and U11278 (N_11278,N_9616,N_8280);
xnor U11279 (N_11279,N_8456,N_8596);
and U11280 (N_11280,N_9799,N_9425);
xnor U11281 (N_11281,N_9478,N_8378);
nor U11282 (N_11282,N_8533,N_8782);
xnor U11283 (N_11283,N_8424,N_9649);
and U11284 (N_11284,N_8906,N_8020);
and U11285 (N_11285,N_8527,N_9441);
and U11286 (N_11286,N_9886,N_9935);
nor U11287 (N_11287,N_9975,N_8068);
and U11288 (N_11288,N_8691,N_9076);
nand U11289 (N_11289,N_8897,N_8608);
xnor U11290 (N_11290,N_8515,N_9156);
nor U11291 (N_11291,N_9446,N_8367);
and U11292 (N_11292,N_9626,N_9282);
nor U11293 (N_11293,N_8529,N_9076);
nand U11294 (N_11294,N_8534,N_9655);
nand U11295 (N_11295,N_9696,N_9105);
nand U11296 (N_11296,N_8559,N_9362);
xor U11297 (N_11297,N_8563,N_8182);
nand U11298 (N_11298,N_9526,N_9916);
or U11299 (N_11299,N_8013,N_9575);
nand U11300 (N_11300,N_8054,N_8311);
nor U11301 (N_11301,N_9350,N_8549);
nor U11302 (N_11302,N_8421,N_8670);
xnor U11303 (N_11303,N_9540,N_8483);
nand U11304 (N_11304,N_9805,N_9638);
nor U11305 (N_11305,N_8537,N_9200);
or U11306 (N_11306,N_8057,N_9368);
and U11307 (N_11307,N_9779,N_9712);
nand U11308 (N_11308,N_8650,N_9181);
and U11309 (N_11309,N_8244,N_9711);
and U11310 (N_11310,N_8468,N_9978);
xnor U11311 (N_11311,N_9473,N_9269);
and U11312 (N_11312,N_8173,N_9483);
or U11313 (N_11313,N_9150,N_9003);
and U11314 (N_11314,N_9034,N_8871);
and U11315 (N_11315,N_8571,N_8380);
nand U11316 (N_11316,N_8878,N_8110);
nand U11317 (N_11317,N_8463,N_8667);
xor U11318 (N_11318,N_8019,N_9434);
nor U11319 (N_11319,N_8370,N_8813);
xor U11320 (N_11320,N_8556,N_8869);
xor U11321 (N_11321,N_9688,N_8940);
and U11322 (N_11322,N_8849,N_9574);
nand U11323 (N_11323,N_9167,N_9830);
xor U11324 (N_11324,N_9270,N_8927);
nor U11325 (N_11325,N_9235,N_9940);
nand U11326 (N_11326,N_8905,N_9926);
xnor U11327 (N_11327,N_8377,N_9562);
nand U11328 (N_11328,N_8909,N_9844);
xnor U11329 (N_11329,N_8307,N_9674);
nor U11330 (N_11330,N_8363,N_9673);
nand U11331 (N_11331,N_8768,N_8373);
xor U11332 (N_11332,N_9303,N_9889);
and U11333 (N_11333,N_8825,N_9717);
xnor U11334 (N_11334,N_8373,N_8697);
nor U11335 (N_11335,N_8858,N_9808);
nand U11336 (N_11336,N_9960,N_9702);
nand U11337 (N_11337,N_9559,N_9620);
xnor U11338 (N_11338,N_9399,N_9105);
nand U11339 (N_11339,N_9829,N_8324);
nor U11340 (N_11340,N_9081,N_9424);
nand U11341 (N_11341,N_8041,N_8455);
nor U11342 (N_11342,N_8211,N_9785);
and U11343 (N_11343,N_9340,N_8872);
nand U11344 (N_11344,N_8207,N_9244);
nand U11345 (N_11345,N_9583,N_8631);
nand U11346 (N_11346,N_9990,N_8559);
nand U11347 (N_11347,N_8993,N_8644);
nor U11348 (N_11348,N_9212,N_9994);
or U11349 (N_11349,N_9619,N_8130);
nor U11350 (N_11350,N_8265,N_9527);
and U11351 (N_11351,N_9107,N_8177);
xor U11352 (N_11352,N_9659,N_9000);
nor U11353 (N_11353,N_8384,N_9966);
nand U11354 (N_11354,N_9696,N_9613);
and U11355 (N_11355,N_9203,N_9914);
or U11356 (N_11356,N_8019,N_9273);
nor U11357 (N_11357,N_9473,N_8058);
nand U11358 (N_11358,N_8102,N_9191);
nand U11359 (N_11359,N_8332,N_8270);
nor U11360 (N_11360,N_8295,N_8253);
and U11361 (N_11361,N_8366,N_9656);
nand U11362 (N_11362,N_9293,N_8391);
xnor U11363 (N_11363,N_9273,N_9423);
xor U11364 (N_11364,N_9616,N_9393);
nand U11365 (N_11365,N_9625,N_8687);
nand U11366 (N_11366,N_9047,N_9803);
and U11367 (N_11367,N_8869,N_9209);
or U11368 (N_11368,N_9644,N_8738);
nor U11369 (N_11369,N_9145,N_9979);
xor U11370 (N_11370,N_8720,N_8776);
xor U11371 (N_11371,N_8205,N_9549);
nor U11372 (N_11372,N_8141,N_9771);
nor U11373 (N_11373,N_9862,N_9924);
or U11374 (N_11374,N_9049,N_9436);
nor U11375 (N_11375,N_9570,N_9805);
or U11376 (N_11376,N_9460,N_8551);
nor U11377 (N_11377,N_8103,N_8993);
xor U11378 (N_11378,N_9450,N_9934);
nand U11379 (N_11379,N_9727,N_9622);
nor U11380 (N_11380,N_8197,N_9162);
xor U11381 (N_11381,N_9115,N_8829);
or U11382 (N_11382,N_8331,N_8516);
nor U11383 (N_11383,N_9771,N_9715);
xnor U11384 (N_11384,N_9564,N_8431);
or U11385 (N_11385,N_8967,N_8987);
and U11386 (N_11386,N_9411,N_8618);
and U11387 (N_11387,N_9626,N_9432);
xor U11388 (N_11388,N_8604,N_8691);
xor U11389 (N_11389,N_9113,N_8974);
or U11390 (N_11390,N_9613,N_8263);
or U11391 (N_11391,N_9613,N_9452);
or U11392 (N_11392,N_9322,N_9131);
or U11393 (N_11393,N_8688,N_9384);
and U11394 (N_11394,N_9562,N_8637);
and U11395 (N_11395,N_8120,N_8815);
and U11396 (N_11396,N_8128,N_9451);
or U11397 (N_11397,N_8942,N_9977);
nand U11398 (N_11398,N_8376,N_8415);
or U11399 (N_11399,N_9059,N_9345);
and U11400 (N_11400,N_8877,N_9955);
nand U11401 (N_11401,N_8063,N_8689);
nor U11402 (N_11402,N_9477,N_8339);
xnor U11403 (N_11403,N_9330,N_8633);
and U11404 (N_11404,N_8432,N_9098);
nand U11405 (N_11405,N_9442,N_9846);
xor U11406 (N_11406,N_9751,N_9385);
nor U11407 (N_11407,N_9018,N_8471);
nand U11408 (N_11408,N_9985,N_8481);
or U11409 (N_11409,N_8934,N_9014);
xor U11410 (N_11410,N_9026,N_8584);
or U11411 (N_11411,N_9244,N_9090);
nor U11412 (N_11412,N_8891,N_9504);
nand U11413 (N_11413,N_8130,N_8653);
or U11414 (N_11414,N_9275,N_9439);
xor U11415 (N_11415,N_8915,N_9254);
or U11416 (N_11416,N_8534,N_9410);
or U11417 (N_11417,N_9394,N_8882);
or U11418 (N_11418,N_9872,N_9927);
nor U11419 (N_11419,N_9616,N_9042);
nand U11420 (N_11420,N_9171,N_8551);
xnor U11421 (N_11421,N_9762,N_8568);
xor U11422 (N_11422,N_8208,N_8254);
or U11423 (N_11423,N_8390,N_9274);
or U11424 (N_11424,N_8787,N_9493);
and U11425 (N_11425,N_8821,N_8908);
nor U11426 (N_11426,N_9554,N_9868);
nor U11427 (N_11427,N_9217,N_9776);
and U11428 (N_11428,N_9136,N_9087);
or U11429 (N_11429,N_9477,N_8171);
xnor U11430 (N_11430,N_9886,N_8608);
nand U11431 (N_11431,N_8283,N_8235);
xnor U11432 (N_11432,N_8502,N_8193);
or U11433 (N_11433,N_9160,N_8508);
xor U11434 (N_11434,N_8814,N_9934);
nor U11435 (N_11435,N_9522,N_8953);
xor U11436 (N_11436,N_9809,N_8433);
and U11437 (N_11437,N_9540,N_9579);
nand U11438 (N_11438,N_8149,N_8220);
xor U11439 (N_11439,N_8831,N_9972);
or U11440 (N_11440,N_8333,N_8970);
nand U11441 (N_11441,N_8461,N_8861);
or U11442 (N_11442,N_9096,N_9195);
nor U11443 (N_11443,N_9082,N_8447);
nand U11444 (N_11444,N_9584,N_9974);
nand U11445 (N_11445,N_9283,N_8303);
nand U11446 (N_11446,N_8298,N_9651);
or U11447 (N_11447,N_9354,N_8760);
xnor U11448 (N_11448,N_9080,N_8279);
nand U11449 (N_11449,N_9142,N_9303);
nor U11450 (N_11450,N_9857,N_9158);
xnor U11451 (N_11451,N_9866,N_8037);
nor U11452 (N_11452,N_8832,N_9375);
xnor U11453 (N_11453,N_9549,N_9257);
nor U11454 (N_11454,N_9438,N_9112);
and U11455 (N_11455,N_9420,N_8983);
or U11456 (N_11456,N_8321,N_8985);
nand U11457 (N_11457,N_8451,N_9891);
or U11458 (N_11458,N_9441,N_8299);
xor U11459 (N_11459,N_8145,N_8420);
xnor U11460 (N_11460,N_9080,N_9299);
or U11461 (N_11461,N_9299,N_8386);
and U11462 (N_11462,N_8802,N_9446);
xor U11463 (N_11463,N_9904,N_8970);
nand U11464 (N_11464,N_9204,N_8172);
nand U11465 (N_11465,N_9231,N_9767);
or U11466 (N_11466,N_8751,N_9379);
nand U11467 (N_11467,N_8678,N_9139);
nand U11468 (N_11468,N_9097,N_8291);
and U11469 (N_11469,N_8651,N_8523);
nand U11470 (N_11470,N_9355,N_9782);
nand U11471 (N_11471,N_9134,N_9038);
or U11472 (N_11472,N_9723,N_9880);
xnor U11473 (N_11473,N_8306,N_9637);
nor U11474 (N_11474,N_8209,N_8746);
xor U11475 (N_11475,N_9743,N_8272);
and U11476 (N_11476,N_9252,N_8093);
xor U11477 (N_11477,N_8380,N_9973);
or U11478 (N_11478,N_9804,N_8659);
or U11479 (N_11479,N_8800,N_8705);
and U11480 (N_11480,N_8552,N_9664);
nand U11481 (N_11481,N_9256,N_8920);
nor U11482 (N_11482,N_8005,N_8711);
and U11483 (N_11483,N_9675,N_9998);
and U11484 (N_11484,N_9658,N_9217);
nand U11485 (N_11485,N_8264,N_8581);
nand U11486 (N_11486,N_9306,N_9396);
nand U11487 (N_11487,N_8088,N_9970);
and U11488 (N_11488,N_8334,N_8545);
nor U11489 (N_11489,N_9949,N_8532);
nor U11490 (N_11490,N_8887,N_9815);
and U11491 (N_11491,N_9020,N_8349);
and U11492 (N_11492,N_8676,N_8439);
nor U11493 (N_11493,N_9025,N_8569);
or U11494 (N_11494,N_9113,N_9204);
and U11495 (N_11495,N_8116,N_9611);
nor U11496 (N_11496,N_8143,N_9595);
and U11497 (N_11497,N_9818,N_8942);
xnor U11498 (N_11498,N_9741,N_8502);
xnor U11499 (N_11499,N_8574,N_8690);
nor U11500 (N_11500,N_9647,N_9503);
nor U11501 (N_11501,N_9064,N_9897);
or U11502 (N_11502,N_9546,N_9175);
nor U11503 (N_11503,N_8441,N_9259);
nor U11504 (N_11504,N_8777,N_9130);
nand U11505 (N_11505,N_9396,N_9911);
nor U11506 (N_11506,N_9664,N_8283);
or U11507 (N_11507,N_9287,N_8788);
or U11508 (N_11508,N_9935,N_9208);
or U11509 (N_11509,N_9651,N_9331);
and U11510 (N_11510,N_9691,N_9201);
and U11511 (N_11511,N_8162,N_8115);
or U11512 (N_11512,N_8821,N_9531);
nand U11513 (N_11513,N_8511,N_9313);
nor U11514 (N_11514,N_8308,N_9133);
nand U11515 (N_11515,N_9802,N_9114);
and U11516 (N_11516,N_8150,N_9315);
nand U11517 (N_11517,N_9336,N_8248);
nor U11518 (N_11518,N_9306,N_9251);
nor U11519 (N_11519,N_9293,N_9576);
and U11520 (N_11520,N_9932,N_8163);
nand U11521 (N_11521,N_9808,N_9049);
xnor U11522 (N_11522,N_9836,N_9113);
nor U11523 (N_11523,N_9660,N_8382);
and U11524 (N_11524,N_9478,N_8783);
or U11525 (N_11525,N_8753,N_8575);
nand U11526 (N_11526,N_9101,N_9793);
nor U11527 (N_11527,N_9957,N_9805);
and U11528 (N_11528,N_8869,N_8344);
xor U11529 (N_11529,N_8984,N_9716);
nor U11530 (N_11530,N_8682,N_9015);
nor U11531 (N_11531,N_8208,N_8627);
and U11532 (N_11532,N_8108,N_9470);
nor U11533 (N_11533,N_9908,N_8344);
and U11534 (N_11534,N_8198,N_9573);
and U11535 (N_11535,N_8740,N_8269);
and U11536 (N_11536,N_8887,N_8172);
and U11537 (N_11537,N_8927,N_9838);
nor U11538 (N_11538,N_8408,N_8470);
nand U11539 (N_11539,N_8787,N_8690);
nand U11540 (N_11540,N_8543,N_9691);
xnor U11541 (N_11541,N_9099,N_9734);
or U11542 (N_11542,N_9434,N_8601);
nand U11543 (N_11543,N_9428,N_8738);
nand U11544 (N_11544,N_8310,N_9289);
nand U11545 (N_11545,N_9799,N_9072);
or U11546 (N_11546,N_9764,N_9604);
or U11547 (N_11547,N_8793,N_8445);
and U11548 (N_11548,N_8910,N_9658);
or U11549 (N_11549,N_8997,N_8025);
nor U11550 (N_11550,N_8183,N_9712);
nor U11551 (N_11551,N_8611,N_8204);
and U11552 (N_11552,N_8633,N_9252);
or U11553 (N_11553,N_8455,N_8707);
nand U11554 (N_11554,N_9655,N_9761);
and U11555 (N_11555,N_8498,N_9086);
xor U11556 (N_11556,N_8391,N_9678);
and U11557 (N_11557,N_8180,N_9681);
xnor U11558 (N_11558,N_8098,N_9608);
nor U11559 (N_11559,N_8186,N_9807);
nand U11560 (N_11560,N_8358,N_8731);
or U11561 (N_11561,N_8426,N_9785);
nand U11562 (N_11562,N_8477,N_9870);
or U11563 (N_11563,N_8919,N_9918);
nor U11564 (N_11564,N_8129,N_8164);
nor U11565 (N_11565,N_9980,N_9864);
nor U11566 (N_11566,N_9520,N_8432);
nor U11567 (N_11567,N_9540,N_9442);
xnor U11568 (N_11568,N_8999,N_9754);
nor U11569 (N_11569,N_8733,N_9965);
xor U11570 (N_11570,N_8755,N_9993);
nand U11571 (N_11571,N_8997,N_8401);
or U11572 (N_11572,N_8986,N_9536);
nor U11573 (N_11573,N_8827,N_8635);
xnor U11574 (N_11574,N_9943,N_9864);
or U11575 (N_11575,N_9589,N_8397);
or U11576 (N_11576,N_9161,N_8576);
or U11577 (N_11577,N_9766,N_9357);
and U11578 (N_11578,N_9372,N_9753);
nand U11579 (N_11579,N_8235,N_9423);
and U11580 (N_11580,N_8853,N_8527);
or U11581 (N_11581,N_9236,N_9597);
nor U11582 (N_11582,N_9426,N_9590);
nor U11583 (N_11583,N_9798,N_9240);
or U11584 (N_11584,N_8495,N_8180);
nor U11585 (N_11585,N_9602,N_9411);
nor U11586 (N_11586,N_9601,N_9487);
or U11587 (N_11587,N_9172,N_9838);
xnor U11588 (N_11588,N_9558,N_9750);
and U11589 (N_11589,N_8573,N_9888);
or U11590 (N_11590,N_9939,N_9899);
nor U11591 (N_11591,N_9005,N_8644);
xor U11592 (N_11592,N_9741,N_8669);
or U11593 (N_11593,N_8335,N_9049);
nor U11594 (N_11594,N_9987,N_9703);
nand U11595 (N_11595,N_8653,N_8028);
xor U11596 (N_11596,N_9781,N_8704);
xor U11597 (N_11597,N_9051,N_9403);
xor U11598 (N_11598,N_9024,N_9723);
and U11599 (N_11599,N_8245,N_8328);
nand U11600 (N_11600,N_9898,N_8440);
nand U11601 (N_11601,N_8475,N_9549);
nor U11602 (N_11602,N_9075,N_8280);
nor U11603 (N_11603,N_9816,N_8645);
nand U11604 (N_11604,N_8013,N_9848);
nor U11605 (N_11605,N_9145,N_8715);
xor U11606 (N_11606,N_8323,N_9465);
xor U11607 (N_11607,N_8427,N_9435);
nand U11608 (N_11608,N_9570,N_9729);
nor U11609 (N_11609,N_9062,N_9409);
and U11610 (N_11610,N_9727,N_8602);
xnor U11611 (N_11611,N_9094,N_9778);
nand U11612 (N_11612,N_8974,N_8259);
xor U11613 (N_11613,N_9273,N_8963);
or U11614 (N_11614,N_9641,N_8987);
and U11615 (N_11615,N_9744,N_8916);
nor U11616 (N_11616,N_9699,N_8039);
nand U11617 (N_11617,N_8357,N_8432);
or U11618 (N_11618,N_8995,N_9187);
or U11619 (N_11619,N_8982,N_8832);
or U11620 (N_11620,N_9692,N_8832);
xnor U11621 (N_11621,N_9056,N_9260);
nor U11622 (N_11622,N_9337,N_8506);
and U11623 (N_11623,N_9398,N_9546);
nor U11624 (N_11624,N_8220,N_9013);
or U11625 (N_11625,N_8325,N_8032);
nor U11626 (N_11626,N_8943,N_9822);
xnor U11627 (N_11627,N_8339,N_8038);
or U11628 (N_11628,N_8093,N_8098);
nor U11629 (N_11629,N_8324,N_8906);
and U11630 (N_11630,N_9574,N_8641);
xor U11631 (N_11631,N_9450,N_8561);
and U11632 (N_11632,N_9858,N_9660);
nand U11633 (N_11633,N_8576,N_8093);
and U11634 (N_11634,N_9326,N_9318);
nand U11635 (N_11635,N_9481,N_9230);
and U11636 (N_11636,N_9692,N_9646);
and U11637 (N_11637,N_8445,N_8219);
nand U11638 (N_11638,N_9146,N_8114);
and U11639 (N_11639,N_9847,N_8833);
nand U11640 (N_11640,N_8950,N_8311);
nand U11641 (N_11641,N_9270,N_9089);
nor U11642 (N_11642,N_9554,N_8805);
nand U11643 (N_11643,N_9118,N_8293);
nand U11644 (N_11644,N_8922,N_8657);
and U11645 (N_11645,N_8923,N_9883);
nor U11646 (N_11646,N_8577,N_8101);
and U11647 (N_11647,N_9584,N_9412);
nor U11648 (N_11648,N_8953,N_9153);
and U11649 (N_11649,N_8599,N_8966);
xor U11650 (N_11650,N_8072,N_9252);
xor U11651 (N_11651,N_9752,N_8342);
or U11652 (N_11652,N_9459,N_8968);
or U11653 (N_11653,N_8849,N_9794);
nand U11654 (N_11654,N_8136,N_9813);
and U11655 (N_11655,N_9356,N_8056);
nor U11656 (N_11656,N_8843,N_9523);
nand U11657 (N_11657,N_9421,N_9891);
xnor U11658 (N_11658,N_9789,N_8387);
nand U11659 (N_11659,N_9957,N_9030);
xnor U11660 (N_11660,N_9887,N_8072);
xnor U11661 (N_11661,N_8355,N_9397);
nand U11662 (N_11662,N_8165,N_9071);
nor U11663 (N_11663,N_8313,N_8384);
or U11664 (N_11664,N_8729,N_9589);
or U11665 (N_11665,N_9962,N_9816);
nand U11666 (N_11666,N_9068,N_8708);
and U11667 (N_11667,N_8092,N_8814);
or U11668 (N_11668,N_8699,N_9900);
xor U11669 (N_11669,N_8827,N_8893);
xnor U11670 (N_11670,N_9727,N_9408);
xor U11671 (N_11671,N_8264,N_9262);
nor U11672 (N_11672,N_8437,N_8088);
and U11673 (N_11673,N_9188,N_9119);
nor U11674 (N_11674,N_8538,N_8556);
and U11675 (N_11675,N_8982,N_8477);
or U11676 (N_11676,N_8018,N_8527);
nor U11677 (N_11677,N_8548,N_8206);
xnor U11678 (N_11678,N_9412,N_8914);
xnor U11679 (N_11679,N_8078,N_9362);
and U11680 (N_11680,N_8024,N_9004);
nand U11681 (N_11681,N_9544,N_9668);
and U11682 (N_11682,N_9277,N_8257);
nor U11683 (N_11683,N_9268,N_9935);
and U11684 (N_11684,N_9650,N_8172);
and U11685 (N_11685,N_9056,N_8838);
nor U11686 (N_11686,N_8034,N_8146);
xnor U11687 (N_11687,N_9480,N_9520);
nand U11688 (N_11688,N_8750,N_8415);
nor U11689 (N_11689,N_8887,N_8959);
xnor U11690 (N_11690,N_9687,N_8648);
and U11691 (N_11691,N_9928,N_9450);
xnor U11692 (N_11692,N_8928,N_8439);
xnor U11693 (N_11693,N_9919,N_8062);
or U11694 (N_11694,N_9415,N_9532);
or U11695 (N_11695,N_8195,N_9968);
xor U11696 (N_11696,N_8425,N_8991);
nand U11697 (N_11697,N_8994,N_8428);
or U11698 (N_11698,N_9707,N_9749);
or U11699 (N_11699,N_9167,N_9185);
and U11700 (N_11700,N_8801,N_8237);
or U11701 (N_11701,N_8795,N_9562);
xnor U11702 (N_11702,N_8124,N_9422);
or U11703 (N_11703,N_8648,N_9392);
nand U11704 (N_11704,N_9652,N_9065);
xor U11705 (N_11705,N_8317,N_9218);
nor U11706 (N_11706,N_9592,N_8456);
nor U11707 (N_11707,N_8437,N_8441);
xnor U11708 (N_11708,N_9077,N_9576);
nand U11709 (N_11709,N_9243,N_9307);
and U11710 (N_11710,N_8766,N_9620);
or U11711 (N_11711,N_8449,N_9880);
nor U11712 (N_11712,N_8796,N_9163);
and U11713 (N_11713,N_8270,N_8706);
or U11714 (N_11714,N_8551,N_9368);
nor U11715 (N_11715,N_8361,N_8384);
nand U11716 (N_11716,N_8661,N_8214);
xor U11717 (N_11717,N_8656,N_8339);
and U11718 (N_11718,N_9478,N_9951);
and U11719 (N_11719,N_8662,N_9591);
or U11720 (N_11720,N_8794,N_8915);
nand U11721 (N_11721,N_9409,N_8884);
nor U11722 (N_11722,N_9709,N_8374);
and U11723 (N_11723,N_8614,N_8054);
nand U11724 (N_11724,N_9274,N_9961);
xnor U11725 (N_11725,N_9653,N_8862);
xnor U11726 (N_11726,N_9377,N_8616);
nand U11727 (N_11727,N_9056,N_8289);
and U11728 (N_11728,N_9255,N_9925);
nor U11729 (N_11729,N_8746,N_8988);
nor U11730 (N_11730,N_8919,N_9364);
xnor U11731 (N_11731,N_9459,N_9546);
or U11732 (N_11732,N_9752,N_8056);
nand U11733 (N_11733,N_8140,N_9546);
and U11734 (N_11734,N_9645,N_8199);
or U11735 (N_11735,N_8618,N_9022);
nand U11736 (N_11736,N_9689,N_8948);
xnor U11737 (N_11737,N_9278,N_9842);
nand U11738 (N_11738,N_8107,N_9085);
or U11739 (N_11739,N_9057,N_9341);
nand U11740 (N_11740,N_8337,N_9824);
nand U11741 (N_11741,N_9126,N_9283);
nand U11742 (N_11742,N_9133,N_8758);
nand U11743 (N_11743,N_9949,N_8496);
nand U11744 (N_11744,N_8749,N_8280);
and U11745 (N_11745,N_8159,N_8836);
and U11746 (N_11746,N_8705,N_8238);
or U11747 (N_11747,N_9656,N_8822);
xnor U11748 (N_11748,N_9551,N_8627);
xor U11749 (N_11749,N_9155,N_8360);
nand U11750 (N_11750,N_8877,N_9564);
and U11751 (N_11751,N_8269,N_9246);
nor U11752 (N_11752,N_8072,N_8098);
xnor U11753 (N_11753,N_8427,N_8563);
and U11754 (N_11754,N_8159,N_8271);
and U11755 (N_11755,N_8494,N_9309);
xnor U11756 (N_11756,N_8358,N_9311);
nand U11757 (N_11757,N_9762,N_8356);
nand U11758 (N_11758,N_8579,N_8133);
nand U11759 (N_11759,N_9349,N_9430);
nor U11760 (N_11760,N_8719,N_8145);
xnor U11761 (N_11761,N_8325,N_9547);
xnor U11762 (N_11762,N_8951,N_9623);
nor U11763 (N_11763,N_9604,N_8220);
or U11764 (N_11764,N_8973,N_8696);
or U11765 (N_11765,N_8947,N_9609);
nor U11766 (N_11766,N_8528,N_9888);
and U11767 (N_11767,N_9708,N_9670);
or U11768 (N_11768,N_9491,N_8443);
and U11769 (N_11769,N_9054,N_8298);
nand U11770 (N_11770,N_8065,N_8516);
nand U11771 (N_11771,N_9012,N_8265);
nand U11772 (N_11772,N_8520,N_8566);
nor U11773 (N_11773,N_8079,N_9442);
nor U11774 (N_11774,N_9044,N_8027);
xor U11775 (N_11775,N_9855,N_9443);
nand U11776 (N_11776,N_9123,N_9729);
nor U11777 (N_11777,N_9624,N_9847);
and U11778 (N_11778,N_9343,N_8539);
or U11779 (N_11779,N_9516,N_8461);
nor U11780 (N_11780,N_9735,N_8162);
or U11781 (N_11781,N_9860,N_8199);
xor U11782 (N_11782,N_9291,N_8131);
nand U11783 (N_11783,N_9915,N_9908);
nor U11784 (N_11784,N_9335,N_9437);
xor U11785 (N_11785,N_8284,N_8853);
and U11786 (N_11786,N_9550,N_8322);
xnor U11787 (N_11787,N_9373,N_8450);
or U11788 (N_11788,N_8296,N_9828);
nor U11789 (N_11789,N_9215,N_9937);
xor U11790 (N_11790,N_9479,N_9455);
nor U11791 (N_11791,N_9070,N_9588);
or U11792 (N_11792,N_9425,N_8850);
or U11793 (N_11793,N_8195,N_8601);
and U11794 (N_11794,N_8232,N_9248);
nor U11795 (N_11795,N_8443,N_9852);
or U11796 (N_11796,N_8322,N_8851);
or U11797 (N_11797,N_8668,N_8077);
xnor U11798 (N_11798,N_9451,N_9483);
xnor U11799 (N_11799,N_9579,N_9417);
or U11800 (N_11800,N_8644,N_8871);
xnor U11801 (N_11801,N_9740,N_9237);
and U11802 (N_11802,N_9864,N_8804);
or U11803 (N_11803,N_8689,N_9132);
or U11804 (N_11804,N_8398,N_9173);
nor U11805 (N_11805,N_8595,N_8145);
or U11806 (N_11806,N_8418,N_8742);
or U11807 (N_11807,N_9610,N_8997);
xnor U11808 (N_11808,N_8474,N_8711);
xor U11809 (N_11809,N_9212,N_9867);
nor U11810 (N_11810,N_8570,N_9280);
and U11811 (N_11811,N_9092,N_8131);
nor U11812 (N_11812,N_8131,N_9412);
xnor U11813 (N_11813,N_9749,N_8079);
and U11814 (N_11814,N_9419,N_9065);
nor U11815 (N_11815,N_8860,N_8146);
nor U11816 (N_11816,N_9715,N_8659);
xnor U11817 (N_11817,N_9461,N_9124);
or U11818 (N_11818,N_8362,N_9615);
or U11819 (N_11819,N_8591,N_9329);
xor U11820 (N_11820,N_9597,N_9132);
or U11821 (N_11821,N_8549,N_8267);
or U11822 (N_11822,N_9828,N_9699);
or U11823 (N_11823,N_8344,N_9099);
xor U11824 (N_11824,N_8395,N_8394);
nand U11825 (N_11825,N_8851,N_8623);
xnor U11826 (N_11826,N_8465,N_9648);
nand U11827 (N_11827,N_9903,N_8143);
and U11828 (N_11828,N_9608,N_8026);
or U11829 (N_11829,N_9732,N_8988);
or U11830 (N_11830,N_8005,N_8317);
and U11831 (N_11831,N_8692,N_8309);
nand U11832 (N_11832,N_8982,N_9475);
and U11833 (N_11833,N_9569,N_9882);
nand U11834 (N_11834,N_9021,N_8402);
and U11835 (N_11835,N_8495,N_9740);
and U11836 (N_11836,N_8733,N_9345);
xor U11837 (N_11837,N_8930,N_8949);
xor U11838 (N_11838,N_9758,N_9468);
nand U11839 (N_11839,N_8455,N_9484);
and U11840 (N_11840,N_9561,N_8836);
and U11841 (N_11841,N_9519,N_8237);
nor U11842 (N_11842,N_8108,N_8091);
and U11843 (N_11843,N_8677,N_9349);
and U11844 (N_11844,N_9161,N_8281);
or U11845 (N_11845,N_9878,N_9943);
or U11846 (N_11846,N_9429,N_8668);
nor U11847 (N_11847,N_8021,N_9555);
or U11848 (N_11848,N_9958,N_8631);
xnor U11849 (N_11849,N_9210,N_8838);
and U11850 (N_11850,N_9090,N_9186);
nor U11851 (N_11851,N_9698,N_9481);
nand U11852 (N_11852,N_9906,N_9284);
xnor U11853 (N_11853,N_9001,N_8857);
xnor U11854 (N_11854,N_8570,N_9605);
nor U11855 (N_11855,N_9303,N_8058);
nand U11856 (N_11856,N_8745,N_9401);
and U11857 (N_11857,N_8614,N_9879);
xor U11858 (N_11858,N_8636,N_8439);
xor U11859 (N_11859,N_9972,N_9537);
nor U11860 (N_11860,N_9834,N_8171);
nand U11861 (N_11861,N_9865,N_9439);
nor U11862 (N_11862,N_8737,N_9667);
and U11863 (N_11863,N_9253,N_9307);
nand U11864 (N_11864,N_8692,N_8820);
nor U11865 (N_11865,N_8427,N_9607);
nor U11866 (N_11866,N_8878,N_8921);
nor U11867 (N_11867,N_9505,N_8116);
or U11868 (N_11868,N_9230,N_9959);
nand U11869 (N_11869,N_8810,N_8186);
or U11870 (N_11870,N_8106,N_8055);
nor U11871 (N_11871,N_9886,N_9571);
and U11872 (N_11872,N_9458,N_8933);
or U11873 (N_11873,N_8769,N_9783);
nor U11874 (N_11874,N_9145,N_9774);
or U11875 (N_11875,N_8249,N_9911);
nand U11876 (N_11876,N_9784,N_8458);
nor U11877 (N_11877,N_8751,N_9270);
nand U11878 (N_11878,N_9944,N_8282);
nor U11879 (N_11879,N_9165,N_9608);
xnor U11880 (N_11880,N_8901,N_9261);
nor U11881 (N_11881,N_9916,N_8563);
nor U11882 (N_11882,N_9385,N_8428);
and U11883 (N_11883,N_9754,N_9377);
or U11884 (N_11884,N_8472,N_9511);
and U11885 (N_11885,N_8911,N_8636);
nand U11886 (N_11886,N_9026,N_8003);
nor U11887 (N_11887,N_9353,N_8046);
nand U11888 (N_11888,N_9251,N_8289);
or U11889 (N_11889,N_8624,N_9200);
xnor U11890 (N_11890,N_8094,N_9573);
nand U11891 (N_11891,N_8670,N_9635);
xnor U11892 (N_11892,N_9268,N_8215);
nand U11893 (N_11893,N_8996,N_9932);
nand U11894 (N_11894,N_8109,N_9239);
xor U11895 (N_11895,N_8765,N_8164);
xnor U11896 (N_11896,N_9248,N_9504);
or U11897 (N_11897,N_8574,N_9178);
xor U11898 (N_11898,N_9335,N_8591);
nor U11899 (N_11899,N_9259,N_8841);
xnor U11900 (N_11900,N_8065,N_8148);
xnor U11901 (N_11901,N_9250,N_8484);
xnor U11902 (N_11902,N_8022,N_9814);
and U11903 (N_11903,N_8530,N_8858);
or U11904 (N_11904,N_9967,N_9686);
and U11905 (N_11905,N_9792,N_8528);
and U11906 (N_11906,N_9268,N_8049);
and U11907 (N_11907,N_8072,N_8199);
and U11908 (N_11908,N_8820,N_8867);
nand U11909 (N_11909,N_8087,N_8343);
nor U11910 (N_11910,N_9682,N_8100);
nand U11911 (N_11911,N_8137,N_8606);
and U11912 (N_11912,N_9534,N_8020);
and U11913 (N_11913,N_9486,N_9645);
and U11914 (N_11914,N_8113,N_8854);
and U11915 (N_11915,N_9713,N_8190);
nor U11916 (N_11916,N_8222,N_9436);
or U11917 (N_11917,N_9817,N_8865);
nand U11918 (N_11918,N_8413,N_8915);
xor U11919 (N_11919,N_9596,N_9080);
nor U11920 (N_11920,N_8877,N_9714);
xor U11921 (N_11921,N_9794,N_8189);
nand U11922 (N_11922,N_9774,N_9251);
nor U11923 (N_11923,N_8015,N_8055);
or U11924 (N_11924,N_8704,N_8784);
nor U11925 (N_11925,N_8194,N_9873);
nor U11926 (N_11926,N_8361,N_9982);
nand U11927 (N_11927,N_9647,N_9310);
nand U11928 (N_11928,N_8830,N_8553);
xor U11929 (N_11929,N_9221,N_9250);
xor U11930 (N_11930,N_8490,N_8502);
and U11931 (N_11931,N_9468,N_9860);
or U11932 (N_11932,N_8164,N_8363);
xnor U11933 (N_11933,N_8200,N_9734);
xnor U11934 (N_11934,N_8615,N_9547);
nand U11935 (N_11935,N_9568,N_9214);
nor U11936 (N_11936,N_9438,N_8178);
nand U11937 (N_11937,N_8919,N_8528);
xnor U11938 (N_11938,N_8139,N_9280);
nand U11939 (N_11939,N_9998,N_8032);
and U11940 (N_11940,N_9724,N_8194);
or U11941 (N_11941,N_9933,N_9807);
nand U11942 (N_11942,N_8251,N_9272);
and U11943 (N_11943,N_8326,N_8088);
xnor U11944 (N_11944,N_8826,N_8981);
nor U11945 (N_11945,N_9569,N_9082);
nor U11946 (N_11946,N_8285,N_9256);
and U11947 (N_11947,N_9174,N_9536);
and U11948 (N_11948,N_8833,N_8878);
nand U11949 (N_11949,N_9036,N_8655);
nor U11950 (N_11950,N_8644,N_9159);
nand U11951 (N_11951,N_9728,N_8422);
or U11952 (N_11952,N_8201,N_9819);
xnor U11953 (N_11953,N_8426,N_9489);
xnor U11954 (N_11954,N_8252,N_8135);
nand U11955 (N_11955,N_8582,N_9423);
nor U11956 (N_11956,N_8053,N_9840);
nand U11957 (N_11957,N_8402,N_9838);
and U11958 (N_11958,N_8216,N_9164);
nand U11959 (N_11959,N_9011,N_8592);
or U11960 (N_11960,N_9889,N_9975);
and U11961 (N_11961,N_9351,N_9410);
nand U11962 (N_11962,N_9840,N_9023);
and U11963 (N_11963,N_9195,N_8924);
xor U11964 (N_11964,N_8495,N_8355);
xnor U11965 (N_11965,N_9683,N_9355);
nand U11966 (N_11966,N_8493,N_8944);
and U11967 (N_11967,N_9199,N_8854);
xor U11968 (N_11968,N_8026,N_9809);
nor U11969 (N_11969,N_9355,N_9671);
or U11970 (N_11970,N_9347,N_8565);
xnor U11971 (N_11971,N_8711,N_8456);
or U11972 (N_11972,N_8259,N_9159);
nand U11973 (N_11973,N_8212,N_9808);
nand U11974 (N_11974,N_9714,N_8186);
nor U11975 (N_11975,N_9668,N_9084);
xor U11976 (N_11976,N_9170,N_9999);
xor U11977 (N_11977,N_9753,N_9199);
and U11978 (N_11978,N_9906,N_9374);
nor U11979 (N_11979,N_9537,N_9722);
nor U11980 (N_11980,N_8511,N_9574);
and U11981 (N_11981,N_9742,N_8728);
nand U11982 (N_11982,N_9429,N_8942);
and U11983 (N_11983,N_8433,N_9270);
and U11984 (N_11984,N_8530,N_9724);
nor U11985 (N_11985,N_8805,N_8231);
nor U11986 (N_11986,N_9355,N_8444);
and U11987 (N_11987,N_8003,N_8989);
nor U11988 (N_11988,N_8740,N_9668);
nand U11989 (N_11989,N_8003,N_9260);
and U11990 (N_11990,N_8786,N_8344);
xor U11991 (N_11991,N_8648,N_8092);
or U11992 (N_11992,N_8182,N_8706);
nor U11993 (N_11993,N_8032,N_8301);
and U11994 (N_11994,N_8297,N_8234);
nand U11995 (N_11995,N_9883,N_8500);
xnor U11996 (N_11996,N_8588,N_9202);
nand U11997 (N_11997,N_8536,N_9143);
or U11998 (N_11998,N_8074,N_8446);
nor U11999 (N_11999,N_8361,N_9487);
nor U12000 (N_12000,N_10828,N_10421);
or U12001 (N_12001,N_10170,N_11009);
xor U12002 (N_12002,N_11288,N_10533);
xor U12003 (N_12003,N_11097,N_10371);
or U12004 (N_12004,N_10603,N_11683);
and U12005 (N_12005,N_11643,N_10723);
xor U12006 (N_12006,N_10680,N_11614);
and U12007 (N_12007,N_10472,N_10040);
xor U12008 (N_12008,N_10720,N_10638);
nor U12009 (N_12009,N_11974,N_11223);
or U12010 (N_12010,N_10279,N_11134);
xnor U12011 (N_12011,N_10233,N_11360);
xnor U12012 (N_12012,N_11822,N_11914);
and U12013 (N_12013,N_11273,N_10963);
xor U12014 (N_12014,N_11890,N_10481);
or U12015 (N_12015,N_11606,N_10399);
xnor U12016 (N_12016,N_10731,N_10975);
or U12017 (N_12017,N_10599,N_11029);
and U12018 (N_12018,N_10899,N_11429);
nand U12019 (N_12019,N_11777,N_11850);
xor U12020 (N_12020,N_11151,N_10686);
and U12021 (N_12021,N_10302,N_11607);
nor U12022 (N_12022,N_10778,N_10684);
nand U12023 (N_12023,N_11031,N_11070);
and U12024 (N_12024,N_10570,N_10910);
or U12025 (N_12025,N_11506,N_11855);
and U12026 (N_12026,N_11560,N_11141);
nand U12027 (N_12027,N_11025,N_11576);
nor U12028 (N_12028,N_11086,N_11329);
xor U12029 (N_12029,N_10922,N_10550);
or U12030 (N_12030,N_10206,N_10678);
nor U12031 (N_12031,N_11917,N_10810);
nand U12032 (N_12032,N_10775,N_10500);
or U12033 (N_12033,N_10077,N_10508);
nand U12034 (N_12034,N_10306,N_11509);
nor U12035 (N_12035,N_10955,N_11381);
nor U12036 (N_12036,N_11051,N_11030);
xor U12037 (N_12037,N_10033,N_11886);
xnor U12038 (N_12038,N_10543,N_11748);
nand U12039 (N_12039,N_10613,N_11236);
nor U12040 (N_12040,N_10597,N_10107);
nor U12041 (N_12041,N_11512,N_11922);
xnor U12042 (N_12042,N_11274,N_10877);
or U12043 (N_12043,N_10983,N_10323);
nor U12044 (N_12044,N_11763,N_11037);
and U12045 (N_12045,N_11722,N_10585);
nor U12046 (N_12046,N_11286,N_11148);
nor U12047 (N_12047,N_11760,N_10200);
and U12048 (N_12048,N_11513,N_10735);
nand U12049 (N_12049,N_11658,N_11289);
nor U12050 (N_12050,N_11883,N_11004);
or U12051 (N_12051,N_11552,N_10278);
xor U12052 (N_12052,N_10711,N_10788);
or U12053 (N_12053,N_10820,N_10960);
nand U12054 (N_12054,N_10900,N_10166);
nand U12055 (N_12055,N_11706,N_10795);
xor U12056 (N_12056,N_11965,N_11093);
or U12057 (N_12057,N_10574,N_11232);
nor U12058 (N_12058,N_11282,N_11324);
and U12059 (N_12059,N_11740,N_11448);
xnor U12060 (N_12060,N_11171,N_11889);
or U12061 (N_12061,N_11519,N_10930);
xor U12062 (N_12062,N_10636,N_10458);
xor U12063 (N_12063,N_10642,N_11444);
xnor U12064 (N_12064,N_10477,N_11674);
and U12065 (N_12065,N_10700,N_11712);
nand U12066 (N_12066,N_11612,N_10903);
and U12067 (N_12067,N_10297,N_11830);
nand U12068 (N_12068,N_11986,N_10448);
nor U12069 (N_12069,N_10027,N_10892);
and U12070 (N_12070,N_10282,N_10805);
or U12071 (N_12071,N_10252,N_10881);
xor U12072 (N_12072,N_10016,N_11087);
xnor U12073 (N_12073,N_11348,N_11871);
nand U12074 (N_12074,N_10005,N_11691);
xor U12075 (N_12075,N_11005,N_11493);
or U12076 (N_12076,N_11189,N_11931);
and U12077 (N_12077,N_11632,N_10049);
nor U12078 (N_12078,N_11060,N_11530);
nor U12079 (N_12079,N_10338,N_11131);
nand U12080 (N_12080,N_11563,N_10274);
nor U12081 (N_12081,N_11388,N_11692);
or U12082 (N_12082,N_10014,N_10105);
nand U12083 (N_12083,N_11392,N_11017);
nand U12084 (N_12084,N_11610,N_11019);
and U12085 (N_12085,N_10978,N_11697);
nor U12086 (N_12086,N_10835,N_11230);
nand U12087 (N_12087,N_11210,N_10567);
nand U12088 (N_12088,N_10495,N_11968);
nor U12089 (N_12089,N_10346,N_10093);
and U12090 (N_12090,N_11858,N_10670);
and U12091 (N_12091,N_11000,N_10487);
or U12092 (N_12092,N_10359,N_10773);
and U12093 (N_12093,N_10668,N_11852);
and U12094 (N_12094,N_10406,N_10476);
nor U12095 (N_12095,N_11245,N_11778);
and U12096 (N_12096,N_10794,N_10737);
or U12097 (N_12097,N_11870,N_11417);
or U12098 (N_12098,N_11894,N_10544);
nor U12099 (N_12099,N_10347,N_11196);
and U12100 (N_12100,N_10416,N_10557);
xnor U12101 (N_12101,N_11897,N_11735);
xnor U12102 (N_12102,N_10579,N_10020);
or U12103 (N_12103,N_10609,N_10784);
nand U12104 (N_12104,N_11336,N_10848);
and U12105 (N_12105,N_11895,N_11088);
nor U12106 (N_12106,N_10119,N_10325);
or U12107 (N_12107,N_10473,N_10854);
xor U12108 (N_12108,N_11875,N_10520);
and U12109 (N_12109,N_11995,N_11626);
nor U12110 (N_12110,N_11184,N_10661);
xor U12111 (N_12111,N_10488,N_10867);
nor U12112 (N_12112,N_10149,N_11363);
nor U12113 (N_12113,N_11954,N_10761);
and U12114 (N_12114,N_11075,N_11020);
or U12115 (N_12115,N_10439,N_11385);
nand U12116 (N_12116,N_11755,N_11212);
nand U12117 (N_12117,N_10189,N_11055);
xnor U12118 (N_12118,N_10965,N_10205);
and U12119 (N_12119,N_10808,N_10839);
nand U12120 (N_12120,N_11789,N_11709);
nor U12121 (N_12121,N_10156,N_10845);
nand U12122 (N_12122,N_10202,N_11793);
nand U12123 (N_12123,N_10169,N_10409);
and U12124 (N_12124,N_11843,N_10234);
nand U12125 (N_12125,N_10351,N_11977);
nor U12126 (N_12126,N_10260,N_11222);
and U12127 (N_12127,N_11957,N_10485);
xnor U12128 (N_12128,N_11690,N_11938);
xnor U12129 (N_12129,N_10886,N_11040);
or U12130 (N_12130,N_10130,N_11911);
nor U12131 (N_12131,N_11711,N_11412);
nor U12132 (N_12132,N_11164,N_11350);
or U12133 (N_12133,N_10298,N_10894);
nand U12134 (N_12134,N_10693,N_10694);
xor U12135 (N_12135,N_11540,N_10937);
xor U12136 (N_12136,N_10368,N_11076);
nand U12137 (N_12137,N_11400,N_11034);
and U12138 (N_12138,N_10938,N_11062);
or U12139 (N_12139,N_11061,N_11584);
nand U12140 (N_12140,N_10046,N_11045);
or U12141 (N_12141,N_11090,N_11744);
and U12142 (N_12142,N_10378,N_10531);
xnor U12143 (N_12143,N_11853,N_11701);
nand U12144 (N_12144,N_11165,N_11065);
nand U12145 (N_12145,N_11577,N_10159);
xor U12146 (N_12146,N_11338,N_11963);
xor U12147 (N_12147,N_11550,N_11026);
or U12148 (N_12148,N_10669,N_10022);
and U12149 (N_12149,N_11799,N_10390);
or U12150 (N_12150,N_11473,N_11140);
or U12151 (N_12151,N_10583,N_11564);
xor U12152 (N_12152,N_10984,N_10792);
nand U12153 (N_12153,N_11535,N_10685);
xor U12154 (N_12154,N_11885,N_11556);
nand U12155 (N_12155,N_11526,N_10198);
and U12156 (N_12156,N_11561,N_11152);
and U12157 (N_12157,N_11592,N_11934);
nor U12158 (N_12158,N_11450,N_11228);
or U12159 (N_12159,N_10941,N_10893);
or U12160 (N_12160,N_11961,N_11155);
or U12161 (N_12161,N_11893,N_10836);
nand U12162 (N_12162,N_11107,N_11206);
nor U12163 (N_12163,N_11117,N_11108);
or U12164 (N_12164,N_11868,N_11896);
or U12165 (N_12165,N_10920,N_10499);
nor U12166 (N_12166,N_11100,N_10086);
and U12167 (N_12167,N_10847,N_10355);
or U12168 (N_12168,N_11531,N_11415);
or U12169 (N_12169,N_10629,N_10450);
and U12170 (N_12170,N_11575,N_10092);
xor U12171 (N_12171,N_11379,N_11081);
and U12172 (N_12172,N_11249,N_11723);
and U12173 (N_12173,N_11525,N_10837);
nand U12174 (N_12174,N_11094,N_11546);
nand U12175 (N_12175,N_10729,N_10185);
xnor U12176 (N_12176,N_11772,N_11199);
or U12177 (N_12177,N_10561,N_10463);
nor U12178 (N_12178,N_11484,N_10454);
nand U12179 (N_12179,N_10045,N_10316);
nor U12180 (N_12180,N_10004,N_11605);
xor U12181 (N_12181,N_10687,N_10840);
nand U12182 (N_12182,N_10691,N_10842);
nor U12183 (N_12183,N_10075,N_11826);
xnor U12184 (N_12184,N_11660,N_11817);
xor U12185 (N_12185,N_10326,N_10556);
or U12186 (N_12186,N_11635,N_10709);
and U12187 (N_12187,N_11972,N_11949);
nor U12188 (N_12188,N_10523,N_10770);
and U12189 (N_12189,N_10757,N_10580);
and U12190 (N_12190,N_10374,N_11554);
and U12191 (N_12191,N_11451,N_10021);
nand U12192 (N_12192,N_10857,N_11630);
or U12193 (N_12193,N_10340,N_11290);
and U12194 (N_12194,N_11470,N_11838);
nor U12195 (N_12195,N_11765,N_11064);
and U12196 (N_12196,N_10587,N_11204);
or U12197 (N_12197,N_11686,N_10541);
and U12198 (N_12198,N_11133,N_10428);
nor U12199 (N_12199,N_10874,N_10235);
xor U12200 (N_12200,N_11758,N_10422);
xnor U12201 (N_12201,N_10799,N_10155);
and U12202 (N_12202,N_10578,N_10489);
nand U12203 (N_12203,N_11410,N_10705);
and U12204 (N_12204,N_11042,N_11352);
xnor U12205 (N_12205,N_11035,N_10418);
and U12206 (N_12206,N_10296,N_10214);
and U12207 (N_12207,N_11666,N_11539);
or U12208 (N_12208,N_10446,N_11229);
nand U12209 (N_12209,N_11188,N_11839);
and U12210 (N_12210,N_11437,N_11548);
and U12211 (N_12211,N_10741,N_10364);
xor U12212 (N_12212,N_10644,N_11482);
xor U12213 (N_12213,N_11955,N_11498);
xnor U12214 (N_12214,N_11291,N_11514);
nand U12215 (N_12215,N_10696,N_10436);
xor U12216 (N_12216,N_10923,N_10986);
xnor U12217 (N_12217,N_11559,N_10453);
and U12218 (N_12218,N_10553,N_11021);
or U12219 (N_12219,N_10624,N_11685);
or U12220 (N_12220,N_11303,N_10806);
nand U12221 (N_12221,N_10966,N_10679);
xnor U12222 (N_12222,N_10305,N_10547);
nand U12223 (N_12223,N_10424,N_11589);
and U12224 (N_12224,N_11239,N_10177);
or U12225 (N_12225,N_10209,N_11814);
and U12226 (N_12226,N_10144,N_10442);
nor U12227 (N_12227,N_10562,N_10117);
or U12228 (N_12228,N_11010,N_10370);
nor U12229 (N_12229,N_11840,N_10552);
or U12230 (N_12230,N_11776,N_11447);
xor U12231 (N_12231,N_10250,N_10402);
and U12232 (N_12232,N_11281,N_11664);
nor U12233 (N_12233,N_11816,N_11047);
and U12234 (N_12234,N_10506,N_10315);
nor U12235 (N_12235,N_10514,N_10779);
and U12236 (N_12236,N_11803,N_10431);
nand U12237 (N_12237,N_10111,N_11982);
nand U12238 (N_12238,N_10440,N_11475);
or U12239 (N_12239,N_11594,N_10079);
or U12240 (N_12240,N_11595,N_11295);
xnor U12241 (N_12241,N_11002,N_11497);
or U12242 (N_12242,N_10216,N_10352);
nand U12243 (N_12243,N_11604,N_10755);
nor U12244 (N_12244,N_10878,N_11091);
and U12245 (N_12245,N_11547,N_10555);
or U12246 (N_12246,N_10907,N_11316);
nor U12247 (N_12247,N_11861,N_11203);
nor U12248 (N_12248,N_10611,N_10962);
nand U12249 (N_12249,N_10861,N_10635);
and U12250 (N_12250,N_11993,N_10242);
xnor U12251 (N_12251,N_10362,N_10928);
nand U12252 (N_12252,N_10122,N_10692);
or U12253 (N_12253,N_11636,N_10057);
nand U12254 (N_12254,N_10393,N_10656);
nor U12255 (N_12255,N_11118,N_10262);
or U12256 (N_12256,N_10094,N_10714);
nor U12257 (N_12257,N_11197,N_10002);
or U12258 (N_12258,N_10342,N_11721);
nor U12259 (N_12259,N_11147,N_11537);
nor U12260 (N_12260,N_10558,N_11581);
and U12261 (N_12261,N_11901,N_10379);
nand U12262 (N_12262,N_10645,N_10146);
or U12263 (N_12263,N_10354,N_11084);
and U12264 (N_12264,N_11549,N_11640);
and U12265 (N_12265,N_10751,N_10417);
nor U12266 (N_12266,N_11398,N_10665);
and U12267 (N_12267,N_11714,N_10746);
nor U12268 (N_12268,N_11966,N_11449);
xnor U12269 (N_12269,N_10565,N_10000);
nor U12270 (N_12270,N_10875,N_10754);
or U12271 (N_12271,N_10136,N_11341);
and U12272 (N_12272,N_11695,N_10148);
or U12273 (N_12273,N_11912,N_10332);
xnor U12274 (N_12274,N_11244,N_11737);
nor U12275 (N_12275,N_10151,N_10073);
or U12276 (N_12276,N_10707,N_11041);
nor U12277 (N_12277,N_10162,N_11191);
or U12278 (N_12278,N_10456,N_11225);
nand U12279 (N_12279,N_11616,N_11309);
or U12280 (N_12280,N_11083,N_10249);
and U12281 (N_12281,N_10449,N_10940);
nand U12282 (N_12282,N_10403,N_11728);
nor U12283 (N_12283,N_11190,N_10133);
xor U12284 (N_12284,N_11507,N_11580);
or U12285 (N_12285,N_11574,N_10109);
nand U12286 (N_12286,N_11805,N_10384);
or U12287 (N_12287,N_10138,N_10572);
xor U12288 (N_12288,N_11994,N_10764);
nand U12289 (N_12289,N_10791,N_10884);
and U12290 (N_12290,N_10804,N_10826);
xnor U12291 (N_12291,N_11317,N_11810);
or U12292 (N_12292,N_10267,N_10825);
nand U12293 (N_12293,N_10865,N_10259);
nand U12294 (N_12294,N_11638,N_10116);
and U12295 (N_12295,N_11077,N_10280);
xnor U12296 (N_12296,N_10876,N_10901);
and U12297 (N_12297,N_10082,N_11331);
xnor U12298 (N_12298,N_10108,N_11533);
nor U12299 (N_12299,N_10608,N_11754);
and U12300 (N_12300,N_10942,N_11935);
xnor U12301 (N_12301,N_10672,N_10633);
xor U12302 (N_12302,N_11520,N_10103);
nor U12303 (N_12303,N_11143,N_10659);
xnor U12304 (N_12304,N_10013,N_11371);
xnor U12305 (N_12305,N_10913,N_11058);
and U12306 (N_12306,N_11985,N_10060);
or U12307 (N_12307,N_10433,N_10699);
xor U12308 (N_12308,N_11419,N_10494);
xnor U12309 (N_12309,N_10802,N_11532);
or U12310 (N_12310,N_10927,N_11634);
nor U12311 (N_12311,N_10866,N_11964);
and U12312 (N_12312,N_11434,N_11380);
or U12313 (N_12313,N_10304,N_10361);
or U12314 (N_12314,N_10988,N_11747);
or U12315 (N_12315,N_11401,N_10145);
or U12316 (N_12316,N_11787,N_10977);
nand U12317 (N_12317,N_10911,N_10655);
nor U12318 (N_12318,N_10660,N_11247);
xor U12319 (N_12319,N_11841,N_10382);
nand U12320 (N_12320,N_10733,N_11624);
nor U12321 (N_12321,N_11649,N_10528);
and U12322 (N_12322,N_10841,N_11085);
xnor U12323 (N_12323,N_11168,N_11732);
nand U12324 (N_12324,N_11402,N_11262);
nand U12325 (N_12325,N_11014,N_11794);
nand U12326 (N_12326,N_10851,N_10632);
nor U12327 (N_12327,N_10853,N_11483);
and U12328 (N_12328,N_10178,N_10276);
nor U12329 (N_12329,N_10782,N_10072);
xnor U12330 (N_12330,N_10307,N_11521);
and U12331 (N_12331,N_11588,N_11887);
nor U12332 (N_12332,N_11389,N_10596);
nor U12333 (N_12333,N_10890,N_11137);
xnor U12334 (N_12334,N_10509,N_10657);
nand U12335 (N_12335,N_11569,N_11655);
and U12336 (N_12336,N_11231,N_10623);
or U12337 (N_12337,N_10869,N_11310);
xor U12338 (N_12338,N_10742,N_10879);
xnor U12339 (N_12339,N_11536,N_10519);
nand U12340 (N_12340,N_11491,N_10441);
xor U12341 (N_12341,N_11835,N_11150);
and U12342 (N_12342,N_11541,N_11753);
nor U12343 (N_12343,N_11211,N_10816);
nand U12344 (N_12344,N_10011,N_10760);
or U12345 (N_12345,N_11804,N_11715);
nand U12346 (N_12346,N_10740,N_10525);
nor U12347 (N_12347,N_11471,N_11454);
or U12348 (N_12348,N_10677,N_11718);
or U12349 (N_12349,N_11502,N_10467);
and U12350 (N_12350,N_10465,N_11782);
nand U12351 (N_12351,N_10801,N_10129);
nand U12352 (N_12352,N_11657,N_10445);
nand U12353 (N_12353,N_11725,N_10229);
or U12354 (N_12354,N_10469,N_11136);
nand U12355 (N_12355,N_10211,N_10803);
nor U12356 (N_12356,N_11112,N_11693);
xnor U12357 (N_12357,N_10650,N_10007);
nand U12358 (N_12358,N_10286,N_10386);
nand U12359 (N_12359,N_10993,N_10666);
nor U12360 (N_12360,N_11096,N_10967);
nor U12361 (N_12361,N_10756,N_11662);
nor U12362 (N_12362,N_11873,N_11764);
nand U12363 (N_12363,N_11969,N_10053);
and U12364 (N_12364,N_11233,N_10482);
nand U12365 (N_12365,N_11439,N_11024);
nand U12366 (N_12366,N_11198,N_10961);
xnor U12367 (N_12367,N_10817,N_10154);
xor U12368 (N_12368,N_11499,N_10036);
or U12369 (N_12369,N_11884,N_11611);
or U12370 (N_12370,N_11125,N_10330);
or U12371 (N_12371,N_11749,N_10083);
nor U12372 (N_12372,N_11780,N_10898);
and U12373 (N_12373,N_11771,N_11111);
or U12374 (N_12374,N_10957,N_11302);
or U12375 (N_12375,N_10388,N_10600);
or U12376 (N_12376,N_10947,N_11220);
xnor U12377 (N_12377,N_11330,N_10549);
xnor U12378 (N_12378,N_11266,N_10247);
and U12379 (N_12379,N_10909,N_11218);
or U12380 (N_12380,N_11216,N_11213);
and U12381 (N_12381,N_11393,N_10852);
or U12382 (N_12382,N_11404,N_11932);
nor U12383 (N_12383,N_11105,N_11123);
nor U12384 (N_12384,N_10019,N_11842);
xor U12385 (N_12385,N_10389,N_11790);
and U12386 (N_12386,N_11713,N_11320);
nor U12387 (N_12387,N_11802,N_11877);
or U12388 (N_12388,N_11276,N_11177);
nand U12389 (N_12389,N_10182,N_11593);
xnor U12390 (N_12390,N_10885,N_10979);
xor U12391 (N_12391,N_11242,N_11609);
or U12392 (N_12392,N_10333,N_10767);
nand U12393 (N_12393,N_11347,N_10976);
nand U12394 (N_12394,N_11102,N_10652);
and U12395 (N_12395,N_11126,N_11821);
nand U12396 (N_12396,N_11250,N_10087);
or U12397 (N_12397,N_11494,N_11023);
xnor U12398 (N_12398,N_10241,N_11761);
nand U12399 (N_12399,N_11321,N_10365);
and U12400 (N_12400,N_11261,N_11376);
or U12401 (N_12401,N_11746,N_10532);
nand U12402 (N_12402,N_10176,N_10647);
or U12403 (N_12403,N_11072,N_11872);
and U12404 (N_12404,N_11110,N_10625);
nor U12405 (N_12405,N_11443,N_10950);
xnor U12406 (N_12406,N_11719,N_10998);
or U12407 (N_12407,N_11756,N_10065);
or U12408 (N_12408,N_10524,N_10772);
nor U12409 (N_12409,N_10862,N_10545);
xnor U12410 (N_12410,N_10568,N_11878);
and U12411 (N_12411,N_11903,N_11183);
and U12412 (N_12412,N_10153,N_11620);
or U12413 (N_12413,N_10479,N_10969);
and U12414 (N_12414,N_11278,N_11357);
nor U12415 (N_12415,N_10225,N_10664);
xnor U12416 (N_12416,N_11205,N_11132);
or U12417 (N_12417,N_11708,N_10768);
or U12418 (N_12418,N_11978,N_11488);
nor U12419 (N_12419,N_11054,N_11717);
nand U12420 (N_12420,N_11461,N_10444);
nand U12421 (N_12421,N_11390,N_10777);
xor U12422 (N_12422,N_11769,N_10616);
or U12423 (N_12423,N_11365,N_10595);
nand U12424 (N_12424,N_11166,N_11534);
xor U12425 (N_12425,N_10610,N_10003);
and U12426 (N_12426,N_11435,N_10171);
or U12427 (N_12427,N_11555,N_11775);
and U12428 (N_12428,N_10789,N_11340);
nor U12429 (N_12429,N_10569,N_11372);
xor U12430 (N_12430,N_11207,N_10237);
nor U12431 (N_12431,N_10366,N_11465);
nand U12432 (N_12432,N_10319,N_10023);
xnor U12433 (N_12433,N_11433,N_11059);
and U12434 (N_12434,N_11930,N_11154);
or U12435 (N_12435,N_10367,N_11456);
nor U12436 (N_12436,N_11175,N_11007);
nand U12437 (N_12437,N_11967,N_11268);
nand U12438 (N_12438,N_10673,N_10989);
or U12439 (N_12439,N_11503,N_10968);
nand U12440 (N_12440,N_10076,N_10468);
nand U12441 (N_12441,N_11913,N_10257);
nor U12442 (N_12442,N_10373,N_10098);
and U12443 (N_12443,N_11699,N_11820);
and U12444 (N_12444,N_11163,N_11792);
nor U12445 (N_12445,N_10164,N_11553);
xor U12446 (N_12446,N_11819,N_11335);
xor U12447 (N_12447,N_10486,N_10856);
xnor U12448 (N_12448,N_11436,N_11074);
xor U12449 (N_12449,N_10126,N_10897);
or U12450 (N_12450,N_11867,N_10181);
xnor U12451 (N_12451,N_10201,N_10753);
xnor U12452 (N_12452,N_10849,N_10080);
nor U12453 (N_12453,N_10400,N_11039);
nand U12454 (N_12454,N_11524,N_11353);
and U12455 (N_12455,N_10427,N_11669);
nand U12456 (N_12456,N_11235,N_11384);
or U12457 (N_12457,N_11221,N_11337);
xnor U12458 (N_12458,N_11092,N_11907);
nand U12459 (N_12459,N_11095,N_11022);
nor U12460 (N_12460,N_10415,N_10255);
nor U12461 (N_12461,N_10612,N_10029);
or U12462 (N_12462,N_11418,N_11733);
nor U12463 (N_12463,N_10344,N_10414);
nand U12464 (N_12464,N_11863,N_11325);
nand U12465 (N_12465,N_10398,N_10501);
and U12466 (N_12466,N_10397,N_11891);
and U12467 (N_12467,N_10026,N_10069);
and U12468 (N_12468,N_10478,N_11322);
or U12469 (N_12469,N_10776,N_11496);
xor U12470 (N_12470,N_11942,N_10747);
nand U12471 (N_12471,N_10074,N_10243);
nor U12472 (N_12472,N_11485,N_10762);
nor U12473 (N_12473,N_10648,N_11293);
and U12474 (N_12474,N_11173,N_10534);
nand U12475 (N_12475,N_10739,N_10018);
xor U12476 (N_12476,N_10671,N_11759);
xnor U12477 (N_12477,N_10833,N_10581);
or U12478 (N_12478,N_10999,N_10734);
nand U12479 (N_12479,N_11808,N_11234);
nor U12480 (N_12480,N_10703,N_10576);
xnor U12481 (N_12481,N_10199,N_10459);
or U12482 (N_12482,N_10510,N_11124);
xnor U12483 (N_12483,N_10736,N_10375);
and U12484 (N_12484,N_11675,N_11314);
or U12485 (N_12485,N_10218,N_11921);
xnor U12486 (N_12486,N_10819,N_10035);
and U12487 (N_12487,N_11898,N_10980);
or U12488 (N_12488,N_10091,N_10858);
nor U12489 (N_12489,N_10419,N_10540);
or U12490 (N_12490,N_11187,N_10095);
nand U12491 (N_12491,N_11421,N_10097);
or U12492 (N_12492,N_10443,N_11067);
and U12493 (N_12493,N_10991,N_11424);
and U12494 (N_12494,N_10551,N_11246);
or U12495 (N_12495,N_11343,N_10496);
and U12496 (N_12496,N_11837,N_10724);
and U12497 (N_12497,N_10407,N_10701);
and U12498 (N_12498,N_11618,N_11157);
nand U12499 (N_12499,N_10505,N_10385);
xor U12500 (N_12500,N_11598,N_10051);
xor U12501 (N_12501,N_10193,N_11219);
xor U12502 (N_12502,N_10114,N_10880);
xor U12503 (N_12503,N_10294,N_10815);
nand U12504 (N_12504,N_11926,N_11615);
and U12505 (N_12505,N_11391,N_11694);
or U12506 (N_12506,N_10147,N_11018);
xnor U12507 (N_12507,N_11784,N_10771);
xnor U12508 (N_12508,N_11200,N_10790);
or U12509 (N_12509,N_10032,N_10717);
and U12510 (N_12510,N_11851,N_11573);
xor U12511 (N_12511,N_11720,N_11432);
or U12512 (N_12512,N_11279,N_11215);
and U12513 (N_12513,N_10089,N_11399);
xnor U12514 (N_12514,N_10517,N_11257);
or U12515 (N_12515,N_10589,N_11364);
or U12516 (N_12516,N_10339,N_11910);
nand U12517 (N_12517,N_10504,N_11224);
xor U12518 (N_12518,N_11186,N_10906);
or U12519 (N_12519,N_10824,N_10244);
nand U12520 (N_12520,N_10308,N_10227);
and U12521 (N_12521,N_10377,N_10435);
nand U12522 (N_12522,N_10622,N_10253);
nor U12523 (N_12523,N_10223,N_11989);
or U12524 (N_12524,N_10586,N_10135);
or U12525 (N_12525,N_10059,N_10219);
or U12526 (N_12526,N_11637,N_10123);
nor U12527 (N_12527,N_11752,N_11631);
or U12528 (N_12528,N_11984,N_11710);
nor U12529 (N_12529,N_10827,N_11647);
or U12530 (N_12530,N_10639,N_10598);
nand U12531 (N_12531,N_11738,N_11824);
and U12532 (N_12532,N_10793,N_10522);
nor U12533 (N_12533,N_10285,N_11195);
and U12534 (N_12534,N_10887,N_10264);
or U12535 (N_12535,N_10713,N_11423);
nand U12536 (N_12536,N_11809,N_11676);
xnor U12537 (N_12537,N_11082,N_10704);
nor U12538 (N_12538,N_11900,N_11661);
nor U12539 (N_12539,N_11180,N_10173);
nor U12540 (N_12540,N_10157,N_10337);
nand U12541 (N_12541,N_10054,N_11071);
or U12542 (N_12542,N_10971,N_11476);
nor U12543 (N_12543,N_10100,N_11639);
nor U12544 (N_12544,N_10335,N_11682);
nand U12545 (N_12545,N_11015,N_10240);
or U12546 (N_12546,N_10563,N_11857);
nor U12547 (N_12547,N_10289,N_10743);
nand U12548 (N_12548,N_10959,N_11905);
nor U12549 (N_12549,N_10546,N_10727);
or U12550 (N_12550,N_11142,N_10187);
or U12551 (N_12551,N_10891,N_10321);
or U12552 (N_12552,N_11665,N_11294);
or U12553 (N_12553,N_11796,N_11260);
nor U12554 (N_12554,N_10548,N_10667);
xor U12555 (N_12555,N_11370,N_10646);
xor U12556 (N_12556,N_10873,N_10269);
or U12557 (N_12557,N_11382,N_10012);
nor U12558 (N_12558,N_11726,N_11960);
nor U12559 (N_12559,N_11998,N_11139);
nand U12560 (N_12560,N_10184,N_10626);
nor U12561 (N_12561,N_11162,N_11730);
nor U12562 (N_12562,N_11144,N_11943);
xor U12563 (N_12563,N_10818,N_11312);
nor U12564 (N_12564,N_10931,N_11264);
nand U12565 (N_12565,N_10590,N_11933);
and U12566 (N_12566,N_11120,N_10759);
nor U12567 (N_12567,N_10420,N_11924);
nor U12568 (N_12568,N_10730,N_11651);
or U12569 (N_12569,N_11012,N_11153);
or U12570 (N_12570,N_11823,N_10631);
or U12571 (N_12571,N_10251,N_11464);
nand U12572 (N_12572,N_11477,N_11043);
xor U12573 (N_12573,N_10391,N_11006);
and U12574 (N_12574,N_10662,N_10811);
or U12575 (N_12575,N_11008,N_10141);
nor U12576 (N_12576,N_11505,N_11420);
nand U12577 (N_12577,N_11066,N_10883);
or U12578 (N_12578,N_11255,N_11918);
nor U12579 (N_12579,N_11829,N_11267);
nor U12580 (N_12580,N_11208,N_11779);
nand U12581 (N_12581,N_10239,N_10689);
nor U12582 (N_12582,N_10513,N_11326);
xor U12583 (N_12583,N_10272,N_10408);
xnor U12584 (N_12584,N_11156,N_11413);
xnor U12585 (N_12585,N_10888,N_11241);
nand U12586 (N_12586,N_11226,N_11818);
or U12587 (N_12587,N_11073,N_11904);
nor U12588 (N_12588,N_11979,N_11345);
nor U12589 (N_12589,N_11469,N_10052);
nand U12590 (N_12590,N_10110,N_11860);
and U12591 (N_12591,N_10186,N_11486);
xor U12592 (N_12592,N_11766,N_11386);
or U12593 (N_12593,N_10620,N_11601);
nor U12594 (N_12594,N_11356,N_11256);
nor U12595 (N_12595,N_10112,N_10615);
nor U12596 (N_12596,N_10131,N_10973);
and U12597 (N_12597,N_11367,N_11104);
or U12598 (N_12598,N_10535,N_11844);
xnor U12599 (N_12599,N_11050,N_11625);
and U12600 (N_12600,N_10904,N_10238);
and U12601 (N_12601,N_10217,N_11641);
nor U12602 (N_12602,N_11741,N_11571);
and U12603 (N_12603,N_11416,N_11068);
and U12604 (N_12604,N_10702,N_11916);
nor U12605 (N_12605,N_11248,N_11698);
xor U12606 (N_12606,N_11426,N_10882);
or U12607 (N_12607,N_10946,N_11864);
or U12608 (N_12608,N_10895,N_10412);
nor U12609 (N_12609,N_10474,N_11828);
or U12610 (N_12610,N_11882,N_10676);
or U12611 (N_12611,N_11562,N_11277);
xor U12612 (N_12612,N_11981,N_10380);
and U12613 (N_12613,N_10834,N_10039);
and U12614 (N_12614,N_10266,N_11339);
nand U12615 (N_12615,N_10303,N_10750);
and U12616 (N_12616,N_11292,N_11568);
xnor U12617 (N_12617,N_10030,N_10538);
nand U12618 (N_12618,N_11915,N_11238);
xnor U12619 (N_12619,N_10786,N_10125);
or U12620 (N_12620,N_11510,N_10653);
or U12621 (N_12621,N_11586,N_11462);
or U12622 (N_12622,N_10932,N_11925);
xnor U12623 (N_12623,N_11480,N_11463);
nand U12624 (N_12624,N_10964,N_10594);
xor U12625 (N_12625,N_10024,N_11825);
xnor U12626 (N_12626,N_11185,N_11705);
or U12627 (N_12627,N_10150,N_11349);
xor U12628 (N_12628,N_10542,N_11773);
or U12629 (N_12629,N_11946,N_10034);
xor U12630 (N_12630,N_11254,N_11653);
xor U12631 (N_12631,N_11446,N_11127);
nand U12632 (N_12632,N_11179,N_10798);
or U12633 (N_12633,N_10902,N_10637);
nand U12634 (N_12634,N_11452,N_11848);
and U12635 (N_12635,N_11138,N_10102);
xor U12636 (N_12636,N_11466,N_11801);
and U12637 (N_12637,N_11201,N_11366);
nand U12638 (N_12638,N_11673,N_11599);
xnor U12639 (N_12639,N_10663,N_10683);
or U12640 (N_12640,N_11881,N_11397);
nor U12641 (N_12641,N_11603,N_11313);
nor U12642 (N_12642,N_10763,N_10995);
and U12643 (N_12643,N_10783,N_10607);
and U12644 (N_12644,N_10320,N_11504);
xor U12645 (N_12645,N_10800,N_10716);
xor U12646 (N_12646,N_11578,N_10492);
and U12647 (N_12647,N_10651,N_10273);
or U12648 (N_12648,N_11999,N_11680);
nand U12649 (N_12649,N_10929,N_11284);
xor U12650 (N_12650,N_10605,N_10208);
nand U12651 (N_12651,N_10180,N_10348);
nand U12652 (N_12652,N_10912,N_10071);
nand U12653 (N_12653,N_10328,N_10591);
nor U12654 (N_12654,N_10404,N_11629);
or U12655 (N_12655,N_10015,N_11202);
nor U12656 (N_12656,N_10698,N_10859);
nand U12657 (N_12657,N_10812,N_11959);
xor U12658 (N_12658,N_11768,N_11027);
xor U12659 (N_12659,N_10174,N_10722);
xor U12660 (N_12660,N_10101,N_10744);
and U12661 (N_12661,N_10318,N_11243);
nor U12662 (N_12662,N_11800,N_10006);
nor U12663 (N_12663,N_10601,N_11394);
nor U12664 (N_12664,N_10041,N_11600);
nand U12665 (N_12665,N_11544,N_11160);
nor U12666 (N_12666,N_10058,N_11941);
and U12667 (N_12667,N_10681,N_11308);
xor U12668 (N_12668,N_11996,N_10369);
xnor U12669 (N_12669,N_11596,N_10619);
and U12670 (N_12670,N_10341,N_10275);
and U12671 (N_12671,N_10301,N_11298);
or U12672 (N_12672,N_10823,N_10934);
nor U12673 (N_12673,N_10643,N_10521);
and U12674 (N_12674,N_10192,N_11046);
and U12675 (N_12675,N_10860,N_10426);
or U12676 (N_12676,N_10809,N_11646);
or U12677 (N_12677,N_11159,N_11467);
or U12678 (N_12678,N_11271,N_10844);
and U12679 (N_12679,N_10491,N_11170);
xor U12680 (N_12680,N_11757,N_10028);
nor U12681 (N_12681,N_11135,N_11739);
and U12682 (N_12682,N_11945,N_11269);
or U12683 (N_12683,N_11176,N_11145);
xnor U12684 (N_12684,N_10640,N_10945);
nand U12685 (N_12685,N_10466,N_10787);
nor U12686 (N_12686,N_10868,N_11387);
and U12687 (N_12687,N_11285,N_10256);
xnor U12688 (N_12688,N_11543,N_11888);
and U12689 (N_12689,N_11515,N_11923);
xor U12690 (N_12690,N_10690,N_10728);
or U12691 (N_12691,N_11940,N_10336);
nor U12692 (N_12692,N_10230,N_11259);
nor U12693 (N_12693,N_11407,N_10990);
xor U12694 (N_12694,N_10042,N_11983);
or U12695 (N_12695,N_11570,N_10863);
xor U12696 (N_12696,N_10571,N_11297);
and U12697 (N_12697,N_10025,N_11791);
nand U12698 (N_12698,N_11161,N_10037);
or U12699 (N_12699,N_10392,N_10327);
or U12700 (N_12700,N_10641,N_11178);
or U12701 (N_12701,N_10232,N_11158);
nand U12702 (N_12702,N_11460,N_10405);
and U12703 (N_12703,N_11684,N_11403);
nor U12704 (N_12704,N_10175,N_10291);
nand U12705 (N_12705,N_11597,N_10917);
and U12706 (N_12706,N_11342,N_11847);
nor U12707 (N_12707,N_11272,N_10137);
nor U12708 (N_12708,N_10452,N_10813);
nor U12709 (N_12709,N_10846,N_10674);
xor U12710 (N_12710,N_11368,N_10987);
or U12711 (N_12711,N_10725,N_10807);
nor U12712 (N_12712,N_11323,N_10196);
nand U12713 (N_12713,N_11122,N_10575);
or U12714 (N_12714,N_10924,N_11405);
nor U12715 (N_12715,N_10203,N_10068);
nor U12716 (N_12716,N_11742,N_10451);
nand U12717 (N_12717,N_10220,N_11845);
and U12718 (N_12718,N_10281,N_11987);
or U12719 (N_12719,N_10936,N_10044);
nand U12720 (N_12720,N_11936,N_10953);
and U12721 (N_12721,N_11237,N_11696);
or U12722 (N_12722,N_11583,N_11743);
nor U12723 (N_12723,N_10719,N_11619);
nand U12724 (N_12724,N_10353,N_10952);
nand U12725 (N_12725,N_11587,N_11813);
nor U12726 (N_12726,N_10284,N_10951);
or U12727 (N_12727,N_10067,N_11874);
or U12728 (N_12728,N_11944,N_10958);
or U12729 (N_12729,N_11130,N_10349);
nand U12730 (N_12730,N_11375,N_11032);
nor U12731 (N_12731,N_11627,N_10695);
nand U12732 (N_12732,N_11950,N_10774);
xor U12733 (N_12733,N_11053,N_10322);
nor U12734 (N_12734,N_10309,N_11522);
xnor U12735 (N_12735,N_10821,N_11865);
and U12736 (N_12736,N_10056,N_10566);
nand U12737 (N_12737,N_11859,N_11751);
nand U12738 (N_12738,N_10630,N_11833);
and U12739 (N_12739,N_10283,N_11383);
and U12740 (N_12740,N_10718,N_11468);
nor U12741 (N_12741,N_10152,N_10996);
nor U12742 (N_12742,N_11671,N_11457);
nor U12743 (N_12743,N_11919,N_10483);
xor U12744 (N_12744,N_11762,N_10432);
or U12745 (N_12745,N_11880,N_11253);
nand U12746 (N_12746,N_10158,N_11501);
nor U12747 (N_12747,N_10634,N_10732);
nand U12748 (N_12748,N_10765,N_10314);
nand U12749 (N_12749,N_11306,N_10430);
and U12750 (N_12750,N_10838,N_10604);
or U12751 (N_12751,N_11459,N_11044);
and U12752 (N_12752,N_11724,N_11103);
nor U12753 (N_12753,N_11472,N_10864);
nor U12754 (N_12754,N_10290,N_11217);
and U12755 (N_12755,N_11063,N_11362);
xnor U12756 (N_12756,N_11361,N_10263);
or U12757 (N_12757,N_11962,N_10564);
or U12758 (N_12758,N_11679,N_10047);
or U12759 (N_12759,N_11458,N_10300);
or U12760 (N_12760,N_10994,N_10167);
nand U12761 (N_12761,N_10423,N_11862);
xnor U12762 (N_12762,N_11378,N_11307);
xnor U12763 (N_12763,N_10627,N_11500);
nand U12764 (N_12764,N_11296,N_11172);
or U12765 (N_12765,N_10287,N_10908);
xnor U12766 (N_12766,N_10831,N_10372);
xor U12767 (N_12767,N_11374,N_10277);
nor U12768 (N_12768,N_11304,N_10697);
or U12769 (N_12769,N_10832,N_10437);
or U12770 (N_12770,N_11545,N_11263);
xor U12771 (N_12771,N_11252,N_10484);
nand U12772 (N_12772,N_11395,N_10780);
nand U12773 (N_12773,N_11167,N_11033);
or U12774 (N_12774,N_10288,N_11455);
nor U12775 (N_12775,N_10721,N_11174);
nand U12776 (N_12776,N_10356,N_11908);
xor U12777 (N_12777,N_11668,N_11036);
and U12778 (N_12778,N_10726,N_10190);
and U12779 (N_12779,N_11971,N_11866);
or U12780 (N_12780,N_11734,N_11585);
xnor U12781 (N_12781,N_11411,N_10447);
or U12782 (N_12782,N_10324,N_11644);
and U12783 (N_12783,N_10038,N_11106);
xnor U12784 (N_12784,N_11806,N_10197);
xor U12785 (N_12785,N_10455,N_11952);
and U12786 (N_12786,N_11970,N_10078);
xor U12787 (N_12787,N_10949,N_11089);
xnor U12788 (N_12788,N_10140,N_10829);
nand U12789 (N_12789,N_11902,N_11001);
nor U12790 (N_12790,N_10222,N_11704);
nand U12791 (N_12791,N_10310,N_11591);
or U12792 (N_12792,N_10785,N_10434);
or U12793 (N_12793,N_10096,N_11128);
xor U12794 (N_12794,N_10224,N_11003);
nand U12795 (N_12795,N_10293,N_10139);
nand U12796 (N_12796,N_10331,N_10708);
nor U12797 (N_12797,N_10935,N_10194);
xor U12798 (N_12798,N_11663,N_11240);
nor U12799 (N_12799,N_11052,N_10387);
and U12800 (N_12800,N_10956,N_10972);
or U12801 (N_12801,N_10573,N_10982);
or U12802 (N_12802,N_10118,N_10363);
nand U12803 (N_12803,N_11956,N_11440);
nand U12804 (N_12804,N_10050,N_11146);
nand U12805 (N_12805,N_10425,N_10985);
and U12806 (N_12806,N_10221,N_11929);
nand U12807 (N_12807,N_11689,N_10248);
nand U12808 (N_12808,N_11113,N_10559);
and U12809 (N_12809,N_10916,N_10606);
and U12810 (N_12810,N_10769,N_10475);
and U12811 (N_12811,N_11192,N_10413);
nor U12812 (N_12812,N_11920,N_11750);
xor U12813 (N_12813,N_10464,N_11214);
and U12814 (N_12814,N_11315,N_11508);
xnor U12815 (N_12815,N_11346,N_10749);
and U12816 (N_12816,N_11344,N_10183);
nor U12817 (N_12817,N_11327,N_11788);
and U12818 (N_12818,N_11453,N_11115);
and U12819 (N_12819,N_11869,N_10649);
xnor U12820 (N_12820,N_11258,N_11667);
xor U12821 (N_12821,N_10085,N_10954);
nor U12822 (N_12822,N_11069,N_11892);
and U12823 (N_12823,N_11227,N_11608);
nand U12824 (N_12824,N_10113,N_10334);
and U12825 (N_12825,N_10654,N_10527);
xor U12826 (N_12826,N_10010,N_10539);
or U12827 (N_12827,N_10142,N_10134);
xor U12828 (N_12828,N_10115,N_10621);
and U12829 (N_12829,N_11727,N_11408);
nor U12830 (N_12830,N_10204,N_11566);
or U12831 (N_12831,N_11551,N_10602);
nor U12832 (N_12832,N_11879,N_10165);
nor U12833 (N_12833,N_10870,N_11078);
or U12834 (N_12834,N_10688,N_11038);
nor U12835 (N_12835,N_10896,N_11422);
nor U12836 (N_12836,N_10628,N_10997);
nor U12837 (N_12837,N_11899,N_11856);
xor U12838 (N_12838,N_10758,N_11280);
nor U12839 (N_12839,N_10132,N_10536);
nor U12840 (N_12840,N_11798,N_10682);
and U12841 (N_12841,N_11579,N_10560);
xor U12842 (N_12842,N_11672,N_11182);
xor U12843 (N_12843,N_10343,N_10503);
nand U12844 (N_12844,N_11487,N_10493);
xnor U12845 (N_12845,N_11783,N_11854);
or U12846 (N_12846,N_11849,N_11080);
nand U12847 (N_12847,N_11767,N_11414);
nand U12848 (N_12848,N_10031,N_10511);
xnor U12849 (N_12849,N_10381,N_10161);
xnor U12850 (N_12850,N_11558,N_11702);
or U12851 (N_12851,N_11795,N_10163);
nand U12852 (N_12852,N_11659,N_10925);
and U12853 (N_12853,N_10124,N_10981);
and U12854 (N_12854,N_10710,N_11991);
nand U12855 (N_12855,N_10497,N_10943);
xnor U12856 (N_12856,N_11678,N_10592);
nor U12857 (N_12857,N_11557,N_10706);
or U12858 (N_12858,N_11947,N_11909);
or U12859 (N_12859,N_11193,N_10394);
xnor U12860 (N_12860,N_11906,N_11670);
nand U12861 (N_12861,N_11251,N_11169);
or U12862 (N_12862,N_10350,N_11511);
nor U12863 (N_12863,N_10918,N_10120);
or U12864 (N_12864,N_11359,N_10268);
nand U12865 (N_12865,N_10254,N_11652);
or U12866 (N_12866,N_11567,N_11354);
nand U12867 (N_12867,N_10588,N_11369);
xor U12868 (N_12868,N_11013,N_10429);
nand U12869 (N_12869,N_11319,N_10658);
nor U12870 (N_12870,N_10974,N_11836);
nor U12871 (N_12871,N_11181,N_11707);
or U12872 (N_12872,N_11807,N_10471);
or U12873 (N_12873,N_10715,N_10781);
and U12874 (N_12874,N_10872,N_10617);
nand U12875 (N_12875,N_10172,N_10329);
or U12876 (N_12876,N_11812,N_11351);
nand U12877 (N_12877,N_11270,N_11121);
and U12878 (N_12878,N_10070,N_10797);
nand U12879 (N_12879,N_10933,N_10311);
xnor U12880 (N_12880,N_11528,N_10017);
or U12881 (N_12881,N_11489,N_11028);
and U12882 (N_12882,N_11937,N_11305);
nor U12883 (N_12883,N_11098,N_11927);
nand U12884 (N_12884,N_11687,N_10084);
xor U12885 (N_12885,N_10195,N_11333);
or U12886 (N_12886,N_10299,N_11445);
xnor U12887 (N_12887,N_10516,N_10529);
and U12888 (N_12888,N_10498,N_10062);
and U12889 (N_12889,N_10618,N_11602);
and U12890 (N_12890,N_11396,N_11301);
and U12891 (N_12891,N_10830,N_10009);
nand U12892 (N_12892,N_10914,N_10061);
nand U12893 (N_12893,N_10179,N_11318);
nor U12894 (N_12894,N_10401,N_11431);
nand U12895 (N_12895,N_10822,N_11565);
and U12896 (N_12896,N_11194,N_10295);
or U12897 (N_12897,N_11582,N_11049);
or U12898 (N_12898,N_10921,N_10843);
xnor U12899 (N_12899,N_10358,N_10043);
or U12900 (N_12900,N_11529,N_11628);
nor U12901 (N_12901,N_11654,N_10593);
and U12902 (N_12902,N_11745,N_10480);
xor U12903 (N_12903,N_10889,N_11527);
nor U12904 (N_12904,N_11980,N_10752);
and U12905 (N_12905,N_11016,N_11116);
nand U12906 (N_12906,N_10396,N_10081);
or U12907 (N_12907,N_10515,N_10207);
or U12908 (N_12908,N_10345,N_11516);
nor U12909 (N_12909,N_10063,N_10088);
nor U12910 (N_12910,N_11265,N_10766);
and U12911 (N_12911,N_11797,N_11441);
and U12912 (N_12912,N_11542,N_11774);
xor U12913 (N_12913,N_10213,N_11119);
xor U12914 (N_12914,N_11409,N_10939);
nand U12915 (N_12915,N_11373,N_10160);
and U12916 (N_12916,N_11645,N_10258);
nand U12917 (N_12917,N_11939,N_11988);
nor U12918 (N_12918,N_11048,N_10312);
xor U12919 (N_12919,N_11997,N_11099);
nor U12920 (N_12920,N_10814,N_10128);
and U12921 (N_12921,N_10215,N_10526);
and U12922 (N_12922,N_10871,N_11700);
nand U12923 (N_12923,N_11377,N_10168);
nor U12924 (N_12924,N_10460,N_11427);
nor U12925 (N_12925,N_11975,N_10212);
and U12926 (N_12926,N_11355,N_10313);
nand U12927 (N_12927,N_10360,N_11633);
and U12928 (N_12928,N_10143,N_10490);
nand U12929 (N_12929,N_10104,N_10236);
and U12930 (N_12930,N_11716,N_11832);
nand U12931 (N_12931,N_10554,N_11688);
nor U12932 (N_12932,N_11430,N_10376);
nor U12933 (N_12933,N_10948,N_11428);
or U12934 (N_12934,N_11731,N_10905);
nor U12935 (N_12935,N_10188,N_11621);
or U12936 (N_12936,N_10502,N_10271);
xor U12937 (N_12937,N_10470,N_10614);
nor U12938 (N_12938,N_11334,N_11781);
nand U12939 (N_12939,N_11736,N_10395);
xnor U12940 (N_12940,N_10410,N_11406);
nor U12941 (N_12941,N_10970,N_11283);
and U12942 (N_12942,N_10066,N_10461);
or U12943 (N_12943,N_11275,N_10915);
or U12944 (N_12944,N_11827,N_10231);
nor U12945 (N_12945,N_11948,N_10048);
nand U12946 (N_12946,N_10127,N_11623);
or U12947 (N_12947,N_10210,N_11681);
and U12948 (N_12948,N_11109,N_11538);
or U12949 (N_12949,N_11650,N_11617);
nor U12950 (N_12950,N_11474,N_11729);
and U12951 (N_12951,N_11479,N_10530);
xnor U12952 (N_12952,N_10738,N_11425);
nand U12953 (N_12953,N_10919,N_10462);
or U12954 (N_12954,N_11481,N_11648);
or U12955 (N_12955,N_10855,N_10191);
xor U12956 (N_12956,N_10245,N_11490);
or U12957 (N_12957,N_10228,N_11311);
and U12958 (N_12958,N_10008,N_10748);
nand U12959 (N_12959,N_11951,N_11358);
nor U12960 (N_12960,N_10675,N_11518);
xor U12961 (N_12961,N_11642,N_10518);
nand U12962 (N_12962,N_10457,N_10317);
xor U12963 (N_12963,N_11011,N_10411);
nand U12964 (N_12964,N_10438,N_11492);
or U12965 (N_12965,N_11834,N_11478);
nand U12966 (N_12966,N_11442,N_10745);
or U12967 (N_12967,N_10106,N_10992);
and U12968 (N_12968,N_10064,N_11990);
and U12969 (N_12969,N_11786,N_11770);
or U12970 (N_12970,N_11079,N_10383);
nor U12971 (N_12971,N_10246,N_10850);
or U12972 (N_12972,N_11572,N_11332);
nor U12973 (N_12973,N_10712,N_11287);
and U12974 (N_12974,N_10292,N_10507);
nor U12975 (N_12975,N_11209,N_11613);
and U12976 (N_12976,N_10577,N_10261);
and U12977 (N_12977,N_11129,N_10584);
nand U12978 (N_12978,N_11953,N_10265);
and U12979 (N_12979,N_11495,N_10944);
or U12980 (N_12980,N_11523,N_10090);
or U12981 (N_12981,N_10926,N_10796);
and U12982 (N_12982,N_11992,N_10512);
or U12983 (N_12983,N_10270,N_11590);
nand U12984 (N_12984,N_11056,N_10055);
nor U12985 (N_12985,N_10357,N_11811);
xnor U12986 (N_12986,N_11677,N_10099);
nor U12987 (N_12987,N_11785,N_11846);
or U12988 (N_12988,N_11622,N_10001);
nor U12989 (N_12989,N_11703,N_10582);
or U12990 (N_12990,N_11149,N_10537);
nand U12991 (N_12991,N_11057,N_11517);
xnor U12992 (N_12992,N_11328,N_11101);
xor U12993 (N_12993,N_11973,N_11438);
or U12994 (N_12994,N_11831,N_10121);
nand U12995 (N_12995,N_11656,N_11876);
or U12996 (N_12996,N_11300,N_11114);
nand U12997 (N_12997,N_11976,N_11815);
nand U12998 (N_12998,N_11299,N_11958);
xor U12999 (N_12999,N_11928,N_10226);
or U13000 (N_13000,N_11219,N_10908);
nor U13001 (N_13001,N_10015,N_10594);
xnor U13002 (N_13002,N_11345,N_11607);
xor U13003 (N_13003,N_11312,N_10938);
nand U13004 (N_13004,N_11139,N_10252);
xnor U13005 (N_13005,N_11522,N_11620);
xnor U13006 (N_13006,N_11915,N_11351);
or U13007 (N_13007,N_10197,N_10868);
and U13008 (N_13008,N_11303,N_10755);
nor U13009 (N_13009,N_10205,N_10788);
and U13010 (N_13010,N_11137,N_11436);
nor U13011 (N_13011,N_11879,N_11183);
and U13012 (N_13012,N_10565,N_10514);
nand U13013 (N_13013,N_10706,N_10777);
nor U13014 (N_13014,N_11425,N_10600);
nor U13015 (N_13015,N_10754,N_11084);
xor U13016 (N_13016,N_10734,N_11629);
or U13017 (N_13017,N_11167,N_10701);
xor U13018 (N_13018,N_10697,N_10204);
nor U13019 (N_13019,N_11039,N_11739);
nand U13020 (N_13020,N_11193,N_10026);
xnor U13021 (N_13021,N_10864,N_11541);
nor U13022 (N_13022,N_10228,N_11843);
xnor U13023 (N_13023,N_11068,N_11692);
nor U13024 (N_13024,N_11984,N_11777);
and U13025 (N_13025,N_10340,N_10554);
and U13026 (N_13026,N_10168,N_11776);
nor U13027 (N_13027,N_11345,N_11620);
nand U13028 (N_13028,N_10185,N_10964);
nand U13029 (N_13029,N_11151,N_11004);
or U13030 (N_13030,N_10981,N_11681);
nand U13031 (N_13031,N_10439,N_10212);
nor U13032 (N_13032,N_11990,N_10606);
and U13033 (N_13033,N_11485,N_10517);
xor U13034 (N_13034,N_10721,N_11840);
nor U13035 (N_13035,N_11883,N_10491);
or U13036 (N_13036,N_10102,N_11561);
or U13037 (N_13037,N_11890,N_10215);
and U13038 (N_13038,N_11900,N_11268);
nand U13039 (N_13039,N_10837,N_10641);
or U13040 (N_13040,N_11362,N_11377);
xor U13041 (N_13041,N_10516,N_10622);
and U13042 (N_13042,N_10953,N_10435);
or U13043 (N_13043,N_10718,N_10405);
nand U13044 (N_13044,N_11725,N_11026);
nor U13045 (N_13045,N_10974,N_11940);
nand U13046 (N_13046,N_10165,N_10388);
nand U13047 (N_13047,N_10775,N_11549);
nand U13048 (N_13048,N_11916,N_11303);
xnor U13049 (N_13049,N_10799,N_11437);
or U13050 (N_13050,N_10999,N_10901);
nand U13051 (N_13051,N_10761,N_11361);
or U13052 (N_13052,N_10951,N_11012);
or U13053 (N_13053,N_11933,N_11401);
or U13054 (N_13054,N_10623,N_10490);
xnor U13055 (N_13055,N_10360,N_11852);
or U13056 (N_13056,N_10316,N_11196);
nor U13057 (N_13057,N_10904,N_10691);
nor U13058 (N_13058,N_11700,N_10512);
and U13059 (N_13059,N_10216,N_10493);
nand U13060 (N_13060,N_10411,N_10513);
nor U13061 (N_13061,N_10198,N_10368);
nor U13062 (N_13062,N_10808,N_11791);
and U13063 (N_13063,N_10692,N_10343);
xor U13064 (N_13064,N_10197,N_10824);
xnor U13065 (N_13065,N_10695,N_10954);
and U13066 (N_13066,N_10169,N_10402);
or U13067 (N_13067,N_11893,N_11531);
or U13068 (N_13068,N_10126,N_11757);
nand U13069 (N_13069,N_11088,N_11533);
nor U13070 (N_13070,N_11100,N_11760);
nand U13071 (N_13071,N_10915,N_10239);
xnor U13072 (N_13072,N_11228,N_10921);
nand U13073 (N_13073,N_10694,N_10373);
xnor U13074 (N_13074,N_10887,N_10914);
nand U13075 (N_13075,N_11120,N_10728);
nand U13076 (N_13076,N_10876,N_11259);
and U13077 (N_13077,N_11396,N_10078);
nand U13078 (N_13078,N_11194,N_11391);
and U13079 (N_13079,N_11101,N_11558);
nor U13080 (N_13080,N_10504,N_10031);
nor U13081 (N_13081,N_11708,N_11356);
and U13082 (N_13082,N_11442,N_10037);
or U13083 (N_13083,N_11862,N_11835);
or U13084 (N_13084,N_10376,N_11405);
or U13085 (N_13085,N_10089,N_11758);
and U13086 (N_13086,N_11839,N_11656);
and U13087 (N_13087,N_10806,N_10415);
or U13088 (N_13088,N_10268,N_11328);
xor U13089 (N_13089,N_10174,N_10882);
xnor U13090 (N_13090,N_10325,N_11436);
xor U13091 (N_13091,N_10892,N_10288);
or U13092 (N_13092,N_10014,N_10201);
nand U13093 (N_13093,N_11214,N_11976);
nand U13094 (N_13094,N_11363,N_11190);
nand U13095 (N_13095,N_10107,N_11011);
xor U13096 (N_13096,N_10147,N_11064);
xnor U13097 (N_13097,N_10429,N_11656);
and U13098 (N_13098,N_11747,N_11312);
nand U13099 (N_13099,N_11216,N_11689);
nand U13100 (N_13100,N_10769,N_10376);
nand U13101 (N_13101,N_10520,N_10921);
nand U13102 (N_13102,N_10200,N_10691);
and U13103 (N_13103,N_11738,N_10142);
nand U13104 (N_13104,N_10215,N_11547);
or U13105 (N_13105,N_11325,N_11084);
or U13106 (N_13106,N_10820,N_10308);
nor U13107 (N_13107,N_10603,N_10546);
and U13108 (N_13108,N_10273,N_10048);
xor U13109 (N_13109,N_10908,N_11415);
xnor U13110 (N_13110,N_10401,N_10324);
xor U13111 (N_13111,N_10064,N_10290);
nand U13112 (N_13112,N_10443,N_11934);
nor U13113 (N_13113,N_11326,N_10391);
nor U13114 (N_13114,N_11904,N_11491);
or U13115 (N_13115,N_11528,N_10545);
nand U13116 (N_13116,N_11984,N_11673);
and U13117 (N_13117,N_10674,N_11533);
or U13118 (N_13118,N_10697,N_11081);
nand U13119 (N_13119,N_11876,N_10649);
xnor U13120 (N_13120,N_10937,N_10313);
or U13121 (N_13121,N_11789,N_10265);
and U13122 (N_13122,N_11921,N_11095);
nand U13123 (N_13123,N_10385,N_10970);
or U13124 (N_13124,N_10429,N_10400);
xor U13125 (N_13125,N_11256,N_10512);
nand U13126 (N_13126,N_10379,N_10133);
or U13127 (N_13127,N_10936,N_10118);
and U13128 (N_13128,N_10311,N_10083);
nand U13129 (N_13129,N_11176,N_10862);
and U13130 (N_13130,N_11526,N_10658);
or U13131 (N_13131,N_11214,N_11938);
nand U13132 (N_13132,N_10724,N_11214);
xnor U13133 (N_13133,N_11508,N_10465);
or U13134 (N_13134,N_10565,N_10041);
nor U13135 (N_13135,N_10831,N_11385);
and U13136 (N_13136,N_10027,N_10198);
xnor U13137 (N_13137,N_10075,N_11137);
or U13138 (N_13138,N_10631,N_10149);
or U13139 (N_13139,N_11704,N_11076);
and U13140 (N_13140,N_10659,N_10108);
or U13141 (N_13141,N_11671,N_11360);
nand U13142 (N_13142,N_10921,N_11549);
or U13143 (N_13143,N_11201,N_11856);
xnor U13144 (N_13144,N_11696,N_10006);
xor U13145 (N_13145,N_11257,N_10556);
nor U13146 (N_13146,N_11605,N_11567);
nand U13147 (N_13147,N_10007,N_11010);
and U13148 (N_13148,N_11016,N_10077);
or U13149 (N_13149,N_10357,N_11073);
or U13150 (N_13150,N_11218,N_11286);
nor U13151 (N_13151,N_11568,N_11736);
nor U13152 (N_13152,N_10635,N_11196);
or U13153 (N_13153,N_11227,N_11776);
nor U13154 (N_13154,N_10486,N_10975);
nand U13155 (N_13155,N_10974,N_11532);
xnor U13156 (N_13156,N_10364,N_10619);
nand U13157 (N_13157,N_10505,N_10542);
nor U13158 (N_13158,N_11962,N_11172);
nor U13159 (N_13159,N_10028,N_10587);
or U13160 (N_13160,N_11854,N_11757);
xnor U13161 (N_13161,N_11531,N_11074);
nor U13162 (N_13162,N_10716,N_11376);
and U13163 (N_13163,N_10607,N_11703);
and U13164 (N_13164,N_10236,N_11930);
nor U13165 (N_13165,N_11772,N_11833);
or U13166 (N_13166,N_10329,N_11013);
nand U13167 (N_13167,N_10996,N_10544);
nand U13168 (N_13168,N_11405,N_11244);
nor U13169 (N_13169,N_10518,N_10235);
or U13170 (N_13170,N_10819,N_11875);
and U13171 (N_13171,N_10001,N_10935);
and U13172 (N_13172,N_10046,N_11258);
nor U13173 (N_13173,N_10408,N_11972);
and U13174 (N_13174,N_10254,N_11009);
xnor U13175 (N_13175,N_11279,N_10135);
and U13176 (N_13176,N_11577,N_11419);
or U13177 (N_13177,N_11002,N_10231);
nor U13178 (N_13178,N_10639,N_11363);
or U13179 (N_13179,N_10063,N_11348);
nor U13180 (N_13180,N_10850,N_11717);
or U13181 (N_13181,N_11651,N_10209);
xor U13182 (N_13182,N_11283,N_11094);
or U13183 (N_13183,N_11251,N_11235);
and U13184 (N_13184,N_10734,N_10727);
nor U13185 (N_13185,N_11304,N_10401);
or U13186 (N_13186,N_11632,N_11286);
or U13187 (N_13187,N_11917,N_11770);
and U13188 (N_13188,N_10478,N_11092);
and U13189 (N_13189,N_10544,N_11631);
xor U13190 (N_13190,N_10910,N_11396);
nand U13191 (N_13191,N_11841,N_10779);
nor U13192 (N_13192,N_10653,N_10831);
nor U13193 (N_13193,N_11336,N_11274);
nor U13194 (N_13194,N_11889,N_11957);
nor U13195 (N_13195,N_10439,N_11912);
nand U13196 (N_13196,N_11533,N_11979);
nor U13197 (N_13197,N_11188,N_10258);
or U13198 (N_13198,N_11673,N_10432);
or U13199 (N_13199,N_11962,N_10201);
xor U13200 (N_13200,N_10099,N_11424);
or U13201 (N_13201,N_11295,N_11427);
or U13202 (N_13202,N_11811,N_10324);
or U13203 (N_13203,N_11234,N_11794);
or U13204 (N_13204,N_11484,N_11990);
and U13205 (N_13205,N_10091,N_10309);
xnor U13206 (N_13206,N_10411,N_11307);
xnor U13207 (N_13207,N_11720,N_11855);
or U13208 (N_13208,N_11475,N_11532);
nor U13209 (N_13209,N_11804,N_10793);
nand U13210 (N_13210,N_11989,N_11825);
nor U13211 (N_13211,N_10776,N_10557);
nor U13212 (N_13212,N_11801,N_10451);
xor U13213 (N_13213,N_10453,N_11562);
xor U13214 (N_13214,N_10648,N_11378);
xor U13215 (N_13215,N_11273,N_11122);
nand U13216 (N_13216,N_10282,N_11186);
nand U13217 (N_13217,N_10483,N_11758);
xor U13218 (N_13218,N_11106,N_11978);
or U13219 (N_13219,N_11970,N_10141);
nand U13220 (N_13220,N_10106,N_11995);
or U13221 (N_13221,N_11681,N_10991);
xnor U13222 (N_13222,N_10512,N_10515);
or U13223 (N_13223,N_11880,N_11689);
xor U13224 (N_13224,N_10674,N_11913);
nor U13225 (N_13225,N_11344,N_11687);
nand U13226 (N_13226,N_10583,N_10422);
and U13227 (N_13227,N_10724,N_11805);
nand U13228 (N_13228,N_10512,N_11793);
or U13229 (N_13229,N_11571,N_11590);
or U13230 (N_13230,N_10851,N_10187);
xor U13231 (N_13231,N_10598,N_10355);
and U13232 (N_13232,N_10740,N_10312);
and U13233 (N_13233,N_11875,N_11270);
nor U13234 (N_13234,N_11130,N_10832);
and U13235 (N_13235,N_10606,N_10351);
nor U13236 (N_13236,N_11252,N_11224);
xnor U13237 (N_13237,N_10103,N_11756);
nand U13238 (N_13238,N_11711,N_11353);
xor U13239 (N_13239,N_10696,N_10695);
or U13240 (N_13240,N_11493,N_11548);
nor U13241 (N_13241,N_11543,N_11024);
or U13242 (N_13242,N_10131,N_11038);
nor U13243 (N_13243,N_10382,N_11772);
nor U13244 (N_13244,N_10139,N_10674);
nand U13245 (N_13245,N_11199,N_10639);
or U13246 (N_13246,N_11026,N_11510);
nand U13247 (N_13247,N_10400,N_11957);
nor U13248 (N_13248,N_10422,N_11853);
or U13249 (N_13249,N_10906,N_11826);
nand U13250 (N_13250,N_10174,N_10117);
xnor U13251 (N_13251,N_11653,N_10859);
nor U13252 (N_13252,N_11348,N_11821);
or U13253 (N_13253,N_10065,N_10016);
nor U13254 (N_13254,N_11999,N_10568);
or U13255 (N_13255,N_10468,N_11872);
nor U13256 (N_13256,N_10033,N_11828);
xnor U13257 (N_13257,N_11834,N_10961);
xor U13258 (N_13258,N_10280,N_11570);
nor U13259 (N_13259,N_10296,N_11485);
or U13260 (N_13260,N_10607,N_11422);
xor U13261 (N_13261,N_10480,N_11261);
and U13262 (N_13262,N_11215,N_10370);
nand U13263 (N_13263,N_11193,N_11112);
nand U13264 (N_13264,N_10190,N_10238);
xor U13265 (N_13265,N_11705,N_10617);
and U13266 (N_13266,N_10533,N_11258);
and U13267 (N_13267,N_11161,N_11873);
and U13268 (N_13268,N_11452,N_10932);
nand U13269 (N_13269,N_11833,N_11659);
xnor U13270 (N_13270,N_11768,N_11921);
and U13271 (N_13271,N_11779,N_11060);
nand U13272 (N_13272,N_11920,N_10026);
nand U13273 (N_13273,N_10125,N_11765);
nand U13274 (N_13274,N_10616,N_11511);
nand U13275 (N_13275,N_11486,N_10665);
xnor U13276 (N_13276,N_10758,N_11821);
nor U13277 (N_13277,N_10247,N_11844);
nand U13278 (N_13278,N_11834,N_11152);
nand U13279 (N_13279,N_11353,N_10378);
and U13280 (N_13280,N_10751,N_10438);
xor U13281 (N_13281,N_11693,N_11427);
nor U13282 (N_13282,N_10583,N_11060);
xor U13283 (N_13283,N_11605,N_10487);
or U13284 (N_13284,N_10188,N_10246);
xor U13285 (N_13285,N_10173,N_10450);
or U13286 (N_13286,N_11715,N_10416);
nor U13287 (N_13287,N_11797,N_11932);
xor U13288 (N_13288,N_11027,N_10128);
nor U13289 (N_13289,N_11303,N_10022);
and U13290 (N_13290,N_10830,N_10741);
nand U13291 (N_13291,N_10404,N_11662);
or U13292 (N_13292,N_11185,N_10224);
nand U13293 (N_13293,N_10511,N_10639);
and U13294 (N_13294,N_10095,N_11991);
and U13295 (N_13295,N_11634,N_10090);
nand U13296 (N_13296,N_10592,N_10904);
xnor U13297 (N_13297,N_10185,N_11017);
nand U13298 (N_13298,N_11472,N_11515);
nand U13299 (N_13299,N_11754,N_10851);
nand U13300 (N_13300,N_11161,N_10706);
or U13301 (N_13301,N_10565,N_10118);
or U13302 (N_13302,N_11019,N_11408);
xnor U13303 (N_13303,N_10711,N_11313);
nand U13304 (N_13304,N_10338,N_11399);
and U13305 (N_13305,N_11278,N_11457);
and U13306 (N_13306,N_11893,N_10304);
nor U13307 (N_13307,N_11738,N_10657);
and U13308 (N_13308,N_10181,N_10283);
nor U13309 (N_13309,N_11194,N_11054);
xor U13310 (N_13310,N_11205,N_10160);
nor U13311 (N_13311,N_11740,N_11278);
or U13312 (N_13312,N_11085,N_11595);
xor U13313 (N_13313,N_10164,N_10337);
nor U13314 (N_13314,N_10468,N_11798);
xor U13315 (N_13315,N_11159,N_11005);
nand U13316 (N_13316,N_10855,N_10890);
nand U13317 (N_13317,N_11755,N_11086);
nand U13318 (N_13318,N_10204,N_10619);
nor U13319 (N_13319,N_11666,N_11249);
and U13320 (N_13320,N_11670,N_11657);
and U13321 (N_13321,N_10619,N_11005);
and U13322 (N_13322,N_10800,N_10372);
or U13323 (N_13323,N_11831,N_10656);
nor U13324 (N_13324,N_11121,N_11418);
nor U13325 (N_13325,N_11729,N_11335);
nand U13326 (N_13326,N_11395,N_11105);
and U13327 (N_13327,N_11788,N_11143);
or U13328 (N_13328,N_11831,N_10008);
xnor U13329 (N_13329,N_10491,N_11570);
or U13330 (N_13330,N_10861,N_11395);
nor U13331 (N_13331,N_10586,N_11448);
nand U13332 (N_13332,N_11728,N_10689);
xnor U13333 (N_13333,N_10456,N_11733);
and U13334 (N_13334,N_10525,N_10716);
nand U13335 (N_13335,N_10433,N_11943);
nor U13336 (N_13336,N_11634,N_10583);
or U13337 (N_13337,N_10694,N_11444);
and U13338 (N_13338,N_10902,N_11624);
and U13339 (N_13339,N_11646,N_11520);
xnor U13340 (N_13340,N_11721,N_11236);
nand U13341 (N_13341,N_10780,N_11346);
nor U13342 (N_13342,N_11324,N_11686);
and U13343 (N_13343,N_10240,N_10624);
xnor U13344 (N_13344,N_10140,N_10944);
xnor U13345 (N_13345,N_11524,N_10977);
and U13346 (N_13346,N_11940,N_11938);
nor U13347 (N_13347,N_10506,N_10931);
nand U13348 (N_13348,N_10254,N_10144);
xor U13349 (N_13349,N_11773,N_10644);
nor U13350 (N_13350,N_11940,N_10383);
xnor U13351 (N_13351,N_10615,N_11629);
xor U13352 (N_13352,N_10278,N_10840);
nor U13353 (N_13353,N_10812,N_11235);
or U13354 (N_13354,N_10175,N_11765);
xor U13355 (N_13355,N_11675,N_11031);
xnor U13356 (N_13356,N_11279,N_11081);
xnor U13357 (N_13357,N_11930,N_11749);
or U13358 (N_13358,N_10195,N_11854);
and U13359 (N_13359,N_11662,N_10867);
and U13360 (N_13360,N_11606,N_10123);
and U13361 (N_13361,N_10513,N_10400);
nor U13362 (N_13362,N_10509,N_10794);
or U13363 (N_13363,N_10216,N_11853);
or U13364 (N_13364,N_11882,N_11469);
xor U13365 (N_13365,N_10544,N_10197);
and U13366 (N_13366,N_11854,N_10161);
nor U13367 (N_13367,N_10039,N_11866);
nand U13368 (N_13368,N_11903,N_10995);
nand U13369 (N_13369,N_11156,N_10095);
or U13370 (N_13370,N_10084,N_11677);
nand U13371 (N_13371,N_11076,N_11885);
nor U13372 (N_13372,N_10492,N_10157);
and U13373 (N_13373,N_11111,N_10111);
and U13374 (N_13374,N_10955,N_11516);
nand U13375 (N_13375,N_11343,N_11277);
and U13376 (N_13376,N_10551,N_11196);
or U13377 (N_13377,N_11122,N_10717);
nor U13378 (N_13378,N_10434,N_10411);
xor U13379 (N_13379,N_10038,N_10052);
nand U13380 (N_13380,N_10009,N_10874);
xnor U13381 (N_13381,N_10669,N_10568);
and U13382 (N_13382,N_11756,N_11469);
nor U13383 (N_13383,N_10660,N_11123);
nor U13384 (N_13384,N_11168,N_11282);
or U13385 (N_13385,N_11247,N_10311);
and U13386 (N_13386,N_11398,N_10565);
and U13387 (N_13387,N_11980,N_11613);
nor U13388 (N_13388,N_10798,N_10261);
and U13389 (N_13389,N_11308,N_10056);
or U13390 (N_13390,N_11600,N_10747);
nand U13391 (N_13391,N_11407,N_10021);
nor U13392 (N_13392,N_10804,N_10458);
xnor U13393 (N_13393,N_11802,N_11657);
xnor U13394 (N_13394,N_10213,N_11939);
nand U13395 (N_13395,N_10343,N_11830);
or U13396 (N_13396,N_10674,N_10283);
and U13397 (N_13397,N_10745,N_10332);
or U13398 (N_13398,N_11160,N_10236);
or U13399 (N_13399,N_10020,N_11041);
xor U13400 (N_13400,N_11942,N_10592);
xnor U13401 (N_13401,N_11598,N_10265);
and U13402 (N_13402,N_11202,N_11866);
or U13403 (N_13403,N_10582,N_10021);
and U13404 (N_13404,N_11831,N_11687);
and U13405 (N_13405,N_10397,N_11062);
nand U13406 (N_13406,N_10355,N_11917);
xnor U13407 (N_13407,N_10458,N_11742);
xor U13408 (N_13408,N_11645,N_11680);
xnor U13409 (N_13409,N_10285,N_11002);
or U13410 (N_13410,N_11906,N_10831);
nor U13411 (N_13411,N_11683,N_11062);
xnor U13412 (N_13412,N_10674,N_10932);
nand U13413 (N_13413,N_11070,N_10537);
nor U13414 (N_13414,N_10032,N_11146);
xor U13415 (N_13415,N_10551,N_10472);
and U13416 (N_13416,N_11681,N_11309);
nand U13417 (N_13417,N_10277,N_10998);
nor U13418 (N_13418,N_10551,N_10047);
nor U13419 (N_13419,N_10360,N_10693);
nor U13420 (N_13420,N_11960,N_11731);
xnor U13421 (N_13421,N_11895,N_11180);
nor U13422 (N_13422,N_10363,N_11090);
nand U13423 (N_13423,N_10016,N_11926);
or U13424 (N_13424,N_10595,N_11607);
nand U13425 (N_13425,N_11976,N_11649);
xnor U13426 (N_13426,N_11067,N_11365);
nand U13427 (N_13427,N_11133,N_10426);
nor U13428 (N_13428,N_11820,N_11209);
nor U13429 (N_13429,N_11996,N_10523);
and U13430 (N_13430,N_10219,N_10929);
xor U13431 (N_13431,N_11982,N_11474);
nor U13432 (N_13432,N_11727,N_10042);
nor U13433 (N_13433,N_11325,N_11760);
or U13434 (N_13434,N_11360,N_10624);
or U13435 (N_13435,N_11826,N_10160);
nand U13436 (N_13436,N_10968,N_10672);
and U13437 (N_13437,N_10420,N_10484);
nor U13438 (N_13438,N_10877,N_11568);
and U13439 (N_13439,N_10141,N_10025);
or U13440 (N_13440,N_10386,N_10166);
or U13441 (N_13441,N_10105,N_11801);
or U13442 (N_13442,N_11348,N_10257);
xor U13443 (N_13443,N_11226,N_11822);
nor U13444 (N_13444,N_11209,N_11383);
nand U13445 (N_13445,N_11880,N_10420);
nand U13446 (N_13446,N_11591,N_10294);
and U13447 (N_13447,N_10898,N_11286);
nor U13448 (N_13448,N_11349,N_10370);
or U13449 (N_13449,N_11382,N_10623);
nor U13450 (N_13450,N_11670,N_11593);
and U13451 (N_13451,N_10522,N_10483);
xor U13452 (N_13452,N_10668,N_10879);
or U13453 (N_13453,N_10099,N_10492);
and U13454 (N_13454,N_10136,N_11348);
and U13455 (N_13455,N_10745,N_11680);
nor U13456 (N_13456,N_10663,N_11671);
and U13457 (N_13457,N_11266,N_11923);
xnor U13458 (N_13458,N_10553,N_10335);
nand U13459 (N_13459,N_11057,N_10740);
and U13460 (N_13460,N_10253,N_10560);
xor U13461 (N_13461,N_11972,N_10586);
and U13462 (N_13462,N_10085,N_11759);
xnor U13463 (N_13463,N_11514,N_10252);
xnor U13464 (N_13464,N_10664,N_11455);
nor U13465 (N_13465,N_10543,N_11300);
or U13466 (N_13466,N_10785,N_11334);
or U13467 (N_13467,N_10049,N_11203);
xnor U13468 (N_13468,N_11732,N_10571);
nand U13469 (N_13469,N_10885,N_11586);
and U13470 (N_13470,N_11741,N_10367);
nand U13471 (N_13471,N_11439,N_11487);
xnor U13472 (N_13472,N_11301,N_11489);
nor U13473 (N_13473,N_10067,N_10582);
nand U13474 (N_13474,N_10012,N_11620);
nand U13475 (N_13475,N_10225,N_11783);
xnor U13476 (N_13476,N_11255,N_10592);
or U13477 (N_13477,N_10213,N_10136);
nand U13478 (N_13478,N_11332,N_11877);
and U13479 (N_13479,N_11527,N_11772);
nor U13480 (N_13480,N_10969,N_11942);
and U13481 (N_13481,N_11554,N_10348);
xnor U13482 (N_13482,N_11479,N_11833);
nor U13483 (N_13483,N_11049,N_10098);
and U13484 (N_13484,N_10004,N_10204);
and U13485 (N_13485,N_11181,N_10437);
nand U13486 (N_13486,N_11095,N_11615);
or U13487 (N_13487,N_10231,N_11005);
or U13488 (N_13488,N_11174,N_11826);
xor U13489 (N_13489,N_11566,N_11882);
nor U13490 (N_13490,N_11981,N_10536);
xor U13491 (N_13491,N_11448,N_10350);
nor U13492 (N_13492,N_10187,N_10285);
and U13493 (N_13493,N_11407,N_11637);
nor U13494 (N_13494,N_10087,N_10373);
xor U13495 (N_13495,N_11319,N_10458);
nand U13496 (N_13496,N_11214,N_10810);
nand U13497 (N_13497,N_11581,N_10200);
xnor U13498 (N_13498,N_10365,N_11453);
nor U13499 (N_13499,N_11895,N_11381);
nor U13500 (N_13500,N_10099,N_11834);
nor U13501 (N_13501,N_11615,N_10361);
and U13502 (N_13502,N_10689,N_10609);
nand U13503 (N_13503,N_11272,N_11801);
and U13504 (N_13504,N_11091,N_11916);
nand U13505 (N_13505,N_10118,N_10492);
or U13506 (N_13506,N_10397,N_10842);
nor U13507 (N_13507,N_11708,N_10077);
xnor U13508 (N_13508,N_11799,N_11011);
nand U13509 (N_13509,N_11120,N_10139);
and U13510 (N_13510,N_11168,N_11510);
nor U13511 (N_13511,N_10599,N_10822);
nor U13512 (N_13512,N_11907,N_11258);
and U13513 (N_13513,N_11269,N_10769);
nor U13514 (N_13514,N_11089,N_10190);
nor U13515 (N_13515,N_10826,N_10051);
or U13516 (N_13516,N_11273,N_10299);
and U13517 (N_13517,N_10383,N_11398);
nor U13518 (N_13518,N_10217,N_10145);
xnor U13519 (N_13519,N_11428,N_11013);
xnor U13520 (N_13520,N_11083,N_10977);
nand U13521 (N_13521,N_11395,N_10911);
or U13522 (N_13522,N_10297,N_11114);
xor U13523 (N_13523,N_10571,N_10259);
xor U13524 (N_13524,N_11580,N_10250);
nand U13525 (N_13525,N_10101,N_11085);
and U13526 (N_13526,N_11912,N_10110);
nor U13527 (N_13527,N_11230,N_11246);
or U13528 (N_13528,N_11240,N_10269);
or U13529 (N_13529,N_11378,N_10148);
and U13530 (N_13530,N_11088,N_11616);
xnor U13531 (N_13531,N_11745,N_11954);
and U13532 (N_13532,N_10659,N_10956);
nor U13533 (N_13533,N_11266,N_11133);
nand U13534 (N_13534,N_11340,N_11704);
nor U13535 (N_13535,N_10972,N_10754);
nor U13536 (N_13536,N_11562,N_10629);
nor U13537 (N_13537,N_11974,N_10691);
nor U13538 (N_13538,N_10009,N_10496);
xor U13539 (N_13539,N_11053,N_10796);
nor U13540 (N_13540,N_11618,N_10530);
and U13541 (N_13541,N_11424,N_11582);
nor U13542 (N_13542,N_10484,N_11114);
nand U13543 (N_13543,N_11215,N_10840);
and U13544 (N_13544,N_10530,N_10603);
or U13545 (N_13545,N_11670,N_10548);
xnor U13546 (N_13546,N_10326,N_11728);
or U13547 (N_13547,N_11593,N_10475);
nor U13548 (N_13548,N_10872,N_11857);
and U13549 (N_13549,N_11560,N_11155);
or U13550 (N_13550,N_10566,N_10473);
and U13551 (N_13551,N_11956,N_11044);
or U13552 (N_13552,N_10909,N_11742);
nor U13553 (N_13553,N_11957,N_11477);
nand U13554 (N_13554,N_11086,N_10260);
nor U13555 (N_13555,N_11776,N_11319);
nand U13556 (N_13556,N_10750,N_10716);
nor U13557 (N_13557,N_10782,N_11543);
or U13558 (N_13558,N_11258,N_11597);
nor U13559 (N_13559,N_11936,N_10162);
nor U13560 (N_13560,N_11524,N_11377);
or U13561 (N_13561,N_11889,N_11087);
or U13562 (N_13562,N_10780,N_10243);
nor U13563 (N_13563,N_10291,N_11616);
nor U13564 (N_13564,N_11345,N_10374);
and U13565 (N_13565,N_10647,N_10748);
xnor U13566 (N_13566,N_10526,N_11690);
nor U13567 (N_13567,N_10146,N_11722);
and U13568 (N_13568,N_11492,N_10937);
and U13569 (N_13569,N_10115,N_10834);
xnor U13570 (N_13570,N_11104,N_11574);
xor U13571 (N_13571,N_11090,N_10938);
nand U13572 (N_13572,N_10167,N_11044);
nor U13573 (N_13573,N_11981,N_11169);
xor U13574 (N_13574,N_10096,N_10459);
nor U13575 (N_13575,N_11609,N_11797);
and U13576 (N_13576,N_11490,N_11771);
nor U13577 (N_13577,N_11625,N_10266);
nand U13578 (N_13578,N_10649,N_10719);
nor U13579 (N_13579,N_11410,N_10780);
xor U13580 (N_13580,N_10960,N_10827);
or U13581 (N_13581,N_11886,N_11019);
and U13582 (N_13582,N_10606,N_11760);
xnor U13583 (N_13583,N_10635,N_10955);
xnor U13584 (N_13584,N_10652,N_11213);
and U13585 (N_13585,N_10145,N_11326);
and U13586 (N_13586,N_10562,N_10777);
xor U13587 (N_13587,N_11551,N_10050);
and U13588 (N_13588,N_11654,N_11962);
nor U13589 (N_13589,N_11744,N_11475);
or U13590 (N_13590,N_10793,N_10158);
or U13591 (N_13591,N_10221,N_10889);
nand U13592 (N_13592,N_10605,N_11056);
or U13593 (N_13593,N_11720,N_10016);
nand U13594 (N_13594,N_10805,N_11928);
or U13595 (N_13595,N_11211,N_10220);
xor U13596 (N_13596,N_10657,N_10530);
and U13597 (N_13597,N_11938,N_11772);
and U13598 (N_13598,N_10270,N_10355);
xor U13599 (N_13599,N_10682,N_11395);
xnor U13600 (N_13600,N_10517,N_11146);
and U13601 (N_13601,N_10269,N_10835);
nand U13602 (N_13602,N_10673,N_10913);
nand U13603 (N_13603,N_11709,N_11542);
and U13604 (N_13604,N_10816,N_10982);
and U13605 (N_13605,N_11663,N_11401);
and U13606 (N_13606,N_10303,N_10777);
xnor U13607 (N_13607,N_10966,N_10998);
and U13608 (N_13608,N_10496,N_10044);
xnor U13609 (N_13609,N_10212,N_10732);
or U13610 (N_13610,N_11869,N_10237);
xor U13611 (N_13611,N_10713,N_10346);
or U13612 (N_13612,N_10815,N_11077);
or U13613 (N_13613,N_10867,N_10055);
nand U13614 (N_13614,N_10268,N_11988);
and U13615 (N_13615,N_11843,N_10494);
or U13616 (N_13616,N_11567,N_11579);
or U13617 (N_13617,N_10292,N_10517);
xnor U13618 (N_13618,N_10361,N_10106);
nor U13619 (N_13619,N_11275,N_11315);
xnor U13620 (N_13620,N_11942,N_11804);
xnor U13621 (N_13621,N_10890,N_10720);
and U13622 (N_13622,N_11302,N_11060);
and U13623 (N_13623,N_10758,N_10875);
and U13624 (N_13624,N_11489,N_10883);
xnor U13625 (N_13625,N_10376,N_10123);
and U13626 (N_13626,N_11233,N_11692);
or U13627 (N_13627,N_10328,N_11384);
or U13628 (N_13628,N_10478,N_11001);
nand U13629 (N_13629,N_11519,N_11341);
nor U13630 (N_13630,N_10638,N_11652);
and U13631 (N_13631,N_10249,N_11426);
nand U13632 (N_13632,N_10337,N_11110);
nor U13633 (N_13633,N_11013,N_10822);
or U13634 (N_13634,N_10628,N_10360);
nand U13635 (N_13635,N_11246,N_11981);
xnor U13636 (N_13636,N_11466,N_11514);
and U13637 (N_13637,N_10505,N_10053);
or U13638 (N_13638,N_11731,N_10020);
and U13639 (N_13639,N_10438,N_11613);
xnor U13640 (N_13640,N_11579,N_11481);
or U13641 (N_13641,N_10523,N_10148);
nor U13642 (N_13642,N_11170,N_10052);
xor U13643 (N_13643,N_10951,N_11752);
and U13644 (N_13644,N_11401,N_11633);
and U13645 (N_13645,N_10629,N_11699);
nor U13646 (N_13646,N_10342,N_11269);
and U13647 (N_13647,N_10316,N_10226);
nand U13648 (N_13648,N_11779,N_10833);
nand U13649 (N_13649,N_10022,N_10913);
and U13650 (N_13650,N_10202,N_11925);
nor U13651 (N_13651,N_10529,N_10777);
nor U13652 (N_13652,N_10615,N_11345);
nor U13653 (N_13653,N_11933,N_11177);
or U13654 (N_13654,N_11396,N_11631);
nor U13655 (N_13655,N_10563,N_10690);
or U13656 (N_13656,N_11614,N_11094);
and U13657 (N_13657,N_11727,N_11633);
xor U13658 (N_13658,N_10957,N_11260);
and U13659 (N_13659,N_11259,N_11498);
nor U13660 (N_13660,N_10843,N_10078);
or U13661 (N_13661,N_11696,N_11646);
and U13662 (N_13662,N_10809,N_10444);
and U13663 (N_13663,N_11226,N_11422);
and U13664 (N_13664,N_11695,N_11671);
and U13665 (N_13665,N_10144,N_11801);
xor U13666 (N_13666,N_10789,N_11160);
xor U13667 (N_13667,N_10220,N_10157);
nor U13668 (N_13668,N_11835,N_11782);
nor U13669 (N_13669,N_11690,N_10019);
xnor U13670 (N_13670,N_11431,N_11238);
xor U13671 (N_13671,N_10318,N_11198);
xnor U13672 (N_13672,N_10415,N_10620);
nor U13673 (N_13673,N_11207,N_10556);
nand U13674 (N_13674,N_11348,N_10199);
and U13675 (N_13675,N_10431,N_10469);
nand U13676 (N_13676,N_10445,N_10134);
xor U13677 (N_13677,N_10158,N_11542);
or U13678 (N_13678,N_10787,N_11156);
xnor U13679 (N_13679,N_11484,N_10714);
or U13680 (N_13680,N_10855,N_10087);
nor U13681 (N_13681,N_11933,N_10209);
nor U13682 (N_13682,N_11062,N_10205);
and U13683 (N_13683,N_11349,N_11843);
nand U13684 (N_13684,N_10596,N_11542);
nor U13685 (N_13685,N_10186,N_11527);
xnor U13686 (N_13686,N_11353,N_10237);
and U13687 (N_13687,N_10767,N_11454);
or U13688 (N_13688,N_10449,N_11761);
nor U13689 (N_13689,N_11455,N_11089);
and U13690 (N_13690,N_10203,N_10766);
xnor U13691 (N_13691,N_10526,N_11829);
or U13692 (N_13692,N_10319,N_10327);
or U13693 (N_13693,N_11732,N_11998);
or U13694 (N_13694,N_10231,N_11480);
or U13695 (N_13695,N_11424,N_11880);
nor U13696 (N_13696,N_11706,N_10319);
nor U13697 (N_13697,N_11315,N_10212);
nand U13698 (N_13698,N_11691,N_10290);
or U13699 (N_13699,N_10297,N_10270);
nor U13700 (N_13700,N_11824,N_10096);
xor U13701 (N_13701,N_10172,N_11528);
nor U13702 (N_13702,N_11968,N_11181);
nand U13703 (N_13703,N_11084,N_11562);
or U13704 (N_13704,N_11285,N_10951);
or U13705 (N_13705,N_10708,N_11410);
or U13706 (N_13706,N_10620,N_11292);
and U13707 (N_13707,N_11897,N_10058);
nand U13708 (N_13708,N_11463,N_10690);
and U13709 (N_13709,N_11643,N_11711);
nor U13710 (N_13710,N_11818,N_11098);
or U13711 (N_13711,N_10225,N_10992);
nand U13712 (N_13712,N_10466,N_11268);
or U13713 (N_13713,N_10182,N_10715);
nor U13714 (N_13714,N_11327,N_11892);
nor U13715 (N_13715,N_10622,N_10278);
or U13716 (N_13716,N_11458,N_11751);
nor U13717 (N_13717,N_10389,N_10114);
nor U13718 (N_13718,N_11595,N_10567);
xnor U13719 (N_13719,N_11665,N_11838);
or U13720 (N_13720,N_10460,N_10243);
or U13721 (N_13721,N_11594,N_10565);
and U13722 (N_13722,N_10185,N_10541);
xnor U13723 (N_13723,N_10416,N_11172);
xor U13724 (N_13724,N_10159,N_11205);
or U13725 (N_13725,N_10733,N_10472);
nor U13726 (N_13726,N_11993,N_10310);
nand U13727 (N_13727,N_10853,N_11757);
and U13728 (N_13728,N_11605,N_10815);
nor U13729 (N_13729,N_10822,N_11245);
nand U13730 (N_13730,N_10130,N_11044);
nand U13731 (N_13731,N_10597,N_10342);
and U13732 (N_13732,N_10265,N_11716);
nor U13733 (N_13733,N_11599,N_11873);
nand U13734 (N_13734,N_10847,N_11427);
nor U13735 (N_13735,N_10270,N_11691);
and U13736 (N_13736,N_11549,N_10938);
nor U13737 (N_13737,N_11871,N_10060);
nand U13738 (N_13738,N_11433,N_11925);
or U13739 (N_13739,N_10188,N_11613);
nand U13740 (N_13740,N_11742,N_10331);
xor U13741 (N_13741,N_11218,N_10145);
nand U13742 (N_13742,N_11744,N_10326);
or U13743 (N_13743,N_10515,N_11152);
or U13744 (N_13744,N_11661,N_11654);
xor U13745 (N_13745,N_10373,N_10003);
nand U13746 (N_13746,N_10541,N_10109);
or U13747 (N_13747,N_11733,N_10626);
xnor U13748 (N_13748,N_10901,N_10433);
nand U13749 (N_13749,N_11063,N_10612);
and U13750 (N_13750,N_11730,N_10774);
nor U13751 (N_13751,N_11140,N_11201);
xnor U13752 (N_13752,N_11712,N_10544);
and U13753 (N_13753,N_11650,N_11806);
nor U13754 (N_13754,N_11214,N_11336);
nand U13755 (N_13755,N_10319,N_11055);
xnor U13756 (N_13756,N_10718,N_10750);
xor U13757 (N_13757,N_11129,N_10174);
and U13758 (N_13758,N_10720,N_11010);
or U13759 (N_13759,N_11301,N_10401);
or U13760 (N_13760,N_10748,N_10762);
xnor U13761 (N_13761,N_11262,N_11635);
and U13762 (N_13762,N_11274,N_11382);
xnor U13763 (N_13763,N_10136,N_10338);
nor U13764 (N_13764,N_11333,N_10154);
or U13765 (N_13765,N_11964,N_10363);
nand U13766 (N_13766,N_11696,N_10594);
and U13767 (N_13767,N_11702,N_11637);
xor U13768 (N_13768,N_11484,N_10716);
or U13769 (N_13769,N_10498,N_10662);
nand U13770 (N_13770,N_10865,N_11194);
nor U13771 (N_13771,N_10289,N_11800);
nor U13772 (N_13772,N_10431,N_10917);
and U13773 (N_13773,N_11093,N_11630);
and U13774 (N_13774,N_10974,N_10762);
and U13775 (N_13775,N_11930,N_11431);
and U13776 (N_13776,N_11000,N_11996);
xnor U13777 (N_13777,N_10984,N_11157);
nand U13778 (N_13778,N_11765,N_10340);
xnor U13779 (N_13779,N_10127,N_11052);
and U13780 (N_13780,N_10207,N_10066);
xor U13781 (N_13781,N_11598,N_11721);
nand U13782 (N_13782,N_10023,N_10858);
nand U13783 (N_13783,N_10573,N_11497);
nor U13784 (N_13784,N_10276,N_10581);
nor U13785 (N_13785,N_11106,N_11906);
xnor U13786 (N_13786,N_10761,N_10239);
nor U13787 (N_13787,N_10230,N_11525);
or U13788 (N_13788,N_11174,N_11238);
xor U13789 (N_13789,N_10293,N_11306);
xor U13790 (N_13790,N_10083,N_11389);
and U13791 (N_13791,N_10324,N_11847);
xor U13792 (N_13792,N_11774,N_10204);
nor U13793 (N_13793,N_10444,N_10794);
nor U13794 (N_13794,N_10014,N_11595);
xor U13795 (N_13795,N_11443,N_11869);
or U13796 (N_13796,N_11475,N_11850);
xor U13797 (N_13797,N_11290,N_10478);
xor U13798 (N_13798,N_10802,N_10241);
and U13799 (N_13799,N_10514,N_11556);
xnor U13800 (N_13800,N_10548,N_10212);
and U13801 (N_13801,N_11816,N_10888);
and U13802 (N_13802,N_11586,N_11811);
or U13803 (N_13803,N_10760,N_11362);
and U13804 (N_13804,N_11269,N_10283);
and U13805 (N_13805,N_11693,N_11636);
nand U13806 (N_13806,N_10105,N_10360);
and U13807 (N_13807,N_10018,N_11077);
or U13808 (N_13808,N_10536,N_10632);
or U13809 (N_13809,N_11086,N_11798);
nand U13810 (N_13810,N_11995,N_10501);
and U13811 (N_13811,N_10759,N_10247);
and U13812 (N_13812,N_11816,N_10547);
and U13813 (N_13813,N_10437,N_11449);
nor U13814 (N_13814,N_10090,N_10238);
nor U13815 (N_13815,N_11785,N_11361);
and U13816 (N_13816,N_10215,N_11772);
nor U13817 (N_13817,N_10949,N_10376);
xnor U13818 (N_13818,N_11133,N_10791);
and U13819 (N_13819,N_10436,N_11170);
and U13820 (N_13820,N_10124,N_11514);
nand U13821 (N_13821,N_10578,N_10240);
or U13822 (N_13822,N_10275,N_11445);
or U13823 (N_13823,N_11354,N_11986);
and U13824 (N_13824,N_10632,N_10297);
and U13825 (N_13825,N_11812,N_11517);
nor U13826 (N_13826,N_10565,N_10716);
nor U13827 (N_13827,N_10969,N_11117);
and U13828 (N_13828,N_11026,N_10124);
and U13829 (N_13829,N_10459,N_10195);
xor U13830 (N_13830,N_10594,N_10096);
xnor U13831 (N_13831,N_11455,N_10931);
nand U13832 (N_13832,N_10570,N_10447);
and U13833 (N_13833,N_10573,N_11435);
or U13834 (N_13834,N_11562,N_10835);
and U13835 (N_13835,N_11994,N_11368);
or U13836 (N_13836,N_11658,N_11036);
nor U13837 (N_13837,N_11130,N_10742);
nand U13838 (N_13838,N_10422,N_11141);
xor U13839 (N_13839,N_10903,N_11069);
xnor U13840 (N_13840,N_10564,N_11142);
and U13841 (N_13841,N_11274,N_10137);
and U13842 (N_13842,N_10340,N_11822);
xor U13843 (N_13843,N_10708,N_10055);
xnor U13844 (N_13844,N_11821,N_10406);
xor U13845 (N_13845,N_11847,N_11858);
or U13846 (N_13846,N_10583,N_10667);
or U13847 (N_13847,N_11410,N_11412);
nand U13848 (N_13848,N_11744,N_10583);
nor U13849 (N_13849,N_11952,N_11433);
nand U13850 (N_13850,N_10958,N_11808);
nand U13851 (N_13851,N_11387,N_11381);
nor U13852 (N_13852,N_10228,N_10541);
nor U13853 (N_13853,N_11028,N_10929);
xnor U13854 (N_13854,N_11520,N_11966);
and U13855 (N_13855,N_10781,N_10818);
xnor U13856 (N_13856,N_10765,N_10099);
nor U13857 (N_13857,N_10772,N_10814);
and U13858 (N_13858,N_10542,N_11231);
nor U13859 (N_13859,N_11617,N_10825);
and U13860 (N_13860,N_11777,N_11909);
xnor U13861 (N_13861,N_10698,N_11484);
xnor U13862 (N_13862,N_11618,N_10282);
and U13863 (N_13863,N_11929,N_11827);
or U13864 (N_13864,N_10820,N_11287);
or U13865 (N_13865,N_10000,N_11593);
xnor U13866 (N_13866,N_11680,N_10535);
and U13867 (N_13867,N_10450,N_10719);
xor U13868 (N_13868,N_10206,N_11605);
or U13869 (N_13869,N_10306,N_11231);
nor U13870 (N_13870,N_10181,N_11962);
and U13871 (N_13871,N_10054,N_10700);
xnor U13872 (N_13872,N_11443,N_11597);
or U13873 (N_13873,N_10960,N_11206);
or U13874 (N_13874,N_11807,N_11557);
xor U13875 (N_13875,N_11664,N_10750);
nor U13876 (N_13876,N_11135,N_10122);
nor U13877 (N_13877,N_11679,N_10765);
nand U13878 (N_13878,N_11300,N_10681);
nand U13879 (N_13879,N_10956,N_11285);
or U13880 (N_13880,N_11521,N_10581);
nand U13881 (N_13881,N_11152,N_11581);
nor U13882 (N_13882,N_11632,N_10932);
or U13883 (N_13883,N_11149,N_11481);
xnor U13884 (N_13884,N_10348,N_11393);
nor U13885 (N_13885,N_10242,N_10470);
and U13886 (N_13886,N_10789,N_11902);
or U13887 (N_13887,N_11179,N_11004);
nand U13888 (N_13888,N_10231,N_11620);
xnor U13889 (N_13889,N_11858,N_11443);
nor U13890 (N_13890,N_11580,N_11631);
nor U13891 (N_13891,N_10752,N_10230);
nand U13892 (N_13892,N_10716,N_11868);
xnor U13893 (N_13893,N_10295,N_10063);
nand U13894 (N_13894,N_10742,N_10735);
or U13895 (N_13895,N_11373,N_10126);
xor U13896 (N_13896,N_10131,N_11245);
or U13897 (N_13897,N_11634,N_10341);
or U13898 (N_13898,N_10060,N_11151);
nor U13899 (N_13899,N_11368,N_10508);
nand U13900 (N_13900,N_10024,N_11722);
nand U13901 (N_13901,N_10727,N_10696);
or U13902 (N_13902,N_10565,N_11156);
or U13903 (N_13903,N_10082,N_11133);
nand U13904 (N_13904,N_11369,N_11262);
and U13905 (N_13905,N_10143,N_10589);
xor U13906 (N_13906,N_10806,N_10704);
and U13907 (N_13907,N_11726,N_10596);
or U13908 (N_13908,N_11360,N_11930);
nor U13909 (N_13909,N_10860,N_11616);
nor U13910 (N_13910,N_10357,N_10259);
nor U13911 (N_13911,N_10996,N_10458);
nor U13912 (N_13912,N_10352,N_10584);
or U13913 (N_13913,N_11639,N_11950);
nor U13914 (N_13914,N_10431,N_10730);
or U13915 (N_13915,N_10523,N_11754);
or U13916 (N_13916,N_10321,N_11930);
nor U13917 (N_13917,N_11773,N_10831);
xnor U13918 (N_13918,N_10038,N_11381);
or U13919 (N_13919,N_10836,N_11334);
nor U13920 (N_13920,N_11531,N_10809);
nor U13921 (N_13921,N_11558,N_10295);
or U13922 (N_13922,N_10379,N_10288);
xor U13923 (N_13923,N_11267,N_10131);
nor U13924 (N_13924,N_10062,N_11568);
xor U13925 (N_13925,N_11250,N_11279);
or U13926 (N_13926,N_10245,N_10065);
xor U13927 (N_13927,N_10520,N_10076);
or U13928 (N_13928,N_10720,N_10016);
nor U13929 (N_13929,N_10238,N_11247);
and U13930 (N_13930,N_11991,N_10219);
nor U13931 (N_13931,N_10129,N_10475);
nand U13932 (N_13932,N_11280,N_11895);
xnor U13933 (N_13933,N_11239,N_10058);
nand U13934 (N_13934,N_11884,N_10039);
and U13935 (N_13935,N_10006,N_10593);
xnor U13936 (N_13936,N_10601,N_10565);
or U13937 (N_13937,N_11427,N_10994);
xor U13938 (N_13938,N_11411,N_11061);
or U13939 (N_13939,N_10674,N_11833);
and U13940 (N_13940,N_11547,N_10192);
nand U13941 (N_13941,N_10512,N_11636);
xor U13942 (N_13942,N_11257,N_11873);
and U13943 (N_13943,N_11460,N_10100);
nor U13944 (N_13944,N_11033,N_11487);
nand U13945 (N_13945,N_10511,N_11089);
or U13946 (N_13946,N_11026,N_11012);
and U13947 (N_13947,N_11360,N_11696);
nor U13948 (N_13948,N_10176,N_11590);
xor U13949 (N_13949,N_11612,N_10285);
and U13950 (N_13950,N_10274,N_11874);
or U13951 (N_13951,N_11468,N_11358);
xor U13952 (N_13952,N_10123,N_10418);
nor U13953 (N_13953,N_11400,N_10273);
or U13954 (N_13954,N_11600,N_11690);
nor U13955 (N_13955,N_11502,N_11539);
and U13956 (N_13956,N_10863,N_11925);
and U13957 (N_13957,N_11703,N_10898);
or U13958 (N_13958,N_11899,N_10824);
nor U13959 (N_13959,N_11640,N_10111);
nand U13960 (N_13960,N_11842,N_11899);
or U13961 (N_13961,N_10489,N_10696);
or U13962 (N_13962,N_11666,N_10061);
xnor U13963 (N_13963,N_10986,N_11114);
nand U13964 (N_13964,N_11811,N_10151);
and U13965 (N_13965,N_11896,N_10453);
nand U13966 (N_13966,N_10058,N_11913);
nor U13967 (N_13967,N_11301,N_11537);
nor U13968 (N_13968,N_10611,N_10503);
or U13969 (N_13969,N_10514,N_11640);
xnor U13970 (N_13970,N_10922,N_11163);
or U13971 (N_13971,N_10513,N_11881);
nand U13972 (N_13972,N_11219,N_11589);
nor U13973 (N_13973,N_10288,N_11331);
nor U13974 (N_13974,N_11205,N_10166);
nand U13975 (N_13975,N_11476,N_11799);
and U13976 (N_13976,N_10947,N_11707);
xor U13977 (N_13977,N_11205,N_10161);
nor U13978 (N_13978,N_11669,N_11252);
nor U13979 (N_13979,N_10934,N_11739);
nand U13980 (N_13980,N_10546,N_11440);
and U13981 (N_13981,N_11054,N_11184);
nor U13982 (N_13982,N_10788,N_11168);
nor U13983 (N_13983,N_10074,N_10654);
xnor U13984 (N_13984,N_10056,N_11364);
nand U13985 (N_13985,N_11747,N_11264);
xnor U13986 (N_13986,N_10115,N_10670);
and U13987 (N_13987,N_11660,N_10945);
or U13988 (N_13988,N_10483,N_10278);
nand U13989 (N_13989,N_11823,N_10785);
nor U13990 (N_13990,N_11911,N_11448);
and U13991 (N_13991,N_10517,N_11890);
nor U13992 (N_13992,N_11868,N_11682);
and U13993 (N_13993,N_10378,N_10025);
nor U13994 (N_13994,N_10911,N_11435);
nand U13995 (N_13995,N_11063,N_11585);
and U13996 (N_13996,N_10504,N_10778);
nand U13997 (N_13997,N_11672,N_11700);
xor U13998 (N_13998,N_10249,N_11864);
or U13999 (N_13999,N_10187,N_11771);
xnor U14000 (N_14000,N_13842,N_13920);
nor U14001 (N_14001,N_13848,N_12478);
or U14002 (N_14002,N_12785,N_13200);
xor U14003 (N_14003,N_13273,N_12739);
and U14004 (N_14004,N_12136,N_13220);
nand U14005 (N_14005,N_12466,N_13729);
nand U14006 (N_14006,N_13185,N_13977);
and U14007 (N_14007,N_13858,N_13707);
or U14008 (N_14008,N_12370,N_13950);
or U14009 (N_14009,N_13727,N_13219);
nor U14010 (N_14010,N_12449,N_12199);
nand U14011 (N_14011,N_12640,N_13597);
or U14012 (N_14012,N_13586,N_13009);
or U14013 (N_14013,N_13735,N_12108);
xnor U14014 (N_14014,N_12950,N_13202);
and U14015 (N_14015,N_12653,N_13557);
nand U14016 (N_14016,N_13154,N_13849);
or U14017 (N_14017,N_12485,N_12771);
and U14018 (N_14018,N_13008,N_12876);
and U14019 (N_14019,N_12709,N_12404);
xnor U14020 (N_14020,N_13462,N_12097);
or U14021 (N_14021,N_13109,N_13860);
and U14022 (N_14022,N_13545,N_12407);
or U14023 (N_14023,N_13436,N_13396);
or U14024 (N_14024,N_12593,N_12216);
xnor U14025 (N_14025,N_13603,N_13307);
nand U14026 (N_14026,N_12978,N_12123);
or U14027 (N_14027,N_13825,N_12169);
or U14028 (N_14028,N_12715,N_13136);
xor U14029 (N_14029,N_13286,N_12137);
nand U14030 (N_14030,N_12422,N_13340);
xnor U14031 (N_14031,N_12028,N_13405);
or U14032 (N_14032,N_12489,N_12657);
or U14033 (N_14033,N_13026,N_12079);
nand U14034 (N_14034,N_12113,N_12274);
nand U14035 (N_14035,N_13761,N_13048);
nand U14036 (N_14036,N_13177,N_13425);
or U14037 (N_14037,N_13775,N_13019);
nand U14038 (N_14038,N_13167,N_12026);
nor U14039 (N_14039,N_13995,N_13283);
and U14040 (N_14040,N_13492,N_13041);
and U14041 (N_14041,N_13728,N_13426);
xnor U14042 (N_14042,N_13745,N_13780);
nor U14043 (N_14043,N_13748,N_12387);
nand U14044 (N_14044,N_13631,N_13446);
and U14045 (N_14045,N_12458,N_12580);
or U14046 (N_14046,N_13148,N_13851);
or U14047 (N_14047,N_13166,N_13226);
nor U14048 (N_14048,N_13298,N_13933);
or U14049 (N_14049,N_13108,N_12763);
nor U14050 (N_14050,N_13675,N_13580);
and U14051 (N_14051,N_12822,N_13244);
xnor U14052 (N_14052,N_13990,N_12624);
or U14053 (N_14053,N_13938,N_13218);
xor U14054 (N_14054,N_12804,N_12821);
or U14055 (N_14055,N_12852,N_13628);
nor U14056 (N_14056,N_12985,N_12574);
or U14057 (N_14057,N_12234,N_13269);
or U14058 (N_14058,N_12179,N_13308);
xor U14059 (N_14059,N_13467,N_12164);
nor U14060 (N_14060,N_13355,N_12184);
and U14061 (N_14061,N_13186,N_12486);
and U14062 (N_14062,N_13326,N_13123);
and U14063 (N_14063,N_13310,N_12316);
or U14064 (N_14064,N_12887,N_13043);
xnor U14065 (N_14065,N_13556,N_12359);
nor U14066 (N_14066,N_13841,N_13316);
nor U14067 (N_14067,N_12987,N_13957);
xor U14068 (N_14068,N_12913,N_13481);
nor U14069 (N_14069,N_12718,N_13130);
nor U14070 (N_14070,N_12376,N_13655);
nand U14071 (N_14071,N_13968,N_12322);
nand U14072 (N_14072,N_13353,N_12143);
xor U14073 (N_14073,N_13407,N_12529);
or U14074 (N_14074,N_13335,N_12157);
and U14075 (N_14075,N_12282,N_12459);
xor U14076 (N_14076,N_12608,N_12297);
nor U14077 (N_14077,N_12454,N_13157);
and U14078 (N_14078,N_13179,N_13369);
nand U14079 (N_14079,N_13317,N_13767);
nor U14080 (N_14080,N_13888,N_13739);
xnor U14081 (N_14081,N_13757,N_13807);
xnor U14082 (N_14082,N_12540,N_13480);
and U14083 (N_14083,N_12884,N_12377);
or U14084 (N_14084,N_13502,N_13190);
and U14085 (N_14085,N_13708,N_13459);
nand U14086 (N_14086,N_12443,N_13869);
or U14087 (N_14087,N_13567,N_13354);
xor U14088 (N_14088,N_13798,N_12860);
nor U14089 (N_14089,N_12725,N_12154);
nand U14090 (N_14090,N_13371,N_13223);
and U14091 (N_14091,N_12135,N_13822);
or U14092 (N_14092,N_12545,N_13373);
nor U14093 (N_14093,N_12711,N_12740);
xnor U14094 (N_14094,N_12465,N_13653);
xor U14095 (N_14095,N_12835,N_12922);
nand U14096 (N_14096,N_13583,N_13550);
and U14097 (N_14097,N_13870,N_13656);
and U14098 (N_14098,N_13691,N_12895);
xor U14099 (N_14099,N_12500,N_12346);
nand U14100 (N_14100,N_13195,N_13730);
nor U14101 (N_14101,N_12348,N_13971);
nor U14102 (N_14102,N_13174,N_12746);
nand U14103 (N_14103,N_13922,N_13193);
and U14104 (N_14104,N_12535,N_12463);
nor U14105 (N_14105,N_13828,N_12567);
nand U14106 (N_14106,N_12923,N_12460);
and U14107 (N_14107,N_13051,N_12009);
and U14108 (N_14108,N_12921,N_12498);
xnor U14109 (N_14109,N_13515,N_13954);
nand U14110 (N_14110,N_13619,N_13036);
or U14111 (N_14111,N_12824,N_13577);
nor U14112 (N_14112,N_13855,N_12813);
and U14113 (N_14113,N_13209,N_12298);
or U14114 (N_14114,N_13769,N_12306);
xnor U14115 (N_14115,N_12668,N_13126);
nand U14116 (N_14116,N_13015,N_12770);
nand U14117 (N_14117,N_13912,N_12181);
nor U14118 (N_14118,N_13443,N_12564);
and U14119 (N_14119,N_12305,N_13164);
xor U14120 (N_14120,N_13027,N_13400);
or U14121 (N_14121,N_13958,N_13812);
nor U14122 (N_14122,N_13907,N_12066);
or U14123 (N_14123,N_13596,N_12243);
or U14124 (N_14124,N_12904,N_13790);
or U14125 (N_14125,N_12893,N_13339);
or U14126 (N_14126,N_12089,N_12937);
or U14127 (N_14127,N_13510,N_12111);
nor U14128 (N_14128,N_13948,N_12495);
and U14129 (N_14129,N_12237,N_13225);
and U14130 (N_14130,N_12033,N_12994);
or U14131 (N_14131,N_13248,N_13012);
and U14132 (N_14132,N_13342,N_12627);
nand U14133 (N_14133,N_12991,N_13444);
xor U14134 (N_14134,N_13089,N_12250);
or U14135 (N_14135,N_13584,N_12180);
nand U14136 (N_14136,N_13050,N_12035);
nand U14137 (N_14137,N_13319,N_13721);
xor U14138 (N_14138,N_12319,N_12434);
xor U14139 (N_14139,N_13824,N_12745);
nand U14140 (N_14140,N_12907,N_12114);
nor U14141 (N_14141,N_13724,N_12191);
or U14142 (N_14142,N_13097,N_12122);
nand U14143 (N_14143,N_12712,N_13623);
nor U14144 (N_14144,N_12866,N_12582);
nor U14145 (N_14145,N_13570,N_12132);
nor U14146 (N_14146,N_13213,N_12165);
nand U14147 (N_14147,N_12708,N_12787);
and U14148 (N_14148,N_12690,N_12563);
nor U14149 (N_14149,N_12871,N_13529);
nand U14150 (N_14150,N_13134,N_12816);
nor U14151 (N_14151,N_13093,N_13431);
or U14152 (N_14152,N_13245,N_13695);
and U14153 (N_14153,N_12810,N_12791);
or U14154 (N_14154,N_12431,N_12960);
nand U14155 (N_14155,N_12036,N_13266);
and U14156 (N_14156,N_12554,N_12008);
nor U14157 (N_14157,N_13331,N_13784);
nor U14158 (N_14158,N_13208,N_13676);
nor U14159 (N_14159,N_12899,N_12356);
and U14160 (N_14160,N_12766,N_12491);
nand U14161 (N_14161,N_12508,N_13387);
and U14162 (N_14162,N_12317,N_12217);
nor U14163 (N_14163,N_12772,N_13882);
xor U14164 (N_14164,N_12702,N_12340);
or U14165 (N_14165,N_13936,N_12743);
and U14166 (N_14166,N_13716,N_12192);
nor U14167 (N_14167,N_12286,N_13821);
and U14168 (N_14168,N_12737,N_13427);
xnor U14169 (N_14169,N_12902,N_12230);
and U14170 (N_14170,N_13294,N_13965);
and U14171 (N_14171,N_12476,N_12488);
or U14172 (N_14172,N_12006,N_12834);
or U14173 (N_14173,N_13531,N_13176);
or U14174 (N_14174,N_13081,N_13246);
xor U14175 (N_14175,N_13135,N_13839);
and U14176 (N_14176,N_13483,N_12461);
nor U14177 (N_14177,N_13018,N_12065);
or U14178 (N_14178,N_13474,N_12121);
and U14179 (N_14179,N_13258,N_13559);
xor U14180 (N_14180,N_13599,N_12932);
nand U14181 (N_14181,N_13039,N_12138);
nand U14182 (N_14182,N_13362,N_12717);
nand U14183 (N_14183,N_13463,N_12615);
nand U14184 (N_14184,N_12278,N_12330);
nor U14185 (N_14185,N_12644,N_12038);
or U14186 (N_14186,N_12205,N_13024);
nand U14187 (N_14187,N_12100,N_12981);
and U14188 (N_14188,N_13852,N_12012);
nor U14189 (N_14189,N_13100,N_13376);
or U14190 (N_14190,N_12676,N_12403);
nor U14191 (N_14191,N_13435,N_12856);
nor U14192 (N_14192,N_12505,N_13007);
or U14193 (N_14193,N_13428,N_12974);
nor U14194 (N_14194,N_13025,N_12558);
nand U14195 (N_14195,N_12213,N_12646);
and U14196 (N_14196,N_12185,N_13581);
nor U14197 (N_14197,N_12648,N_12757);
and U14198 (N_14198,N_13595,N_12117);
or U14199 (N_14199,N_12358,N_12130);
nand U14200 (N_14200,N_13891,N_12751);
nor U14201 (N_14201,N_12967,N_12722);
nor U14202 (N_14202,N_13062,N_12954);
nor U14203 (N_14203,N_13921,N_13061);
nand U14204 (N_14204,N_12609,N_12134);
nand U14205 (N_14205,N_13112,N_12936);
nand U14206 (N_14206,N_12384,N_13122);
or U14207 (N_14207,N_12728,N_12539);
xor U14208 (N_14208,N_13911,N_13713);
and U14209 (N_14209,N_13829,N_13890);
nor U14210 (N_14210,N_13830,N_13072);
and U14211 (N_14211,N_12694,N_13471);
or U14212 (N_14212,N_13259,N_12368);
nor U14213 (N_14213,N_12611,N_13329);
and U14214 (N_14214,N_12222,N_12010);
nand U14215 (N_14215,N_12801,N_12769);
nand U14216 (N_14216,N_13982,N_12156);
and U14217 (N_14217,N_12405,N_13189);
or U14218 (N_14218,N_12150,N_12617);
or U14219 (N_14219,N_12200,N_13650);
xor U14220 (N_14220,N_13447,N_12531);
and U14221 (N_14221,N_13408,N_13021);
nand U14222 (N_14222,N_13680,N_13734);
or U14223 (N_14223,N_12504,N_12517);
xor U14224 (N_14224,N_12252,N_12140);
nor U14225 (N_14225,N_12958,N_13278);
nand U14226 (N_14226,N_13850,N_12233);
nand U14227 (N_14227,N_12492,N_13344);
nand U14228 (N_14228,N_13832,N_13931);
and U14229 (N_14229,N_12828,N_13453);
xnor U14230 (N_14230,N_13641,N_13333);
nand U14231 (N_14231,N_12054,N_13605);
and U14232 (N_14232,N_13231,N_13486);
nor U14233 (N_14233,N_12750,N_12139);
nand U14234 (N_14234,N_13993,N_13296);
xnor U14235 (N_14235,N_12515,N_13017);
or U14236 (N_14236,N_13752,N_13658);
and U14237 (N_14237,N_12331,N_12920);
or U14238 (N_14238,N_12050,N_13334);
nand U14239 (N_14239,N_12383,N_13827);
and U14240 (N_14240,N_13667,N_12328);
nor U14241 (N_14241,N_13835,N_13293);
and U14242 (N_14242,N_12998,N_13733);
xor U14243 (N_14243,N_12208,N_12480);
nand U14244 (N_14244,N_13221,N_13366);
nor U14245 (N_14245,N_12326,N_13456);
or U14246 (N_14246,N_13636,N_12897);
xor U14247 (N_14247,N_13925,N_12912);
or U14248 (N_14248,N_13723,N_12170);
xnor U14249 (N_14249,N_12612,N_12968);
or U14250 (N_14250,N_12166,N_13038);
or U14251 (N_14251,N_12031,N_12979);
nor U14252 (N_14252,N_13183,N_12671);
nand U14253 (N_14253,N_12232,N_12412);
nand U14254 (N_14254,N_12736,N_13479);
nand U14255 (N_14255,N_13338,N_13929);
or U14256 (N_14256,N_12865,N_13698);
and U14257 (N_14257,N_13518,N_13146);
or U14258 (N_14258,N_13992,N_13101);
nand U14259 (N_14259,N_13528,N_13624);
or U14260 (N_14260,N_12416,N_13859);
xnor U14261 (N_14261,N_13356,N_13212);
or U14262 (N_14262,N_12837,N_12396);
and U14263 (N_14263,N_12355,N_12919);
nor U14264 (N_14264,N_13493,N_13766);
or U14265 (N_14265,N_13401,N_13254);
nor U14266 (N_14266,N_13924,N_13153);
and U14267 (N_14267,N_12889,N_13845);
nor U14268 (N_14268,N_12879,N_12992);
nand U14269 (N_14269,N_12318,N_13168);
nor U14270 (N_14270,N_12275,N_12613);
and U14271 (N_14271,N_12053,N_13458);
nor U14272 (N_14272,N_13332,N_12586);
and U14273 (N_14273,N_13063,N_12104);
xnor U14274 (N_14274,N_12151,N_12324);
nand U14275 (N_14275,N_12778,N_12189);
or U14276 (N_14276,N_12814,N_13171);
or U14277 (N_14277,N_13881,N_12579);
nand U14278 (N_14278,N_12313,N_12684);
and U14279 (N_14279,N_12691,N_12302);
nand U14280 (N_14280,N_13610,N_13525);
or U14281 (N_14281,N_13074,N_13607);
nor U14282 (N_14282,N_12565,N_13274);
nor U14283 (N_14283,N_13065,N_13934);
and U14284 (N_14284,N_12990,N_12797);
xor U14285 (N_14285,N_12246,N_12409);
or U14286 (N_14286,N_12452,N_12048);
or U14287 (N_14287,N_12490,N_13465);
nand U14288 (N_14288,N_13945,N_13626);
and U14289 (N_14289,N_12367,N_13216);
xor U14290 (N_14290,N_13726,N_13660);
or U14291 (N_14291,N_12872,N_12426);
nand U14292 (N_14292,N_13685,N_12578);
and U14293 (N_14293,N_13546,N_12249);
xor U14294 (N_14294,N_12914,N_12686);
nor U14295 (N_14295,N_12842,N_13141);
and U14296 (N_14296,N_12955,N_13276);
nor U14297 (N_14297,N_13360,N_12072);
or U14298 (N_14298,N_13833,N_13527);
xor U14299 (N_14299,N_13196,N_13969);
nand U14300 (N_14300,N_13256,N_13070);
xnor U14301 (N_14301,N_13406,N_13121);
nand U14302 (N_14302,N_13295,N_13380);
and U14303 (N_14303,N_13511,N_13944);
xor U14304 (N_14304,N_13159,N_13170);
and U14305 (N_14305,N_13949,N_12481);
and U14306 (N_14306,N_12989,N_13238);
nor U14307 (N_14307,N_12850,N_13002);
nor U14308 (N_14308,N_12680,N_13608);
nand U14309 (N_14309,N_12183,N_13395);
or U14310 (N_14310,N_13746,N_13424);
xnor U14311 (N_14311,N_13661,N_12083);
or U14312 (N_14312,N_13306,N_13918);
and U14313 (N_14313,N_12204,N_13811);
or U14314 (N_14314,N_13421,N_12758);
nor U14315 (N_14315,N_12004,N_12647);
xnor U14316 (N_14316,N_13538,N_12716);
nand U14317 (N_14317,N_13184,N_13438);
xor U14318 (N_14318,N_12748,N_13604);
or U14319 (N_14319,N_13322,N_12357);
nand U14320 (N_14320,N_13674,N_13489);
or U14321 (N_14321,N_13782,N_13533);
or U14322 (N_14322,N_12337,N_12524);
and U14323 (N_14323,N_13145,N_13482);
or U14324 (N_14324,N_12174,N_12811);
or U14325 (N_14325,N_12953,N_13302);
nand U14326 (N_14326,N_13020,N_12756);
nor U14327 (N_14327,N_13016,N_12650);
nor U14328 (N_14328,N_12947,N_12543);
and U14329 (N_14329,N_12142,N_12090);
nand U14330 (N_14330,N_12327,N_13037);
xor U14331 (N_14331,N_12765,N_13996);
and U14332 (N_14332,N_13553,N_12941);
xnor U14333 (N_14333,N_13867,N_12501);
and U14334 (N_14334,N_13885,N_13840);
nor U14335 (N_14335,N_13771,N_13098);
nor U14336 (N_14336,N_13499,N_13290);
nand U14337 (N_14337,N_12291,N_12060);
nor U14338 (N_14338,N_12794,N_12528);
xnor U14339 (N_14339,N_13683,N_13067);
nand U14340 (N_14340,N_13336,N_12752);
and U14341 (N_14341,N_13682,N_12323);
xor U14342 (N_14342,N_12670,N_12051);
nor U14343 (N_14343,N_13011,N_13614);
xor U14344 (N_14344,N_12016,N_12020);
and U14345 (N_14345,N_12263,N_13301);
xnor U14346 (N_14346,N_12070,N_13473);
or U14347 (N_14347,N_13742,N_13343);
nor U14348 (N_14348,N_13740,N_12753);
xor U14349 (N_14349,N_13133,N_12632);
or U14350 (N_14350,N_13498,N_13383);
nor U14351 (N_14351,N_13684,N_13455);
and U14352 (N_14352,N_13588,N_13073);
and U14353 (N_14353,N_13536,N_13909);
and U14354 (N_14354,N_12957,N_12497);
or U14355 (N_14355,N_12812,N_13071);
nand U14356 (N_14356,N_12479,N_12602);
or U14357 (N_14357,N_12761,N_12069);
xor U14358 (N_14358,N_12553,N_12639);
or U14359 (N_14359,N_12364,N_13429);
nand U14360 (N_14360,N_13787,N_13388);
xor U14361 (N_14361,N_13468,N_12127);
nand U14362 (N_14362,N_13363,N_13142);
or U14363 (N_14363,N_12862,N_12555);
or U14364 (N_14364,N_12915,N_12710);
and U14365 (N_14365,N_13670,N_13699);
nand U14366 (N_14366,N_13215,N_13994);
and U14367 (N_14367,N_13540,N_12910);
or U14368 (N_14368,N_12583,N_12312);
xor U14369 (N_14369,N_12764,N_13591);
or U14370 (N_14370,N_13928,N_13230);
xor U14371 (N_14371,N_13173,N_12571);
or U14372 (N_14372,N_13242,N_13519);
xor U14373 (N_14373,N_12874,N_12547);
and U14374 (N_14374,N_12663,N_13878);
xnor U14375 (N_14375,N_12456,N_12868);
and U14376 (N_14376,N_13694,N_12848);
or U14377 (N_14377,N_13741,N_12429);
or U14378 (N_14378,N_12264,N_12587);
nand U14379 (N_14379,N_12621,N_12432);
or U14380 (N_14380,N_12641,N_13127);
and U14381 (N_14381,N_13432,N_12982);
nand U14382 (N_14382,N_13495,N_13399);
or U14383 (N_14383,N_13715,N_12858);
or U14384 (N_14384,N_13814,N_13955);
nor U14385 (N_14385,N_12825,N_13114);
xor U14386 (N_14386,N_13714,N_12986);
and U14387 (N_14387,N_12197,N_12017);
nand U14388 (N_14388,N_12148,N_13884);
or U14389 (N_14389,N_13304,N_13198);
xor U14390 (N_14390,N_13485,N_13697);
and U14391 (N_14391,N_13935,N_12883);
nor U14392 (N_14392,N_13454,N_12056);
xor U14393 (N_14393,N_13789,N_13379);
or U14394 (N_14394,N_13452,N_12342);
or U14395 (N_14395,N_13612,N_13594);
xnor U14396 (N_14396,N_12800,N_12839);
xor U14397 (N_14397,N_12354,N_13357);
and U14398 (N_14398,N_13111,N_12236);
and U14399 (N_14399,N_12175,N_12352);
or U14400 (N_14400,N_13629,N_12125);
and U14401 (N_14401,N_13345,N_13253);
or U14402 (N_14402,N_12831,N_12532);
and U14403 (N_14403,N_12229,N_13169);
nand U14404 (N_14404,N_12190,N_13129);
xnor U14405 (N_14405,N_12417,N_13573);
xnor U14406 (N_14406,N_12462,N_13265);
and U14407 (N_14407,N_13564,N_13055);
and U14408 (N_14408,N_12662,N_13664);
or U14409 (N_14409,N_12436,N_12406);
nand U14410 (N_14410,N_12116,N_12043);
and U14411 (N_14411,N_13693,N_12704);
and U14412 (N_14412,N_12546,N_12444);
xnor U14413 (N_14413,N_13116,N_13523);
or U14414 (N_14414,N_13764,N_13854);
nor U14415 (N_14415,N_12254,N_13460);
or U14416 (N_14416,N_13774,N_12413);
nor U14417 (N_14417,N_13252,N_12636);
or U14418 (N_14418,N_13417,N_12258);
and U14419 (N_14419,N_13617,N_13543);
nand U14420 (N_14420,N_13033,N_12167);
or U14421 (N_14421,N_13064,N_13720);
nor U14422 (N_14422,N_13743,N_13625);
or U14423 (N_14423,N_13535,N_12892);
and U14424 (N_14424,N_13413,N_13902);
nand U14425 (N_14425,N_13576,N_13961);
and U14426 (N_14426,N_12000,N_12424);
and U14427 (N_14427,N_12561,N_13908);
or U14428 (N_14428,N_13541,N_12378);
nor U14429 (N_14429,N_12178,N_12956);
and U14430 (N_14430,N_12362,N_12929);
or U14431 (N_14431,N_12988,N_12091);
nor U14432 (N_14432,N_13337,N_13346);
or U14433 (N_14433,N_13005,N_12360);
or U14434 (N_14434,N_13799,N_13967);
xor U14435 (N_14435,N_13781,N_12518);
nor U14436 (N_14436,N_13669,N_12369);
or U14437 (N_14437,N_13754,N_12202);
xnor U14438 (N_14438,N_13247,N_12253);
and U14439 (N_14439,N_12724,N_13505);
or U14440 (N_14440,N_13420,N_12799);
and U14441 (N_14441,N_13937,N_12240);
xnor U14442 (N_14442,N_13770,N_12864);
or U14443 (N_14443,N_12939,N_12300);
and U14444 (N_14444,N_13466,N_13320);
and U14445 (N_14445,N_13192,N_13368);
nor U14446 (N_14446,N_13156,N_13110);
nor U14447 (N_14447,N_12818,N_12102);
or U14448 (N_14448,N_13520,N_12714);
and U14449 (N_14449,N_12503,N_13364);
and U14450 (N_14450,N_13889,N_12059);
nand U14451 (N_14451,N_13046,N_13779);
nand U14452 (N_14452,N_12271,N_13287);
nand U14453 (N_14453,N_12682,N_12350);
and U14454 (N_14454,N_12851,N_12983);
and U14455 (N_14455,N_13914,N_12666);
or U14456 (N_14456,N_12777,N_12141);
nand U14457 (N_14457,N_12610,N_12410);
or U14458 (N_14458,N_13052,N_12194);
nand U14459 (N_14459,N_13834,N_12133);
and U14460 (N_14460,N_12128,N_13214);
nand U14461 (N_14461,N_13386,N_12262);
nor U14462 (N_14462,N_12219,N_12206);
nand U14463 (N_14463,N_13415,N_13088);
or U14464 (N_14464,N_13501,N_13554);
or U14465 (N_14465,N_13987,N_12833);
nor U14466 (N_14466,N_13906,N_13919);
or U14467 (N_14467,N_12341,N_13158);
nor U14468 (N_14468,N_12906,N_13702);
and U14469 (N_14469,N_13517,N_12427);
or U14470 (N_14470,N_13644,N_13497);
nor U14471 (N_14471,N_13140,N_12082);
nor U14472 (N_14472,N_12296,N_13289);
nor U14473 (N_14473,N_12177,N_13989);
and U14474 (N_14474,N_13255,N_12699);
or U14475 (N_14475,N_12293,N_13440);
nor U14476 (N_14476,N_13351,N_12999);
nor U14477 (N_14477,N_13513,N_12373);
and U14478 (N_14478,N_12707,N_12507);
and U14479 (N_14479,N_13817,N_13251);
and U14480 (N_14480,N_12024,N_13117);
xnor U14481 (N_14481,N_13677,N_12599);
nand U14482 (N_14482,N_12701,N_13975);
and U14483 (N_14483,N_12115,N_13374);
nand U14484 (N_14484,N_13392,N_12964);
nor U14485 (N_14485,N_12273,N_13753);
and U14486 (N_14486,N_13946,N_12631);
xnor U14487 (N_14487,N_12329,N_13621);
nor U14488 (N_14488,N_13054,N_12415);
nand U14489 (N_14489,N_13516,N_13325);
nand U14490 (N_14490,N_12677,N_13940);
nand U14491 (N_14491,N_13899,N_12841);
xor U14492 (N_14492,N_12629,N_13942);
or U14493 (N_14493,N_13279,N_12645);
nand U14494 (N_14494,N_12855,N_13657);
and U14495 (N_14495,N_13365,N_12095);
nand U14496 (N_14496,N_12015,N_12391);
nor U14497 (N_14497,N_12103,N_13865);
nor U14498 (N_14498,N_12863,N_13671);
xnor U14499 (N_14499,N_13330,N_13321);
xnor U14500 (N_14500,N_13441,N_12534);
and U14501 (N_14501,N_13563,N_13659);
and U14502 (N_14502,N_13182,N_12487);
and U14503 (N_14503,N_13506,N_12658);
and U14504 (N_14504,N_13926,N_13272);
nor U14505 (N_14505,N_13000,N_13587);
xnor U14506 (N_14506,N_12642,N_12594);
xnor U14507 (N_14507,N_13871,N_12042);
or U14508 (N_14508,N_12592,N_12679);
xor U14509 (N_14509,N_12162,N_12786);
or U14510 (N_14510,N_13512,N_12109);
and U14511 (N_14511,N_12394,N_12651);
xor U14512 (N_14512,N_12533,N_13045);
xnor U14513 (N_14513,N_12802,N_12420);
nand U14514 (N_14514,N_13076,N_13205);
or U14515 (N_14515,N_12457,N_12938);
nor U14516 (N_14516,N_13023,N_12502);
xor U14517 (N_14517,N_12626,N_12309);
nor U14518 (N_14518,N_13470,N_13393);
xnor U14519 (N_14519,N_13795,N_13710);
nand U14520 (N_14520,N_12542,N_12014);
or U14521 (N_14521,N_12965,N_12944);
nand U14522 (N_14522,N_13566,N_13281);
xor U14523 (N_14523,N_12520,N_12926);
nor U14524 (N_14524,N_12093,N_13377);
nand U14525 (N_14525,N_12288,N_12908);
xor U14526 (N_14526,N_12007,N_12361);
nand U14527 (N_14527,N_12073,N_13075);
nor U14528 (N_14528,N_13305,N_12380);
nor U14529 (N_14529,N_13923,N_13616);
xnor U14530 (N_14530,N_12916,N_12187);
nor U14531 (N_14531,N_12519,N_13547);
nand U14532 (N_14532,N_13738,N_13778);
nand U14533 (N_14533,N_13905,N_13391);
nand U14534 (N_14534,N_12898,N_12075);
or U14535 (N_14535,N_13235,N_12727);
nand U14536 (N_14536,N_13143,N_13986);
xor U14537 (N_14537,N_12838,N_12244);
xnor U14538 (N_14538,N_13598,N_12061);
or U14539 (N_14539,N_12159,N_13144);
xor U14540 (N_14540,N_13125,N_13662);
xor U14541 (N_14541,N_12269,N_13652);
nand U14542 (N_14542,N_13261,N_12225);
nand U14543 (N_14543,N_13233,N_12032);
xnor U14544 (N_14544,N_13087,N_13791);
and U14545 (N_14545,N_13537,N_13763);
or U14546 (N_14546,N_13194,N_13115);
and U14547 (N_14547,N_12857,N_12210);
nor U14548 (N_14548,N_13758,N_12685);
nor U14549 (N_14549,N_13705,N_13032);
xor U14550 (N_14550,N_12146,N_13894);
nand U14551 (N_14551,N_12656,N_13224);
xnor U14552 (N_14552,N_12793,N_13375);
nor U14553 (N_14553,N_12451,N_12438);
and U14554 (N_14554,N_12019,N_12034);
and U14555 (N_14555,N_12667,N_12976);
or U14556 (N_14556,N_13551,N_13820);
and U14557 (N_14557,N_12966,N_12696);
xor U14558 (N_14558,N_12847,N_13382);
nand U14559 (N_14559,N_12226,N_13359);
or U14560 (N_14560,N_12882,N_12675);
and U14561 (N_14561,N_12755,N_12849);
nand U14562 (N_14562,N_12803,N_13056);
or U14563 (N_14563,N_12430,N_12112);
or U14564 (N_14564,N_13449,N_12759);
or U14565 (N_14565,N_13574,N_13737);
or U14566 (N_14566,N_12314,N_12596);
nand U14567 (N_14567,N_12266,N_13347);
nand U14568 (N_14568,N_12484,N_13491);
or U14569 (N_14569,N_12927,N_12494);
or U14570 (N_14570,N_12347,N_13999);
and U14571 (N_14571,N_13084,N_13010);
xnor U14572 (N_14572,N_12940,N_13836);
or U14573 (N_14573,N_13309,N_12468);
nor U14574 (N_14574,N_12760,N_13507);
nor U14575 (N_14575,N_12762,N_12683);
xor U14576 (N_14576,N_13217,N_12975);
nor U14577 (N_14577,N_13947,N_13119);
xor U14578 (N_14578,N_12301,N_13750);
nand U14579 (N_14579,N_12493,N_12562);
nand U14580 (N_14580,N_12344,N_13423);
nor U14581 (N_14581,N_12076,N_12723);
nor U14582 (N_14582,N_13718,N_12094);
xor U14583 (N_14583,N_13719,N_13409);
nand U14584 (N_14584,N_13679,N_13262);
or U14585 (N_14585,N_13606,N_12623);
and U14586 (N_14586,N_12315,N_12078);
xor U14587 (N_14587,N_12238,N_13916);
and U14588 (N_14588,N_13412,N_12455);
and U14589 (N_14589,N_12351,N_12211);
nand U14590 (N_14590,N_12550,N_13856);
or U14591 (N_14591,N_13910,N_12433);
nand U14592 (N_14592,N_13210,N_13068);
or U14593 (N_14593,N_13096,N_13260);
or U14594 (N_14594,N_13701,N_12823);
or U14595 (N_14595,N_13128,N_13956);
and U14596 (N_14596,N_12290,N_12124);
or U14597 (N_14597,N_12209,N_13418);
nor U14598 (N_14598,N_13837,N_13029);
or U14599 (N_14599,N_12055,N_13901);
and U14600 (N_14600,N_12446,N_12721);
nor U14601 (N_14601,N_13241,N_13651);
nand U14602 (N_14602,N_12276,N_12660);
xnor U14603 (N_14603,N_13349,N_13264);
and U14604 (N_14604,N_12552,N_13285);
or U14605 (N_14605,N_13288,N_12730);
and U14606 (N_14606,N_13756,N_13542);
xor U14607 (N_14607,N_12633,N_12447);
and U14608 (N_14608,N_13804,N_12603);
xnor U14609 (N_14609,N_13149,N_13960);
xor U14610 (N_14610,N_13280,N_12654);
and U14611 (N_14611,N_12469,N_13561);
and U14612 (N_14612,N_12379,N_12227);
xor U14613 (N_14613,N_12005,N_12310);
xor U14614 (N_14614,N_13985,N_13138);
nand U14615 (N_14615,N_12840,N_13654);
nand U14616 (N_14616,N_12414,N_13549);
or U14617 (N_14617,N_13451,N_13951);
nand U14618 (N_14618,N_13430,N_13323);
xnor U14619 (N_14619,N_13797,N_13736);
xnor U14620 (N_14620,N_12098,N_13042);
nand U14621 (N_14621,N_13866,N_13394);
xor U14622 (N_14622,N_12477,N_12577);
and U14623 (N_14623,N_13139,N_12689);
nor U14624 (N_14624,N_13411,N_12706);
or U14625 (N_14625,N_12375,N_12581);
nor U14626 (N_14626,N_13469,N_12106);
or U14627 (N_14627,N_13303,N_13777);
or U14628 (N_14628,N_13952,N_12516);
nor U14629 (N_14629,N_13892,N_12788);
nand U14630 (N_14630,N_12289,N_13284);
nor U14631 (N_14631,N_13297,N_13900);
nand U14632 (N_14632,N_13978,N_13530);
xor U14633 (N_14633,N_12147,N_13378);
and U14634 (N_14634,N_12513,N_13979);
xnor U14635 (N_14635,N_13991,N_12203);
or U14636 (N_14636,N_12129,N_13861);
or U14637 (N_14637,N_12619,N_13234);
and U14638 (N_14638,N_13700,N_12280);
or U14639 (N_14639,N_12092,N_13472);
nor U14640 (N_14640,N_12742,N_12620);
nor U14641 (N_14641,N_12248,N_12172);
or U14642 (N_14642,N_13592,N_12638);
or U14643 (N_14643,N_12809,N_13602);
nand U14644 (N_14644,N_13282,N_12120);
or U14645 (N_14645,N_12844,N_12928);
or U14646 (N_14646,N_12040,N_12901);
xor U14647 (N_14647,N_12635,N_12085);
nor U14648 (N_14648,N_13959,N_13092);
nand U14649 (N_14649,N_12836,N_12984);
nor U14650 (N_14650,N_13001,N_12496);
and U14651 (N_14651,N_13877,N_13893);
xnor U14652 (N_14652,N_12107,N_12002);
and U14653 (N_14653,N_13800,N_13204);
nor U14654 (N_14654,N_13494,N_13161);
nor U14655 (N_14655,N_12784,N_12946);
nor U14656 (N_14656,N_12559,N_12652);
and U14657 (N_14657,N_12437,N_12925);
nor U14658 (N_14658,N_13620,N_12399);
or U14659 (N_14659,N_12891,N_13786);
or U14660 (N_14660,N_12201,N_13448);
nand U14661 (N_14661,N_12163,N_12338);
or U14662 (N_14662,N_12086,N_13103);
and U14663 (N_14663,N_13270,N_13639);
xor U14664 (N_14664,N_12397,N_13666);
and U14665 (N_14665,N_12080,N_13083);
nand U14666 (N_14666,N_13590,N_13402);
xor U14667 (N_14667,N_12597,N_12931);
xor U14668 (N_14668,N_12972,N_13299);
or U14669 (N_14669,N_13095,N_13222);
xnor U14670 (N_14670,N_13291,N_12295);
nand U14671 (N_14671,N_12118,N_12695);
and U14672 (N_14672,N_12817,N_12470);
or U14673 (N_14673,N_12713,N_13521);
xnor U14674 (N_14674,N_12428,N_12256);
nand U14675 (N_14675,N_12336,N_12158);
and U14676 (N_14676,N_13328,N_13105);
or U14677 (N_14677,N_13793,N_12659);
and U14678 (N_14678,N_13014,N_13783);
nand U14679 (N_14679,N_13404,N_12917);
and U14680 (N_14680,N_13818,N_12467);
nand U14681 (N_14681,N_13348,N_12588);
nand U14682 (N_14682,N_13410,N_13381);
xor U14683 (N_14683,N_12726,N_12231);
or U14684 (N_14684,N_13803,N_12569);
nand U14685 (N_14685,N_13689,N_13953);
xnor U14686 (N_14686,N_12214,N_12285);
nand U14687 (N_14687,N_13484,N_13751);
and U14688 (N_14688,N_12768,N_12830);
xnor U14689 (N_14689,N_12870,N_13846);
nand U14690 (N_14690,N_13227,N_13663);
xor U14691 (N_14691,N_12149,N_12145);
xnor U14692 (N_14692,N_13648,N_12933);
nand U14693 (N_14693,N_13236,N_13090);
nor U14694 (N_14694,N_13981,N_12307);
and U14695 (N_14695,N_13006,N_12353);
nor U14696 (N_14696,N_12071,N_12930);
nor U14697 (N_14697,N_13106,N_13647);
or U14698 (N_14698,N_12995,N_12924);
xnor U14699 (N_14699,N_12464,N_13600);
xor U14700 (N_14700,N_12997,N_13522);
and U14701 (N_14701,N_12678,N_12267);
or U14702 (N_14702,N_12119,N_13880);
nor U14703 (N_14703,N_12993,N_13998);
or U14704 (N_14704,N_12780,N_13532);
xnor U14705 (N_14705,N_12512,N_12945);
xor U14706 (N_14706,N_12909,N_12698);
or U14707 (N_14707,N_13450,N_13500);
and U14708 (N_14708,N_13589,N_12084);
nand U14709 (N_14709,N_12962,N_12747);
nor U14710 (N_14710,N_12025,N_13257);
and U14711 (N_14711,N_13442,N_13915);
and U14712 (N_14712,N_13988,N_12029);
and U14713 (N_14713,N_12700,N_13028);
and U14714 (N_14714,N_13311,N_12789);
and U14715 (N_14715,N_12959,N_12878);
and U14716 (N_14716,N_13579,N_13895);
and U14717 (N_14717,N_13147,N_13477);
or U14718 (N_14718,N_13197,N_13461);
nor U14719 (N_14719,N_13414,N_13731);
or U14720 (N_14720,N_12027,N_13879);
nor U14721 (N_14721,N_12257,N_13524);
xor U14722 (N_14722,N_12215,N_12845);
nor U14723 (N_14723,N_13886,N_13646);
xor U14724 (N_14724,N_12160,N_12198);
nand U14725 (N_14725,N_12510,N_12400);
or U14726 (N_14726,N_13358,N_12536);
nor U14727 (N_14727,N_13060,N_12819);
or U14728 (N_14728,N_12905,N_12401);
nand U14729 (N_14729,N_13815,N_13180);
nand U14730 (N_14730,N_12475,N_12692);
or U14731 (N_14731,N_12894,N_12411);
or U14732 (N_14732,N_12506,N_12212);
xor U14733 (N_14733,N_13372,N_12321);
nor U14734 (N_14734,N_13904,N_13615);
nor U14735 (N_14735,N_12885,N_12294);
and U14736 (N_14736,N_13160,N_13044);
nand U14737 (N_14737,N_13792,N_13268);
and U14738 (N_14738,N_12445,N_13030);
xor U14739 (N_14739,N_12473,N_13571);
and U14740 (N_14740,N_12221,N_12873);
or U14741 (N_14741,N_13047,N_13941);
nand U14742 (N_14742,N_13562,N_13250);
and U14743 (N_14743,N_12105,N_12441);
xor U14744 (N_14744,N_12022,N_13678);
and U14745 (N_14745,N_13565,N_13984);
nand U14746 (N_14746,N_12688,N_12886);
or U14747 (N_14747,N_12334,N_13609);
xnor U14748 (N_14748,N_13434,N_12349);
xor U14749 (N_14749,N_12176,N_12585);
nor U14750 (N_14750,N_12182,N_12733);
or U14751 (N_14751,N_12074,N_13178);
xor U14752 (N_14752,N_12731,N_12013);
xnor U14753 (N_14753,N_12867,N_12241);
and U14754 (N_14754,N_12021,N_12283);
and U14755 (N_14755,N_13749,N_13802);
nand U14756 (N_14756,N_13099,N_13082);
xor U14757 (N_14757,N_13843,N_13643);
nand U14758 (N_14758,N_12796,N_12365);
nor U14759 (N_14759,N_12661,N_12807);
or U14760 (N_14760,N_12570,N_13640);
and U14761 (N_14761,N_13318,N_13022);
and U14762 (N_14762,N_13514,N_13341);
nor U14763 (N_14763,N_13077,N_12573);
or U14764 (N_14764,N_13898,N_13544);
xnor U14765 (N_14765,N_13788,N_13690);
xor U14766 (N_14766,N_13091,N_13124);
nor U14767 (N_14767,N_12062,N_13352);
xnor U14768 (N_14768,N_13172,N_12186);
or U14769 (N_14769,N_12450,N_12284);
nor U14770 (N_14770,N_13973,N_12792);
or U14771 (N_14771,N_12511,N_13211);
nor U14772 (N_14772,N_12228,N_13903);
xnor U14773 (N_14773,N_13635,N_13887);
xnor U14774 (N_14774,N_12382,N_13243);
or U14775 (N_14775,N_12096,N_13593);
xor U14776 (N_14776,N_13131,N_13004);
and U14777 (N_14777,N_12265,N_13107);
and U14778 (N_14778,N_12155,N_13206);
or U14779 (N_14779,N_12260,N_12538);
nand U14780 (N_14780,N_13873,N_13805);
xnor U14781 (N_14781,N_13162,N_12499);
nor U14782 (N_14782,N_13966,N_12077);
nand U14783 (N_14783,N_12196,N_13709);
or U14784 (N_14784,N_12223,N_13712);
nor U14785 (N_14785,N_12372,N_12308);
nand U14786 (N_14786,N_13367,N_13229);
and U14787 (N_14787,N_13203,N_13872);
nand U14788 (N_14788,N_13445,N_12859);
nor U14789 (N_14789,N_13085,N_12977);
nor U14790 (N_14790,N_13575,N_12669);
xnor U14791 (N_14791,N_13181,N_13132);
or U14792 (N_14792,N_12598,N_12037);
xor U14793 (N_14793,N_13692,N_13673);
xor U14794 (N_14794,N_13155,N_13104);
nand U14795 (N_14795,N_12949,N_12101);
nor U14796 (N_14796,N_13275,N_12744);
xor U14797 (N_14797,N_12418,N_12600);
and U14798 (N_14798,N_12943,N_13526);
and U14799 (N_14799,N_13207,N_12398);
nand U14800 (N_14800,N_13534,N_12846);
nor U14801 (N_14801,N_13943,N_12948);
nor U14802 (N_14802,N_13686,N_12126);
xor U14803 (N_14803,N_12903,N_13040);
or U14804 (N_14804,N_12687,N_13853);
or U14805 (N_14805,N_13237,N_12299);
nor U14806 (N_14806,N_12934,N_12333);
and U14807 (N_14807,N_13755,N_12734);
nor U14808 (N_14808,N_12729,N_12058);
nand U14809 (N_14809,N_12530,N_12435);
nor U14810 (N_14810,N_13403,N_12408);
xor U14811 (N_14811,N_12390,N_13964);
and U14812 (N_14812,N_12767,N_12325);
and U14813 (N_14813,N_13794,N_12442);
or U14814 (N_14814,N_12649,N_13188);
and U14815 (N_14815,N_13863,N_12952);
xor U14816 (N_14816,N_13582,N_12514);
and U14817 (N_14817,N_12808,N_13416);
nor U14818 (N_14818,N_13725,N_12402);
xnor U14819 (N_14819,N_12595,N_13503);
xor U14820 (N_14820,N_13831,N_13927);
nor U14821 (N_14821,N_13560,N_13312);
nand U14822 (N_14822,N_13118,N_12281);
xnor U14823 (N_14823,N_12386,N_13370);
and U14824 (N_14824,N_13199,N_13816);
nor U14825 (N_14825,N_13810,N_12173);
nor U14826 (N_14826,N_12526,N_13476);
nor U14827 (N_14827,N_13972,N_13475);
nor U14828 (N_14828,N_12047,N_12311);
xnor U14829 (N_14829,N_12782,N_13433);
xnor U14830 (N_14830,N_12332,N_12052);
nand U14831 (N_14831,N_13496,N_12820);
or U14832 (N_14832,N_13398,N_13747);
xnor U14833 (N_14833,N_13706,N_12614);
nand U14834 (N_14834,N_12601,N_12371);
or U14835 (N_14835,N_12239,N_12970);
nor U14836 (N_14836,N_13760,N_13630);
and U14837 (N_14837,N_13868,N_12969);
or U14838 (N_14838,N_12279,N_12393);
nor U14839 (N_14839,N_13759,N_13315);
nor U14840 (N_14840,N_13552,N_12888);
or U14841 (N_14841,N_13437,N_13585);
and U14842 (N_14842,N_13883,N_12440);
or U14843 (N_14843,N_12754,N_13696);
nand U14844 (N_14844,N_12935,N_12732);
xor U14845 (N_14845,N_12735,N_13645);
or U14846 (N_14846,N_12703,N_12087);
or U14847 (N_14847,N_12277,N_12423);
and U14848 (N_14848,N_12951,N_13980);
nor U14849 (N_14849,N_13249,N_12304);
or U14850 (N_14850,N_12011,N_13508);
nand U14851 (N_14851,N_13069,N_13053);
nand U14852 (N_14852,N_12374,N_13102);
or U14853 (N_14853,N_13930,N_13151);
or U14854 (N_14854,N_12303,N_13031);
nand U14855 (N_14855,N_12591,N_13704);
nand U14856 (N_14856,N_12483,N_12131);
nor U14857 (N_14857,N_13819,N_12551);
xnor U14858 (N_14858,N_12245,N_12673);
and U14859 (N_14859,N_13913,N_13633);
nor U14860 (N_14860,N_13490,N_12590);
or U14861 (N_14861,N_12247,N_13847);
nand U14862 (N_14862,N_12482,N_12693);
xnor U14863 (N_14863,N_12439,N_13801);
nand U14864 (N_14864,N_13773,N_13113);
and U14865 (N_14865,N_13478,N_13634);
xnor U14866 (N_14866,N_13240,N_12081);
and U14867 (N_14867,N_12161,N_12068);
nand U14868 (N_14868,N_12171,N_13876);
or U14869 (N_14869,N_12971,N_12544);
or U14870 (N_14870,N_12890,N_13300);
and U14871 (N_14871,N_12815,N_12843);
xor U14872 (N_14872,N_13711,N_13613);
nand U14873 (N_14873,N_13350,N_13917);
nor U14874 (N_14874,N_12541,N_13385);
nor U14875 (N_14875,N_13687,N_12255);
and U14876 (N_14876,N_13601,N_12790);
xnor U14877 (N_14877,N_12207,N_13638);
nor U14878 (N_14878,N_12144,N_12057);
or U14879 (N_14879,N_12572,N_13267);
nor U14880 (N_14880,N_13163,N_12041);
or U14881 (N_14881,N_12618,N_12655);
and U14882 (N_14882,N_12522,N_13120);
and U14883 (N_14883,N_12001,N_12634);
xor U14884 (N_14884,N_13397,N_13997);
nor U14885 (N_14885,N_12474,N_12749);
nor U14886 (N_14886,N_12900,N_12388);
nor U14887 (N_14887,N_13569,N_13717);
or U14888 (N_14888,N_12272,N_12829);
xor U14889 (N_14889,N_13013,N_12425);
nand U14890 (N_14890,N_12681,N_12854);
or U14891 (N_14891,N_13578,N_12044);
or U14892 (N_14892,N_12259,N_13419);
nor U14893 (N_14893,N_12911,N_13049);
xnor U14894 (N_14894,N_13324,N_13744);
nor U14895 (N_14895,N_12039,N_12616);
nand U14896 (N_14896,N_12576,N_12099);
xor U14897 (N_14897,N_13983,N_13384);
nand U14898 (N_14898,N_12339,N_12381);
nor U14899 (N_14899,N_13932,N_13703);
and U14900 (N_14900,N_13313,N_13539);
nand U14901 (N_14901,N_13642,N_12063);
nor U14902 (N_14902,N_12973,N_12881);
nor U14903 (N_14903,N_12861,N_13504);
or U14904 (N_14904,N_13080,N_12509);
and U14905 (N_14905,N_13875,N_13813);
nand U14906 (N_14906,N_12961,N_13035);
or U14907 (N_14907,N_12674,N_13864);
nand U14908 (N_14908,N_12049,N_13732);
nand U14909 (N_14909,N_13962,N_12775);
and U14910 (N_14910,N_12385,N_12018);
and U14911 (N_14911,N_12918,N_12896);
or U14912 (N_14912,N_12607,N_12548);
nor U14913 (N_14913,N_12575,N_12235);
xor U14914 (N_14914,N_13826,N_13137);
nand U14915 (N_14915,N_13232,N_12523);
nor U14916 (N_14916,N_13390,N_13672);
or U14917 (N_14917,N_12023,N_13823);
nand U14918 (N_14918,N_12152,N_12343);
xnor U14919 (N_14919,N_12193,N_12472);
nand U14920 (N_14920,N_13263,N_12453);
nor U14921 (N_14921,N_13555,N_13558);
nand U14922 (N_14922,N_12389,N_12335);
nor U14923 (N_14923,N_13785,N_13765);
and U14924 (N_14924,N_12345,N_12877);
nand U14925 (N_14925,N_12251,N_12697);
or U14926 (N_14926,N_12664,N_12220);
or U14927 (N_14927,N_13688,N_12774);
nor U14928 (N_14928,N_13034,N_12045);
or U14929 (N_14929,N_13796,N_12320);
or U14930 (N_14930,N_12153,N_13897);
nand U14931 (N_14931,N_13003,N_12363);
nand U14932 (N_14932,N_12195,N_12448);
nand U14933 (N_14933,N_13632,N_13422);
and U14934 (N_14934,N_12287,N_12292);
xnor U14935 (N_14935,N_12261,N_13809);
xnor U14936 (N_14936,N_13457,N_13722);
xnor U14937 (N_14937,N_12779,N_13057);
nand U14938 (N_14938,N_12705,N_12366);
nor U14939 (N_14939,N_13896,N_12421);
nand U14940 (N_14940,N_12392,N_13649);
xnor U14941 (N_14941,N_13776,N_13201);
and U14942 (N_14942,N_13094,N_12521);
nand U14943 (N_14943,N_13488,N_13618);
nor U14944 (N_14944,N_12980,N_12776);
xor U14945 (N_14945,N_12270,N_13239);
and U14946 (N_14946,N_13568,N_12806);
nand U14947 (N_14947,N_12798,N_13389);
nor U14948 (N_14948,N_12637,N_13058);
nor U14949 (N_14949,N_12067,N_13939);
nand U14950 (N_14950,N_12605,N_12853);
xor U14951 (N_14951,N_12419,N_12942);
nand U14952 (N_14952,N_13762,N_12672);
nand U14953 (N_14953,N_13874,N_12568);
nor U14954 (N_14954,N_13681,N_13059);
or U14955 (N_14955,N_13187,N_12556);
nor U14956 (N_14956,N_13509,N_12584);
and U14957 (N_14957,N_13078,N_12242);
xor U14958 (N_14958,N_12783,N_13066);
and U14959 (N_14959,N_12805,N_13572);
nand U14960 (N_14960,N_12549,N_12773);
nor U14961 (N_14961,N_13439,N_12630);
xnor U14962 (N_14962,N_13150,N_13970);
or U14963 (N_14963,N_13191,N_13665);
or U14964 (N_14964,N_13086,N_13808);
nor U14965 (N_14965,N_12525,N_13768);
or U14966 (N_14966,N_12064,N_12003);
xor U14967 (N_14967,N_13627,N_12643);
and U14968 (N_14968,N_13963,N_13228);
and U14969 (N_14969,N_12224,N_12527);
xor U14970 (N_14970,N_12795,N_12088);
nor U14971 (N_14971,N_12395,N_12826);
xor U14972 (N_14972,N_12110,N_12996);
or U14973 (N_14973,N_12781,N_13622);
nand U14974 (N_14974,N_12720,N_13079);
nor U14975 (N_14975,N_13862,N_12827);
nor U14976 (N_14976,N_12665,N_12589);
nor U14977 (N_14977,N_12738,N_12030);
nand U14978 (N_14978,N_12869,N_12557);
nand U14979 (N_14979,N_12963,N_12537);
nand U14980 (N_14980,N_13292,N_12832);
nand U14981 (N_14981,N_13806,N_12741);
xor U14982 (N_14982,N_12560,N_12188);
or U14983 (N_14983,N_13271,N_12628);
nand U14984 (N_14984,N_12268,N_12218);
or U14985 (N_14985,N_13844,N_13361);
nand U14986 (N_14986,N_13974,N_13152);
nor U14987 (N_14987,N_12719,N_12604);
and U14988 (N_14988,N_13611,N_13772);
and U14989 (N_14989,N_12566,N_13487);
or U14990 (N_14990,N_13165,N_12625);
or U14991 (N_14991,N_12168,N_12046);
and U14992 (N_14992,N_13277,N_13976);
and U14993 (N_14993,N_13175,N_13464);
and U14994 (N_14994,N_13857,N_13668);
xnor U14995 (N_14995,N_13314,N_12471);
nor U14996 (N_14996,N_13637,N_12606);
or U14997 (N_14997,N_12875,N_12622);
nor U14998 (N_14998,N_13327,N_12880);
nor U14999 (N_14999,N_13548,N_13838);
and U15000 (N_15000,N_13249,N_13622);
or U15001 (N_15001,N_12200,N_12095);
xor U15002 (N_15002,N_13531,N_12858);
or U15003 (N_15003,N_12584,N_13504);
nand U15004 (N_15004,N_13106,N_13167);
or U15005 (N_15005,N_13381,N_12131);
nor U15006 (N_15006,N_13748,N_12208);
and U15007 (N_15007,N_13266,N_13414);
and U15008 (N_15008,N_12866,N_13722);
and U15009 (N_15009,N_13971,N_13411);
nand U15010 (N_15010,N_13959,N_12224);
and U15011 (N_15011,N_13790,N_13468);
nand U15012 (N_15012,N_12169,N_12373);
nor U15013 (N_15013,N_12378,N_13772);
and U15014 (N_15014,N_13756,N_12761);
xor U15015 (N_15015,N_12945,N_13171);
xnor U15016 (N_15016,N_12562,N_12949);
xor U15017 (N_15017,N_12794,N_13238);
xor U15018 (N_15018,N_13852,N_12836);
nor U15019 (N_15019,N_13221,N_12215);
nand U15020 (N_15020,N_13742,N_12813);
xor U15021 (N_15021,N_13178,N_13787);
xor U15022 (N_15022,N_13634,N_12811);
nand U15023 (N_15023,N_12874,N_12773);
and U15024 (N_15024,N_12537,N_13772);
or U15025 (N_15025,N_13154,N_12109);
or U15026 (N_15026,N_12712,N_12458);
nor U15027 (N_15027,N_13778,N_13954);
nor U15028 (N_15028,N_13693,N_12358);
and U15029 (N_15029,N_13463,N_12360);
xor U15030 (N_15030,N_13093,N_12889);
xor U15031 (N_15031,N_13583,N_12533);
and U15032 (N_15032,N_12506,N_13751);
nand U15033 (N_15033,N_13756,N_12731);
and U15034 (N_15034,N_12245,N_13965);
or U15035 (N_15035,N_13099,N_13818);
and U15036 (N_15036,N_13218,N_12907);
and U15037 (N_15037,N_13703,N_13423);
nor U15038 (N_15038,N_13999,N_12752);
or U15039 (N_15039,N_13289,N_12702);
xnor U15040 (N_15040,N_13260,N_13651);
or U15041 (N_15041,N_13018,N_13005);
or U15042 (N_15042,N_12956,N_12218);
or U15043 (N_15043,N_12315,N_12633);
nand U15044 (N_15044,N_13207,N_13846);
nand U15045 (N_15045,N_13050,N_13446);
nor U15046 (N_15046,N_12181,N_12945);
or U15047 (N_15047,N_12792,N_12166);
and U15048 (N_15048,N_12722,N_13066);
nand U15049 (N_15049,N_12903,N_13257);
and U15050 (N_15050,N_13560,N_12746);
nor U15051 (N_15051,N_13635,N_13421);
or U15052 (N_15052,N_13646,N_12437);
nor U15053 (N_15053,N_13889,N_12428);
nand U15054 (N_15054,N_13928,N_12838);
xor U15055 (N_15055,N_12786,N_12830);
nand U15056 (N_15056,N_13412,N_12205);
or U15057 (N_15057,N_12697,N_13911);
xnor U15058 (N_15058,N_12483,N_12743);
nand U15059 (N_15059,N_13229,N_13461);
and U15060 (N_15060,N_13754,N_13537);
xnor U15061 (N_15061,N_12203,N_13760);
nand U15062 (N_15062,N_12181,N_12097);
nand U15063 (N_15063,N_12773,N_13258);
xor U15064 (N_15064,N_12430,N_13253);
and U15065 (N_15065,N_13188,N_12611);
nand U15066 (N_15066,N_13151,N_13964);
and U15067 (N_15067,N_13047,N_12122);
and U15068 (N_15068,N_13738,N_12620);
and U15069 (N_15069,N_12147,N_13246);
or U15070 (N_15070,N_12392,N_13498);
and U15071 (N_15071,N_12599,N_13024);
nor U15072 (N_15072,N_12229,N_12589);
nor U15073 (N_15073,N_12602,N_12525);
and U15074 (N_15074,N_12262,N_12373);
and U15075 (N_15075,N_13918,N_12908);
or U15076 (N_15076,N_12134,N_13840);
nor U15077 (N_15077,N_12099,N_12258);
xor U15078 (N_15078,N_12764,N_13037);
nand U15079 (N_15079,N_12647,N_13921);
and U15080 (N_15080,N_13316,N_13341);
xor U15081 (N_15081,N_12031,N_13627);
nor U15082 (N_15082,N_12591,N_12321);
xnor U15083 (N_15083,N_13632,N_12054);
or U15084 (N_15084,N_12543,N_13767);
and U15085 (N_15085,N_13540,N_12542);
xor U15086 (N_15086,N_12915,N_13013);
xnor U15087 (N_15087,N_13324,N_12734);
nor U15088 (N_15088,N_12200,N_13425);
nand U15089 (N_15089,N_13568,N_13796);
nor U15090 (N_15090,N_13983,N_13843);
nor U15091 (N_15091,N_12233,N_13800);
nor U15092 (N_15092,N_12134,N_13405);
and U15093 (N_15093,N_13770,N_13577);
nor U15094 (N_15094,N_13426,N_13620);
nand U15095 (N_15095,N_13463,N_12752);
nand U15096 (N_15096,N_12331,N_12804);
nand U15097 (N_15097,N_13801,N_13726);
and U15098 (N_15098,N_12585,N_12995);
and U15099 (N_15099,N_12698,N_12588);
nand U15100 (N_15100,N_12196,N_12479);
nand U15101 (N_15101,N_13202,N_13365);
and U15102 (N_15102,N_12613,N_13438);
nand U15103 (N_15103,N_13386,N_13688);
or U15104 (N_15104,N_13671,N_13262);
xnor U15105 (N_15105,N_12082,N_12355);
nor U15106 (N_15106,N_13770,N_13823);
nand U15107 (N_15107,N_12499,N_13071);
nor U15108 (N_15108,N_12064,N_12321);
nand U15109 (N_15109,N_13534,N_13373);
or U15110 (N_15110,N_12425,N_13008);
nor U15111 (N_15111,N_13667,N_13463);
or U15112 (N_15112,N_13520,N_12017);
and U15113 (N_15113,N_12125,N_12725);
nand U15114 (N_15114,N_13486,N_13541);
and U15115 (N_15115,N_13144,N_12604);
and U15116 (N_15116,N_13495,N_12381);
and U15117 (N_15117,N_13717,N_12859);
and U15118 (N_15118,N_12872,N_12202);
xor U15119 (N_15119,N_13381,N_13326);
nor U15120 (N_15120,N_12683,N_13231);
nand U15121 (N_15121,N_13132,N_13041);
xor U15122 (N_15122,N_13833,N_12569);
and U15123 (N_15123,N_12464,N_13714);
and U15124 (N_15124,N_12246,N_12558);
or U15125 (N_15125,N_13605,N_13763);
nor U15126 (N_15126,N_13452,N_13333);
nand U15127 (N_15127,N_12881,N_12870);
nand U15128 (N_15128,N_13266,N_13409);
xnor U15129 (N_15129,N_13158,N_13027);
xnor U15130 (N_15130,N_13029,N_13541);
and U15131 (N_15131,N_12804,N_13868);
nand U15132 (N_15132,N_13602,N_13997);
or U15133 (N_15133,N_13901,N_12160);
nand U15134 (N_15134,N_12422,N_13089);
or U15135 (N_15135,N_13032,N_12424);
nor U15136 (N_15136,N_13532,N_13353);
nor U15137 (N_15137,N_13813,N_13925);
xor U15138 (N_15138,N_13345,N_12817);
nor U15139 (N_15139,N_12553,N_12799);
xor U15140 (N_15140,N_13199,N_13800);
nand U15141 (N_15141,N_12106,N_12826);
nor U15142 (N_15142,N_13818,N_12919);
xor U15143 (N_15143,N_13841,N_13063);
or U15144 (N_15144,N_13965,N_12071);
nand U15145 (N_15145,N_13072,N_13899);
nand U15146 (N_15146,N_13899,N_13732);
and U15147 (N_15147,N_12277,N_12600);
nor U15148 (N_15148,N_13572,N_12803);
xnor U15149 (N_15149,N_13780,N_13672);
xor U15150 (N_15150,N_13448,N_13913);
xnor U15151 (N_15151,N_12316,N_12270);
and U15152 (N_15152,N_13853,N_12229);
and U15153 (N_15153,N_12176,N_12558);
xor U15154 (N_15154,N_12202,N_12722);
xnor U15155 (N_15155,N_13428,N_12087);
and U15156 (N_15156,N_12484,N_13258);
nand U15157 (N_15157,N_13312,N_12510);
xor U15158 (N_15158,N_13576,N_13287);
xnor U15159 (N_15159,N_12352,N_12357);
or U15160 (N_15160,N_13807,N_12464);
and U15161 (N_15161,N_12688,N_12681);
xnor U15162 (N_15162,N_13482,N_12138);
nor U15163 (N_15163,N_13475,N_12765);
nor U15164 (N_15164,N_12397,N_13098);
or U15165 (N_15165,N_13174,N_12844);
nor U15166 (N_15166,N_13881,N_12529);
and U15167 (N_15167,N_13887,N_13122);
nand U15168 (N_15168,N_12928,N_12600);
xor U15169 (N_15169,N_12882,N_13927);
nor U15170 (N_15170,N_12798,N_12837);
nor U15171 (N_15171,N_12076,N_12509);
or U15172 (N_15172,N_13061,N_12334);
nand U15173 (N_15173,N_13065,N_12708);
xor U15174 (N_15174,N_13750,N_12836);
and U15175 (N_15175,N_12611,N_12577);
or U15176 (N_15176,N_13398,N_12861);
or U15177 (N_15177,N_13876,N_12841);
and U15178 (N_15178,N_12651,N_12419);
nand U15179 (N_15179,N_12708,N_13644);
nor U15180 (N_15180,N_12375,N_13164);
xnor U15181 (N_15181,N_13026,N_13516);
or U15182 (N_15182,N_13158,N_13372);
nor U15183 (N_15183,N_12494,N_13905);
xnor U15184 (N_15184,N_12645,N_12456);
nor U15185 (N_15185,N_13905,N_12083);
xnor U15186 (N_15186,N_13159,N_12694);
and U15187 (N_15187,N_12027,N_13280);
and U15188 (N_15188,N_12480,N_12452);
nor U15189 (N_15189,N_12388,N_12412);
nand U15190 (N_15190,N_12430,N_13746);
nor U15191 (N_15191,N_12292,N_13216);
or U15192 (N_15192,N_13252,N_13966);
nand U15193 (N_15193,N_13682,N_13763);
or U15194 (N_15194,N_12736,N_12342);
and U15195 (N_15195,N_13296,N_12908);
nor U15196 (N_15196,N_12973,N_12889);
nand U15197 (N_15197,N_12212,N_13987);
xnor U15198 (N_15198,N_12954,N_13388);
nand U15199 (N_15199,N_13236,N_13197);
nor U15200 (N_15200,N_12515,N_12058);
nand U15201 (N_15201,N_13594,N_13371);
nor U15202 (N_15202,N_13098,N_12840);
or U15203 (N_15203,N_12248,N_13749);
xnor U15204 (N_15204,N_13029,N_13222);
xor U15205 (N_15205,N_13995,N_13497);
and U15206 (N_15206,N_13947,N_12741);
xnor U15207 (N_15207,N_12200,N_12520);
nor U15208 (N_15208,N_13819,N_12240);
and U15209 (N_15209,N_12972,N_12895);
or U15210 (N_15210,N_12321,N_13018);
nand U15211 (N_15211,N_12061,N_13537);
nand U15212 (N_15212,N_13871,N_13612);
nor U15213 (N_15213,N_13188,N_13713);
nor U15214 (N_15214,N_12468,N_12430);
or U15215 (N_15215,N_12552,N_13021);
or U15216 (N_15216,N_12566,N_12637);
or U15217 (N_15217,N_13257,N_12258);
and U15218 (N_15218,N_12824,N_13181);
or U15219 (N_15219,N_12949,N_12557);
or U15220 (N_15220,N_13482,N_12774);
or U15221 (N_15221,N_12070,N_12943);
xnor U15222 (N_15222,N_12843,N_12471);
nand U15223 (N_15223,N_13994,N_13205);
nor U15224 (N_15224,N_13979,N_12246);
xor U15225 (N_15225,N_13296,N_13880);
or U15226 (N_15226,N_12832,N_12175);
or U15227 (N_15227,N_12399,N_13015);
nor U15228 (N_15228,N_13570,N_13269);
xor U15229 (N_15229,N_13136,N_12450);
or U15230 (N_15230,N_12746,N_12679);
xor U15231 (N_15231,N_13341,N_12401);
nand U15232 (N_15232,N_13513,N_13524);
xnor U15233 (N_15233,N_13808,N_12074);
nor U15234 (N_15234,N_12279,N_13450);
xnor U15235 (N_15235,N_12390,N_12667);
or U15236 (N_15236,N_13588,N_13793);
xnor U15237 (N_15237,N_12421,N_13010);
nor U15238 (N_15238,N_13690,N_12217);
xor U15239 (N_15239,N_12967,N_12969);
xor U15240 (N_15240,N_13032,N_13092);
nand U15241 (N_15241,N_12505,N_12297);
nor U15242 (N_15242,N_13280,N_12723);
xnor U15243 (N_15243,N_12266,N_13140);
nor U15244 (N_15244,N_12321,N_13985);
or U15245 (N_15245,N_12921,N_13760);
or U15246 (N_15246,N_13248,N_12546);
nand U15247 (N_15247,N_13635,N_13409);
nand U15248 (N_15248,N_13627,N_13501);
xor U15249 (N_15249,N_13471,N_12712);
xnor U15250 (N_15250,N_12911,N_13617);
xor U15251 (N_15251,N_13062,N_12656);
or U15252 (N_15252,N_13150,N_12474);
or U15253 (N_15253,N_12072,N_13392);
and U15254 (N_15254,N_13053,N_12203);
nor U15255 (N_15255,N_13030,N_13073);
nand U15256 (N_15256,N_13904,N_13784);
and U15257 (N_15257,N_13835,N_12133);
nor U15258 (N_15258,N_12782,N_12218);
nand U15259 (N_15259,N_13427,N_12411);
xnor U15260 (N_15260,N_12124,N_13644);
nor U15261 (N_15261,N_13137,N_12882);
nand U15262 (N_15262,N_12640,N_13415);
and U15263 (N_15263,N_13878,N_13402);
and U15264 (N_15264,N_12258,N_13106);
nor U15265 (N_15265,N_12748,N_12546);
and U15266 (N_15266,N_12333,N_12492);
nor U15267 (N_15267,N_13558,N_12724);
xor U15268 (N_15268,N_12936,N_12760);
xnor U15269 (N_15269,N_12949,N_12539);
or U15270 (N_15270,N_13866,N_13376);
nor U15271 (N_15271,N_12261,N_12371);
and U15272 (N_15272,N_12862,N_13162);
nor U15273 (N_15273,N_12752,N_12030);
xor U15274 (N_15274,N_13879,N_12011);
or U15275 (N_15275,N_13917,N_12823);
nand U15276 (N_15276,N_12086,N_12287);
or U15277 (N_15277,N_12006,N_12628);
nand U15278 (N_15278,N_12831,N_12416);
xor U15279 (N_15279,N_12878,N_12330);
nor U15280 (N_15280,N_13310,N_12054);
and U15281 (N_15281,N_13730,N_12834);
xor U15282 (N_15282,N_12382,N_13623);
and U15283 (N_15283,N_13883,N_13944);
and U15284 (N_15284,N_13677,N_13102);
nor U15285 (N_15285,N_12459,N_13361);
or U15286 (N_15286,N_13098,N_12608);
and U15287 (N_15287,N_13730,N_13862);
nor U15288 (N_15288,N_13880,N_13017);
nor U15289 (N_15289,N_12505,N_12894);
or U15290 (N_15290,N_12569,N_12576);
nand U15291 (N_15291,N_12822,N_13883);
nor U15292 (N_15292,N_13866,N_12075);
and U15293 (N_15293,N_12656,N_13337);
or U15294 (N_15294,N_13698,N_13951);
or U15295 (N_15295,N_12155,N_12166);
xnor U15296 (N_15296,N_13006,N_12839);
nor U15297 (N_15297,N_12932,N_13969);
and U15298 (N_15298,N_12892,N_13461);
nand U15299 (N_15299,N_12410,N_12211);
and U15300 (N_15300,N_13994,N_13819);
nor U15301 (N_15301,N_13203,N_13359);
or U15302 (N_15302,N_12049,N_12222);
and U15303 (N_15303,N_13592,N_12963);
nor U15304 (N_15304,N_13502,N_12257);
nor U15305 (N_15305,N_12544,N_13679);
nand U15306 (N_15306,N_13896,N_12624);
and U15307 (N_15307,N_13194,N_13590);
xor U15308 (N_15308,N_13965,N_13763);
nand U15309 (N_15309,N_12881,N_13260);
nand U15310 (N_15310,N_12084,N_12628);
nand U15311 (N_15311,N_13089,N_12531);
xnor U15312 (N_15312,N_12462,N_13193);
xnor U15313 (N_15313,N_12541,N_12900);
nor U15314 (N_15314,N_13192,N_12878);
or U15315 (N_15315,N_13650,N_12091);
or U15316 (N_15316,N_13180,N_12776);
and U15317 (N_15317,N_12959,N_13834);
nand U15318 (N_15318,N_13978,N_12161);
nor U15319 (N_15319,N_13116,N_13009);
nand U15320 (N_15320,N_12353,N_13476);
nand U15321 (N_15321,N_12216,N_12312);
and U15322 (N_15322,N_12127,N_13867);
and U15323 (N_15323,N_13946,N_13345);
nor U15324 (N_15324,N_13723,N_13782);
nor U15325 (N_15325,N_13898,N_13643);
nand U15326 (N_15326,N_13390,N_13739);
and U15327 (N_15327,N_12193,N_12915);
and U15328 (N_15328,N_12867,N_12686);
nor U15329 (N_15329,N_12339,N_12085);
nor U15330 (N_15330,N_12378,N_12071);
nand U15331 (N_15331,N_12917,N_13515);
and U15332 (N_15332,N_12292,N_12886);
or U15333 (N_15333,N_13152,N_12409);
or U15334 (N_15334,N_12923,N_12627);
xor U15335 (N_15335,N_12991,N_13903);
or U15336 (N_15336,N_12184,N_12674);
nor U15337 (N_15337,N_13951,N_13535);
nand U15338 (N_15338,N_13730,N_13937);
xnor U15339 (N_15339,N_13743,N_12878);
or U15340 (N_15340,N_13278,N_13529);
nor U15341 (N_15341,N_13204,N_13233);
nand U15342 (N_15342,N_12311,N_13374);
and U15343 (N_15343,N_13057,N_12490);
nand U15344 (N_15344,N_13048,N_13871);
nand U15345 (N_15345,N_13350,N_13112);
nand U15346 (N_15346,N_13004,N_12932);
nand U15347 (N_15347,N_12081,N_12041);
xnor U15348 (N_15348,N_12011,N_13371);
and U15349 (N_15349,N_13433,N_13867);
and U15350 (N_15350,N_13421,N_12287);
xnor U15351 (N_15351,N_13381,N_13720);
or U15352 (N_15352,N_13276,N_12787);
nand U15353 (N_15353,N_13952,N_12471);
nor U15354 (N_15354,N_12557,N_12560);
xor U15355 (N_15355,N_12066,N_12207);
nand U15356 (N_15356,N_13967,N_12557);
or U15357 (N_15357,N_12252,N_13603);
nor U15358 (N_15358,N_13395,N_13459);
xnor U15359 (N_15359,N_13689,N_12079);
nor U15360 (N_15360,N_13229,N_12269);
xnor U15361 (N_15361,N_12940,N_13993);
or U15362 (N_15362,N_13023,N_13968);
xor U15363 (N_15363,N_13149,N_13209);
or U15364 (N_15364,N_12861,N_13029);
nand U15365 (N_15365,N_12023,N_12619);
and U15366 (N_15366,N_12311,N_12912);
nor U15367 (N_15367,N_13691,N_13970);
nor U15368 (N_15368,N_12760,N_13080);
or U15369 (N_15369,N_12867,N_13743);
or U15370 (N_15370,N_12449,N_13583);
nand U15371 (N_15371,N_12397,N_13064);
nand U15372 (N_15372,N_12870,N_13529);
and U15373 (N_15373,N_13416,N_13955);
nand U15374 (N_15374,N_13641,N_13258);
and U15375 (N_15375,N_12562,N_12644);
xor U15376 (N_15376,N_13900,N_13954);
nor U15377 (N_15377,N_12900,N_12668);
or U15378 (N_15378,N_12707,N_13035);
or U15379 (N_15379,N_12173,N_13898);
nand U15380 (N_15380,N_13034,N_13172);
or U15381 (N_15381,N_12455,N_13851);
nand U15382 (N_15382,N_12472,N_12349);
and U15383 (N_15383,N_12039,N_13257);
or U15384 (N_15384,N_12614,N_12046);
xnor U15385 (N_15385,N_13747,N_13195);
or U15386 (N_15386,N_12347,N_12874);
xor U15387 (N_15387,N_12645,N_13084);
nor U15388 (N_15388,N_13522,N_13343);
xor U15389 (N_15389,N_13917,N_13973);
or U15390 (N_15390,N_12516,N_12028);
or U15391 (N_15391,N_13563,N_13109);
and U15392 (N_15392,N_13600,N_12269);
nor U15393 (N_15393,N_13869,N_13534);
nor U15394 (N_15394,N_12984,N_12974);
nor U15395 (N_15395,N_13073,N_12883);
nand U15396 (N_15396,N_12632,N_12669);
or U15397 (N_15397,N_13535,N_12298);
nor U15398 (N_15398,N_13869,N_13703);
xor U15399 (N_15399,N_12070,N_12693);
or U15400 (N_15400,N_13012,N_12299);
or U15401 (N_15401,N_13011,N_12583);
xor U15402 (N_15402,N_12075,N_12077);
nand U15403 (N_15403,N_12934,N_12160);
nor U15404 (N_15404,N_13703,N_12059);
or U15405 (N_15405,N_12890,N_13989);
xnor U15406 (N_15406,N_12691,N_13388);
and U15407 (N_15407,N_12699,N_12553);
or U15408 (N_15408,N_12008,N_12081);
nand U15409 (N_15409,N_13438,N_13876);
nand U15410 (N_15410,N_12763,N_12870);
and U15411 (N_15411,N_12495,N_13056);
nand U15412 (N_15412,N_13189,N_13167);
nor U15413 (N_15413,N_12683,N_12225);
xnor U15414 (N_15414,N_13154,N_13451);
and U15415 (N_15415,N_12790,N_12158);
nand U15416 (N_15416,N_12327,N_12927);
and U15417 (N_15417,N_12197,N_12413);
or U15418 (N_15418,N_12418,N_13721);
nor U15419 (N_15419,N_12654,N_13983);
xor U15420 (N_15420,N_12300,N_13445);
or U15421 (N_15421,N_12667,N_12232);
xnor U15422 (N_15422,N_13909,N_13059);
nand U15423 (N_15423,N_13141,N_12950);
xor U15424 (N_15424,N_13086,N_12898);
and U15425 (N_15425,N_12747,N_13795);
and U15426 (N_15426,N_12518,N_12030);
xor U15427 (N_15427,N_12334,N_13834);
or U15428 (N_15428,N_12456,N_13742);
nand U15429 (N_15429,N_12855,N_12597);
nand U15430 (N_15430,N_12548,N_12340);
nand U15431 (N_15431,N_13209,N_12739);
or U15432 (N_15432,N_13267,N_12510);
nand U15433 (N_15433,N_13454,N_13366);
or U15434 (N_15434,N_13202,N_12043);
and U15435 (N_15435,N_13263,N_13429);
or U15436 (N_15436,N_12255,N_12273);
xnor U15437 (N_15437,N_13517,N_12495);
and U15438 (N_15438,N_12221,N_12332);
nor U15439 (N_15439,N_12043,N_13817);
or U15440 (N_15440,N_13190,N_13287);
nor U15441 (N_15441,N_13593,N_12352);
xnor U15442 (N_15442,N_12759,N_13593);
nor U15443 (N_15443,N_12872,N_13990);
nor U15444 (N_15444,N_13435,N_13867);
or U15445 (N_15445,N_12078,N_12772);
nor U15446 (N_15446,N_12466,N_12442);
or U15447 (N_15447,N_13168,N_12848);
xor U15448 (N_15448,N_13097,N_13142);
nor U15449 (N_15449,N_12531,N_12460);
xnor U15450 (N_15450,N_13883,N_12835);
or U15451 (N_15451,N_12639,N_13697);
or U15452 (N_15452,N_12806,N_13682);
and U15453 (N_15453,N_12026,N_12867);
nand U15454 (N_15454,N_12079,N_12322);
or U15455 (N_15455,N_13970,N_13945);
nor U15456 (N_15456,N_12258,N_12973);
xnor U15457 (N_15457,N_13920,N_12549);
xor U15458 (N_15458,N_13714,N_13785);
nor U15459 (N_15459,N_12354,N_12144);
and U15460 (N_15460,N_13486,N_13156);
xnor U15461 (N_15461,N_12170,N_12475);
and U15462 (N_15462,N_13300,N_12361);
nor U15463 (N_15463,N_12231,N_13274);
nand U15464 (N_15464,N_12829,N_13772);
or U15465 (N_15465,N_12425,N_12397);
nand U15466 (N_15466,N_12419,N_13183);
nor U15467 (N_15467,N_13412,N_13543);
and U15468 (N_15468,N_13084,N_12037);
xnor U15469 (N_15469,N_12012,N_12473);
nor U15470 (N_15470,N_13763,N_12214);
and U15471 (N_15471,N_12005,N_13154);
xnor U15472 (N_15472,N_12062,N_13364);
nand U15473 (N_15473,N_12990,N_13129);
or U15474 (N_15474,N_13543,N_12718);
nand U15475 (N_15475,N_13381,N_13798);
or U15476 (N_15476,N_12654,N_12522);
nand U15477 (N_15477,N_13246,N_12106);
and U15478 (N_15478,N_12182,N_13913);
and U15479 (N_15479,N_12619,N_12860);
nand U15480 (N_15480,N_12859,N_13704);
nand U15481 (N_15481,N_12400,N_12087);
nand U15482 (N_15482,N_12101,N_12701);
xor U15483 (N_15483,N_12907,N_12736);
nor U15484 (N_15484,N_13266,N_13767);
and U15485 (N_15485,N_13456,N_13676);
nand U15486 (N_15486,N_13439,N_12441);
nand U15487 (N_15487,N_12099,N_12884);
xnor U15488 (N_15488,N_12981,N_12323);
xor U15489 (N_15489,N_12427,N_12175);
and U15490 (N_15490,N_12716,N_13531);
or U15491 (N_15491,N_12194,N_12852);
nand U15492 (N_15492,N_12269,N_13658);
and U15493 (N_15493,N_13637,N_12272);
and U15494 (N_15494,N_13659,N_13349);
or U15495 (N_15495,N_13561,N_13391);
or U15496 (N_15496,N_12504,N_12110);
nor U15497 (N_15497,N_12766,N_13007);
nor U15498 (N_15498,N_12092,N_13293);
nor U15499 (N_15499,N_13453,N_12354);
and U15500 (N_15500,N_13849,N_13095);
nand U15501 (N_15501,N_13014,N_13450);
nand U15502 (N_15502,N_12483,N_13191);
or U15503 (N_15503,N_12401,N_12670);
nor U15504 (N_15504,N_13053,N_12724);
nand U15505 (N_15505,N_13205,N_12626);
and U15506 (N_15506,N_13572,N_13554);
nand U15507 (N_15507,N_12460,N_12820);
xor U15508 (N_15508,N_12959,N_13840);
xor U15509 (N_15509,N_13024,N_12803);
xnor U15510 (N_15510,N_13725,N_12092);
xor U15511 (N_15511,N_12694,N_13919);
or U15512 (N_15512,N_13822,N_13065);
or U15513 (N_15513,N_12804,N_12702);
and U15514 (N_15514,N_12756,N_13357);
nand U15515 (N_15515,N_12079,N_12885);
xor U15516 (N_15516,N_13853,N_12760);
nand U15517 (N_15517,N_13348,N_13255);
or U15518 (N_15518,N_13757,N_13349);
and U15519 (N_15519,N_12945,N_13091);
and U15520 (N_15520,N_13823,N_13327);
nand U15521 (N_15521,N_13703,N_12359);
xnor U15522 (N_15522,N_13451,N_13044);
nor U15523 (N_15523,N_12894,N_12488);
nor U15524 (N_15524,N_12917,N_12916);
nand U15525 (N_15525,N_12008,N_13555);
or U15526 (N_15526,N_13800,N_13234);
xnor U15527 (N_15527,N_13750,N_12561);
and U15528 (N_15528,N_13537,N_13576);
xnor U15529 (N_15529,N_13191,N_13433);
nor U15530 (N_15530,N_12043,N_12253);
or U15531 (N_15531,N_13638,N_12392);
and U15532 (N_15532,N_12789,N_12244);
or U15533 (N_15533,N_12124,N_13489);
or U15534 (N_15534,N_12968,N_12714);
or U15535 (N_15535,N_13390,N_12805);
nand U15536 (N_15536,N_13247,N_12271);
nor U15537 (N_15537,N_13967,N_12985);
or U15538 (N_15538,N_13621,N_13524);
and U15539 (N_15539,N_13595,N_13105);
nand U15540 (N_15540,N_12562,N_13776);
nor U15541 (N_15541,N_13577,N_13781);
xor U15542 (N_15542,N_13454,N_13737);
xnor U15543 (N_15543,N_13392,N_13092);
and U15544 (N_15544,N_12496,N_13973);
nand U15545 (N_15545,N_13125,N_12781);
and U15546 (N_15546,N_13817,N_13031);
nand U15547 (N_15547,N_13695,N_13266);
or U15548 (N_15548,N_13683,N_13639);
and U15549 (N_15549,N_13016,N_12557);
xnor U15550 (N_15550,N_13702,N_13979);
xnor U15551 (N_15551,N_12070,N_12833);
nor U15552 (N_15552,N_13259,N_12754);
or U15553 (N_15553,N_12805,N_13755);
and U15554 (N_15554,N_13021,N_12827);
and U15555 (N_15555,N_12893,N_13489);
xnor U15556 (N_15556,N_12349,N_12057);
nor U15557 (N_15557,N_12612,N_13667);
nor U15558 (N_15558,N_13823,N_13982);
and U15559 (N_15559,N_12326,N_12210);
and U15560 (N_15560,N_12585,N_12947);
nand U15561 (N_15561,N_13652,N_12743);
xnor U15562 (N_15562,N_13173,N_12624);
or U15563 (N_15563,N_12272,N_12515);
nand U15564 (N_15564,N_13742,N_12672);
or U15565 (N_15565,N_12114,N_13236);
or U15566 (N_15566,N_12112,N_12021);
or U15567 (N_15567,N_13567,N_12187);
nor U15568 (N_15568,N_13776,N_13930);
or U15569 (N_15569,N_12475,N_12855);
nor U15570 (N_15570,N_12725,N_12326);
nand U15571 (N_15571,N_13966,N_12217);
and U15572 (N_15572,N_12946,N_12081);
and U15573 (N_15573,N_13376,N_12740);
and U15574 (N_15574,N_12487,N_13346);
and U15575 (N_15575,N_13797,N_13281);
xor U15576 (N_15576,N_13269,N_12311);
nand U15577 (N_15577,N_12115,N_12554);
nand U15578 (N_15578,N_13610,N_12137);
nand U15579 (N_15579,N_12598,N_12105);
and U15580 (N_15580,N_13081,N_12535);
or U15581 (N_15581,N_12543,N_12472);
nor U15582 (N_15582,N_12977,N_12546);
nor U15583 (N_15583,N_13085,N_12337);
nor U15584 (N_15584,N_13021,N_12177);
or U15585 (N_15585,N_12169,N_13611);
nand U15586 (N_15586,N_13841,N_13011);
and U15587 (N_15587,N_13554,N_13635);
xnor U15588 (N_15588,N_13255,N_12177);
xor U15589 (N_15589,N_12235,N_12813);
and U15590 (N_15590,N_12977,N_13498);
nor U15591 (N_15591,N_13823,N_13909);
or U15592 (N_15592,N_13866,N_12169);
or U15593 (N_15593,N_12185,N_12054);
or U15594 (N_15594,N_13852,N_12645);
nor U15595 (N_15595,N_12863,N_13687);
nor U15596 (N_15596,N_13563,N_12352);
or U15597 (N_15597,N_13499,N_12282);
xnor U15598 (N_15598,N_13863,N_12667);
xor U15599 (N_15599,N_13483,N_12978);
or U15600 (N_15600,N_12390,N_13599);
xor U15601 (N_15601,N_13430,N_13206);
xor U15602 (N_15602,N_13941,N_12403);
or U15603 (N_15603,N_13087,N_12708);
nor U15604 (N_15604,N_13466,N_12090);
and U15605 (N_15605,N_13943,N_12166);
and U15606 (N_15606,N_13810,N_13470);
and U15607 (N_15607,N_13755,N_12628);
xnor U15608 (N_15608,N_12071,N_12627);
nor U15609 (N_15609,N_13766,N_13725);
nand U15610 (N_15610,N_13564,N_12269);
and U15611 (N_15611,N_12590,N_13071);
nand U15612 (N_15612,N_13612,N_13691);
nor U15613 (N_15613,N_13192,N_12518);
and U15614 (N_15614,N_12232,N_13968);
nand U15615 (N_15615,N_12268,N_12032);
or U15616 (N_15616,N_13116,N_13900);
xor U15617 (N_15617,N_13903,N_13406);
and U15618 (N_15618,N_12646,N_12491);
nor U15619 (N_15619,N_13753,N_13327);
nor U15620 (N_15620,N_12356,N_13234);
nor U15621 (N_15621,N_12292,N_13568);
or U15622 (N_15622,N_12198,N_13300);
nor U15623 (N_15623,N_13800,N_13701);
or U15624 (N_15624,N_12918,N_13576);
xnor U15625 (N_15625,N_12841,N_12032);
and U15626 (N_15626,N_13393,N_13642);
nor U15627 (N_15627,N_12635,N_13357);
nor U15628 (N_15628,N_12349,N_13591);
and U15629 (N_15629,N_12505,N_13082);
nand U15630 (N_15630,N_12371,N_13047);
and U15631 (N_15631,N_12633,N_12661);
nand U15632 (N_15632,N_12887,N_12858);
nand U15633 (N_15633,N_13239,N_12707);
xor U15634 (N_15634,N_13153,N_13443);
or U15635 (N_15635,N_13438,N_13305);
or U15636 (N_15636,N_13788,N_12956);
nand U15637 (N_15637,N_12755,N_12345);
xor U15638 (N_15638,N_13417,N_12326);
or U15639 (N_15639,N_13822,N_13882);
nand U15640 (N_15640,N_13529,N_12058);
nand U15641 (N_15641,N_12226,N_13424);
or U15642 (N_15642,N_13584,N_12324);
xnor U15643 (N_15643,N_13085,N_12473);
nor U15644 (N_15644,N_12049,N_13462);
nand U15645 (N_15645,N_13569,N_13566);
nor U15646 (N_15646,N_12483,N_13998);
nor U15647 (N_15647,N_12633,N_12230);
nand U15648 (N_15648,N_13764,N_13356);
and U15649 (N_15649,N_12109,N_13522);
nand U15650 (N_15650,N_12950,N_13891);
and U15651 (N_15651,N_13699,N_12588);
xnor U15652 (N_15652,N_13390,N_12955);
nand U15653 (N_15653,N_12991,N_13790);
nor U15654 (N_15654,N_13413,N_12484);
or U15655 (N_15655,N_12717,N_13829);
and U15656 (N_15656,N_12290,N_13510);
nor U15657 (N_15657,N_13131,N_12506);
xnor U15658 (N_15658,N_13026,N_13711);
xor U15659 (N_15659,N_13367,N_12273);
nand U15660 (N_15660,N_12060,N_13576);
and U15661 (N_15661,N_13195,N_13464);
xor U15662 (N_15662,N_12079,N_13766);
nor U15663 (N_15663,N_13948,N_13117);
nand U15664 (N_15664,N_13397,N_13164);
nor U15665 (N_15665,N_13317,N_12670);
nor U15666 (N_15666,N_12033,N_13065);
xnor U15667 (N_15667,N_12798,N_13798);
or U15668 (N_15668,N_12915,N_13885);
xnor U15669 (N_15669,N_12770,N_12531);
and U15670 (N_15670,N_13102,N_12594);
nand U15671 (N_15671,N_12056,N_12283);
nand U15672 (N_15672,N_13147,N_12656);
nor U15673 (N_15673,N_13310,N_13080);
and U15674 (N_15674,N_12967,N_13197);
nor U15675 (N_15675,N_13466,N_12449);
nor U15676 (N_15676,N_13379,N_12854);
or U15677 (N_15677,N_12145,N_12536);
nor U15678 (N_15678,N_12785,N_12990);
and U15679 (N_15679,N_12754,N_13264);
xor U15680 (N_15680,N_12202,N_12754);
and U15681 (N_15681,N_13448,N_12591);
or U15682 (N_15682,N_13529,N_12574);
nor U15683 (N_15683,N_12308,N_12829);
nand U15684 (N_15684,N_13799,N_13924);
nand U15685 (N_15685,N_13894,N_13886);
nor U15686 (N_15686,N_13812,N_12744);
nand U15687 (N_15687,N_13410,N_13826);
or U15688 (N_15688,N_12594,N_13021);
nor U15689 (N_15689,N_12641,N_13689);
nor U15690 (N_15690,N_13813,N_12347);
xnor U15691 (N_15691,N_12196,N_13192);
nand U15692 (N_15692,N_12818,N_13983);
or U15693 (N_15693,N_12105,N_13254);
or U15694 (N_15694,N_13466,N_12648);
nand U15695 (N_15695,N_12007,N_12705);
xor U15696 (N_15696,N_12758,N_12349);
nand U15697 (N_15697,N_12538,N_12976);
nand U15698 (N_15698,N_12737,N_13651);
nand U15699 (N_15699,N_13859,N_13599);
xor U15700 (N_15700,N_13789,N_13772);
nor U15701 (N_15701,N_13643,N_12635);
and U15702 (N_15702,N_13576,N_12205);
nor U15703 (N_15703,N_13197,N_13338);
xnor U15704 (N_15704,N_12935,N_12642);
and U15705 (N_15705,N_13863,N_12206);
or U15706 (N_15706,N_12951,N_12677);
nor U15707 (N_15707,N_12612,N_12534);
or U15708 (N_15708,N_12889,N_13418);
nand U15709 (N_15709,N_13045,N_12912);
xor U15710 (N_15710,N_13733,N_13013);
nand U15711 (N_15711,N_13135,N_12908);
xor U15712 (N_15712,N_12497,N_13366);
xnor U15713 (N_15713,N_13829,N_12775);
nand U15714 (N_15714,N_12928,N_12560);
or U15715 (N_15715,N_12041,N_12589);
nor U15716 (N_15716,N_13350,N_13633);
nor U15717 (N_15717,N_12745,N_13726);
xor U15718 (N_15718,N_12240,N_12656);
xnor U15719 (N_15719,N_13158,N_13507);
nand U15720 (N_15720,N_13936,N_12702);
nand U15721 (N_15721,N_13715,N_13614);
xnor U15722 (N_15722,N_12890,N_12102);
or U15723 (N_15723,N_12462,N_13081);
and U15724 (N_15724,N_12906,N_12460);
xnor U15725 (N_15725,N_12221,N_12416);
xnor U15726 (N_15726,N_12336,N_12961);
and U15727 (N_15727,N_13796,N_12008);
nand U15728 (N_15728,N_13645,N_13634);
nand U15729 (N_15729,N_12796,N_13554);
and U15730 (N_15730,N_12706,N_12971);
or U15731 (N_15731,N_13120,N_12154);
nor U15732 (N_15732,N_12087,N_12097);
nand U15733 (N_15733,N_13972,N_12817);
and U15734 (N_15734,N_13201,N_13954);
nor U15735 (N_15735,N_13858,N_12178);
or U15736 (N_15736,N_13662,N_12455);
xnor U15737 (N_15737,N_12733,N_12177);
or U15738 (N_15738,N_13163,N_12118);
and U15739 (N_15739,N_12998,N_12350);
nand U15740 (N_15740,N_12468,N_12470);
and U15741 (N_15741,N_12384,N_13135);
nand U15742 (N_15742,N_13989,N_12880);
xor U15743 (N_15743,N_12058,N_13387);
xor U15744 (N_15744,N_13312,N_12308);
nor U15745 (N_15745,N_12253,N_12113);
and U15746 (N_15746,N_12053,N_12684);
or U15747 (N_15747,N_13808,N_12472);
xnor U15748 (N_15748,N_13024,N_13397);
nand U15749 (N_15749,N_13041,N_12392);
nor U15750 (N_15750,N_13030,N_13992);
nand U15751 (N_15751,N_13953,N_13976);
xnor U15752 (N_15752,N_13928,N_12833);
or U15753 (N_15753,N_12383,N_13342);
nand U15754 (N_15754,N_12123,N_12940);
or U15755 (N_15755,N_13484,N_12880);
nand U15756 (N_15756,N_12279,N_13540);
or U15757 (N_15757,N_13723,N_13792);
nor U15758 (N_15758,N_12322,N_12999);
nand U15759 (N_15759,N_12703,N_13915);
or U15760 (N_15760,N_12817,N_12813);
or U15761 (N_15761,N_13349,N_13918);
or U15762 (N_15762,N_13273,N_13135);
nor U15763 (N_15763,N_12356,N_12504);
nor U15764 (N_15764,N_12461,N_12152);
or U15765 (N_15765,N_13944,N_12923);
nor U15766 (N_15766,N_13163,N_13539);
and U15767 (N_15767,N_12285,N_13659);
nand U15768 (N_15768,N_13023,N_13622);
xor U15769 (N_15769,N_12759,N_12064);
and U15770 (N_15770,N_13995,N_12487);
xnor U15771 (N_15771,N_13532,N_13516);
nand U15772 (N_15772,N_13729,N_13672);
and U15773 (N_15773,N_12635,N_12038);
xor U15774 (N_15774,N_12512,N_13157);
nand U15775 (N_15775,N_13623,N_12308);
and U15776 (N_15776,N_12320,N_13138);
xor U15777 (N_15777,N_12980,N_13405);
and U15778 (N_15778,N_13223,N_13660);
xor U15779 (N_15779,N_12258,N_12800);
and U15780 (N_15780,N_13583,N_13308);
nor U15781 (N_15781,N_13264,N_12035);
nor U15782 (N_15782,N_13142,N_12779);
nor U15783 (N_15783,N_12422,N_13100);
or U15784 (N_15784,N_12916,N_13123);
nor U15785 (N_15785,N_13101,N_12074);
nand U15786 (N_15786,N_13105,N_13508);
nor U15787 (N_15787,N_12359,N_12493);
and U15788 (N_15788,N_12133,N_12572);
and U15789 (N_15789,N_12850,N_12603);
nand U15790 (N_15790,N_13074,N_12019);
and U15791 (N_15791,N_12358,N_12525);
nand U15792 (N_15792,N_12144,N_13784);
and U15793 (N_15793,N_13016,N_12996);
nor U15794 (N_15794,N_12273,N_13546);
nand U15795 (N_15795,N_13667,N_12486);
nor U15796 (N_15796,N_13474,N_12754);
nand U15797 (N_15797,N_13524,N_12389);
nor U15798 (N_15798,N_13643,N_12238);
xnor U15799 (N_15799,N_13652,N_13981);
and U15800 (N_15800,N_13921,N_12908);
or U15801 (N_15801,N_13804,N_12585);
xor U15802 (N_15802,N_12332,N_13929);
nand U15803 (N_15803,N_13738,N_13197);
and U15804 (N_15804,N_12067,N_13280);
xor U15805 (N_15805,N_13333,N_12903);
xnor U15806 (N_15806,N_12087,N_12839);
xnor U15807 (N_15807,N_12868,N_12679);
and U15808 (N_15808,N_12646,N_12731);
xor U15809 (N_15809,N_12133,N_13080);
nor U15810 (N_15810,N_13031,N_13747);
and U15811 (N_15811,N_12488,N_12327);
or U15812 (N_15812,N_12340,N_13124);
xnor U15813 (N_15813,N_12002,N_12350);
nand U15814 (N_15814,N_12044,N_12583);
nand U15815 (N_15815,N_13559,N_13141);
xor U15816 (N_15816,N_12461,N_12019);
or U15817 (N_15817,N_12779,N_12894);
nand U15818 (N_15818,N_13272,N_13550);
xnor U15819 (N_15819,N_13778,N_13514);
nor U15820 (N_15820,N_12487,N_12207);
or U15821 (N_15821,N_12591,N_13671);
nand U15822 (N_15822,N_13046,N_12071);
or U15823 (N_15823,N_12284,N_13931);
xor U15824 (N_15824,N_13357,N_12712);
nand U15825 (N_15825,N_13332,N_12451);
or U15826 (N_15826,N_13775,N_12648);
and U15827 (N_15827,N_12305,N_13806);
nor U15828 (N_15828,N_13525,N_12746);
nand U15829 (N_15829,N_12854,N_13844);
nand U15830 (N_15830,N_12184,N_13925);
xnor U15831 (N_15831,N_13754,N_12671);
xnor U15832 (N_15832,N_13652,N_12012);
xnor U15833 (N_15833,N_13257,N_12753);
or U15834 (N_15834,N_13565,N_13026);
xor U15835 (N_15835,N_12568,N_13136);
or U15836 (N_15836,N_12431,N_13334);
or U15837 (N_15837,N_12611,N_13897);
nand U15838 (N_15838,N_13485,N_13778);
nand U15839 (N_15839,N_12426,N_12359);
and U15840 (N_15840,N_12368,N_12578);
or U15841 (N_15841,N_12252,N_12097);
nor U15842 (N_15842,N_12435,N_12067);
nand U15843 (N_15843,N_12654,N_12131);
nand U15844 (N_15844,N_13130,N_12700);
nand U15845 (N_15845,N_12778,N_13734);
nand U15846 (N_15846,N_13949,N_12847);
nor U15847 (N_15847,N_13299,N_13330);
xnor U15848 (N_15848,N_12286,N_12534);
or U15849 (N_15849,N_12269,N_12277);
xnor U15850 (N_15850,N_13197,N_13432);
xnor U15851 (N_15851,N_13479,N_12441);
and U15852 (N_15852,N_13150,N_13307);
and U15853 (N_15853,N_13450,N_12615);
and U15854 (N_15854,N_13956,N_12264);
nor U15855 (N_15855,N_12052,N_13254);
nand U15856 (N_15856,N_13069,N_12542);
nor U15857 (N_15857,N_13081,N_12663);
nor U15858 (N_15858,N_13471,N_12196);
nor U15859 (N_15859,N_13753,N_12197);
nor U15860 (N_15860,N_12001,N_13058);
xor U15861 (N_15861,N_12921,N_12043);
and U15862 (N_15862,N_12147,N_12309);
nor U15863 (N_15863,N_12962,N_12556);
nor U15864 (N_15864,N_12880,N_13797);
or U15865 (N_15865,N_13224,N_13487);
nor U15866 (N_15866,N_12027,N_13151);
nor U15867 (N_15867,N_12529,N_13495);
or U15868 (N_15868,N_12629,N_13229);
nor U15869 (N_15869,N_12313,N_12173);
xor U15870 (N_15870,N_13570,N_13120);
xor U15871 (N_15871,N_13617,N_13917);
xor U15872 (N_15872,N_12672,N_13772);
nand U15873 (N_15873,N_13838,N_13916);
nand U15874 (N_15874,N_13938,N_13557);
nor U15875 (N_15875,N_13312,N_12353);
nand U15876 (N_15876,N_12336,N_13313);
xnor U15877 (N_15877,N_12573,N_13264);
xor U15878 (N_15878,N_13113,N_12688);
nor U15879 (N_15879,N_12990,N_12722);
or U15880 (N_15880,N_13510,N_12179);
nand U15881 (N_15881,N_12115,N_12599);
or U15882 (N_15882,N_12918,N_12307);
or U15883 (N_15883,N_12931,N_13767);
xor U15884 (N_15884,N_12843,N_13092);
nor U15885 (N_15885,N_12878,N_12571);
and U15886 (N_15886,N_12790,N_13695);
and U15887 (N_15887,N_12354,N_13198);
or U15888 (N_15888,N_12788,N_12335);
nor U15889 (N_15889,N_13111,N_12905);
nand U15890 (N_15890,N_13083,N_12474);
and U15891 (N_15891,N_13506,N_12574);
and U15892 (N_15892,N_12298,N_12873);
nor U15893 (N_15893,N_13893,N_12174);
and U15894 (N_15894,N_13704,N_13354);
nor U15895 (N_15895,N_13523,N_13536);
nor U15896 (N_15896,N_13314,N_13217);
and U15897 (N_15897,N_13983,N_13725);
or U15898 (N_15898,N_12650,N_12908);
and U15899 (N_15899,N_13947,N_12302);
nand U15900 (N_15900,N_12817,N_12006);
or U15901 (N_15901,N_13529,N_12312);
and U15902 (N_15902,N_12063,N_13496);
nor U15903 (N_15903,N_13949,N_12176);
nand U15904 (N_15904,N_13878,N_13205);
xor U15905 (N_15905,N_12514,N_13710);
nor U15906 (N_15906,N_12026,N_12134);
nor U15907 (N_15907,N_12976,N_12710);
xnor U15908 (N_15908,N_13702,N_12781);
and U15909 (N_15909,N_13981,N_12891);
nand U15910 (N_15910,N_12307,N_12242);
or U15911 (N_15911,N_12024,N_13884);
and U15912 (N_15912,N_13774,N_12897);
and U15913 (N_15913,N_12852,N_12271);
nor U15914 (N_15914,N_13354,N_13110);
and U15915 (N_15915,N_12155,N_12385);
or U15916 (N_15916,N_13091,N_12680);
xor U15917 (N_15917,N_13366,N_12625);
or U15918 (N_15918,N_13476,N_12462);
and U15919 (N_15919,N_13042,N_12762);
nand U15920 (N_15920,N_12695,N_12085);
nand U15921 (N_15921,N_13208,N_12148);
nor U15922 (N_15922,N_13901,N_12477);
and U15923 (N_15923,N_12201,N_12526);
and U15924 (N_15924,N_13040,N_13648);
and U15925 (N_15925,N_13997,N_12836);
nor U15926 (N_15926,N_12160,N_13630);
nor U15927 (N_15927,N_13566,N_13004);
xor U15928 (N_15928,N_12413,N_12566);
nor U15929 (N_15929,N_13176,N_13363);
nand U15930 (N_15930,N_12738,N_12728);
xnor U15931 (N_15931,N_12336,N_12223);
or U15932 (N_15932,N_13739,N_12379);
nand U15933 (N_15933,N_12569,N_12734);
and U15934 (N_15934,N_13700,N_12241);
and U15935 (N_15935,N_13533,N_13759);
nor U15936 (N_15936,N_13062,N_13594);
nor U15937 (N_15937,N_12876,N_13676);
nor U15938 (N_15938,N_12854,N_13928);
nand U15939 (N_15939,N_13109,N_12825);
or U15940 (N_15940,N_13548,N_12691);
nand U15941 (N_15941,N_13011,N_12139);
nand U15942 (N_15942,N_12723,N_13687);
nand U15943 (N_15943,N_13103,N_13367);
xor U15944 (N_15944,N_13744,N_12552);
nand U15945 (N_15945,N_13383,N_12534);
xor U15946 (N_15946,N_12155,N_12762);
nand U15947 (N_15947,N_13942,N_13596);
nor U15948 (N_15948,N_12468,N_12638);
or U15949 (N_15949,N_12176,N_12139);
and U15950 (N_15950,N_13073,N_12907);
xor U15951 (N_15951,N_12363,N_12209);
or U15952 (N_15952,N_13963,N_13775);
and U15953 (N_15953,N_13330,N_12107);
or U15954 (N_15954,N_12050,N_12852);
nand U15955 (N_15955,N_13765,N_12181);
xnor U15956 (N_15956,N_13800,N_12398);
or U15957 (N_15957,N_12794,N_13877);
nand U15958 (N_15958,N_13933,N_12938);
xnor U15959 (N_15959,N_12748,N_13098);
xor U15960 (N_15960,N_13558,N_13814);
nand U15961 (N_15961,N_12221,N_12684);
or U15962 (N_15962,N_13882,N_13687);
nor U15963 (N_15963,N_13695,N_12728);
nand U15964 (N_15964,N_13496,N_13882);
xnor U15965 (N_15965,N_12897,N_12288);
and U15966 (N_15966,N_13210,N_12049);
nor U15967 (N_15967,N_13178,N_13799);
xor U15968 (N_15968,N_12377,N_13854);
or U15969 (N_15969,N_13473,N_13329);
xor U15970 (N_15970,N_12731,N_13005);
or U15971 (N_15971,N_13584,N_12759);
nand U15972 (N_15972,N_13598,N_13300);
or U15973 (N_15973,N_13981,N_13501);
xor U15974 (N_15974,N_13407,N_12143);
nor U15975 (N_15975,N_12679,N_12321);
and U15976 (N_15976,N_12962,N_13475);
nor U15977 (N_15977,N_12715,N_12436);
or U15978 (N_15978,N_13014,N_12046);
xnor U15979 (N_15979,N_13027,N_12430);
nor U15980 (N_15980,N_12455,N_12325);
and U15981 (N_15981,N_13458,N_13128);
nor U15982 (N_15982,N_12060,N_13812);
and U15983 (N_15983,N_13779,N_12847);
or U15984 (N_15984,N_12999,N_12219);
xnor U15985 (N_15985,N_12712,N_12338);
xor U15986 (N_15986,N_12378,N_13068);
nand U15987 (N_15987,N_12068,N_12750);
nand U15988 (N_15988,N_12776,N_12628);
and U15989 (N_15989,N_13638,N_13323);
nor U15990 (N_15990,N_13187,N_13601);
nand U15991 (N_15991,N_12708,N_12213);
and U15992 (N_15992,N_13154,N_13823);
or U15993 (N_15993,N_12114,N_13342);
and U15994 (N_15994,N_13465,N_13365);
nand U15995 (N_15995,N_12770,N_12884);
nand U15996 (N_15996,N_13307,N_13804);
and U15997 (N_15997,N_12596,N_13157);
nor U15998 (N_15998,N_13927,N_13690);
nand U15999 (N_15999,N_12939,N_13364);
nor U16000 (N_16000,N_14582,N_15239);
xnor U16001 (N_16001,N_14639,N_15642);
or U16002 (N_16002,N_15110,N_14179);
xor U16003 (N_16003,N_15391,N_14903);
nor U16004 (N_16004,N_14596,N_15418);
xor U16005 (N_16005,N_15376,N_14560);
nand U16006 (N_16006,N_14211,N_14021);
and U16007 (N_16007,N_15645,N_15848);
nor U16008 (N_16008,N_15030,N_14273);
and U16009 (N_16009,N_14876,N_14991);
nand U16010 (N_16010,N_15345,N_15143);
or U16011 (N_16011,N_15728,N_14270);
nor U16012 (N_16012,N_14241,N_14906);
nor U16013 (N_16013,N_15495,N_15254);
nor U16014 (N_16014,N_15475,N_15086);
nand U16015 (N_16015,N_15516,N_14282);
nand U16016 (N_16016,N_15730,N_15206);
xnor U16017 (N_16017,N_15936,N_14435);
xnor U16018 (N_16018,N_15320,N_15613);
nand U16019 (N_16019,N_14386,N_15287);
or U16020 (N_16020,N_15546,N_15330);
or U16021 (N_16021,N_14061,N_15713);
nor U16022 (N_16022,N_15149,N_14075);
nor U16023 (N_16023,N_14234,N_15091);
xnor U16024 (N_16024,N_15170,N_15069);
or U16025 (N_16025,N_15009,N_15465);
nand U16026 (N_16026,N_15694,N_14620);
nand U16027 (N_16027,N_15103,N_14455);
xor U16028 (N_16028,N_14709,N_15035);
and U16029 (N_16029,N_14520,N_14786);
and U16030 (N_16030,N_14653,N_14664);
or U16031 (N_16031,N_14100,N_14073);
xnor U16032 (N_16032,N_14819,N_15467);
nor U16033 (N_16033,N_14918,N_14603);
or U16034 (N_16034,N_14841,N_14838);
xor U16035 (N_16035,N_15136,N_14099);
or U16036 (N_16036,N_15357,N_14087);
xnor U16037 (N_16037,N_15138,N_15273);
or U16038 (N_16038,N_15839,N_15162);
or U16039 (N_16039,N_15702,N_15359);
or U16040 (N_16040,N_14816,N_15837);
nor U16041 (N_16041,N_15981,N_14464);
and U16042 (N_16042,N_14152,N_14198);
or U16043 (N_16043,N_14562,N_15854);
or U16044 (N_16044,N_14742,N_15466);
and U16045 (N_16045,N_14243,N_14064);
nor U16046 (N_16046,N_15260,N_14964);
nor U16047 (N_16047,N_15530,N_14122);
xnor U16048 (N_16048,N_14005,N_14388);
and U16049 (N_16049,N_15844,N_15064);
and U16050 (N_16050,N_14200,N_15797);
nor U16051 (N_16051,N_15288,N_15807);
and U16052 (N_16052,N_14264,N_15571);
nor U16053 (N_16053,N_15010,N_15439);
nor U16054 (N_16054,N_14377,N_14412);
or U16055 (N_16055,N_14789,N_14533);
and U16056 (N_16056,N_14269,N_15248);
nand U16057 (N_16057,N_15880,N_14083);
nor U16058 (N_16058,N_14111,N_14765);
and U16059 (N_16059,N_14602,N_15887);
xor U16060 (N_16060,N_15251,N_14513);
nand U16061 (N_16061,N_15502,N_15884);
or U16062 (N_16062,N_15696,N_14683);
nor U16063 (N_16063,N_14424,N_15105);
nand U16064 (N_16064,N_15974,N_14660);
xor U16065 (N_16065,N_15434,N_14298);
nor U16066 (N_16066,N_14728,N_15099);
nor U16067 (N_16067,N_15169,N_15209);
nor U16068 (N_16068,N_15553,N_15435);
xnor U16069 (N_16069,N_14946,N_14313);
xnor U16070 (N_16070,N_14842,N_15322);
xor U16071 (N_16071,N_15698,N_15221);
xnor U16072 (N_16072,N_14440,N_14771);
nor U16073 (N_16073,N_15924,N_14693);
or U16074 (N_16074,N_14778,N_15021);
nor U16075 (N_16075,N_15853,N_15646);
nor U16076 (N_16076,N_14724,N_15501);
nor U16077 (N_16077,N_14535,N_14416);
nor U16078 (N_16078,N_14925,N_15449);
nand U16079 (N_16079,N_14894,N_14400);
and U16080 (N_16080,N_15392,N_15044);
nor U16081 (N_16081,N_15405,N_14407);
or U16082 (N_16082,N_15989,N_14672);
and U16083 (N_16083,N_15472,N_15255);
and U16084 (N_16084,N_15775,N_15908);
or U16085 (N_16085,N_15963,N_14038);
and U16086 (N_16086,N_15205,N_14056);
or U16087 (N_16087,N_14125,N_15343);
and U16088 (N_16088,N_14248,N_14626);
nand U16089 (N_16089,N_15722,N_14352);
and U16090 (N_16090,N_14833,N_15999);
xor U16091 (N_16091,N_15212,N_14402);
or U16092 (N_16092,N_14847,N_15005);
nand U16093 (N_16093,N_15835,N_15686);
or U16094 (N_16094,N_14315,N_15972);
nor U16095 (N_16095,N_14357,N_14525);
or U16096 (N_16096,N_14527,N_14580);
or U16097 (N_16097,N_15047,N_15580);
xnor U16098 (N_16098,N_15671,N_15036);
nor U16099 (N_16099,N_14654,N_14265);
nor U16100 (N_16100,N_15760,N_14851);
xor U16101 (N_16101,N_15609,N_15590);
xnor U16102 (N_16102,N_14929,N_15558);
nor U16103 (N_16103,N_15046,N_14034);
nand U16104 (N_16104,N_14036,N_14170);
nand U16105 (N_16105,N_14204,N_15290);
or U16106 (N_16106,N_14066,N_15709);
nand U16107 (N_16107,N_14290,N_14237);
xor U16108 (N_16108,N_14011,N_15117);
nor U16109 (N_16109,N_14104,N_14342);
xor U16110 (N_16110,N_15457,N_15104);
nand U16111 (N_16111,N_15125,N_14578);
nor U16112 (N_16112,N_15937,N_15406);
nand U16113 (N_16113,N_14961,N_14311);
and U16114 (N_16114,N_14356,N_15902);
nor U16115 (N_16115,N_14803,N_15802);
nand U16116 (N_16116,N_14835,N_15689);
nand U16117 (N_16117,N_14935,N_15390);
nor U16118 (N_16118,N_14216,N_14589);
xnor U16119 (N_16119,N_15876,N_14146);
or U16120 (N_16120,N_15267,N_15443);
or U16121 (N_16121,N_14327,N_14768);
or U16122 (N_16122,N_14340,N_15763);
xor U16123 (N_16123,N_14249,N_14538);
and U16124 (N_16124,N_14442,N_14246);
nand U16125 (N_16125,N_15263,N_14516);
nand U16126 (N_16126,N_14740,N_14809);
or U16127 (N_16127,N_15824,N_14031);
nor U16128 (N_16128,N_15218,N_14868);
nor U16129 (N_16129,N_14697,N_14871);
nand U16130 (N_16130,N_14700,N_15121);
nand U16131 (N_16131,N_14799,N_15675);
nand U16132 (N_16132,N_14648,N_14201);
nor U16133 (N_16133,N_15300,N_15274);
or U16134 (N_16134,N_15424,N_15393);
and U16135 (N_16135,N_15993,N_14254);
and U16136 (N_16136,N_14154,N_14158);
nor U16137 (N_16137,N_14606,N_14458);
or U16138 (N_16138,N_15083,N_15333);
nor U16139 (N_16139,N_15409,N_14877);
and U16140 (N_16140,N_15298,N_14539);
xnor U16141 (N_16141,N_14554,N_14556);
nor U16142 (N_16142,N_15624,N_14757);
nand U16143 (N_16143,N_15102,N_14611);
nand U16144 (N_16144,N_15517,N_15473);
or U16145 (N_16145,N_15991,N_15574);
and U16146 (N_16146,N_14632,N_15822);
or U16147 (N_16147,N_15183,N_15308);
xor U16148 (N_16148,N_14601,N_15244);
xnor U16149 (N_16149,N_15454,N_15953);
nand U16150 (N_16150,N_15348,N_15327);
or U16151 (N_16151,N_15804,N_14511);
nand U16152 (N_16152,N_14526,N_14820);
xor U16153 (N_16153,N_14225,N_15794);
and U16154 (N_16154,N_14504,N_15927);
nand U16155 (N_16155,N_14451,N_14659);
or U16156 (N_16156,N_14532,N_15858);
xnor U16157 (N_16157,N_15758,N_14780);
or U16158 (N_16158,N_15237,N_15626);
xor U16159 (N_16159,N_14414,N_14177);
and U16160 (N_16160,N_14908,N_15331);
nor U16161 (N_16161,N_15378,N_15453);
or U16162 (N_16162,N_15695,N_14937);
and U16163 (N_16163,N_14755,N_14756);
xnor U16164 (N_16164,N_15965,N_15707);
or U16165 (N_16165,N_15592,N_15855);
or U16166 (N_16166,N_14068,N_15401);
and U16167 (N_16167,N_14597,N_15762);
xnor U16168 (N_16168,N_14323,N_14507);
xnor U16169 (N_16169,N_14297,N_14845);
and U16170 (N_16170,N_15129,N_15124);
and U16171 (N_16171,N_15411,N_15485);
or U16172 (N_16172,N_15353,N_15647);
xor U16173 (N_16173,N_14354,N_14174);
or U16174 (N_16174,N_14417,N_15422);
or U16175 (N_16175,N_14930,N_14167);
nor U16176 (N_16176,N_14370,N_15544);
or U16177 (N_16177,N_14879,N_14481);
nor U16178 (N_16178,N_14896,N_14694);
and U16179 (N_16179,N_15634,N_15177);
nand U16180 (N_16180,N_14529,N_15076);
and U16181 (N_16181,N_14522,N_14921);
or U16182 (N_16182,N_14128,N_14848);
or U16183 (N_16183,N_14067,N_14832);
or U16184 (N_16184,N_15753,N_14643);
nand U16185 (N_16185,N_15190,N_14957);
or U16186 (N_16186,N_14677,N_14818);
and U16187 (N_16187,N_15909,N_15447);
nor U16188 (N_16188,N_15635,N_14897);
nor U16189 (N_16189,N_15875,N_15564);
nand U16190 (N_16190,N_14114,N_15342);
xnor U16191 (N_16191,N_14119,N_14625);
xnor U16192 (N_16192,N_15795,N_14934);
nand U16193 (N_16193,N_15660,N_15462);
and U16194 (N_16194,N_14893,N_14762);
and U16195 (N_16195,N_15982,N_14014);
or U16196 (N_16196,N_14536,N_15662);
xnor U16197 (N_16197,N_14194,N_15264);
and U16198 (N_16198,N_15524,N_15400);
or U16199 (N_16199,N_14493,N_15396);
or U16200 (N_16200,N_14055,N_14076);
nand U16201 (N_16201,N_14227,N_15643);
or U16202 (N_16202,N_15305,N_15262);
or U16203 (N_16203,N_15856,N_14191);
nand U16204 (N_16204,N_14239,N_15432);
xor U16205 (N_16205,N_14035,N_14737);
xor U16206 (N_16206,N_15810,N_15040);
or U16207 (N_16207,N_15368,N_14182);
and U16208 (N_16208,N_15633,N_14524);
xnor U16209 (N_16209,N_15610,N_15277);
xnor U16210 (N_16210,N_15976,N_14051);
and U16211 (N_16211,N_14115,N_14716);
xor U16212 (N_16212,N_15898,N_15120);
nand U16213 (N_16213,N_14463,N_15967);
or U16214 (N_16214,N_15606,N_14749);
nand U16215 (N_16215,N_14380,N_14362);
or U16216 (N_16216,N_15764,N_14149);
and U16217 (N_16217,N_15272,N_14886);
nor U16218 (N_16218,N_15257,N_15559);
or U16219 (N_16219,N_14423,N_15754);
or U16220 (N_16220,N_14595,N_14806);
nor U16221 (N_16221,N_15868,N_14408);
nand U16222 (N_16222,N_15388,N_14272);
or U16223 (N_16223,N_14502,N_14418);
nand U16224 (N_16224,N_15509,N_14633);
nor U16225 (N_16225,N_14523,N_14199);
or U16226 (N_16226,N_15903,N_14397);
and U16227 (N_16227,N_15906,N_15625);
or U16228 (N_16228,N_14292,N_14287);
and U16229 (N_16229,N_15828,N_14245);
xnor U16230 (N_16230,N_14193,N_15302);
nor U16231 (N_16231,N_14118,N_14624);
xnor U16232 (N_16232,N_15446,N_14933);
or U16233 (N_16233,N_14656,N_14053);
xor U16234 (N_16234,N_14341,N_15072);
and U16235 (N_16235,N_15483,N_15594);
nor U16236 (N_16236,N_15293,N_15080);
xnor U16237 (N_16237,N_15245,N_14283);
or U16238 (N_16238,N_14263,N_15106);
xor U16239 (N_16239,N_14781,N_14884);
xor U16240 (N_16240,N_15334,N_14593);
and U16241 (N_16241,N_14004,N_15360);
and U16242 (N_16242,N_15512,N_15441);
nor U16243 (N_16243,N_15088,N_15479);
or U16244 (N_16244,N_14049,N_15510);
nand U16245 (N_16245,N_15112,N_15744);
or U16246 (N_16246,N_15377,N_14289);
nor U16247 (N_16247,N_14967,N_14197);
xor U16248 (N_16248,N_14276,N_14404);
xor U16249 (N_16249,N_14092,N_14202);
nor U16250 (N_16250,N_14133,N_15496);
xnor U16251 (N_16251,N_14782,N_15486);
nor U16252 (N_16252,N_15039,N_15017);
nand U16253 (N_16253,N_15407,N_14218);
or U16254 (N_16254,N_14175,N_14647);
xnor U16255 (N_16255,N_14666,N_14013);
or U16256 (N_16256,N_15202,N_15242);
nor U16257 (N_16257,N_14837,N_14293);
xor U16258 (N_16258,N_15195,N_14335);
and U16259 (N_16259,N_15881,N_14102);
xnor U16260 (N_16260,N_14376,N_15016);
xor U16261 (N_16261,N_15618,N_14856);
or U16262 (N_16262,N_15291,N_15975);
xor U16263 (N_16263,N_15068,N_14079);
nor U16264 (N_16264,N_14394,N_15787);
nand U16265 (N_16265,N_14576,N_15135);
and U16266 (N_16266,N_14337,N_15816);
xor U16267 (N_16267,N_15374,N_14547);
nor U16268 (N_16268,N_15065,N_14044);
nand U16269 (N_16269,N_15949,N_15750);
and U16270 (N_16270,N_15012,N_14718);
and U16271 (N_16271,N_14431,N_15830);
or U16272 (N_16272,N_15751,N_14330);
nand U16273 (N_16273,N_15747,N_14622);
or U16274 (N_16274,N_15523,N_14326);
xnor U16275 (N_16275,N_15598,N_15299);
xnor U16276 (N_16276,N_14347,N_14579);
nand U16277 (N_16277,N_14301,N_15285);
xor U16278 (N_16278,N_14508,N_15167);
xnor U16279 (N_16279,N_15600,N_15281);
nor U16280 (N_16280,N_15180,N_15387);
or U16281 (N_16281,N_14396,N_15301);
nand U16282 (N_16282,N_15629,N_14453);
xor U16283 (N_16283,N_15476,N_15737);
nor U16284 (N_16284,N_15096,N_15872);
and U16285 (N_16285,N_14260,N_15528);
or U16286 (N_16286,N_15535,N_14528);
or U16287 (N_16287,N_14422,N_15061);
xor U16288 (N_16288,N_14678,N_14911);
nand U16289 (N_16289,N_14085,N_14325);
xor U16290 (N_16290,N_14040,N_15361);
or U16291 (N_16291,N_15402,N_15961);
and U16292 (N_16292,N_15461,N_15259);
xor U16293 (N_16293,N_15394,N_15160);
or U16294 (N_16294,N_15504,N_14619);
or U16295 (N_16295,N_15507,N_15211);
or U16296 (N_16296,N_15605,N_14302);
and U16297 (N_16297,N_14558,N_15716);
nor U16298 (N_16298,N_15265,N_15951);
or U16299 (N_16299,N_14178,N_14753);
nand U16300 (N_16300,N_15790,N_14738);
and U16301 (N_16301,N_15131,N_15986);
nand U16302 (N_16302,N_15860,N_15018);
xnor U16303 (N_16303,N_15042,N_14120);
nor U16304 (N_16304,N_14881,N_14669);
xor U16305 (N_16305,N_15720,N_15670);
and U16306 (N_16306,N_14153,N_14494);
or U16307 (N_16307,N_15210,N_15907);
xnor U16308 (N_16308,N_15997,N_14888);
nand U16309 (N_16309,N_15203,N_15487);
nor U16310 (N_16310,N_14534,N_15664);
and U16311 (N_16311,N_15778,N_14452);
xnor U16312 (N_16312,N_15819,N_15352);
nand U16313 (N_16313,N_15998,N_14996);
or U16314 (N_16314,N_14696,N_15591);
nand U16315 (N_16315,N_15630,N_15307);
or U16316 (N_16316,N_14584,N_15252);
nor U16317 (N_16317,N_15452,N_14018);
xor U16318 (N_16318,N_14989,N_15770);
nand U16319 (N_16319,N_14460,N_15145);
and U16320 (N_16320,N_14480,N_15870);
nand U16321 (N_16321,N_14438,N_15782);
and U16322 (N_16322,N_15067,N_15513);
or U16323 (N_16323,N_14016,N_15236);
and U16324 (N_16324,N_14634,N_14932);
xnor U16325 (N_16325,N_15692,N_14971);
nor U16326 (N_16326,N_14675,N_14462);
xor U16327 (N_16327,N_14710,N_15988);
or U16328 (N_16328,N_15745,N_15712);
nand U16329 (N_16329,N_14434,N_15231);
or U16330 (N_16330,N_15756,N_14840);
or U16331 (N_16331,N_14296,N_14505);
xnor U16332 (N_16332,N_14566,N_15531);
nand U16333 (N_16333,N_14256,N_15585);
xnor U16334 (N_16334,N_15289,N_14640);
nor U16335 (N_16335,N_14430,N_15929);
or U16336 (N_16336,N_14637,N_14873);
nor U16337 (N_16337,N_14086,N_15187);
and U16338 (N_16338,N_14486,N_15958);
and U16339 (N_16339,N_15911,N_14735);
and U16340 (N_16340,N_14895,N_14349);
xnor U16341 (N_16341,N_14824,N_14890);
and U16342 (N_16342,N_15074,N_14096);
nor U16343 (N_16343,N_14915,N_15777);
nor U16344 (N_16344,N_14854,N_15148);
nand U16345 (N_16345,N_14332,N_15666);
or U16346 (N_16346,N_15776,N_15247);
nand U16347 (N_16347,N_15832,N_14145);
and U16348 (N_16348,N_14047,N_14926);
nor U16349 (N_16349,N_15404,N_14324);
and U16350 (N_16350,N_14108,N_14319);
nand U16351 (N_16351,N_15771,N_15413);
nand U16352 (N_16352,N_15621,N_15749);
or U16353 (N_16353,N_14711,N_15948);
nor U16354 (N_16354,N_14846,N_15878);
or U16355 (N_16355,N_15139,N_14081);
or U16356 (N_16356,N_15155,N_15834);
or U16357 (N_16357,N_14155,N_14322);
or U16358 (N_16358,N_15415,N_14131);
and U16359 (N_16359,N_15679,N_15176);
xor U16360 (N_16360,N_15324,N_15107);
or U16361 (N_16361,N_14413,N_14392);
nor U16362 (N_16362,N_15164,N_15665);
nor U16363 (N_16363,N_15078,N_15286);
or U16364 (N_16364,N_14927,N_14224);
nor U16365 (N_16365,N_14776,N_15056);
or U16366 (N_16366,N_14623,N_15850);
nand U16367 (N_16367,N_15372,N_14148);
and U16368 (N_16368,N_14057,N_15426);
xnor U16369 (N_16369,N_15674,N_14823);
nor U16370 (N_16370,N_15623,N_15026);
or U16371 (N_16371,N_14232,N_15450);
nand U16372 (N_16372,N_14746,N_14215);
nor U16373 (N_16373,N_15494,N_15442);
nand U16374 (N_16374,N_14866,N_14787);
xnor U16375 (N_16375,N_15081,N_14106);
nor U16376 (N_16376,N_15229,N_15650);
nand U16377 (N_16377,N_14891,N_14110);
and U16378 (N_16378,N_15410,N_15539);
xor U16379 (N_16379,N_14280,N_15736);
nor U16380 (N_16380,N_15729,N_15704);
or U16381 (N_16381,N_15966,N_14981);
or U16382 (N_16382,N_14288,N_14207);
and U16383 (N_16383,N_14985,N_15383);
or U16384 (N_16384,N_15556,N_14844);
and U16385 (N_16385,N_14450,N_14229);
nor U16386 (N_16386,N_15367,N_15134);
xnor U16387 (N_16387,N_14387,N_14140);
and U16388 (N_16388,N_14600,N_14317);
nor U16389 (N_16389,N_15395,N_14609);
nor U16390 (N_16390,N_15885,N_15208);
nand U16391 (N_16391,N_14630,N_14503);
nor U16392 (N_16392,N_14271,N_15332);
xnor U16393 (N_16393,N_14752,N_15693);
nor U16394 (N_16394,N_14939,N_15188);
nor U16395 (N_16395,N_15586,N_15127);
and U16396 (N_16396,N_14267,N_15799);
xnor U16397 (N_16397,N_15869,N_15701);
nand U16398 (N_16398,N_15784,N_14261);
and U16399 (N_16399,N_14112,N_15216);
and U16400 (N_16400,N_15962,N_14121);
and U16401 (N_16401,N_15493,N_15817);
nor U16402 (N_16402,N_14334,N_14468);
nand U16403 (N_16403,N_14770,N_15399);
or U16404 (N_16404,N_15873,N_15358);
and U16405 (N_16405,N_15258,N_14238);
nor U16406 (N_16406,N_14938,N_14855);
and U16407 (N_16407,N_15373,N_15841);
or U16408 (N_16408,N_15077,N_15891);
xnor U16409 (N_16409,N_15888,N_15964);
or U16410 (N_16410,N_14421,N_15339);
nor U16411 (N_16411,N_14916,N_14138);
and U16412 (N_16412,N_15969,N_15901);
nand U16413 (N_16413,N_14321,N_14590);
xnor U16414 (N_16414,N_15651,N_14312);
nand U16415 (N_16415,N_14371,N_14763);
or U16416 (N_16416,N_14466,N_14975);
xnor U16417 (N_16417,N_14251,N_14180);
nor U16418 (N_16418,N_15939,N_14613);
or U16419 (N_16419,N_15719,N_14429);
xnor U16420 (N_16420,N_14320,N_15992);
xor U16421 (N_16421,N_14344,N_14492);
nand U16422 (N_16422,N_15561,N_14472);
xor U16423 (N_16423,N_15057,N_15282);
nand U16424 (N_16424,N_14567,N_14807);
nor U16425 (N_16425,N_14682,N_15551);
nor U16426 (N_16426,N_14266,N_15738);
xor U16427 (N_16427,N_14420,N_15836);
nand U16428 (N_16428,N_15568,N_14662);
nor U16429 (N_16429,N_15349,N_15217);
xor U16430 (N_16430,N_15363,N_15726);
nand U16431 (N_16431,N_14834,N_14253);
nand U16432 (N_16432,N_14875,N_15604);
or U16433 (N_16433,N_15011,N_14954);
xnor U16434 (N_16434,N_15655,N_14439);
xor U16435 (N_16435,N_15224,N_14947);
nand U16436 (N_16436,N_14960,N_14427);
or U16437 (N_16437,N_14867,N_14316);
nor U16438 (N_16438,N_15663,N_14974);
or U16439 (N_16439,N_15329,N_15806);
xnor U16440 (N_16440,N_14808,N_14663);
xor U16441 (N_16441,N_14722,N_14258);
xnor U16442 (N_16442,N_15996,N_15573);
nand U16443 (N_16443,N_15041,N_15550);
and U16444 (N_16444,N_14754,N_15978);
and U16445 (N_16445,N_14374,N_15004);
nor U16446 (N_16446,N_14173,N_14655);
and U16447 (N_16447,N_14052,N_14779);
xor U16448 (N_16448,N_14428,N_15230);
xor U16449 (N_16449,N_15567,N_14684);
and U16450 (N_16450,N_15708,N_14113);
or U16451 (N_16451,N_14644,N_14491);
and U16452 (N_16452,N_14457,N_14210);
nor U16453 (N_16453,N_15984,N_15350);
or U16454 (N_16454,N_14046,N_15788);
xnor U16455 (N_16455,N_15542,N_14990);
nor U16456 (N_16456,N_14360,N_15168);
or U16457 (N_16457,N_14994,N_15137);
and U16458 (N_16458,N_14591,N_14060);
or U16459 (N_16459,N_14409,N_14432);
and U16460 (N_16460,N_15603,N_14187);
or U16461 (N_16461,N_14236,N_14213);
xor U16462 (N_16462,N_15470,N_15488);
and U16463 (N_16463,N_15700,N_14163);
nand U16464 (N_16464,N_14708,N_15612);
and U16465 (N_16465,N_14817,N_15656);
nor U16466 (N_16466,N_15825,N_15781);
nand U16467 (N_16467,N_15191,N_14345);
or U16468 (N_16468,N_15222,N_15882);
and U16469 (N_16469,N_15667,N_15566);
and U16470 (N_16470,N_14869,N_14375);
nor U16471 (N_16471,N_14605,N_14403);
nand U16472 (N_16472,N_14917,N_15514);
nand U16473 (N_16473,N_14949,N_14476);
nor U16474 (N_16474,N_15464,N_14515);
nor U16475 (N_16475,N_14030,N_15182);
nor U16476 (N_16476,N_15955,N_15007);
nand U16477 (N_16477,N_14661,N_14758);
and U16478 (N_16478,N_15685,N_14736);
nor U16479 (N_16479,N_14367,N_14530);
xor U16480 (N_16480,N_15743,N_14594);
nand U16481 (N_16481,N_14080,N_15602);
or U16482 (N_16482,N_14945,N_15283);
or U16483 (N_16483,N_14156,N_14471);
xor U16484 (N_16484,N_14278,N_14565);
nor U16485 (N_16485,N_15555,N_15628);
nor U16486 (N_16486,N_14039,N_14901);
and U16487 (N_16487,N_14310,N_14027);
xor U16488 (N_16488,N_14902,N_14761);
and U16489 (N_16489,N_14373,N_15582);
xor U16490 (N_16490,N_14006,N_15150);
nand U16491 (N_16491,N_15108,N_15027);
and U16492 (N_16492,N_15431,N_15351);
nand U16493 (N_16493,N_14727,N_15022);
nand U16494 (N_16494,N_15680,N_15940);
xnor U16495 (N_16495,N_14037,N_14725);
nor U16496 (N_16496,N_14563,N_14222);
nand U16497 (N_16497,N_15721,N_15425);
nor U16498 (N_16498,N_15115,N_14348);
xor U16499 (N_16499,N_15611,N_14226);
or U16500 (N_16500,N_14559,N_14825);
xor U16501 (N_16501,N_14262,N_15589);
or U16502 (N_16502,N_15920,N_15658);
nand U16503 (N_16503,N_14998,N_15774);
nand U16504 (N_16504,N_15627,N_15877);
and U16505 (N_16505,N_15673,N_14135);
or U16506 (N_16506,N_14003,N_14168);
or U16507 (N_16507,N_15430,N_14023);
nand U16508 (N_16508,N_15968,N_14510);
and U16509 (N_16509,N_15956,N_15805);
or U16510 (N_16510,N_15003,N_14892);
or U16511 (N_16511,N_14343,N_14361);
nor U16512 (N_16512,N_15499,N_14864);
and U16513 (N_16513,N_15196,N_15250);
or U16514 (N_16514,N_15101,N_14368);
nor U16515 (N_16515,N_15560,N_15733);
and U16516 (N_16516,N_15639,N_14446);
nand U16517 (N_16517,N_14720,N_14859);
and U16518 (N_16518,N_14870,N_15140);
xor U16519 (N_16519,N_14733,N_15020);
and U16520 (N_16520,N_14285,N_15313);
or U16521 (N_16521,N_14936,N_15468);
xor U16522 (N_16522,N_14105,N_15172);
or U16523 (N_16523,N_15883,N_14924);
nor U16524 (N_16524,N_15050,N_15380);
xnor U16525 (N_16525,N_14699,N_15809);
nand U16526 (N_16526,N_15938,N_14483);
and U16527 (N_16527,N_14689,N_14351);
or U16528 (N_16528,N_14797,N_14642);
xor U16529 (N_16529,N_15829,N_15100);
nand U16530 (N_16530,N_15279,N_15318);
nand U16531 (N_16531,N_14043,N_15641);
xor U16532 (N_16532,N_15717,N_15356);
xnor U16533 (N_16533,N_15532,N_15607);
xor U16534 (N_16534,N_15142,N_14355);
nand U16535 (N_16535,N_14557,N_14062);
nand U16536 (N_16536,N_14872,N_15033);
nand U16537 (N_16537,N_15654,N_15079);
nor U16538 (N_16538,N_14958,N_15718);
nand U16539 (N_16539,N_15581,N_15175);
xnor U16540 (N_16540,N_14860,N_14717);
and U16541 (N_16541,N_14764,N_14747);
or U16542 (N_16542,N_15979,N_14090);
xor U16543 (N_16543,N_15133,N_14657);
xnor U16544 (N_16544,N_15147,N_15306);
xnor U16545 (N_16545,N_15253,N_15173);
nand U16546 (N_16546,N_15522,N_15636);
and U16547 (N_16547,N_14127,N_15793);
and U16548 (N_16548,N_15798,N_14604);
nor U16549 (N_16549,N_14792,N_14001);
and U16550 (N_16550,N_14788,N_14801);
nand U16551 (N_16551,N_14495,N_15119);
nand U16552 (N_16552,N_14072,N_15386);
nor U16553 (N_16553,N_14955,N_15058);
and U16554 (N_16554,N_15132,N_14517);
nor U16555 (N_16555,N_14790,N_15015);
xnor U16556 (N_16556,N_15765,N_15292);
or U16557 (N_16557,N_15772,N_15543);
or U16558 (N_16558,N_14688,N_14705);
or U16559 (N_16559,N_15894,N_15918);
and U16560 (N_16560,N_15688,N_14071);
xor U16561 (N_16561,N_15648,N_14116);
and U16562 (N_16562,N_15294,N_15225);
nand U16563 (N_16563,N_14369,N_15821);
and U16564 (N_16564,N_14714,N_15497);
and U16565 (N_16565,N_14988,N_14544);
nor U16566 (N_16566,N_15595,N_15631);
xor U16567 (N_16567,N_15826,N_14305);
and U16568 (N_16568,N_15326,N_15480);
nand U16569 (N_16569,N_14134,N_14189);
xor U16570 (N_16570,N_15928,N_15013);
nor U16571 (N_16571,N_14521,N_15536);
xnor U16572 (N_16572,N_15866,N_14658);
nand U16573 (N_16573,N_14772,N_15416);
nand U16574 (N_16574,N_14058,N_15917);
or U16575 (N_16575,N_15093,N_15228);
xor U16576 (N_16576,N_14196,N_15128);
or U16577 (N_16577,N_14217,N_15319);
nand U16578 (N_16578,N_14759,N_15214);
nand U16579 (N_16579,N_14015,N_14309);
xor U16580 (N_16580,N_14564,N_15703);
nand U16581 (N_16581,N_15970,N_14910);
and U16582 (N_16582,N_14953,N_15491);
xor U16583 (N_16583,N_15682,N_14931);
nor U16584 (N_16584,N_15001,N_14461);
nor U16585 (N_16585,N_14542,N_15316);
xor U16586 (N_16586,N_14951,N_15786);
xor U16587 (N_16587,N_15570,N_14028);
or U16588 (N_16588,N_14997,N_15240);
and U16589 (N_16589,N_15219,N_14865);
xnor U16590 (N_16590,N_14497,N_14117);
and U16591 (N_16591,N_15932,N_15490);
xor U16592 (N_16592,N_14509,N_14398);
or U16593 (N_16593,N_14952,N_14674);
nand U16594 (N_16594,N_14089,N_14235);
xnor U16595 (N_16595,N_14691,N_15525);
xor U16596 (N_16596,N_14275,N_14443);
nand U16597 (N_16597,N_14889,N_14598);
or U16598 (N_16598,N_14830,N_14880);
xnor U16599 (N_16599,N_15921,N_14793);
nor U16600 (N_16600,N_15616,N_15983);
xor U16601 (N_16601,N_15699,N_15608);
xnor U16602 (N_16602,N_14706,N_14702);
and U16603 (N_16603,N_15533,N_14069);
nand U16604 (N_16604,N_14181,N_15934);
or U16605 (N_16605,N_14569,N_14905);
and U16606 (N_16606,N_14704,N_14009);
nor U16607 (N_16607,N_15095,N_14571);
nand U16608 (N_16608,N_15249,N_14393);
and U16609 (N_16609,N_14732,N_15896);
nor U16610 (N_16610,N_14208,N_14979);
or U16611 (N_16611,N_14853,N_14852);
xor U16612 (N_16612,N_14795,N_15233);
nor U16613 (N_16613,N_14192,N_14922);
nor U16614 (N_16614,N_14032,N_14339);
xor U16615 (N_16615,N_15842,N_15547);
or U16616 (N_16616,N_15460,N_15597);
and U16617 (N_16617,N_15813,N_14157);
nor U16618 (N_16618,N_14615,N_15672);
xnor U16619 (N_16619,N_15448,N_15960);
nor U16620 (N_16620,N_14641,N_15181);
nor U16621 (N_16621,N_14353,N_15534);
nand U16622 (N_16622,N_15537,N_14518);
or U16623 (N_16623,N_15584,N_14415);
or U16624 (N_16624,N_14000,N_14804);
xor U16625 (N_16625,N_15159,N_15098);
xor U16626 (N_16626,N_14712,N_15583);
xnor U16627 (N_16627,N_15846,N_15375);
nand U16628 (N_16628,N_14585,N_15735);
nor U16629 (N_16629,N_14631,N_14328);
or U16630 (N_16630,N_15803,N_14381);
nand U16631 (N_16631,N_14449,N_15433);
and U16632 (N_16632,N_15614,N_15029);
nor U16633 (N_16633,N_15578,N_15243);
or U16634 (N_16634,N_15893,N_15311);
xor U16635 (N_16635,N_14426,N_14383);
or U16636 (N_16636,N_14745,N_15904);
xor U16637 (N_16637,N_14652,N_15801);
nor U16638 (N_16638,N_14454,N_14882);
nor U16639 (N_16639,N_14791,N_15575);
xnor U16640 (N_16640,N_15840,N_15122);
or U16641 (N_16641,N_15994,N_14977);
or U16642 (N_16642,N_15032,N_15985);
and U16643 (N_16643,N_15498,N_14912);
or U16644 (N_16644,N_15779,N_14101);
and U16645 (N_16645,N_14231,N_15347);
nor U16646 (N_16646,N_15838,N_14940);
or U16647 (N_16647,N_15508,N_15062);
and U16648 (N_16648,N_14618,N_14599);
xor U16649 (N_16649,N_15238,N_15959);
xor U16650 (N_16650,N_14065,N_15849);
and U16651 (N_16651,N_14378,N_15820);
xnor U16652 (N_16652,N_14822,N_14874);
xnor U16653 (N_16653,N_14406,N_14959);
nor U16654 (N_16654,N_15505,N_15773);
nand U16655 (N_16655,N_15711,N_14195);
and U16656 (N_16656,N_15678,N_15995);
and U16657 (N_16657,N_14751,N_14166);
and U16658 (N_16658,N_15922,N_14329);
or U16659 (N_16659,N_15303,N_15739);
and U16660 (N_16660,N_14577,N_15266);
xnor U16661 (N_16661,N_15545,N_14350);
nor U16662 (N_16662,N_14548,N_14022);
nand U16663 (N_16663,N_14151,N_15905);
xnor U16664 (N_16664,N_14448,N_15914);
nor U16665 (N_16665,N_15028,N_14794);
or U16666 (N_16666,N_15066,N_14255);
xor U16667 (N_16667,N_15362,N_14496);
nand U16668 (N_16668,N_15034,N_14665);
or U16669 (N_16669,N_15220,N_15766);
or U16670 (N_16670,N_15338,N_14479);
or U16671 (N_16671,N_15370,N_14963);
nand U16672 (N_16672,N_14919,N_15178);
or U16673 (N_16673,N_14411,N_14303);
or U16674 (N_16674,N_14966,N_15006);
xnor U16675 (N_16675,N_15576,N_15500);
nor U16676 (N_16676,N_14673,N_14074);
xor U16677 (N_16677,N_14379,N_15389);
and U16678 (N_16678,N_14007,N_15084);
nor U16679 (N_16679,N_15049,N_14171);
and U16680 (N_16680,N_15785,N_14815);
or U16681 (N_16681,N_15075,N_14487);
or U16682 (N_16682,N_15000,N_15163);
or U16683 (N_16683,N_14190,N_14813);
xor U16684 (N_16684,N_14646,N_14729);
xor U16685 (N_16685,N_15557,N_15890);
nand U16686 (N_16686,N_14132,N_14686);
and U16687 (N_16687,N_15827,N_15601);
xnor U16688 (N_16688,N_15193,N_14731);
nand U16689 (N_16689,N_15146,N_14827);
nor U16690 (N_16690,N_14063,N_15463);
and U16691 (N_16691,N_15429,N_15270);
xor U16692 (N_16692,N_15861,N_14026);
nor U16693 (N_16693,N_15144,N_14206);
nor U16694 (N_16694,N_15746,N_14690);
nor U16695 (N_16695,N_14048,N_15954);
and U16696 (N_16696,N_14250,N_15053);
or U16697 (N_16697,N_15328,N_14465);
or U16698 (N_16698,N_15089,N_15458);
xnor U16699 (N_16699,N_14010,N_14553);
and U16700 (N_16700,N_14359,N_15166);
or U16701 (N_16701,N_15622,N_14670);
or U16702 (N_16702,N_15048,N_14968);
and U16703 (N_16703,N_15185,N_15198);
nor U16704 (N_16704,N_14291,N_14221);
xnor U16705 (N_16705,N_14800,N_15973);
xnor U16706 (N_16706,N_15977,N_14364);
or U16707 (N_16707,N_14760,N_14980);
nor U16708 (N_16708,N_15436,N_14441);
xor U16709 (N_16709,N_14723,N_14410);
xor U16710 (N_16710,N_15538,N_14574);
nor U16711 (N_16711,N_14501,N_15895);
or U16712 (N_16712,N_14984,N_15354);
nor U16713 (N_16713,N_15620,N_14734);
or U16714 (N_16714,N_15572,N_14887);
and U16715 (N_16715,N_15755,N_14839);
nand U16716 (N_16716,N_15925,N_14017);
and U16717 (N_16717,N_14203,N_14220);
nor U16718 (N_16718,N_15569,N_14572);
nand U16719 (N_16719,N_15097,N_15130);
or U16720 (N_16720,N_15831,N_15451);
nor U16721 (N_16721,N_15725,N_15280);
xor U16722 (N_16722,N_14144,N_14995);
nand U16723 (N_16723,N_14774,N_15867);
nor U16724 (N_16724,N_14103,N_15661);
or U16725 (N_16725,N_14484,N_15019);
xnor U16726 (N_16726,N_14913,N_14172);
or U16727 (N_16727,N_15037,N_14685);
nor U16728 (N_16728,N_15278,N_15950);
nor U16729 (N_16729,N_15085,N_14469);
xnor U16730 (N_16730,N_14907,N_15577);
or U16731 (N_16731,N_15833,N_15926);
nand U16732 (N_16732,N_14259,N_15412);
nand U16733 (N_16733,N_14695,N_14233);
nand U16734 (N_16734,N_15268,N_15070);
nor U16735 (N_16735,N_14136,N_14671);
and U16736 (N_16736,N_15506,N_15800);
nand U16737 (N_16737,N_15579,N_15296);
xnor U16738 (N_16738,N_14545,N_14812);
or U16739 (N_16739,N_14970,N_15269);
xnor U16740 (N_16740,N_14651,N_15141);
nand U16741 (N_16741,N_15640,N_15847);
xnor U16742 (N_16742,N_15593,N_14008);
and U16743 (N_16743,N_15731,N_15596);
nor U16744 (N_16744,N_15420,N_14987);
or U16745 (N_16745,N_15477,N_15060);
or U16746 (N_16746,N_15456,N_14920);
or U16747 (N_16747,N_14537,N_15687);
nand U16748 (N_16748,N_15340,N_15653);
nand U16749 (N_16749,N_15520,N_15549);
nand U16750 (N_16750,N_15706,N_14284);
and U16751 (N_16751,N_15227,N_14419);
and U16752 (N_16752,N_14552,N_14811);
nand U16753 (N_16753,N_14054,N_15174);
and U16754 (N_16754,N_15123,N_14923);
nand U16755 (N_16755,N_15478,N_15541);
and U16756 (N_16756,N_15474,N_15864);
or U16757 (N_16757,N_14095,N_15059);
and U16758 (N_16758,N_14719,N_15043);
xnor U16759 (N_16759,N_15444,N_14898);
nand U16760 (N_16760,N_15428,N_14474);
and U16761 (N_16761,N_14561,N_14617);
xor U16762 (N_16762,N_15179,N_15371);
and U16763 (N_16763,N_15789,N_15152);
xor U16764 (N_16764,N_14878,N_15369);
nor U16765 (N_16765,N_15341,N_15638);
nand U16766 (N_16766,N_14176,N_15489);
nor U16767 (N_16767,N_15304,N_15200);
nor U16768 (N_16768,N_14904,N_14286);
or U16769 (N_16769,N_15052,N_15082);
xor U16770 (N_16770,N_15649,N_15957);
and U16771 (N_16771,N_15197,N_14425);
and U16772 (N_16772,N_15857,N_14242);
nand U16773 (N_16773,N_15714,N_15683);
and U16774 (N_16774,N_15421,N_15644);
nand U16775 (N_16775,N_15379,N_14628);
nor U16776 (N_16776,N_15808,N_15364);
xor U16777 (N_16777,N_15886,N_14078);
nor U16778 (N_16778,N_14586,N_15438);
xor U16779 (N_16779,N_15768,N_14391);
xor U16780 (N_16780,N_14459,N_15309);
nand U16781 (N_16781,N_15023,N_15892);
or U16782 (N_16782,N_15599,N_14721);
and U16783 (N_16783,N_15054,N_14581);
xor U16784 (N_16784,N_15910,N_14214);
xnor U16785 (N_16785,N_14247,N_15796);
nand U16786 (N_16786,N_14785,N_14050);
xnor U16787 (N_16787,N_14300,N_14540);
nor U16788 (N_16788,N_15859,N_14713);
nand U16789 (N_16789,N_14676,N_14992);
xnor U16790 (N_16790,N_14024,N_15382);
nand U16791 (N_16791,N_15156,N_14703);
and U16792 (N_16792,N_15346,N_14485);
nand U16793 (N_16793,N_15271,N_14636);
and U16794 (N_16794,N_15780,N_15710);
nand U16795 (N_16795,N_14784,N_14956);
nor U16796 (N_16796,N_15529,N_14976);
nand U16797 (N_16797,N_15915,N_14549);
nand U16798 (N_16798,N_14186,N_14307);
nor U16799 (N_16799,N_14775,N_15715);
nand U16800 (N_16800,N_14543,N_14783);
xnor U16801 (N_16801,N_15310,N_14109);
nor U16802 (N_16802,N_15090,N_15863);
xnor U16803 (N_16803,N_14318,N_15677);
and U16804 (N_16804,N_15912,N_14928);
or U16805 (N_16805,N_15862,N_15153);
nor U16806 (N_16806,N_15384,N_14070);
and U16807 (N_16807,N_15323,N_15843);
nand U16808 (N_16808,N_14831,N_15192);
xor U16809 (N_16809,N_14629,N_15365);
nand U16810 (N_16810,N_14899,N_15171);
xnor U16811 (N_16811,N_14650,N_14436);
or U16812 (N_16812,N_15851,N_14978);
or U16813 (N_16813,N_14858,N_14739);
and U16814 (N_16814,N_15705,N_14094);
xnor U16815 (N_16815,N_15038,N_15109);
nand U16816 (N_16816,N_15414,N_15727);
or U16817 (N_16817,N_14943,N_14333);
nor U16818 (N_16818,N_15741,N_14482);
nor U16819 (N_16819,N_14228,N_15511);
xor U16820 (N_16820,N_15337,N_14730);
nand U16821 (N_16821,N_15469,N_14777);
or U16822 (N_16822,N_14372,N_14942);
nor U16823 (N_16823,N_14230,N_14948);
and U16824 (N_16824,N_14627,N_15945);
xnor U16825 (N_16825,N_15314,N_14909);
nand U16826 (N_16826,N_15874,N_15503);
and U16827 (N_16827,N_14240,N_15092);
xnor U16828 (N_16828,N_15814,N_15423);
nor U16829 (N_16829,N_14219,N_15275);
nor U16830 (N_16830,N_15668,N_15923);
nand U16831 (N_16831,N_14033,N_15235);
xnor U16832 (N_16832,N_15812,N_15740);
or U16833 (N_16833,N_14142,N_15742);
xnor U16834 (N_16834,N_15199,N_15919);
and U16835 (N_16835,N_14583,N_15397);
and U16836 (N_16836,N_14531,N_15930);
or U16837 (N_16837,N_15652,N_14012);
xnor U16838 (N_16838,N_15657,N_14857);
or U16839 (N_16839,N_15845,N_15031);
or U16840 (N_16840,N_15521,N_14382);
and U16841 (N_16841,N_15344,N_14701);
xor U16842 (N_16842,N_15669,N_14680);
or U16843 (N_16843,N_14137,N_14437);
or U16844 (N_16844,N_14614,N_15697);
and U16845 (N_16845,N_14478,N_14541);
nand U16846 (N_16846,N_14467,N_14395);
xor U16847 (N_16847,N_15317,N_14308);
nand U16848 (N_16848,N_15158,N_14274);
nand U16849 (N_16849,N_14826,N_14849);
xnor U16850 (N_16850,N_14088,N_15154);
or U16851 (N_16851,N_15659,N_15312);
or U16852 (N_16852,N_15732,N_15990);
nor U16853 (N_16853,N_14972,N_15899);
or U16854 (N_16854,N_15234,N_15767);
nor U16855 (N_16855,N_15223,N_14029);
or U16856 (N_16856,N_14477,N_15201);
and U16857 (N_16857,N_14829,N_15818);
and U16858 (N_16858,N_15315,N_14456);
or U16859 (N_16859,N_14973,N_14962);
nor U16860 (N_16860,N_14570,N_14999);
xor U16861 (N_16861,N_14944,N_15724);
nand U16862 (N_16862,N_14098,N_15437);
nand U16863 (N_16863,N_14850,N_14045);
nor U16864 (N_16864,N_15684,N_14025);
nor U16865 (N_16865,N_14470,N_14750);
and U16866 (N_16866,N_14314,N_14185);
and U16867 (N_16867,N_15515,N_15941);
or U16868 (N_16868,N_14766,N_15051);
nand U16869 (N_16869,N_15871,N_15459);
nor U16870 (N_16870,N_14512,N_15207);
or U16871 (N_16871,N_14645,N_14743);
xor U16872 (N_16872,N_14592,N_14707);
xor U16873 (N_16873,N_14223,N_15261);
nor U16874 (N_16874,N_15114,N_14687);
nor U16875 (N_16875,N_14519,N_14124);
or U16876 (N_16876,N_15482,N_15094);
nor U16877 (N_16877,N_14810,N_14399);
nand U16878 (N_16878,N_14002,N_15943);
nand U16879 (N_16879,N_15637,N_14366);
nand U16880 (N_16880,N_15913,N_15757);
and U16881 (N_16881,N_14741,N_14506);
nand U16882 (N_16882,N_14331,N_15355);
or U16883 (N_16883,N_15184,N_15025);
nand U16884 (N_16884,N_15366,N_14059);
nor U16885 (N_16885,N_14097,N_15471);
or U16886 (N_16886,N_15276,N_14162);
nand U16887 (N_16887,N_15204,N_14159);
or U16888 (N_16888,N_14295,N_15518);
or U16889 (N_16889,N_14621,N_15748);
nand U16890 (N_16890,N_14160,N_14304);
and U16891 (N_16891,N_15295,N_14941);
nor U16892 (N_16892,N_15073,N_15865);
nor U16893 (N_16893,N_14914,N_15615);
or U16894 (N_16894,N_14802,N_15947);
nor U16895 (N_16895,N_14698,N_14401);
nor U16896 (N_16896,N_14635,N_15165);
or U16897 (N_16897,N_15759,N_14500);
nand U16898 (N_16898,N_14141,N_14183);
xnor U16899 (N_16899,N_14798,N_14363);
xor U16900 (N_16900,N_15445,N_14546);
and U16901 (N_16901,N_14184,N_14550);
and U16902 (N_16902,N_14139,N_15381);
nor U16903 (N_16903,N_15232,N_15226);
and U16904 (N_16904,N_14638,N_14205);
nand U16905 (N_16905,N_15690,N_15408);
nor U16906 (N_16906,N_14129,N_14965);
nor U16907 (N_16907,N_14077,N_15946);
xor U16908 (N_16908,N_14130,N_15256);
xor U16909 (N_16909,N_14390,N_14294);
or U16910 (N_16910,N_14123,N_14473);
xnor U16911 (N_16911,N_15935,N_14475);
nor U16912 (N_16912,N_14821,N_14188);
xnor U16913 (N_16913,N_15944,N_14444);
and U16914 (N_16914,N_14209,N_14365);
or U16915 (N_16915,N_15879,N_15897);
or U16916 (N_16916,N_15087,N_15055);
nor U16917 (N_16917,N_15617,N_15157);
nor U16918 (N_16918,N_14551,N_14161);
xnor U16919 (N_16919,N_15151,N_15540);
nor U16920 (N_16920,N_15024,N_14982);
xnor U16921 (N_16921,N_14405,N_14950);
nand U16922 (N_16922,N_15527,N_15111);
nor U16923 (N_16923,N_15823,N_14336);
or U16924 (N_16924,N_14306,N_15723);
nand U16925 (N_16925,N_14692,N_14885);
xnor U16926 (N_16926,N_14796,N_15194);
or U16927 (N_16927,N_14608,N_15417);
nand U16928 (N_16928,N_14126,N_14499);
nand U16929 (N_16929,N_15045,N_15761);
nand U16930 (N_16930,N_14863,N_15071);
xnor U16931 (N_16931,N_14993,N_15419);
xnor U16932 (N_16932,N_14490,N_15933);
nand U16933 (N_16933,N_14244,N_15971);
and U16934 (N_16934,N_14883,N_15014);
or U16935 (N_16935,N_15403,N_15161);
nand U16936 (N_16936,N_15791,N_15189);
xnor U16937 (N_16937,N_15335,N_14082);
xor U16938 (N_16938,N_14433,N_15931);
nand U16939 (N_16939,N_15297,N_14607);
nand U16940 (N_16940,N_15002,N_14612);
and U16941 (N_16941,N_15734,N_14573);
nand U16942 (N_16942,N_14715,N_15980);
and U16943 (N_16943,N_14836,N_14555);
xor U16944 (N_16944,N_15284,N_14252);
or U16945 (N_16945,N_15676,N_15213);
and U16946 (N_16946,N_14042,N_14169);
xnor U16947 (N_16947,N_14862,N_14091);
or U16948 (N_16948,N_15691,N_14588);
nor U16949 (N_16949,N_15552,N_14861);
and U16950 (N_16950,N_14358,N_14767);
xor U16951 (N_16951,N_15455,N_14681);
nand U16952 (N_16952,N_14093,N_14610);
xor U16953 (N_16953,N_15681,N_15427);
nand U16954 (N_16954,N_15126,N_14257);
and U16955 (N_16955,N_15554,N_14587);
nor U16956 (N_16956,N_15241,N_14445);
and U16957 (N_16957,N_15562,N_15484);
and U16958 (N_16958,N_14488,N_14384);
xnor U16959 (N_16959,N_15565,N_15916);
or U16960 (N_16960,N_14389,N_14150);
nor U16961 (N_16961,N_15952,N_14385);
and U16962 (N_16962,N_14165,N_14212);
nand U16963 (N_16963,N_14084,N_14805);
xnor U16964 (N_16964,N_15769,N_15563);
or U16965 (N_16965,N_15063,N_14299);
and U16966 (N_16966,N_14147,N_14575);
nand U16967 (N_16967,N_15811,N_14019);
xnor U16968 (N_16968,N_15325,N_15118);
or U16969 (N_16969,N_15385,N_15752);
nor U16970 (N_16970,N_14814,N_14107);
nand U16971 (N_16971,N_14568,N_14726);
and U16972 (N_16972,N_15548,N_14649);
nand U16973 (N_16973,N_15783,N_14667);
xnor U16974 (N_16974,N_15008,N_14828);
and U16975 (N_16975,N_15588,N_15336);
and U16976 (N_16976,N_14346,N_14986);
and U16977 (N_16977,N_14679,N_14900);
nand U16978 (N_16978,N_15587,N_14020);
and U16979 (N_16979,N_15815,N_15792);
and U16980 (N_16980,N_14277,N_15321);
or U16981 (N_16981,N_15987,N_15440);
xnor U16982 (N_16982,N_14748,N_14773);
and U16983 (N_16983,N_15113,N_14616);
nor U16984 (N_16984,N_14041,N_15519);
xnor U16985 (N_16985,N_15619,N_15398);
and U16986 (N_16986,N_14143,N_14769);
and U16987 (N_16987,N_14983,N_14281);
nor U16988 (N_16988,N_15186,N_15481);
nor U16989 (N_16989,N_14268,N_14489);
nor U16990 (N_16990,N_14843,N_15889);
nand U16991 (N_16991,N_15215,N_15942);
nor U16992 (N_16992,N_15526,N_14498);
and U16993 (N_16993,N_14338,N_14447);
xor U16994 (N_16994,N_14969,N_15852);
nand U16995 (N_16995,N_14164,N_14668);
xnor U16996 (N_16996,N_15116,N_14279);
nand U16997 (N_16997,N_14744,N_15632);
nor U16998 (N_16998,N_15492,N_15900);
nand U16999 (N_16999,N_14514,N_15246);
nor U17000 (N_17000,N_15155,N_15550);
nor U17001 (N_17001,N_15334,N_15690);
xor U17002 (N_17002,N_14151,N_14081);
or U17003 (N_17003,N_15028,N_14201);
or U17004 (N_17004,N_14889,N_14812);
and U17005 (N_17005,N_15474,N_15756);
and U17006 (N_17006,N_15697,N_15942);
or U17007 (N_17007,N_14707,N_14227);
or U17008 (N_17008,N_14674,N_15864);
and U17009 (N_17009,N_14950,N_15423);
nor U17010 (N_17010,N_14365,N_14457);
and U17011 (N_17011,N_15158,N_15623);
nand U17012 (N_17012,N_14851,N_15830);
and U17013 (N_17013,N_14513,N_14567);
xnor U17014 (N_17014,N_14612,N_15991);
and U17015 (N_17015,N_14466,N_15739);
nor U17016 (N_17016,N_14854,N_15252);
nand U17017 (N_17017,N_15026,N_15620);
and U17018 (N_17018,N_15706,N_14060);
or U17019 (N_17019,N_14127,N_15260);
or U17020 (N_17020,N_15603,N_14732);
xor U17021 (N_17021,N_15306,N_15455);
xor U17022 (N_17022,N_14437,N_15117);
nand U17023 (N_17023,N_15963,N_15616);
nand U17024 (N_17024,N_14008,N_14683);
xnor U17025 (N_17025,N_15976,N_15736);
xor U17026 (N_17026,N_14161,N_15032);
or U17027 (N_17027,N_15041,N_15672);
nand U17028 (N_17028,N_14530,N_15456);
xor U17029 (N_17029,N_14973,N_14535);
nand U17030 (N_17030,N_14149,N_15808);
xor U17031 (N_17031,N_15701,N_15353);
and U17032 (N_17032,N_15770,N_14658);
or U17033 (N_17033,N_14131,N_15856);
nand U17034 (N_17034,N_14383,N_15897);
nor U17035 (N_17035,N_14799,N_15546);
xnor U17036 (N_17036,N_14572,N_14310);
or U17037 (N_17037,N_14437,N_14652);
xor U17038 (N_17038,N_14163,N_15079);
and U17039 (N_17039,N_14885,N_15941);
and U17040 (N_17040,N_14724,N_14263);
nor U17041 (N_17041,N_14539,N_14150);
or U17042 (N_17042,N_14275,N_14863);
or U17043 (N_17043,N_14215,N_14071);
nor U17044 (N_17044,N_15168,N_15680);
and U17045 (N_17045,N_14772,N_15348);
xor U17046 (N_17046,N_15143,N_14515);
nand U17047 (N_17047,N_15906,N_15223);
and U17048 (N_17048,N_14507,N_15653);
and U17049 (N_17049,N_15958,N_14601);
nor U17050 (N_17050,N_14895,N_14460);
and U17051 (N_17051,N_14860,N_14792);
and U17052 (N_17052,N_14674,N_14429);
nor U17053 (N_17053,N_14081,N_15766);
nor U17054 (N_17054,N_14324,N_15754);
nand U17055 (N_17055,N_15921,N_14898);
xor U17056 (N_17056,N_14041,N_14225);
nor U17057 (N_17057,N_15720,N_15028);
or U17058 (N_17058,N_14778,N_15810);
or U17059 (N_17059,N_14561,N_15459);
or U17060 (N_17060,N_14793,N_14733);
nand U17061 (N_17061,N_15179,N_15753);
nand U17062 (N_17062,N_15371,N_14476);
or U17063 (N_17063,N_15887,N_15895);
or U17064 (N_17064,N_15908,N_15854);
nor U17065 (N_17065,N_15690,N_15970);
xor U17066 (N_17066,N_15594,N_15165);
xor U17067 (N_17067,N_14109,N_15065);
nand U17068 (N_17068,N_14080,N_14971);
nor U17069 (N_17069,N_14204,N_15356);
xor U17070 (N_17070,N_14530,N_14123);
nand U17071 (N_17071,N_15783,N_15457);
xnor U17072 (N_17072,N_15397,N_15372);
xor U17073 (N_17073,N_14444,N_14325);
and U17074 (N_17074,N_14710,N_14664);
and U17075 (N_17075,N_15095,N_15765);
or U17076 (N_17076,N_15692,N_15548);
nor U17077 (N_17077,N_14086,N_15218);
nand U17078 (N_17078,N_14869,N_14608);
and U17079 (N_17079,N_15108,N_15382);
or U17080 (N_17080,N_15294,N_15205);
or U17081 (N_17081,N_14827,N_14292);
nand U17082 (N_17082,N_14563,N_15252);
xnor U17083 (N_17083,N_15562,N_15910);
and U17084 (N_17084,N_15554,N_14574);
nor U17085 (N_17085,N_14880,N_15088);
nor U17086 (N_17086,N_14723,N_15909);
or U17087 (N_17087,N_14875,N_15046);
nand U17088 (N_17088,N_14738,N_15105);
nand U17089 (N_17089,N_14398,N_15970);
or U17090 (N_17090,N_15267,N_15713);
nand U17091 (N_17091,N_14475,N_15853);
nand U17092 (N_17092,N_14400,N_14016);
nand U17093 (N_17093,N_14740,N_14994);
xor U17094 (N_17094,N_14760,N_14589);
or U17095 (N_17095,N_15121,N_14392);
and U17096 (N_17096,N_14516,N_15401);
or U17097 (N_17097,N_15809,N_14246);
xnor U17098 (N_17098,N_15377,N_14802);
and U17099 (N_17099,N_15942,N_15887);
and U17100 (N_17100,N_15438,N_15305);
xor U17101 (N_17101,N_15309,N_15986);
or U17102 (N_17102,N_15882,N_14581);
xnor U17103 (N_17103,N_14055,N_14682);
xnor U17104 (N_17104,N_14142,N_14488);
xnor U17105 (N_17105,N_15516,N_14943);
or U17106 (N_17106,N_14120,N_15809);
xnor U17107 (N_17107,N_15959,N_14522);
nand U17108 (N_17108,N_15444,N_14908);
nor U17109 (N_17109,N_15992,N_15555);
xnor U17110 (N_17110,N_15123,N_15098);
xor U17111 (N_17111,N_15511,N_15294);
xnor U17112 (N_17112,N_15452,N_14133);
nand U17113 (N_17113,N_15317,N_15835);
nor U17114 (N_17114,N_14140,N_14639);
xor U17115 (N_17115,N_15688,N_14673);
and U17116 (N_17116,N_14077,N_14648);
or U17117 (N_17117,N_14297,N_14803);
nor U17118 (N_17118,N_15026,N_15181);
and U17119 (N_17119,N_14755,N_14403);
or U17120 (N_17120,N_15172,N_14062);
xor U17121 (N_17121,N_15134,N_14157);
or U17122 (N_17122,N_14452,N_15088);
nor U17123 (N_17123,N_14893,N_15650);
or U17124 (N_17124,N_14978,N_15579);
or U17125 (N_17125,N_15622,N_15514);
xor U17126 (N_17126,N_14852,N_14618);
nor U17127 (N_17127,N_15089,N_15352);
and U17128 (N_17128,N_14159,N_15824);
or U17129 (N_17129,N_14221,N_14339);
xnor U17130 (N_17130,N_14028,N_14008);
nor U17131 (N_17131,N_14874,N_14879);
nand U17132 (N_17132,N_15959,N_14489);
and U17133 (N_17133,N_14607,N_15442);
nor U17134 (N_17134,N_14363,N_15979);
or U17135 (N_17135,N_14273,N_14511);
xnor U17136 (N_17136,N_15175,N_15066);
or U17137 (N_17137,N_15943,N_15550);
xor U17138 (N_17138,N_15698,N_15909);
nor U17139 (N_17139,N_14398,N_14019);
nor U17140 (N_17140,N_15910,N_15524);
and U17141 (N_17141,N_14221,N_14074);
and U17142 (N_17142,N_15665,N_14974);
nor U17143 (N_17143,N_15447,N_14384);
or U17144 (N_17144,N_15267,N_15585);
and U17145 (N_17145,N_14747,N_15073);
and U17146 (N_17146,N_14525,N_15430);
nand U17147 (N_17147,N_15789,N_15991);
xnor U17148 (N_17148,N_14570,N_14284);
nand U17149 (N_17149,N_14573,N_15998);
nand U17150 (N_17150,N_14610,N_15267);
xnor U17151 (N_17151,N_15957,N_14307);
or U17152 (N_17152,N_14196,N_14889);
xnor U17153 (N_17153,N_14264,N_14365);
xnor U17154 (N_17154,N_14396,N_14110);
nor U17155 (N_17155,N_14179,N_15233);
nor U17156 (N_17156,N_15895,N_15751);
nand U17157 (N_17157,N_15617,N_15201);
nor U17158 (N_17158,N_14176,N_14539);
xor U17159 (N_17159,N_15602,N_15148);
and U17160 (N_17160,N_15136,N_14833);
xnor U17161 (N_17161,N_14108,N_14096);
or U17162 (N_17162,N_14892,N_15215);
xnor U17163 (N_17163,N_14003,N_15281);
xor U17164 (N_17164,N_14831,N_15044);
or U17165 (N_17165,N_14262,N_15067);
nand U17166 (N_17166,N_15392,N_15716);
nor U17167 (N_17167,N_15770,N_15116);
and U17168 (N_17168,N_15201,N_15697);
nor U17169 (N_17169,N_14343,N_15743);
nand U17170 (N_17170,N_15444,N_15079);
or U17171 (N_17171,N_15466,N_14490);
and U17172 (N_17172,N_15920,N_15191);
or U17173 (N_17173,N_14791,N_14063);
xor U17174 (N_17174,N_14850,N_15148);
or U17175 (N_17175,N_14999,N_14794);
nand U17176 (N_17176,N_14516,N_15476);
nand U17177 (N_17177,N_14766,N_14411);
and U17178 (N_17178,N_15944,N_14976);
nor U17179 (N_17179,N_15693,N_15665);
xnor U17180 (N_17180,N_14945,N_15222);
nand U17181 (N_17181,N_14736,N_15493);
or U17182 (N_17182,N_15242,N_15520);
nor U17183 (N_17183,N_14094,N_14140);
nor U17184 (N_17184,N_14632,N_14121);
nand U17185 (N_17185,N_14783,N_15413);
xnor U17186 (N_17186,N_15812,N_14395);
xor U17187 (N_17187,N_14472,N_15293);
and U17188 (N_17188,N_14200,N_15744);
and U17189 (N_17189,N_14915,N_14572);
nor U17190 (N_17190,N_14694,N_14164);
nor U17191 (N_17191,N_15525,N_15049);
xnor U17192 (N_17192,N_15442,N_15731);
and U17193 (N_17193,N_15636,N_15394);
nand U17194 (N_17194,N_15328,N_15127);
and U17195 (N_17195,N_14190,N_14524);
nand U17196 (N_17196,N_14898,N_15668);
or U17197 (N_17197,N_14553,N_15067);
nand U17198 (N_17198,N_15896,N_15847);
nor U17199 (N_17199,N_14787,N_15064);
xnor U17200 (N_17200,N_15719,N_14181);
or U17201 (N_17201,N_15901,N_15419);
nand U17202 (N_17202,N_14645,N_14070);
nor U17203 (N_17203,N_14686,N_14024);
nor U17204 (N_17204,N_15199,N_14134);
or U17205 (N_17205,N_14660,N_14652);
nand U17206 (N_17206,N_14174,N_14042);
nor U17207 (N_17207,N_15759,N_14930);
nor U17208 (N_17208,N_15825,N_14952);
or U17209 (N_17209,N_15153,N_14698);
and U17210 (N_17210,N_14298,N_14959);
and U17211 (N_17211,N_15742,N_15979);
and U17212 (N_17212,N_14943,N_15172);
xor U17213 (N_17213,N_15826,N_14793);
nand U17214 (N_17214,N_15894,N_14227);
nor U17215 (N_17215,N_14799,N_15708);
and U17216 (N_17216,N_14374,N_15609);
and U17217 (N_17217,N_15712,N_14455);
nor U17218 (N_17218,N_15582,N_15640);
xor U17219 (N_17219,N_14195,N_15277);
and U17220 (N_17220,N_15243,N_15702);
xnor U17221 (N_17221,N_15053,N_14025);
xnor U17222 (N_17222,N_14944,N_14089);
nor U17223 (N_17223,N_15386,N_15713);
or U17224 (N_17224,N_14636,N_14263);
nor U17225 (N_17225,N_14918,N_14443);
and U17226 (N_17226,N_14395,N_14688);
xor U17227 (N_17227,N_14214,N_14097);
nor U17228 (N_17228,N_15027,N_15689);
and U17229 (N_17229,N_15607,N_15621);
nand U17230 (N_17230,N_15672,N_15131);
or U17231 (N_17231,N_14157,N_15681);
and U17232 (N_17232,N_14588,N_15498);
xor U17233 (N_17233,N_14128,N_14751);
or U17234 (N_17234,N_14915,N_15092);
xor U17235 (N_17235,N_15227,N_14589);
nor U17236 (N_17236,N_15941,N_14104);
xnor U17237 (N_17237,N_14408,N_14830);
xor U17238 (N_17238,N_15691,N_15918);
nand U17239 (N_17239,N_15500,N_14515);
or U17240 (N_17240,N_15729,N_14724);
nor U17241 (N_17241,N_15175,N_15250);
nand U17242 (N_17242,N_15479,N_14057);
or U17243 (N_17243,N_15293,N_15665);
and U17244 (N_17244,N_14557,N_14076);
nand U17245 (N_17245,N_14227,N_14857);
xor U17246 (N_17246,N_14685,N_15274);
xor U17247 (N_17247,N_15607,N_14709);
or U17248 (N_17248,N_14256,N_14833);
nand U17249 (N_17249,N_15404,N_14918);
xnor U17250 (N_17250,N_14260,N_14083);
nor U17251 (N_17251,N_15838,N_14664);
nor U17252 (N_17252,N_14169,N_15257);
nor U17253 (N_17253,N_15403,N_15260);
nor U17254 (N_17254,N_14004,N_15868);
nand U17255 (N_17255,N_15404,N_14383);
nand U17256 (N_17256,N_14166,N_15499);
or U17257 (N_17257,N_15094,N_14640);
nor U17258 (N_17258,N_15264,N_15382);
nand U17259 (N_17259,N_14952,N_14080);
nor U17260 (N_17260,N_14069,N_15923);
xnor U17261 (N_17261,N_15836,N_15578);
xor U17262 (N_17262,N_14406,N_14945);
nor U17263 (N_17263,N_14270,N_15189);
or U17264 (N_17264,N_14001,N_15100);
or U17265 (N_17265,N_14265,N_14671);
and U17266 (N_17266,N_14174,N_14464);
nand U17267 (N_17267,N_15027,N_15165);
nor U17268 (N_17268,N_14911,N_14029);
xnor U17269 (N_17269,N_14208,N_15770);
xnor U17270 (N_17270,N_15264,N_15736);
and U17271 (N_17271,N_14022,N_15059);
nand U17272 (N_17272,N_14434,N_15581);
nor U17273 (N_17273,N_15957,N_15604);
or U17274 (N_17274,N_15081,N_14412);
or U17275 (N_17275,N_14077,N_15939);
xor U17276 (N_17276,N_15216,N_14568);
nor U17277 (N_17277,N_14679,N_14233);
nor U17278 (N_17278,N_14604,N_15294);
nor U17279 (N_17279,N_15237,N_14111);
nand U17280 (N_17280,N_15060,N_14697);
nand U17281 (N_17281,N_15481,N_14156);
or U17282 (N_17282,N_14193,N_14197);
and U17283 (N_17283,N_15646,N_15193);
nand U17284 (N_17284,N_14175,N_15445);
and U17285 (N_17285,N_15140,N_15292);
nor U17286 (N_17286,N_14742,N_14648);
xor U17287 (N_17287,N_14691,N_15228);
nor U17288 (N_17288,N_14151,N_14124);
xnor U17289 (N_17289,N_14328,N_14353);
nor U17290 (N_17290,N_15274,N_15793);
nor U17291 (N_17291,N_14770,N_14500);
or U17292 (N_17292,N_15951,N_15395);
nand U17293 (N_17293,N_14521,N_14350);
and U17294 (N_17294,N_15840,N_14759);
nand U17295 (N_17295,N_15522,N_14468);
xnor U17296 (N_17296,N_14846,N_15571);
nand U17297 (N_17297,N_14280,N_14840);
nand U17298 (N_17298,N_15111,N_15840);
xnor U17299 (N_17299,N_14689,N_15483);
or U17300 (N_17300,N_14043,N_14243);
and U17301 (N_17301,N_15355,N_15562);
and U17302 (N_17302,N_14124,N_15510);
nand U17303 (N_17303,N_15982,N_15339);
or U17304 (N_17304,N_15972,N_14010);
xor U17305 (N_17305,N_14062,N_14455);
nor U17306 (N_17306,N_14590,N_15415);
nand U17307 (N_17307,N_14498,N_14565);
and U17308 (N_17308,N_14293,N_15992);
and U17309 (N_17309,N_15211,N_15541);
nand U17310 (N_17310,N_14486,N_14518);
or U17311 (N_17311,N_15483,N_14581);
nand U17312 (N_17312,N_15505,N_14865);
or U17313 (N_17313,N_15015,N_15571);
nand U17314 (N_17314,N_14921,N_15900);
xnor U17315 (N_17315,N_15112,N_15902);
or U17316 (N_17316,N_14356,N_15653);
and U17317 (N_17317,N_14950,N_14475);
nor U17318 (N_17318,N_14685,N_15017);
or U17319 (N_17319,N_15501,N_15285);
and U17320 (N_17320,N_15589,N_14882);
xnor U17321 (N_17321,N_14183,N_15429);
and U17322 (N_17322,N_15462,N_14365);
xnor U17323 (N_17323,N_15110,N_15350);
nor U17324 (N_17324,N_15576,N_15558);
and U17325 (N_17325,N_15321,N_15729);
nand U17326 (N_17326,N_14876,N_15309);
or U17327 (N_17327,N_14287,N_15428);
nor U17328 (N_17328,N_15633,N_14659);
nand U17329 (N_17329,N_14017,N_14028);
or U17330 (N_17330,N_15393,N_15735);
xnor U17331 (N_17331,N_14082,N_14297);
nor U17332 (N_17332,N_14346,N_14373);
nand U17333 (N_17333,N_15715,N_15490);
nor U17334 (N_17334,N_15637,N_15934);
nor U17335 (N_17335,N_15413,N_14444);
nor U17336 (N_17336,N_14600,N_14768);
nor U17337 (N_17337,N_15841,N_14429);
xor U17338 (N_17338,N_15334,N_14470);
nand U17339 (N_17339,N_15864,N_15681);
nand U17340 (N_17340,N_15479,N_14436);
or U17341 (N_17341,N_14294,N_15012);
and U17342 (N_17342,N_14926,N_14498);
nor U17343 (N_17343,N_14640,N_14790);
and U17344 (N_17344,N_14394,N_15937);
and U17345 (N_17345,N_14374,N_15277);
nand U17346 (N_17346,N_14577,N_15850);
nor U17347 (N_17347,N_15836,N_14288);
nand U17348 (N_17348,N_14545,N_14993);
or U17349 (N_17349,N_15128,N_15802);
xor U17350 (N_17350,N_15519,N_15069);
or U17351 (N_17351,N_15467,N_14244);
xnor U17352 (N_17352,N_14615,N_15410);
xnor U17353 (N_17353,N_15217,N_15684);
or U17354 (N_17354,N_15175,N_14913);
and U17355 (N_17355,N_15725,N_15567);
nor U17356 (N_17356,N_14823,N_15470);
and U17357 (N_17357,N_14118,N_15146);
nor U17358 (N_17358,N_14968,N_15906);
or U17359 (N_17359,N_14463,N_14214);
xor U17360 (N_17360,N_15123,N_15990);
or U17361 (N_17361,N_14768,N_15313);
nor U17362 (N_17362,N_14464,N_15124);
and U17363 (N_17363,N_15271,N_15470);
nand U17364 (N_17364,N_14276,N_15497);
or U17365 (N_17365,N_14669,N_14004);
and U17366 (N_17366,N_15902,N_15194);
xnor U17367 (N_17367,N_14957,N_14511);
nor U17368 (N_17368,N_15974,N_14469);
and U17369 (N_17369,N_15123,N_15942);
nand U17370 (N_17370,N_14473,N_15015);
and U17371 (N_17371,N_15174,N_14414);
nand U17372 (N_17372,N_14193,N_14692);
nor U17373 (N_17373,N_14083,N_14048);
nand U17374 (N_17374,N_14139,N_14755);
or U17375 (N_17375,N_15160,N_14235);
nor U17376 (N_17376,N_14466,N_14800);
nand U17377 (N_17377,N_14985,N_15179);
and U17378 (N_17378,N_15783,N_15242);
and U17379 (N_17379,N_14495,N_14319);
nand U17380 (N_17380,N_14248,N_14510);
or U17381 (N_17381,N_14226,N_15589);
nand U17382 (N_17382,N_14914,N_14899);
or U17383 (N_17383,N_14238,N_14344);
or U17384 (N_17384,N_15667,N_14542);
nor U17385 (N_17385,N_15497,N_15588);
nor U17386 (N_17386,N_15723,N_15101);
or U17387 (N_17387,N_15459,N_14942);
xor U17388 (N_17388,N_15028,N_14446);
xnor U17389 (N_17389,N_14799,N_14707);
xnor U17390 (N_17390,N_14658,N_14396);
nor U17391 (N_17391,N_14743,N_14909);
nor U17392 (N_17392,N_15913,N_15502);
xnor U17393 (N_17393,N_15416,N_15497);
nor U17394 (N_17394,N_14291,N_15463);
nand U17395 (N_17395,N_14673,N_15614);
or U17396 (N_17396,N_14496,N_14574);
nand U17397 (N_17397,N_15213,N_15175);
nand U17398 (N_17398,N_15513,N_14915);
nor U17399 (N_17399,N_14496,N_14690);
nand U17400 (N_17400,N_15632,N_15056);
and U17401 (N_17401,N_14600,N_14666);
or U17402 (N_17402,N_14206,N_14999);
or U17403 (N_17403,N_15068,N_14006);
nand U17404 (N_17404,N_14595,N_15492);
xnor U17405 (N_17405,N_14436,N_15385);
nor U17406 (N_17406,N_15818,N_14684);
nor U17407 (N_17407,N_14913,N_15235);
nand U17408 (N_17408,N_15488,N_15837);
nor U17409 (N_17409,N_14088,N_14920);
or U17410 (N_17410,N_15391,N_14301);
or U17411 (N_17411,N_14525,N_14726);
and U17412 (N_17412,N_15991,N_14494);
or U17413 (N_17413,N_15082,N_14516);
xor U17414 (N_17414,N_15306,N_14005);
nand U17415 (N_17415,N_15171,N_14174);
xnor U17416 (N_17416,N_15581,N_14996);
xor U17417 (N_17417,N_15268,N_15397);
or U17418 (N_17418,N_14594,N_15435);
or U17419 (N_17419,N_15917,N_15621);
and U17420 (N_17420,N_15815,N_14561);
and U17421 (N_17421,N_15770,N_14787);
and U17422 (N_17422,N_14177,N_15599);
or U17423 (N_17423,N_15913,N_14223);
xnor U17424 (N_17424,N_15508,N_15219);
or U17425 (N_17425,N_14280,N_15567);
nand U17426 (N_17426,N_14457,N_14822);
nand U17427 (N_17427,N_14867,N_14818);
xor U17428 (N_17428,N_15340,N_15263);
or U17429 (N_17429,N_15173,N_15532);
or U17430 (N_17430,N_14352,N_15975);
xnor U17431 (N_17431,N_15715,N_15095);
nor U17432 (N_17432,N_15880,N_14922);
or U17433 (N_17433,N_15968,N_14805);
or U17434 (N_17434,N_14935,N_15133);
or U17435 (N_17435,N_14633,N_14936);
or U17436 (N_17436,N_14764,N_15000);
or U17437 (N_17437,N_14151,N_15334);
or U17438 (N_17438,N_14652,N_15487);
or U17439 (N_17439,N_14947,N_15589);
or U17440 (N_17440,N_15353,N_15136);
and U17441 (N_17441,N_14868,N_15549);
xnor U17442 (N_17442,N_15518,N_14526);
xor U17443 (N_17443,N_14346,N_15464);
or U17444 (N_17444,N_14524,N_14197);
or U17445 (N_17445,N_15703,N_15013);
xnor U17446 (N_17446,N_14390,N_15572);
and U17447 (N_17447,N_14174,N_15443);
xor U17448 (N_17448,N_15926,N_14672);
and U17449 (N_17449,N_14963,N_14603);
and U17450 (N_17450,N_14183,N_15865);
and U17451 (N_17451,N_14488,N_14227);
nand U17452 (N_17452,N_15510,N_14694);
xor U17453 (N_17453,N_14037,N_14284);
nor U17454 (N_17454,N_14748,N_15043);
nor U17455 (N_17455,N_15783,N_14274);
nand U17456 (N_17456,N_14338,N_15371);
nor U17457 (N_17457,N_14723,N_15203);
nor U17458 (N_17458,N_14042,N_15110);
nor U17459 (N_17459,N_14017,N_14394);
nand U17460 (N_17460,N_15432,N_15974);
nand U17461 (N_17461,N_15522,N_15766);
nor U17462 (N_17462,N_14207,N_14469);
nand U17463 (N_17463,N_14745,N_14530);
and U17464 (N_17464,N_15493,N_14755);
nor U17465 (N_17465,N_14696,N_15458);
nor U17466 (N_17466,N_14067,N_14866);
xnor U17467 (N_17467,N_14131,N_14509);
and U17468 (N_17468,N_15937,N_15192);
or U17469 (N_17469,N_15622,N_15262);
nor U17470 (N_17470,N_15190,N_15660);
nand U17471 (N_17471,N_15730,N_14679);
and U17472 (N_17472,N_15824,N_14821);
xor U17473 (N_17473,N_15128,N_14260);
nor U17474 (N_17474,N_14482,N_14234);
or U17475 (N_17475,N_15962,N_14660);
nand U17476 (N_17476,N_14056,N_14355);
nand U17477 (N_17477,N_15828,N_14863);
or U17478 (N_17478,N_14695,N_14401);
nor U17479 (N_17479,N_15704,N_15414);
xor U17480 (N_17480,N_15043,N_15136);
and U17481 (N_17481,N_15811,N_15447);
and U17482 (N_17482,N_14046,N_15129);
and U17483 (N_17483,N_15243,N_15937);
or U17484 (N_17484,N_15955,N_15286);
nand U17485 (N_17485,N_15278,N_15371);
and U17486 (N_17486,N_15854,N_15820);
or U17487 (N_17487,N_14849,N_14853);
nand U17488 (N_17488,N_14293,N_14520);
and U17489 (N_17489,N_14609,N_15139);
nand U17490 (N_17490,N_15022,N_14004);
and U17491 (N_17491,N_15178,N_14943);
nand U17492 (N_17492,N_14132,N_14158);
nor U17493 (N_17493,N_15267,N_15229);
nor U17494 (N_17494,N_15421,N_14450);
and U17495 (N_17495,N_15257,N_14822);
or U17496 (N_17496,N_15416,N_14159);
and U17497 (N_17497,N_14230,N_15816);
nor U17498 (N_17498,N_15186,N_15701);
or U17499 (N_17499,N_14628,N_15829);
and U17500 (N_17500,N_14875,N_14044);
xor U17501 (N_17501,N_15230,N_15702);
and U17502 (N_17502,N_15824,N_14117);
nand U17503 (N_17503,N_15987,N_15826);
nor U17504 (N_17504,N_14313,N_14227);
nand U17505 (N_17505,N_14286,N_15526);
or U17506 (N_17506,N_15784,N_14718);
xnor U17507 (N_17507,N_14635,N_15629);
and U17508 (N_17508,N_14075,N_15119);
nand U17509 (N_17509,N_14682,N_15498);
and U17510 (N_17510,N_15074,N_14082);
nand U17511 (N_17511,N_15584,N_14299);
nor U17512 (N_17512,N_15098,N_14853);
nor U17513 (N_17513,N_15494,N_15926);
nor U17514 (N_17514,N_14871,N_14613);
or U17515 (N_17515,N_14176,N_14579);
nor U17516 (N_17516,N_14417,N_14250);
nor U17517 (N_17517,N_15147,N_14050);
and U17518 (N_17518,N_14264,N_15741);
xor U17519 (N_17519,N_14869,N_14192);
nor U17520 (N_17520,N_14185,N_15020);
nor U17521 (N_17521,N_14735,N_14738);
nor U17522 (N_17522,N_14108,N_15952);
nor U17523 (N_17523,N_14831,N_14083);
nand U17524 (N_17524,N_14708,N_15190);
nand U17525 (N_17525,N_15301,N_14037);
nand U17526 (N_17526,N_15562,N_14798);
nor U17527 (N_17527,N_15509,N_14764);
or U17528 (N_17528,N_15188,N_15418);
nand U17529 (N_17529,N_15085,N_14406);
and U17530 (N_17530,N_15275,N_14958);
nor U17531 (N_17531,N_14124,N_14803);
xor U17532 (N_17532,N_14038,N_14238);
nand U17533 (N_17533,N_15471,N_15517);
and U17534 (N_17534,N_15670,N_15535);
xnor U17535 (N_17535,N_14719,N_14831);
and U17536 (N_17536,N_14925,N_15194);
and U17537 (N_17537,N_14380,N_14113);
nand U17538 (N_17538,N_15612,N_15994);
nand U17539 (N_17539,N_14837,N_14798);
or U17540 (N_17540,N_15404,N_15006);
xor U17541 (N_17541,N_15784,N_15481);
or U17542 (N_17542,N_15359,N_15157);
and U17543 (N_17543,N_14954,N_14664);
xnor U17544 (N_17544,N_14309,N_14340);
nand U17545 (N_17545,N_14155,N_14170);
nand U17546 (N_17546,N_15340,N_15686);
or U17547 (N_17547,N_15148,N_15532);
and U17548 (N_17548,N_14753,N_15378);
and U17549 (N_17549,N_15776,N_15235);
nand U17550 (N_17550,N_15905,N_15817);
or U17551 (N_17551,N_15513,N_15846);
and U17552 (N_17552,N_15632,N_14419);
nand U17553 (N_17553,N_14538,N_14271);
xnor U17554 (N_17554,N_15040,N_15404);
nand U17555 (N_17555,N_14739,N_15501);
nor U17556 (N_17556,N_15533,N_14077);
xnor U17557 (N_17557,N_15715,N_15390);
nand U17558 (N_17558,N_14565,N_14258);
nand U17559 (N_17559,N_15185,N_14526);
xor U17560 (N_17560,N_14320,N_15531);
or U17561 (N_17561,N_15774,N_15329);
nand U17562 (N_17562,N_14135,N_15949);
nand U17563 (N_17563,N_15066,N_14967);
or U17564 (N_17564,N_15217,N_15829);
nand U17565 (N_17565,N_14911,N_15067);
and U17566 (N_17566,N_14916,N_14012);
and U17567 (N_17567,N_15492,N_14778);
or U17568 (N_17568,N_15981,N_15737);
nor U17569 (N_17569,N_15292,N_14718);
xor U17570 (N_17570,N_15949,N_14230);
and U17571 (N_17571,N_15968,N_15137);
or U17572 (N_17572,N_15588,N_14145);
nor U17573 (N_17573,N_15326,N_14549);
xnor U17574 (N_17574,N_15660,N_14509);
nor U17575 (N_17575,N_15443,N_15035);
or U17576 (N_17576,N_14587,N_14879);
or U17577 (N_17577,N_14591,N_15620);
or U17578 (N_17578,N_14849,N_14846);
and U17579 (N_17579,N_14121,N_15912);
nand U17580 (N_17580,N_14000,N_14838);
or U17581 (N_17581,N_14927,N_15172);
or U17582 (N_17582,N_14357,N_15584);
and U17583 (N_17583,N_15420,N_15497);
nand U17584 (N_17584,N_14013,N_14394);
or U17585 (N_17585,N_14228,N_14975);
xnor U17586 (N_17586,N_14431,N_15340);
nor U17587 (N_17587,N_15955,N_14708);
or U17588 (N_17588,N_14040,N_14789);
and U17589 (N_17589,N_15467,N_15173);
and U17590 (N_17590,N_15833,N_14119);
xor U17591 (N_17591,N_15446,N_15527);
nor U17592 (N_17592,N_14111,N_15181);
or U17593 (N_17593,N_15729,N_14989);
xor U17594 (N_17594,N_15916,N_15880);
or U17595 (N_17595,N_14623,N_14384);
xor U17596 (N_17596,N_14386,N_14847);
or U17597 (N_17597,N_14375,N_15996);
xnor U17598 (N_17598,N_14730,N_15891);
xnor U17599 (N_17599,N_14677,N_15650);
and U17600 (N_17600,N_14532,N_15250);
xor U17601 (N_17601,N_14775,N_14148);
nor U17602 (N_17602,N_15186,N_14027);
or U17603 (N_17603,N_15461,N_14926);
or U17604 (N_17604,N_14128,N_14559);
xor U17605 (N_17605,N_15291,N_14553);
and U17606 (N_17606,N_15486,N_15190);
nand U17607 (N_17607,N_14091,N_15065);
nand U17608 (N_17608,N_14593,N_14955);
nor U17609 (N_17609,N_15854,N_14899);
xor U17610 (N_17610,N_14370,N_15374);
nand U17611 (N_17611,N_14922,N_14146);
and U17612 (N_17612,N_14635,N_15688);
or U17613 (N_17613,N_15670,N_14591);
and U17614 (N_17614,N_15119,N_15510);
xnor U17615 (N_17615,N_14349,N_14464);
or U17616 (N_17616,N_15688,N_14052);
nand U17617 (N_17617,N_15151,N_15026);
and U17618 (N_17618,N_15457,N_14403);
and U17619 (N_17619,N_14468,N_15696);
and U17620 (N_17620,N_14696,N_15231);
and U17621 (N_17621,N_14819,N_14199);
nor U17622 (N_17622,N_14383,N_15804);
xor U17623 (N_17623,N_15614,N_15415);
nor U17624 (N_17624,N_14130,N_15661);
nand U17625 (N_17625,N_15188,N_15149);
and U17626 (N_17626,N_14696,N_14851);
nand U17627 (N_17627,N_14796,N_14498);
nand U17628 (N_17628,N_15263,N_14400);
and U17629 (N_17629,N_15932,N_14658);
nor U17630 (N_17630,N_14610,N_15081);
and U17631 (N_17631,N_14343,N_15998);
nand U17632 (N_17632,N_14555,N_15576);
and U17633 (N_17633,N_14089,N_15591);
or U17634 (N_17634,N_15060,N_14755);
xor U17635 (N_17635,N_14821,N_14442);
nand U17636 (N_17636,N_14121,N_15518);
nor U17637 (N_17637,N_15217,N_15298);
or U17638 (N_17638,N_15626,N_14010);
or U17639 (N_17639,N_14935,N_15931);
nor U17640 (N_17640,N_14893,N_15128);
or U17641 (N_17641,N_15502,N_14261);
or U17642 (N_17642,N_14366,N_15194);
or U17643 (N_17643,N_15632,N_15316);
or U17644 (N_17644,N_14534,N_14360);
xnor U17645 (N_17645,N_15701,N_14597);
xor U17646 (N_17646,N_14427,N_15743);
nand U17647 (N_17647,N_15515,N_15446);
and U17648 (N_17648,N_15713,N_15920);
xor U17649 (N_17649,N_14591,N_15887);
nor U17650 (N_17650,N_14156,N_14671);
xor U17651 (N_17651,N_14148,N_14882);
nand U17652 (N_17652,N_15832,N_14620);
or U17653 (N_17653,N_14932,N_15610);
or U17654 (N_17654,N_14774,N_15245);
xor U17655 (N_17655,N_15825,N_15725);
or U17656 (N_17656,N_14374,N_15991);
xnor U17657 (N_17657,N_14118,N_14147);
nand U17658 (N_17658,N_15107,N_14210);
nor U17659 (N_17659,N_15903,N_15248);
nor U17660 (N_17660,N_14599,N_14075);
and U17661 (N_17661,N_15672,N_14376);
xor U17662 (N_17662,N_14802,N_14507);
or U17663 (N_17663,N_14228,N_14686);
or U17664 (N_17664,N_14485,N_15630);
and U17665 (N_17665,N_14199,N_15304);
xor U17666 (N_17666,N_15888,N_14092);
and U17667 (N_17667,N_15276,N_15568);
or U17668 (N_17668,N_15496,N_15212);
nand U17669 (N_17669,N_15540,N_15843);
nor U17670 (N_17670,N_15631,N_14037);
nand U17671 (N_17671,N_15831,N_15601);
nor U17672 (N_17672,N_14819,N_14142);
nand U17673 (N_17673,N_14713,N_15548);
nand U17674 (N_17674,N_15060,N_15144);
and U17675 (N_17675,N_15108,N_15069);
xnor U17676 (N_17676,N_15927,N_14771);
nor U17677 (N_17677,N_15114,N_15290);
nand U17678 (N_17678,N_14575,N_14549);
nor U17679 (N_17679,N_14580,N_15398);
xnor U17680 (N_17680,N_14536,N_15752);
nand U17681 (N_17681,N_15907,N_15750);
xnor U17682 (N_17682,N_14942,N_15082);
nand U17683 (N_17683,N_14612,N_15686);
nor U17684 (N_17684,N_14533,N_15413);
or U17685 (N_17685,N_14530,N_15758);
xnor U17686 (N_17686,N_15074,N_15257);
nor U17687 (N_17687,N_15468,N_14448);
and U17688 (N_17688,N_14766,N_14601);
and U17689 (N_17689,N_14617,N_15465);
and U17690 (N_17690,N_14437,N_14481);
xnor U17691 (N_17691,N_15390,N_15908);
nor U17692 (N_17692,N_14962,N_14243);
nor U17693 (N_17693,N_14759,N_15897);
nor U17694 (N_17694,N_14417,N_14508);
and U17695 (N_17695,N_15361,N_15969);
or U17696 (N_17696,N_14622,N_15656);
xor U17697 (N_17697,N_15640,N_15679);
nor U17698 (N_17698,N_15456,N_15237);
nor U17699 (N_17699,N_14522,N_14101);
xnor U17700 (N_17700,N_15805,N_14192);
or U17701 (N_17701,N_14443,N_14904);
or U17702 (N_17702,N_14461,N_14543);
or U17703 (N_17703,N_15256,N_15747);
and U17704 (N_17704,N_14076,N_15764);
nor U17705 (N_17705,N_14324,N_15391);
nor U17706 (N_17706,N_15176,N_14936);
nand U17707 (N_17707,N_14210,N_14292);
nor U17708 (N_17708,N_14638,N_14106);
xor U17709 (N_17709,N_15954,N_14394);
or U17710 (N_17710,N_14539,N_14653);
and U17711 (N_17711,N_15205,N_14299);
nor U17712 (N_17712,N_15067,N_14447);
nor U17713 (N_17713,N_14478,N_14057);
nand U17714 (N_17714,N_14152,N_14060);
and U17715 (N_17715,N_15941,N_15999);
nor U17716 (N_17716,N_14767,N_14022);
and U17717 (N_17717,N_14957,N_15405);
and U17718 (N_17718,N_15151,N_14558);
and U17719 (N_17719,N_14468,N_14476);
or U17720 (N_17720,N_15604,N_15295);
xor U17721 (N_17721,N_15592,N_14705);
and U17722 (N_17722,N_14397,N_14433);
xor U17723 (N_17723,N_15486,N_15340);
nor U17724 (N_17724,N_14730,N_14079);
nand U17725 (N_17725,N_15106,N_14161);
xor U17726 (N_17726,N_14428,N_14683);
and U17727 (N_17727,N_15559,N_15905);
or U17728 (N_17728,N_14070,N_15297);
xor U17729 (N_17729,N_14022,N_15611);
and U17730 (N_17730,N_14332,N_14963);
or U17731 (N_17731,N_14833,N_15088);
xnor U17732 (N_17732,N_14471,N_15519);
nand U17733 (N_17733,N_15709,N_15058);
xor U17734 (N_17734,N_15302,N_14727);
and U17735 (N_17735,N_14436,N_15690);
nand U17736 (N_17736,N_15406,N_15218);
nand U17737 (N_17737,N_15343,N_14524);
nand U17738 (N_17738,N_14116,N_14718);
and U17739 (N_17739,N_14438,N_15526);
nand U17740 (N_17740,N_15466,N_14743);
nor U17741 (N_17741,N_15374,N_14197);
or U17742 (N_17742,N_15231,N_15580);
or U17743 (N_17743,N_15104,N_14246);
or U17744 (N_17744,N_15634,N_14460);
nand U17745 (N_17745,N_14021,N_14697);
nor U17746 (N_17746,N_14638,N_15007);
xor U17747 (N_17747,N_14243,N_15118);
or U17748 (N_17748,N_14961,N_15812);
nor U17749 (N_17749,N_14419,N_14522);
xnor U17750 (N_17750,N_15919,N_15528);
or U17751 (N_17751,N_14661,N_14457);
and U17752 (N_17752,N_15093,N_15393);
nor U17753 (N_17753,N_14801,N_14796);
xor U17754 (N_17754,N_15605,N_15963);
and U17755 (N_17755,N_14009,N_14487);
and U17756 (N_17756,N_15263,N_15106);
or U17757 (N_17757,N_15334,N_15400);
xnor U17758 (N_17758,N_15772,N_15643);
or U17759 (N_17759,N_15342,N_14080);
and U17760 (N_17760,N_14881,N_14978);
or U17761 (N_17761,N_14326,N_15304);
and U17762 (N_17762,N_15941,N_15921);
nor U17763 (N_17763,N_14023,N_15310);
nor U17764 (N_17764,N_15045,N_15708);
nand U17765 (N_17765,N_14312,N_14848);
nand U17766 (N_17766,N_15126,N_14399);
nor U17767 (N_17767,N_14789,N_15142);
xor U17768 (N_17768,N_15348,N_14707);
nor U17769 (N_17769,N_14639,N_15839);
or U17770 (N_17770,N_14244,N_15465);
and U17771 (N_17771,N_14260,N_14688);
and U17772 (N_17772,N_14131,N_15374);
nand U17773 (N_17773,N_15845,N_14183);
or U17774 (N_17774,N_14652,N_14707);
and U17775 (N_17775,N_14105,N_15822);
nor U17776 (N_17776,N_15825,N_14805);
nor U17777 (N_17777,N_14915,N_14891);
xnor U17778 (N_17778,N_14659,N_15854);
or U17779 (N_17779,N_14559,N_14312);
or U17780 (N_17780,N_15111,N_14444);
and U17781 (N_17781,N_15305,N_14497);
or U17782 (N_17782,N_14481,N_15260);
xor U17783 (N_17783,N_14241,N_15427);
nand U17784 (N_17784,N_15913,N_15950);
and U17785 (N_17785,N_15651,N_14065);
nor U17786 (N_17786,N_14484,N_15050);
or U17787 (N_17787,N_14126,N_14511);
and U17788 (N_17788,N_14485,N_15610);
nand U17789 (N_17789,N_15651,N_14732);
or U17790 (N_17790,N_15559,N_15642);
or U17791 (N_17791,N_14180,N_15464);
xor U17792 (N_17792,N_14215,N_15442);
and U17793 (N_17793,N_14590,N_15109);
nor U17794 (N_17794,N_14781,N_15420);
and U17795 (N_17795,N_15331,N_15628);
nand U17796 (N_17796,N_14034,N_15051);
or U17797 (N_17797,N_15665,N_14084);
and U17798 (N_17798,N_14576,N_15748);
or U17799 (N_17799,N_14845,N_15884);
or U17800 (N_17800,N_15607,N_15427);
xnor U17801 (N_17801,N_15016,N_15787);
or U17802 (N_17802,N_14288,N_15362);
nor U17803 (N_17803,N_15907,N_14555);
or U17804 (N_17804,N_14646,N_14801);
nand U17805 (N_17805,N_14373,N_14875);
or U17806 (N_17806,N_14738,N_15410);
and U17807 (N_17807,N_14556,N_15046);
nand U17808 (N_17808,N_15681,N_14910);
nor U17809 (N_17809,N_14464,N_15278);
nor U17810 (N_17810,N_14359,N_15741);
nor U17811 (N_17811,N_15666,N_15251);
nor U17812 (N_17812,N_15335,N_14374);
or U17813 (N_17813,N_14507,N_15568);
and U17814 (N_17814,N_14368,N_15998);
nand U17815 (N_17815,N_15517,N_15484);
xor U17816 (N_17816,N_14760,N_14146);
xor U17817 (N_17817,N_14421,N_15737);
xnor U17818 (N_17818,N_14462,N_15381);
nand U17819 (N_17819,N_15005,N_15912);
xnor U17820 (N_17820,N_14037,N_15747);
or U17821 (N_17821,N_14993,N_15826);
nor U17822 (N_17822,N_14703,N_14207);
nor U17823 (N_17823,N_15778,N_14584);
nor U17824 (N_17824,N_15080,N_14901);
or U17825 (N_17825,N_15594,N_14510);
xnor U17826 (N_17826,N_15765,N_14585);
nor U17827 (N_17827,N_15998,N_14844);
nand U17828 (N_17828,N_14381,N_15345);
xor U17829 (N_17829,N_15420,N_14771);
nor U17830 (N_17830,N_15320,N_15570);
and U17831 (N_17831,N_15614,N_15046);
xor U17832 (N_17832,N_14675,N_14093);
nor U17833 (N_17833,N_14749,N_14600);
or U17834 (N_17834,N_14162,N_14395);
nand U17835 (N_17835,N_15108,N_14787);
nor U17836 (N_17836,N_14960,N_15450);
xnor U17837 (N_17837,N_14239,N_14223);
xnor U17838 (N_17838,N_15506,N_14435);
or U17839 (N_17839,N_15097,N_15362);
or U17840 (N_17840,N_14185,N_14391);
or U17841 (N_17841,N_15179,N_15976);
nand U17842 (N_17842,N_15934,N_15457);
or U17843 (N_17843,N_14204,N_14881);
or U17844 (N_17844,N_14015,N_15012);
or U17845 (N_17845,N_15260,N_15671);
and U17846 (N_17846,N_15490,N_15708);
and U17847 (N_17847,N_15897,N_14548);
nor U17848 (N_17848,N_14604,N_15242);
and U17849 (N_17849,N_15890,N_14784);
nor U17850 (N_17850,N_14786,N_14587);
or U17851 (N_17851,N_14584,N_14439);
nand U17852 (N_17852,N_14911,N_14872);
xor U17853 (N_17853,N_14046,N_14083);
and U17854 (N_17854,N_15111,N_14602);
and U17855 (N_17855,N_14232,N_15861);
nor U17856 (N_17856,N_15349,N_14361);
xor U17857 (N_17857,N_14076,N_15688);
or U17858 (N_17858,N_14210,N_15607);
or U17859 (N_17859,N_14475,N_14325);
xnor U17860 (N_17860,N_14427,N_15436);
xor U17861 (N_17861,N_14098,N_14500);
xor U17862 (N_17862,N_15115,N_14737);
and U17863 (N_17863,N_15085,N_14306);
and U17864 (N_17864,N_14860,N_14033);
xor U17865 (N_17865,N_15714,N_14064);
or U17866 (N_17866,N_14149,N_15855);
and U17867 (N_17867,N_14674,N_15493);
xnor U17868 (N_17868,N_15260,N_14090);
nand U17869 (N_17869,N_14736,N_14396);
xor U17870 (N_17870,N_14148,N_14600);
xor U17871 (N_17871,N_14266,N_15599);
nor U17872 (N_17872,N_14906,N_14587);
or U17873 (N_17873,N_14360,N_14177);
and U17874 (N_17874,N_14239,N_15771);
xor U17875 (N_17875,N_15990,N_14981);
nor U17876 (N_17876,N_15553,N_15811);
nand U17877 (N_17877,N_14394,N_14554);
or U17878 (N_17878,N_15456,N_14396);
and U17879 (N_17879,N_15732,N_15006);
xnor U17880 (N_17880,N_15407,N_14106);
nor U17881 (N_17881,N_14061,N_15216);
nand U17882 (N_17882,N_14218,N_14588);
and U17883 (N_17883,N_15902,N_14716);
xor U17884 (N_17884,N_14811,N_14326);
nor U17885 (N_17885,N_15106,N_14398);
nor U17886 (N_17886,N_14397,N_14812);
nand U17887 (N_17887,N_15018,N_15799);
or U17888 (N_17888,N_15934,N_15075);
nor U17889 (N_17889,N_14283,N_15936);
xnor U17890 (N_17890,N_15877,N_14666);
nand U17891 (N_17891,N_14651,N_14052);
nand U17892 (N_17892,N_15980,N_14801);
xor U17893 (N_17893,N_15395,N_14878);
and U17894 (N_17894,N_15945,N_15421);
nand U17895 (N_17895,N_15234,N_14838);
nor U17896 (N_17896,N_15421,N_14464);
and U17897 (N_17897,N_14650,N_14832);
nand U17898 (N_17898,N_14368,N_14477);
nor U17899 (N_17899,N_14134,N_14173);
or U17900 (N_17900,N_14889,N_15331);
or U17901 (N_17901,N_14009,N_14871);
and U17902 (N_17902,N_15702,N_15597);
nor U17903 (N_17903,N_14300,N_14046);
and U17904 (N_17904,N_14870,N_15995);
and U17905 (N_17905,N_14291,N_14016);
and U17906 (N_17906,N_15547,N_15786);
nand U17907 (N_17907,N_14404,N_14768);
and U17908 (N_17908,N_15163,N_15877);
xnor U17909 (N_17909,N_15904,N_14467);
nand U17910 (N_17910,N_15875,N_14452);
nor U17911 (N_17911,N_14730,N_15811);
xor U17912 (N_17912,N_14094,N_15623);
or U17913 (N_17913,N_15348,N_15589);
nand U17914 (N_17914,N_14677,N_15161);
xnor U17915 (N_17915,N_15232,N_14266);
and U17916 (N_17916,N_14480,N_14231);
or U17917 (N_17917,N_15772,N_15235);
nor U17918 (N_17918,N_15101,N_15277);
and U17919 (N_17919,N_15651,N_15680);
and U17920 (N_17920,N_15633,N_14104);
and U17921 (N_17921,N_15332,N_15121);
and U17922 (N_17922,N_14478,N_14520);
nand U17923 (N_17923,N_14215,N_15399);
xnor U17924 (N_17924,N_15130,N_15302);
and U17925 (N_17925,N_14788,N_14150);
or U17926 (N_17926,N_14074,N_14216);
xor U17927 (N_17927,N_14921,N_14564);
or U17928 (N_17928,N_15230,N_14143);
nor U17929 (N_17929,N_15468,N_15566);
or U17930 (N_17930,N_15689,N_15628);
or U17931 (N_17931,N_15301,N_15624);
nor U17932 (N_17932,N_14262,N_15399);
nand U17933 (N_17933,N_15137,N_15825);
nand U17934 (N_17934,N_15179,N_15820);
and U17935 (N_17935,N_15383,N_15750);
or U17936 (N_17936,N_14324,N_15331);
and U17937 (N_17937,N_14222,N_15207);
and U17938 (N_17938,N_15949,N_15146);
or U17939 (N_17939,N_15761,N_15411);
nor U17940 (N_17940,N_15507,N_15936);
nand U17941 (N_17941,N_15097,N_15840);
and U17942 (N_17942,N_14209,N_14139);
nor U17943 (N_17943,N_14782,N_14312);
or U17944 (N_17944,N_15039,N_15976);
nor U17945 (N_17945,N_14018,N_15633);
xnor U17946 (N_17946,N_15937,N_15586);
nand U17947 (N_17947,N_14826,N_14811);
xnor U17948 (N_17948,N_15347,N_14910);
nor U17949 (N_17949,N_15646,N_15865);
nor U17950 (N_17950,N_15667,N_14259);
nand U17951 (N_17951,N_14002,N_14888);
nor U17952 (N_17952,N_15463,N_15792);
or U17953 (N_17953,N_14952,N_14393);
nand U17954 (N_17954,N_15988,N_15322);
and U17955 (N_17955,N_15517,N_14794);
xor U17956 (N_17956,N_15449,N_14254);
xor U17957 (N_17957,N_14173,N_14423);
xor U17958 (N_17958,N_15335,N_15144);
or U17959 (N_17959,N_15398,N_14145);
nand U17960 (N_17960,N_15297,N_14738);
xor U17961 (N_17961,N_14062,N_14667);
nor U17962 (N_17962,N_14281,N_15250);
nor U17963 (N_17963,N_15949,N_14388);
nor U17964 (N_17964,N_15993,N_14529);
nor U17965 (N_17965,N_15808,N_14553);
and U17966 (N_17966,N_15163,N_14161);
or U17967 (N_17967,N_14158,N_15704);
nand U17968 (N_17968,N_14825,N_14383);
xnor U17969 (N_17969,N_14704,N_14203);
nor U17970 (N_17970,N_15139,N_15582);
or U17971 (N_17971,N_15337,N_15631);
xor U17972 (N_17972,N_15524,N_15022);
or U17973 (N_17973,N_15833,N_15381);
nand U17974 (N_17974,N_14380,N_14594);
and U17975 (N_17975,N_15273,N_14515);
and U17976 (N_17976,N_15559,N_15142);
nand U17977 (N_17977,N_14640,N_14510);
xor U17978 (N_17978,N_14867,N_15296);
xnor U17979 (N_17979,N_15144,N_15653);
nand U17980 (N_17980,N_14432,N_15750);
nand U17981 (N_17981,N_15331,N_15618);
nand U17982 (N_17982,N_15067,N_15663);
xnor U17983 (N_17983,N_14943,N_15379);
xnor U17984 (N_17984,N_15050,N_14501);
and U17985 (N_17985,N_14450,N_14335);
or U17986 (N_17986,N_15870,N_15900);
xor U17987 (N_17987,N_14733,N_15065);
xnor U17988 (N_17988,N_15732,N_15474);
xor U17989 (N_17989,N_15483,N_14087);
xnor U17990 (N_17990,N_14533,N_14556);
nor U17991 (N_17991,N_14760,N_15502);
nor U17992 (N_17992,N_15761,N_14637);
nor U17993 (N_17993,N_14989,N_14284);
nor U17994 (N_17994,N_14936,N_14224);
xnor U17995 (N_17995,N_15687,N_15997);
nor U17996 (N_17996,N_15240,N_15362);
and U17997 (N_17997,N_14642,N_15513);
or U17998 (N_17998,N_15662,N_14193);
or U17999 (N_17999,N_14799,N_14889);
and U18000 (N_18000,N_17549,N_17151);
xor U18001 (N_18001,N_16917,N_17082);
nor U18002 (N_18002,N_17351,N_17315);
xnor U18003 (N_18003,N_16536,N_16648);
and U18004 (N_18004,N_17334,N_17579);
and U18005 (N_18005,N_17058,N_17123);
or U18006 (N_18006,N_16188,N_16570);
xnor U18007 (N_18007,N_16098,N_17721);
nor U18008 (N_18008,N_17087,N_16320);
or U18009 (N_18009,N_17956,N_16706);
nand U18010 (N_18010,N_17968,N_17517);
nor U18011 (N_18011,N_16768,N_16685);
xor U18012 (N_18012,N_17659,N_17905);
nand U18013 (N_18013,N_16093,N_16091);
or U18014 (N_18014,N_17491,N_16013);
and U18015 (N_18015,N_17642,N_16951);
nand U18016 (N_18016,N_16425,N_16177);
nor U18017 (N_18017,N_16781,N_16112);
and U18018 (N_18018,N_16046,N_16563);
xnor U18019 (N_18019,N_17568,N_16383);
or U18020 (N_18020,N_17886,N_16861);
nor U18021 (N_18021,N_17432,N_17969);
nor U18022 (N_18022,N_17394,N_17006);
nor U18023 (N_18023,N_17373,N_17484);
and U18024 (N_18024,N_17786,N_16345);
nor U18025 (N_18025,N_16612,N_16272);
and U18026 (N_18026,N_16457,N_16025);
nor U18027 (N_18027,N_17388,N_17486);
nand U18028 (N_18028,N_16749,N_17652);
xor U18029 (N_18029,N_17881,N_16171);
nor U18030 (N_18030,N_17530,N_16634);
nor U18031 (N_18031,N_16059,N_16035);
xor U18032 (N_18032,N_17555,N_17331);
nand U18033 (N_18033,N_16722,N_17272);
nor U18034 (N_18034,N_16762,N_17858);
or U18035 (N_18035,N_17892,N_17092);
nor U18036 (N_18036,N_16974,N_17931);
xor U18037 (N_18037,N_17333,N_17499);
or U18038 (N_18038,N_17975,N_16387);
and U18039 (N_18039,N_17026,N_16018);
and U18040 (N_18040,N_16785,N_16080);
nand U18041 (N_18041,N_17241,N_16022);
and U18042 (N_18042,N_16438,N_16089);
nand U18043 (N_18043,N_17581,N_16693);
xnor U18044 (N_18044,N_16099,N_17984);
or U18045 (N_18045,N_16740,N_16359);
xnor U18046 (N_18046,N_16194,N_17698);
or U18047 (N_18047,N_17164,N_17749);
and U18048 (N_18048,N_16114,N_16213);
and U18049 (N_18049,N_16637,N_16314);
or U18050 (N_18050,N_17547,N_16560);
nand U18051 (N_18051,N_16829,N_16006);
xnor U18052 (N_18052,N_17622,N_17165);
and U18053 (N_18053,N_16282,N_16190);
and U18054 (N_18054,N_17426,N_17929);
nand U18055 (N_18055,N_16849,N_17071);
and U18056 (N_18056,N_17500,N_16931);
and U18057 (N_18057,N_16632,N_17531);
nand U18058 (N_18058,N_17512,N_17002);
or U18059 (N_18059,N_17270,N_16290);
nand U18060 (N_18060,N_16330,N_16718);
nor U18061 (N_18061,N_17212,N_17306);
nor U18062 (N_18062,N_16423,N_16441);
xor U18063 (N_18063,N_16057,N_16586);
nand U18064 (N_18064,N_16010,N_17717);
nor U18065 (N_18065,N_17086,N_17494);
nand U18066 (N_18066,N_16890,N_17247);
nor U18067 (N_18067,N_17218,N_16110);
xor U18068 (N_18068,N_16280,N_17941);
and U18069 (N_18069,N_17601,N_16253);
nor U18070 (N_18070,N_16831,N_16975);
nor U18071 (N_18071,N_17224,N_16809);
nand U18072 (N_18072,N_17016,N_17485);
or U18073 (N_18073,N_16381,N_17391);
and U18074 (N_18074,N_17636,N_17940);
or U18075 (N_18075,N_17299,N_16716);
xor U18076 (N_18076,N_16893,N_16606);
xor U18077 (N_18077,N_16262,N_17365);
and U18078 (N_18078,N_17758,N_17357);
or U18079 (N_18079,N_16851,N_16689);
or U18080 (N_18080,N_16588,N_16494);
xnor U18081 (N_18081,N_16406,N_17310);
nand U18082 (N_18082,N_16531,N_17945);
nand U18083 (N_18083,N_16147,N_17809);
xnor U18084 (N_18084,N_17837,N_17609);
nor U18085 (N_18085,N_16968,N_16552);
nor U18086 (N_18086,N_17489,N_17671);
xor U18087 (N_18087,N_16357,N_17267);
and U18088 (N_18088,N_17197,N_17669);
nor U18089 (N_18089,N_17480,N_16187);
xor U18090 (N_18090,N_16132,N_17222);
nor U18091 (N_18091,N_16976,N_16780);
or U18092 (N_18092,N_17187,N_16611);
and U18093 (N_18093,N_17115,N_16503);
nor U18094 (N_18094,N_16125,N_17116);
or U18095 (N_18095,N_16230,N_16541);
and U18096 (N_18096,N_16720,N_16141);
or U18097 (N_18097,N_16196,N_16622);
nor U18098 (N_18098,N_16602,N_16452);
xnor U18099 (N_18099,N_17126,N_16555);
nand U18100 (N_18100,N_17204,N_16767);
nor U18101 (N_18101,N_16614,N_17346);
and U18102 (N_18102,N_16240,N_17577);
nor U18103 (N_18103,N_16300,N_17600);
xor U18104 (N_18104,N_17050,N_16859);
nand U18105 (N_18105,N_16769,N_17643);
nor U18106 (N_18106,N_17979,N_17064);
nand U18107 (N_18107,N_17768,N_17751);
and U18108 (N_18108,N_17487,N_16543);
or U18109 (N_18109,N_16542,N_16286);
xnor U18110 (N_18110,N_17295,N_17850);
nor U18111 (N_18111,N_16987,N_16942);
and U18112 (N_18112,N_16398,N_16283);
xnor U18113 (N_18113,N_17313,N_16327);
xnor U18114 (N_18114,N_16812,N_17043);
nor U18115 (N_18115,N_17830,N_17580);
xnor U18116 (N_18116,N_17651,N_16770);
xor U18117 (N_18117,N_16549,N_16910);
and U18118 (N_18118,N_17863,N_16579);
and U18119 (N_18119,N_16894,N_16468);
xnor U18120 (N_18120,N_16649,N_17475);
or U18121 (N_18121,N_16391,N_17469);
nand U18122 (N_18122,N_17720,N_16002);
and U18123 (N_18123,N_16538,N_16958);
and U18124 (N_18124,N_16568,N_17181);
nand U18125 (N_18125,N_16003,N_16094);
nor U18126 (N_18126,N_16318,N_17390);
and U18127 (N_18127,N_16410,N_16642);
xor U18128 (N_18128,N_17702,N_17067);
or U18129 (N_18129,N_16741,N_17807);
xor U18130 (N_18130,N_16683,N_17178);
xor U18131 (N_18131,N_17788,N_16673);
and U18132 (N_18132,N_16823,N_16313);
xor U18133 (N_18133,N_16402,N_17081);
nand U18134 (N_18134,N_17845,N_17149);
and U18135 (N_18135,N_17454,N_16553);
or U18136 (N_18136,N_16260,N_17019);
or U18137 (N_18137,N_16412,N_17121);
nand U18138 (N_18138,N_17102,N_17311);
nor U18139 (N_18139,N_16090,N_16507);
nand U18140 (N_18140,N_17550,N_16928);
and U18141 (N_18141,N_17192,N_17632);
nand U18142 (N_18142,N_17034,N_16226);
nor U18143 (N_18143,N_17157,N_17705);
and U18144 (N_18144,N_16984,N_17562);
or U18145 (N_18145,N_17833,N_17235);
and U18146 (N_18146,N_16498,N_16730);
and U18147 (N_18147,N_16615,N_16192);
nor U18148 (N_18148,N_16523,N_16078);
nor U18149 (N_18149,N_17456,N_17857);
xor U18150 (N_18150,N_16103,N_17183);
nand U18151 (N_18151,N_16651,N_16437);
and U18152 (N_18152,N_17118,N_16454);
nor U18153 (N_18153,N_16252,N_17701);
xnor U18154 (N_18154,N_16800,N_17106);
nor U18155 (N_18155,N_17629,N_17281);
nand U18156 (N_18156,N_17173,N_17817);
or U18157 (N_18157,N_16058,N_16775);
or U18158 (N_18158,N_16645,N_17099);
xnor U18159 (N_18159,N_17909,N_16191);
and U18160 (N_18160,N_16932,N_17777);
and U18161 (N_18161,N_16004,N_17022);
and U18162 (N_18162,N_16640,N_17784);
and U18163 (N_18163,N_16265,N_16604);
or U18164 (N_18164,N_16447,N_17997);
nor U18165 (N_18165,N_16639,N_17757);
and U18166 (N_18166,N_16550,N_16569);
or U18167 (N_18167,N_16742,N_16040);
and U18168 (N_18168,N_17623,N_16599);
or U18169 (N_18169,N_16895,N_16212);
and U18170 (N_18170,N_16126,N_17927);
or U18171 (N_18171,N_17389,N_17190);
and U18172 (N_18172,N_16765,N_16348);
xnor U18173 (N_18173,N_16519,N_16292);
or U18174 (N_18174,N_17936,N_17482);
xnor U18175 (N_18175,N_16424,N_17774);
or U18176 (N_18176,N_16941,N_16053);
or U18177 (N_18177,N_16295,N_17011);
nand U18178 (N_18178,N_16178,N_16514);
nand U18179 (N_18179,N_17298,N_16723);
nand U18180 (N_18180,N_17048,N_16774);
or U18181 (N_18181,N_17505,N_16909);
or U18182 (N_18182,N_17556,N_17185);
xor U18183 (N_18183,N_16308,N_17041);
nand U18184 (N_18184,N_17551,N_16624);
nor U18185 (N_18185,N_17226,N_17981);
and U18186 (N_18186,N_17410,N_16060);
nor U18187 (N_18187,N_16985,N_16826);
or U18188 (N_18188,N_16729,N_16376);
nand U18189 (N_18189,N_16021,N_16745);
nor U18190 (N_18190,N_16778,N_16176);
nand U18191 (N_18191,N_17603,N_17473);
xor U18192 (N_18192,N_17982,N_16956);
nand U18193 (N_18193,N_17278,N_16486);
and U18194 (N_18194,N_16827,N_17534);
nand U18195 (N_18195,N_16241,N_17887);
and U18196 (N_18196,N_16900,N_17209);
and U18197 (N_18197,N_17619,N_17096);
or U18198 (N_18198,N_17266,N_16635);
nor U18199 (N_18199,N_16015,N_17742);
xnor U18200 (N_18200,N_16458,N_17282);
and U18201 (N_18201,N_17472,N_16734);
nand U18202 (N_18202,N_17498,N_17253);
nand U18203 (N_18203,N_17347,N_17465);
and U18204 (N_18204,N_17894,N_16721);
or U18205 (N_18205,N_16118,N_17668);
and U18206 (N_18206,N_16166,N_16480);
or U18207 (N_18207,N_17177,N_17436);
and U18208 (N_18208,N_17591,N_17802);
nand U18209 (N_18209,N_17220,N_17162);
xor U18210 (N_18210,N_16150,N_16613);
xnor U18211 (N_18211,N_16964,N_17934);
nand U18212 (N_18212,N_17951,N_16940);
and U18213 (N_18213,N_17640,N_17663);
and U18214 (N_18214,N_17535,N_17678);
xor U18215 (N_18215,N_17841,N_16001);
nor U18216 (N_18216,N_16411,N_16955);
or U18217 (N_18217,N_17168,N_17312);
nand U18218 (N_18218,N_16317,N_17359);
xnor U18219 (N_18219,N_17888,N_17345);
or U18220 (N_18220,N_16807,N_16527);
or U18221 (N_18221,N_16771,N_16609);
or U18222 (N_18222,N_16218,N_16083);
or U18223 (N_18223,N_16914,N_16596);
xor U18224 (N_18224,N_17477,N_16845);
nor U18225 (N_18225,N_16195,N_17964);
nand U18226 (N_18226,N_16735,N_17854);
or U18227 (N_18227,N_16291,N_16878);
xor U18228 (N_18228,N_16165,N_16456);
nor U18229 (N_18229,N_16788,N_16705);
xor U18230 (N_18230,N_17908,N_16920);
xnor U18231 (N_18231,N_17324,N_16972);
nand U18232 (N_18232,N_16344,N_16045);
nor U18233 (N_18233,N_17152,N_16268);
nor U18234 (N_18234,N_16281,N_17385);
nor U18235 (N_18235,N_17458,N_17166);
nand U18236 (N_18236,N_16202,N_16752);
and U18237 (N_18237,N_17319,N_16173);
xnor U18238 (N_18238,N_17593,N_16853);
nand U18239 (N_18239,N_17508,N_16312);
or U18240 (N_18240,N_17649,N_17821);
nand U18241 (N_18241,N_17061,N_17153);
or U18242 (N_18242,N_16016,N_17748);
or U18243 (N_18243,N_17844,N_16136);
nand U18244 (N_18244,N_17504,N_17100);
xor U18245 (N_18245,N_17617,N_16353);
or U18246 (N_18246,N_17033,N_16911);
xor U18247 (N_18247,N_17793,N_17262);
xnor U18248 (N_18248,N_17925,N_16181);
nand U18249 (N_18249,N_16279,N_17159);
nor U18250 (N_18250,N_17348,N_17978);
xnor U18251 (N_18251,N_16821,N_16075);
xor U18252 (N_18252,N_16855,N_16032);
xnor U18253 (N_18253,N_17873,N_16031);
and U18254 (N_18254,N_16062,N_17274);
or U18255 (N_18255,N_17570,N_16760);
nor U18256 (N_18256,N_16077,N_17805);
or U18257 (N_18257,N_17259,N_17077);
nand U18258 (N_18258,N_17406,N_17397);
or U18259 (N_18259,N_17912,N_17367);
nand U18260 (N_18260,N_17297,N_17852);
xor U18261 (N_18261,N_16284,N_16990);
nand U18262 (N_18262,N_17571,N_16336);
or U18263 (N_18263,N_17032,N_17878);
nand U18264 (N_18264,N_16200,N_16786);
nor U18265 (N_18265,N_16688,N_17003);
or U18266 (N_18266,N_16419,N_16051);
and U18267 (N_18267,N_16309,N_16847);
or U18268 (N_18268,N_17957,N_17434);
nor U18269 (N_18269,N_16816,N_17386);
and U18270 (N_18270,N_17366,N_16631);
nand U18271 (N_18271,N_17248,N_16205);
nand U18272 (N_18272,N_17587,N_17239);
or U18273 (N_18273,N_16794,N_17765);
or U18274 (N_18274,N_16719,N_16048);
and U18275 (N_18275,N_16652,N_17402);
nand U18276 (N_18276,N_17725,N_17735);
nor U18277 (N_18277,N_17815,N_16085);
and U18278 (N_18278,N_16506,N_17599);
and U18279 (N_18279,N_17690,N_16669);
and U18280 (N_18280,N_17935,N_17287);
nor U18281 (N_18281,N_17814,N_17094);
xnor U18282 (N_18282,N_17740,N_16427);
xnor U18283 (N_18283,N_17417,N_16843);
nand U18284 (N_18284,N_17481,N_17378);
and U18285 (N_18285,N_17303,N_16872);
or U18286 (N_18286,N_16332,N_17136);
and U18287 (N_18287,N_17362,N_16009);
nand U18288 (N_18288,N_17179,N_17163);
nand U18289 (N_18289,N_16977,N_16193);
xor U18290 (N_18290,N_16271,N_16540);
nand U18291 (N_18291,N_16127,N_16222);
and U18292 (N_18292,N_16228,N_16203);
xor U18293 (N_18293,N_16483,N_17066);
or U18294 (N_18294,N_17588,N_16619);
xnor U18295 (N_18295,N_17503,N_16758);
or U18296 (N_18296,N_16180,N_17686);
nor U18297 (N_18297,N_17810,N_16727);
nor U18298 (N_18298,N_17679,N_17342);
xnor U18299 (N_18299,N_17670,N_17418);
nor U18300 (N_18300,N_17132,N_16443);
and U18301 (N_18301,N_17114,N_17618);
nor U18302 (N_18302,N_16838,N_16858);
or U18303 (N_18303,N_16516,N_17200);
or U18304 (N_18304,N_16802,N_17021);
nor U18305 (N_18305,N_16469,N_16736);
xnor U18306 (N_18306,N_16938,N_17730);
nand U18307 (N_18307,N_17488,N_17910);
nor U18308 (N_18308,N_17953,N_17990);
nand U18309 (N_18309,N_16375,N_17903);
or U18310 (N_18310,N_16636,N_16577);
and U18311 (N_18311,N_17037,N_17523);
or U18312 (N_18312,N_17608,N_17943);
nand U18313 (N_18313,N_17884,N_17620);
nand U18314 (N_18314,N_16160,N_17685);
or U18315 (N_18315,N_16811,N_17726);
or U18316 (N_18316,N_17741,N_17724);
nor U18317 (N_18317,N_17921,N_17464);
xor U18318 (N_18318,N_16369,N_16813);
nand U18319 (N_18319,N_16933,N_16607);
nor U18320 (N_18320,N_17545,N_17352);
or U18321 (N_18321,N_16436,N_17400);
nand U18322 (N_18322,N_17667,N_17231);
and U18323 (N_18323,N_16426,N_16902);
xor U18324 (N_18324,N_17137,N_17761);
nor U18325 (N_18325,N_17072,N_17614);
nor U18326 (N_18326,N_17461,N_16333);
or U18327 (N_18327,N_17332,N_17329);
xor U18328 (N_18328,N_17513,N_17683);
nand U18329 (N_18329,N_17875,N_17383);
nand U18330 (N_18330,N_17973,N_16287);
and U18331 (N_18331,N_17752,N_17896);
nor U18332 (N_18332,N_17760,N_16086);
or U18333 (N_18333,N_16310,N_17891);
or U18334 (N_18334,N_17384,N_17012);
xor U18335 (N_18335,N_16473,N_16824);
or U18336 (N_18336,N_16717,N_17519);
or U18337 (N_18337,N_16403,N_17895);
or U18338 (N_18338,N_17130,N_17506);
and U18339 (N_18339,N_17950,N_16764);
and U18340 (N_18340,N_17425,N_17502);
nand U18341 (N_18341,N_16491,N_17057);
xor U18342 (N_18342,N_17405,N_17198);
or U18343 (N_18343,N_16998,N_16581);
or U18344 (N_18344,N_16365,N_16535);
and U18345 (N_18345,N_17343,N_16466);
and U18346 (N_18346,N_17368,N_17996);
or U18347 (N_18347,N_17290,N_17284);
nor U18348 (N_18348,N_16589,N_17864);
nand U18349 (N_18349,N_16929,N_16061);
xnor U18350 (N_18350,N_17897,N_17129);
and U18351 (N_18351,N_16208,N_17899);
nor U18352 (N_18352,N_16948,N_16533);
nor U18353 (N_18353,N_16474,N_17928);
or U18354 (N_18354,N_17855,N_16965);
or U18355 (N_18355,N_16499,N_16791);
nor U18356 (N_18356,N_17662,N_17732);
nor U18357 (N_18357,N_17687,N_16065);
xor U18358 (N_18358,N_17540,N_17230);
nor U18359 (N_18359,N_16445,N_16924);
nor U18360 (N_18360,N_17052,N_17635);
xnor U18361 (N_18361,N_17219,N_16695);
nand U18362 (N_18362,N_17654,N_16960);
xnor U18363 (N_18363,N_16041,N_17103);
and U18364 (N_18364,N_17017,N_17630);
nand U18365 (N_18365,N_16743,N_16747);
or U18366 (N_18366,N_16905,N_16700);
xor U18367 (N_18367,N_17089,N_16784);
nand U18368 (N_18368,N_16687,N_17452);
and U18369 (N_18369,N_17144,N_17337);
nand U18370 (N_18370,N_16037,N_17713);
or U18371 (N_18371,N_17699,N_16346);
or U18372 (N_18372,N_17776,N_17328);
and U18373 (N_18373,N_16294,N_16414);
and U18374 (N_18374,N_17769,N_16963);
nand U18375 (N_18375,N_16121,N_16834);
nand U18376 (N_18376,N_16329,N_17798);
nand U18377 (N_18377,N_17141,N_16017);
nor U18378 (N_18378,N_17869,N_16701);
xnor U18379 (N_18379,N_17370,N_16019);
or U18380 (N_18380,N_16565,N_17291);
xnor U18381 (N_18381,N_16113,N_16405);
and U18382 (N_18382,N_16039,N_17898);
and U18383 (N_18383,N_16131,N_16850);
nand U18384 (N_18384,N_16580,N_17576);
and U18385 (N_18385,N_16509,N_17195);
nand U18386 (N_18386,N_16149,N_17327);
xor U18387 (N_18387,N_16275,N_17803);
and U18388 (N_18388,N_16899,N_17318);
xor U18389 (N_18389,N_16880,N_17339);
xnor U18390 (N_18390,N_17656,N_16751);
and U18391 (N_18391,N_16707,N_16655);
nand U18392 (N_18392,N_16777,N_17381);
and U18393 (N_18393,N_17279,N_16216);
xnor U18394 (N_18394,N_17451,N_17321);
or U18395 (N_18395,N_17341,N_17242);
nand U18396 (N_18396,N_16638,N_17215);
nor U18397 (N_18397,N_17778,N_17246);
nor U18398 (N_18398,N_16368,N_17589);
and U18399 (N_18399,N_17420,N_16168);
or U18400 (N_18400,N_16799,N_17790);
xnor U18401 (N_18401,N_17107,N_16351);
and U18402 (N_18402,N_17360,N_16879);
and U18403 (N_18403,N_16460,N_17439);
and U18404 (N_18404,N_17992,N_17201);
xor U18405 (N_18405,N_16140,N_16626);
and U18406 (N_18406,N_17411,N_16641);
nand U18407 (N_18407,N_17572,N_17866);
and U18408 (N_18408,N_17148,N_17785);
nor U18409 (N_18409,N_17915,N_16795);
xnor U18410 (N_18410,N_16134,N_17257);
and U18411 (N_18411,N_16374,N_16959);
and U18412 (N_18412,N_16597,N_16378);
nand U18413 (N_18413,N_17254,N_17971);
nor U18414 (N_18414,N_17084,N_17316);
xor U18415 (N_18415,N_16420,N_17001);
xor U18416 (N_18416,N_17024,N_16887);
or U18417 (N_18417,N_17827,N_16817);
nor U18418 (N_18418,N_17079,N_17661);
xor U18419 (N_18419,N_17447,N_17967);
or U18420 (N_18420,N_17093,N_16366);
or U18421 (N_18421,N_17182,N_16819);
and U18422 (N_18422,N_17792,N_17574);
or U18423 (N_18423,N_16501,N_16341);
and U18424 (N_18424,N_17675,N_16027);
nor U18425 (N_18425,N_17650,N_16529);
nand U18426 (N_18426,N_16571,N_17697);
nand U18427 (N_18427,N_17233,N_16201);
or U18428 (N_18428,N_17972,N_16302);
xor U18429 (N_18429,N_16392,N_17926);
xor U18430 (N_18430,N_16724,N_17688);
nor U18431 (N_18431,N_16682,N_16029);
xor U18432 (N_18432,N_16528,N_16926);
and U18433 (N_18433,N_17441,N_17541);
nor U18434 (N_18434,N_16559,N_16444);
and U18435 (N_18435,N_16066,N_17354);
xnor U18436 (N_18436,N_16884,N_16750);
or U18437 (N_18437,N_16070,N_17638);
and U18438 (N_18438,N_16674,N_17628);
and U18439 (N_18439,N_16143,N_16726);
nand U18440 (N_18440,N_17710,N_17853);
and U18441 (N_18441,N_17020,N_16304);
nand U18442 (N_18442,N_16756,N_16810);
and U18443 (N_18443,N_16145,N_16908);
nor U18444 (N_18444,N_16835,N_16979);
nor U18445 (N_18445,N_16556,N_17419);
nand U18446 (N_18446,N_16906,N_17265);
xnor U18447 (N_18447,N_16199,N_17801);
or U18448 (N_18448,N_17756,N_17573);
or U18449 (N_18449,N_16014,N_16477);
nand U18450 (N_18450,N_16513,N_16630);
and U18451 (N_18451,N_16647,N_17446);
and U18452 (N_18452,N_17435,N_16792);
xnor U18453 (N_18453,N_17787,N_17133);
nand U18454 (N_18454,N_17323,N_17569);
xor U18455 (N_18455,N_16583,N_16482);
xor U18456 (N_18456,N_16343,N_17322);
xor U18457 (N_18457,N_17229,N_17772);
nand U18458 (N_18458,N_16081,N_16593);
or U18459 (N_18459,N_16231,N_17091);
and U18460 (N_18460,N_17120,N_17216);
or U18461 (N_18461,N_17703,N_16363);
nand U18462 (N_18462,N_17154,N_17559);
or U18463 (N_18463,N_17946,N_17509);
and U18464 (N_18464,N_17958,N_16882);
and U18465 (N_18465,N_17677,N_16625);
nor U18466 (N_18466,N_16898,N_17010);
xor U18467 (N_18467,N_16892,N_17719);
or U18468 (N_18468,N_17186,N_16805);
and U18469 (N_18469,N_17736,N_16746);
xor U18470 (N_18470,N_17062,N_17715);
nand U18471 (N_18471,N_16105,N_17812);
nor U18472 (N_18472,N_17789,N_17538);
or U18473 (N_18473,N_16912,N_17042);
nor U18474 (N_18474,N_17849,N_17544);
nand U18475 (N_18475,N_16856,N_17408);
nor U18476 (N_18476,N_16221,N_17380);
nor U18477 (N_18477,N_17528,N_16415);
and U18478 (N_18478,N_17770,N_17263);
nor U18479 (N_18479,N_16907,N_17516);
and U18480 (N_18480,N_16511,N_17135);
nand U18481 (N_18481,N_17271,N_16434);
nor U18482 (N_18482,N_17681,N_17819);
xor U18483 (N_18483,N_16227,N_16670);
nor U18484 (N_18484,N_17169,N_16573);
or U18485 (N_18485,N_17644,N_16159);
nand U18486 (N_18486,N_16500,N_16453);
or U18487 (N_18487,N_17566,N_16833);
nand U18488 (N_18488,N_17913,N_17914);
xnor U18489 (N_18489,N_17073,N_16169);
and U18490 (N_18490,N_17515,N_16120);
and U18491 (N_18491,N_17966,N_17529);
and U18492 (N_18492,N_16980,N_16508);
xor U18493 (N_18493,N_17111,N_17918);
and U18494 (N_18494,N_17542,N_16023);
and U18495 (N_18495,N_16818,N_16534);
nand U18496 (N_18496,N_16495,N_17470);
or U18497 (N_18497,N_16303,N_17949);
nor U18498 (N_18498,N_17797,N_17302);
or U18499 (N_18499,N_16479,N_17796);
and U18500 (N_18500,N_16863,N_16471);
and U18501 (N_18501,N_17009,N_17522);
and U18502 (N_18502,N_17336,N_17917);
or U18503 (N_18503,N_16422,N_17870);
and U18504 (N_18504,N_16796,N_16372);
nand U18505 (N_18505,N_16656,N_17208);
nand U18506 (N_18506,N_16243,N_16921);
nor U18507 (N_18507,N_16144,N_17744);
nor U18508 (N_18508,N_16259,N_17754);
or U18509 (N_18509,N_16493,N_16459);
xor U18510 (N_18510,N_16367,N_16184);
nand U18511 (N_18511,N_16867,N_16922);
xnor U18512 (N_18512,N_16961,N_17521);
or U18513 (N_18513,N_16012,N_17563);
nand U18514 (N_18514,N_16595,N_16711);
nor U18515 (N_18515,N_16148,N_16020);
nand U18516 (N_18516,N_16151,N_17848);
or U18517 (N_18517,N_17080,N_16904);
nor U18518 (N_18518,N_16755,N_17101);
and U18519 (N_18519,N_17142,N_16119);
nor U18520 (N_18520,N_17054,N_17363);
or U18521 (N_18521,N_17963,N_17606);
and U18522 (N_18522,N_16484,N_16950);
or U18523 (N_18523,N_17110,N_17404);
and U18524 (N_18524,N_17031,N_17412);
xnor U18525 (N_18525,N_17139,N_16876);
and U18526 (N_18526,N_17694,N_16146);
and U18527 (N_18527,N_16311,N_17199);
xor U18528 (N_18528,N_17700,N_16525);
and U18529 (N_18529,N_17592,N_17586);
or U18530 (N_18530,N_17249,N_16323);
or U18531 (N_18531,N_17483,N_16334);
nor U18532 (N_18532,N_17561,N_16219);
xor U18533 (N_18533,N_16174,N_17867);
nor U18534 (N_18534,N_17727,N_16923);
nor U18535 (N_18535,N_16076,N_16305);
xor U18536 (N_18536,N_17762,N_16744);
nor U18537 (N_18537,N_16680,N_16617);
and U18538 (N_18538,N_17743,N_17273);
nand U18539 (N_18539,N_16666,N_17738);
nor U18540 (N_18540,N_17922,N_16024);
xor U18541 (N_18541,N_17783,N_16844);
nand U18542 (N_18542,N_17444,N_17214);
or U18543 (N_18543,N_16505,N_17564);
nand U18544 (N_18544,N_16633,N_16697);
nand U18545 (N_18545,N_17847,N_16590);
xnor U18546 (N_18546,N_16355,N_17714);
or U18547 (N_18547,N_16623,N_16874);
nand U18548 (N_18548,N_16970,N_16733);
and U18549 (N_18549,N_16815,N_16164);
or U18550 (N_18550,N_17206,N_17427);
nand U18551 (N_18551,N_17307,N_17074);
or U18552 (N_18552,N_17904,N_17065);
xor U18553 (N_18553,N_17836,N_16797);
xor U18554 (N_18554,N_17666,N_16049);
or U18555 (N_18555,N_17145,N_17430);
or U18556 (N_18556,N_17974,N_17860);
and U18557 (N_18557,N_16175,N_17739);
nor U18558 (N_18558,N_17877,N_16214);
and U18559 (N_18559,N_16273,N_16936);
and U18560 (N_18560,N_16481,N_16738);
xnor U18561 (N_18561,N_16510,N_17952);
xnor U18562 (N_18562,N_17525,N_17511);
nor U18563 (N_18563,N_16067,N_16830);
nor U18564 (N_18564,N_16671,N_16832);
xnor U18565 (N_18565,N_17989,N_17376);
xor U18566 (N_18566,N_16836,N_17474);
xnor U18567 (N_18567,N_16518,N_17015);
xnor U18568 (N_18568,N_17143,N_16981);
nand U18569 (N_18569,N_16601,N_16034);
and U18570 (N_18570,N_17260,N_17055);
or U18571 (N_18571,N_17184,N_17938);
xor U18572 (N_18572,N_16757,N_16913);
and U18573 (N_18573,N_17285,N_17122);
nand U18574 (N_18574,N_17314,N_16301);
or U18575 (N_18575,N_16448,N_17546);
nand U18576 (N_18576,N_17839,N_16574);
or U18577 (N_18577,N_17851,N_16207);
nor U18578 (N_18578,N_17040,N_17961);
nor U18579 (N_18579,N_16385,N_16446);
nand U18580 (N_18580,N_17308,N_17075);
xor U18581 (N_18581,N_17453,N_16567);
nor U18582 (N_18582,N_17030,N_16660);
nand U18583 (N_18583,N_16661,N_16088);
or U18584 (N_18584,N_16229,N_16440);
xor U18585 (N_18585,N_17944,N_16274);
nand U18586 (N_18586,N_16306,N_17407);
xnor U18587 (N_18587,N_16714,N_17393);
or U18588 (N_18588,N_17170,N_16450);
nand U18589 (N_18589,N_16071,N_16397);
xnor U18590 (N_18590,N_17495,N_17293);
nor U18591 (N_18591,N_16954,N_16658);
or U18592 (N_18592,N_17471,N_16934);
xnor U18593 (N_18593,N_16564,N_16881);
and U18594 (N_18594,N_16261,N_16248);
or U18595 (N_18595,N_16044,N_17044);
xor U18596 (N_18596,N_17256,N_17942);
or U18597 (N_18597,N_17237,N_16517);
nor U18598 (N_18598,N_16096,N_16704);
nand U18599 (N_18599,N_17364,N_16901);
xor U18600 (N_18600,N_16587,N_17180);
nor U18601 (N_18601,N_16915,N_16038);
nor U18602 (N_18602,N_16407,N_16047);
xnor U18603 (N_18603,N_16395,N_16852);
nand U18604 (N_18604,N_17994,N_17134);
or U18605 (N_18605,N_17585,N_16100);
nand U18606 (N_18606,N_17673,N_17900);
or U18607 (N_18607,N_17865,N_16944);
or U18608 (N_18608,N_16582,N_16686);
nor U18609 (N_18609,N_16490,N_17578);
and U18610 (N_18610,N_16699,N_17046);
or U18611 (N_18611,N_16873,N_16713);
xor U18612 (N_18612,N_17289,N_17317);
nand U18613 (N_18613,N_17320,N_17880);
or U18614 (N_18614,N_16715,N_16739);
nor U18615 (N_18615,N_17999,N_16991);
or U18616 (N_18616,N_17988,N_16042);
and U18617 (N_18617,N_17005,N_17047);
nand U18618 (N_18618,N_16254,N_16008);
or U18619 (N_18619,N_16325,N_16316);
xor U18620 (N_18620,N_16978,N_17059);
and U18621 (N_18621,N_16702,N_17188);
nor U18622 (N_18622,N_17369,N_16598);
and U18623 (N_18623,N_16352,N_17128);
or U18624 (N_18624,N_17292,N_17639);
or U18625 (N_18625,N_17755,N_17029);
nand U18626 (N_18626,N_17095,N_16496);
nor U18627 (N_18627,N_16137,N_17076);
nor U18628 (N_18628,N_17025,N_17172);
and U18629 (N_18629,N_16322,N_17804);
xnor U18630 (N_18630,N_16937,N_17871);
nand U18631 (N_18631,N_17816,N_16354);
nand U18632 (N_18632,N_17492,N_17882);
xor U18633 (N_18633,N_16592,N_17510);
and U18634 (N_18634,N_17746,N_17083);
xor U18635 (N_18635,N_16183,N_17403);
or U18636 (N_18636,N_17038,N_17027);
nand U18637 (N_18637,N_17211,N_16935);
or U18638 (N_18638,N_16837,N_16783);
nand U18639 (N_18639,N_16868,N_17560);
xor U18640 (N_18640,N_17879,N_17063);
and U18641 (N_18641,N_16866,N_17460);
and U18642 (N_18642,N_16875,N_17954);
nor U18643 (N_18643,N_16953,N_17476);
and U18644 (N_18644,N_16416,N_17227);
nor U18645 (N_18645,N_17131,N_17962);
xnor U18646 (N_18646,N_16945,N_17349);
and U18647 (N_18647,N_16677,N_16382);
nand U18648 (N_18648,N_16130,N_17440);
and U18649 (N_18649,N_17747,N_17532);
or U18650 (N_18650,N_17467,N_17117);
or U18651 (N_18651,N_17023,N_17998);
xor U18652 (N_18652,N_16947,N_17109);
xnor U18653 (N_18653,N_17893,N_16896);
nand U18654 (N_18654,N_17497,N_16331);
or U18655 (N_18655,N_17907,N_16449);
nor U18656 (N_18656,N_17955,N_16285);
and U18657 (N_18657,N_17202,N_16465);
and U18658 (N_18658,N_16708,N_17301);
xnor U18659 (N_18659,N_17602,N_16430);
or U18660 (N_18660,N_17286,N_17965);
xor U18661 (N_18661,N_17243,N_16999);
nor U18662 (N_18662,N_17085,N_17060);
nand U18663 (N_18663,N_16011,N_16725);
nor U18664 (N_18664,N_16591,N_17340);
or U18665 (N_18665,N_17842,N_17693);
and U18666 (N_18666,N_17832,N_16663);
or U18667 (N_18667,N_17799,N_17834);
nand U18668 (N_18668,N_17653,N_16782);
nand U18669 (N_18669,N_16753,N_16054);
xnor U18670 (N_18670,N_16249,N_17416);
or U18671 (N_18671,N_16710,N_17859);
or U18672 (N_18672,N_17358,N_16995);
nand U18673 (N_18673,N_16801,N_16798);
and U18674 (N_18674,N_16298,N_17734);
nand U18675 (N_18675,N_17993,N_16115);
or U18676 (N_18676,N_16326,N_16239);
nand U18677 (N_18677,N_17174,N_16703);
nand U18678 (N_18678,N_16530,N_17146);
nand U18679 (N_18679,N_17462,N_17377);
xnor U18680 (N_18680,N_16885,N_16278);
or U18681 (N_18681,N_16545,N_17035);
and U18682 (N_18682,N_16839,N_16497);
nor U18683 (N_18683,N_17078,N_16521);
and U18684 (N_18684,N_17150,N_17876);
nor U18685 (N_18685,N_16429,N_17750);
nand U18686 (N_18686,N_17228,N_17433);
or U18687 (N_18687,N_17674,N_16247);
and U18688 (N_18688,N_16432,N_16170);
or U18689 (N_18689,N_17737,N_16198);
nor U18690 (N_18690,N_16277,N_16224);
nand U18691 (N_18691,N_17627,N_16594);
xor U18692 (N_18692,N_17616,N_17463);
and U18693 (N_18693,N_17238,N_16846);
xnor U18694 (N_18694,N_17223,N_17478);
xor U18695 (N_18695,N_17709,N_16000);
nand U18696 (N_18696,N_16056,N_16966);
and U18697 (N_18697,N_16512,N_17621);
or U18698 (N_18698,N_16918,N_17995);
or U18699 (N_18699,N_16028,N_17811);
or U18700 (N_18700,N_16237,N_17794);
nand U18701 (N_18701,N_17014,N_16475);
xnor U18702 (N_18702,N_17007,N_16242);
nand U18703 (N_18703,N_17775,N_17959);
nor U18704 (N_18704,N_16220,N_17647);
xnor U18705 (N_18705,N_17507,N_17655);
nor U18706 (N_18706,N_16650,N_16772);
xor U18707 (N_18707,N_16319,N_17696);
and U18708 (N_18708,N_17533,N_17782);
nand U18709 (N_18709,N_17911,N_16197);
or U18710 (N_18710,N_17119,N_17947);
nand U18711 (N_18711,N_17916,N_17582);
and U18712 (N_18712,N_16748,N_17553);
nor U18713 (N_18713,N_16842,N_16916);
nor U18714 (N_18714,N_16478,N_17097);
nor U18715 (N_18715,N_17791,N_17902);
nor U18716 (N_18716,N_17070,N_17413);
and U18717 (N_18717,N_17013,N_17140);
nor U18718 (N_18718,N_17872,N_16139);
nor U18719 (N_18719,N_16996,N_16324);
nand U18720 (N_18720,N_16236,N_16074);
and U18721 (N_18721,N_16244,N_17196);
and U18722 (N_18722,N_16665,N_17932);
or U18723 (N_18723,N_16266,N_17862);
or U18724 (N_18724,N_16117,N_16779);
nor U18725 (N_18725,N_16558,N_16957);
xor U18726 (N_18726,N_17325,N_16186);
and U18727 (N_18727,N_17933,N_17712);
nand U18728 (N_18728,N_17258,N_17300);
nand U18729 (N_18729,N_17824,N_17889);
nor U18730 (N_18730,N_16886,N_17217);
nor U18731 (N_18731,N_17275,N_17840);
and U18732 (N_18732,N_16467,N_17689);
and U18733 (N_18733,N_16211,N_16167);
nor U18734 (N_18734,N_17004,N_17537);
nor U18735 (N_18735,N_17401,N_16264);
nor U18736 (N_18736,N_16492,N_16854);
or U18737 (N_18737,N_16206,N_17442);
nor U18738 (N_18738,N_17594,N_16654);
xor U18739 (N_18739,N_16554,N_17379);
nor U18740 (N_18740,N_16223,N_17806);
or U18741 (N_18741,N_16547,N_17112);
xnor U18742 (N_18742,N_17890,N_17808);
xor U18743 (N_18743,N_16349,N_16256);
nand U18744 (N_18744,N_17795,N_17008);
nor U18745 (N_18745,N_16084,N_16690);
nor U18746 (N_18746,N_16653,N_17053);
nand U18747 (N_18747,N_16949,N_17398);
nand U18748 (N_18748,N_16296,N_16043);
nor U18749 (N_18749,N_17203,N_16712);
nand U18750 (N_18750,N_16400,N_16939);
nor U18751 (N_18751,N_16128,N_16408);
and U18752 (N_18752,N_17457,N_16919);
xor U18753 (N_18753,N_17773,N_16161);
nand U18754 (N_18754,N_17780,N_17641);
xnor U18755 (N_18755,N_16575,N_16989);
and U18756 (N_18756,N_16502,N_17160);
nor U18757 (N_18757,N_17088,N_16225);
or U18758 (N_18758,N_16644,N_17948);
nand U18759 (N_18759,N_17596,N_16162);
or U18760 (N_18760,N_16551,N_16731);
or U18761 (N_18761,N_17045,N_16488);
nor U18762 (N_18762,N_16621,N_16828);
nor U18763 (N_18763,N_16421,N_17234);
xnor U18764 (N_18764,N_16158,N_16288);
or U18765 (N_18765,N_17069,N_16664);
nor U18766 (N_18766,N_17856,N_17923);
and U18767 (N_18767,N_17374,N_17213);
or U18768 (N_18768,N_17193,N_17449);
and U18769 (N_18769,N_17098,N_16092);
xnor U18770 (N_18770,N_17976,N_16888);
nand U18771 (N_18771,N_16871,N_16362);
xnor U18772 (N_18772,N_16258,N_17448);
or U18773 (N_18773,N_17176,N_16364);
xor U18774 (N_18774,N_16463,N_16869);
nand U18775 (N_18775,N_16627,N_17036);
nand U18776 (N_18776,N_16399,N_17822);
nand U18777 (N_18777,N_17548,N_16620);
or U18778 (N_18778,N_16217,N_17684);
nor U18779 (N_18779,N_16073,N_16903);
xor U18780 (N_18780,N_16315,N_17826);
and U18781 (N_18781,N_17707,N_17729);
nor U18782 (N_18782,N_17191,N_17987);
xnor U18783 (N_18783,N_16806,N_17236);
nand U18784 (N_18784,N_16215,N_17423);
and U18785 (N_18785,N_17356,N_17610);
or U18786 (N_18786,N_17906,N_17501);
nor U18787 (N_18787,N_17733,N_16848);
nand U18788 (N_18788,N_16925,N_16562);
nor U18789 (N_18789,N_17104,N_17983);
nor U18790 (N_18790,N_16897,N_17028);
and U18791 (N_18791,N_17818,N_16584);
or U18792 (N_18792,N_17781,N_17985);
or U18793 (N_18793,N_17283,N_16339);
nand U18794 (N_18794,N_16433,N_17350);
xnor U18795 (N_18795,N_16373,N_16557);
xnor U18796 (N_18796,N_16431,N_17437);
or U18797 (N_18797,N_17210,N_16967);
or U18798 (N_18798,N_17147,N_17680);
or U18799 (N_18799,N_17846,N_17396);
nor U18800 (N_18800,N_17108,N_16026);
and U18801 (N_18801,N_16413,N_17625);
xnor U18802 (N_18802,N_17304,N_16870);
and U18803 (N_18803,N_16461,N_17167);
and U18804 (N_18804,N_16210,N_17338);
or U18805 (N_18805,N_17450,N_17676);
nor U18806 (N_18806,N_16052,N_17597);
nand U18807 (N_18807,N_17455,N_16616);
or U18808 (N_18808,N_17459,N_17225);
and U18809 (N_18809,N_17825,N_16684);
nor U18810 (N_18810,N_16370,N_17800);
xnor U18811 (N_18811,N_16676,N_16263);
nand U18812 (N_18812,N_16153,N_16087);
and U18813 (N_18813,N_16943,N_17353);
nor U18814 (N_18814,N_16154,N_17392);
nand U18815 (N_18815,N_17874,N_16860);
or U18816 (N_18816,N_17838,N_17704);
or U18817 (N_18817,N_16814,N_17613);
xor U18818 (N_18818,N_16737,N_16520);
nor U18819 (N_18819,N_16992,N_17125);
nor U18820 (N_18820,N_16504,N_17245);
and U18821 (N_18821,N_17682,N_17646);
xor U18822 (N_18822,N_16111,N_16728);
nor U18823 (N_18823,N_16585,N_17443);
or U18824 (N_18824,N_16255,N_17883);
or U18825 (N_18825,N_16124,N_16546);
xnor U18826 (N_18826,N_17375,N_16335);
nand U18827 (N_18827,N_16050,N_16185);
nand U18828 (N_18828,N_17718,N_16340);
xnor U18829 (N_18829,N_16610,N_17557);
xor U18830 (N_18830,N_16793,N_16276);
xnor U18831 (N_18831,N_17829,N_16068);
and U18832 (N_18832,N_16347,N_16360);
nor U18833 (N_18833,N_17624,N_16293);
xnor U18834 (N_18834,N_17920,N_16646);
and U18835 (N_18835,N_17251,N_16790);
and U18836 (N_18836,N_16393,N_17280);
nor U18837 (N_18837,N_17335,N_17382);
nor U18838 (N_18838,N_17524,N_16993);
or U18839 (N_18839,N_16548,N_16377);
xnor U18840 (N_18840,N_16578,N_16971);
and U18841 (N_18841,N_17438,N_17607);
nand U18842 (N_18842,N_16969,N_16063);
nand U18843 (N_18843,N_17445,N_17355);
nor U18844 (N_18844,N_17708,N_16122);
nor U18845 (N_18845,N_16328,N_17692);
xor U18846 (N_18846,N_17520,N_17039);
xnor U18847 (N_18847,N_17155,N_17722);
or U18848 (N_18848,N_16997,N_17766);
and U18849 (N_18849,N_16079,N_17660);
nand U18850 (N_18850,N_17584,N_17414);
nand U18851 (N_18851,N_16390,N_17490);
or U18852 (N_18852,N_16101,N_16489);
and U18853 (N_18853,N_16116,N_16234);
or U18854 (N_18854,N_16250,N_16055);
xor U18855 (N_18855,N_16107,N_16104);
or U18856 (N_18856,N_16307,N_16732);
or U18857 (N_18857,N_16952,N_16603);
xor U18858 (N_18858,N_17496,N_16787);
nor U18859 (N_18859,N_16841,N_16618);
and U18860 (N_18860,N_17731,N_16152);
nand U18861 (N_18861,N_16235,N_16251);
xnor U18862 (N_18862,N_16539,N_17479);
nand U18863 (N_18863,N_17664,N_17372);
nand U18864 (N_18864,N_17612,N_16396);
xor U18865 (N_18865,N_17049,N_16672);
xor U18866 (N_18866,N_17861,N_17626);
or U18867 (N_18867,N_16072,N_17543);
and U18868 (N_18868,N_17631,N_17431);
or U18869 (N_18869,N_16973,N_16401);
nor U18870 (N_18870,N_16379,N_17138);
xnor U18871 (N_18871,N_17706,N_17831);
or U18872 (N_18872,N_17753,N_17615);
nor U18873 (N_18873,N_16544,N_16643);
or U18874 (N_18874,N_16384,N_17960);
nand U18875 (N_18875,N_17565,N_17068);
nor U18876 (N_18876,N_16442,N_16464);
nand U18877 (N_18877,N_17930,N_16526);
nand U18878 (N_18878,N_17105,N_17415);
xnor U18879 (N_18879,N_17371,N_17723);
nand U18880 (N_18880,N_17294,N_16389);
nor U18881 (N_18881,N_16204,N_16386);
nand U18882 (N_18882,N_16182,N_16803);
nand U18883 (N_18883,N_16069,N_16696);
xor U18884 (N_18884,N_16455,N_17745);
and U18885 (N_18885,N_17637,N_17567);
nor U18886 (N_18886,N_16033,N_16988);
or U18887 (N_18887,N_17244,N_17657);
or U18888 (N_18888,N_17645,N_16629);
and U18889 (N_18889,N_17648,N_16342);
or U18890 (N_18890,N_16409,N_16692);
xor U18891 (N_18891,N_17658,N_16246);
and U18892 (N_18892,N_17526,N_17158);
or U18893 (N_18893,N_16524,N_17605);
or U18894 (N_18894,N_17395,N_16946);
or U18895 (N_18895,N_17189,N_16189);
and U18896 (N_18896,N_17527,N_16857);
and U18897 (N_18897,N_17835,N_16532);
nand U18898 (N_18898,N_17221,N_17728);
and U18899 (N_18899,N_16163,N_16804);
and U18900 (N_18900,N_17468,N_16337);
xnor U18901 (N_18901,N_16108,N_17691);
and U18902 (N_18902,N_16930,N_16889);
or U18903 (N_18903,N_17261,N_16761);
and U18904 (N_18904,N_17828,N_16417);
nor U18905 (N_18905,N_16709,N_17575);
nor U18906 (N_18906,N_17558,N_17255);
xor U18907 (N_18907,N_17813,N_17277);
and U18908 (N_18908,N_16679,N_17611);
and U18909 (N_18909,N_16822,N_17264);
or U18910 (N_18910,N_17634,N_16404);
nor U18911 (N_18911,N_16605,N_17466);
and U18912 (N_18912,N_16109,N_16156);
and U18913 (N_18913,N_16005,N_16129);
and U18914 (N_18914,N_17090,N_17595);
nand U18915 (N_18915,N_16269,N_17161);
or U18916 (N_18916,N_17232,N_17604);
and U18917 (N_18917,N_16883,N_16394);
nand U18918 (N_18918,N_17924,N_16338);
nand U18919 (N_18919,N_16877,N_16289);
and U18920 (N_18920,N_17127,N_16825);
and U18921 (N_18921,N_17672,N_17590);
and U18922 (N_18922,N_16862,N_16388);
xnor U18923 (N_18923,N_16361,N_16808);
nor U18924 (N_18924,N_17552,N_16668);
and U18925 (N_18925,N_17885,N_17991);
or U18926 (N_18926,N_16157,N_16608);
and U18927 (N_18927,N_16566,N_16297);
nor U18928 (N_18928,N_17296,N_16030);
xor U18929 (N_18929,N_17422,N_17518);
and U18930 (N_18930,N_16675,N_16462);
or U18931 (N_18931,N_17759,N_17399);
and U18932 (N_18932,N_16064,N_17056);
and U18933 (N_18933,N_17428,N_17633);
nor U18934 (N_18934,N_17539,N_16865);
and U18935 (N_18935,N_16097,N_16358);
nor U18936 (N_18936,N_17305,N_16659);
nor U18937 (N_18937,N_17330,N_16102);
xor U18938 (N_18938,N_16840,N_16350);
and U18939 (N_18939,N_17771,N_16470);
and U18940 (N_18940,N_16257,N_16600);
or U18941 (N_18941,N_16371,N_16138);
or U18942 (N_18942,N_17493,N_17763);
nor U18943 (N_18943,N_16356,N_16561);
and U18944 (N_18944,N_17421,N_17939);
nor U18945 (N_18945,N_17124,N_17665);
or U18946 (N_18946,N_17554,N_17868);
or U18947 (N_18947,N_16891,N_16628);
or U18948 (N_18948,N_17820,N_17424);
nor U18949 (N_18949,N_16678,N_16657);
nor U18950 (N_18950,N_17194,N_16820);
nand U18951 (N_18951,N_16789,N_17937);
xnor U18952 (N_18952,N_16172,N_17309);
nor U18953 (N_18953,N_16238,N_16209);
nor U18954 (N_18954,N_16321,N_17711);
nor U18955 (N_18955,N_16036,N_17409);
xnor U18956 (N_18956,N_17207,N_16773);
and U18957 (N_18957,N_16694,N_17205);
xor U18958 (N_18958,N_17268,N_16299);
or U18959 (N_18959,N_17288,N_16451);
and U18960 (N_18960,N_16986,N_16418);
nor U18961 (N_18961,N_17977,N_16007);
or U18962 (N_18962,N_16270,N_17767);
and U18963 (N_18963,N_17764,N_16994);
xor U18964 (N_18964,N_17276,N_17980);
and U18965 (N_18965,N_16576,N_16123);
and U18966 (N_18966,N_16380,N_16082);
xor U18967 (N_18967,N_17901,N_16435);
xor U18968 (N_18968,N_17051,N_17250);
xor U18969 (N_18969,N_17175,N_17695);
and U18970 (N_18970,N_16142,N_16232);
nand U18971 (N_18971,N_17823,N_16428);
nor U18972 (N_18972,N_17113,N_17344);
xnor U18973 (N_18973,N_16472,N_17429);
and U18974 (N_18974,N_16962,N_17843);
xor U18975 (N_18975,N_16245,N_17986);
xor U18976 (N_18976,N_16572,N_16982);
xor U18977 (N_18977,N_16515,N_16662);
xnor U18978 (N_18978,N_16754,N_16095);
nor U18979 (N_18979,N_17716,N_16439);
nand U18980 (N_18980,N_16267,N_16179);
or U18981 (N_18981,N_16681,N_16766);
nand U18982 (N_18982,N_16133,N_17171);
nor U18983 (N_18983,N_17583,N_17240);
or U18984 (N_18984,N_17387,N_16537);
xor U18985 (N_18985,N_17919,N_17514);
nor U18986 (N_18986,N_16759,N_16983);
nor U18987 (N_18987,N_17598,N_17018);
nor U18988 (N_18988,N_17156,N_17970);
and U18989 (N_18989,N_17252,N_17269);
nand U18990 (N_18990,N_17361,N_16476);
or U18991 (N_18991,N_17000,N_16691);
and U18992 (N_18992,N_16135,N_17536);
nand U18993 (N_18993,N_17779,N_16667);
nand U18994 (N_18994,N_16927,N_16155);
and U18995 (N_18995,N_16763,N_16864);
nand U18996 (N_18996,N_17326,N_16233);
and U18997 (N_18997,N_16698,N_16776);
xor U18998 (N_18998,N_16485,N_16106);
and U18999 (N_18999,N_16487,N_16522);
or U19000 (N_19000,N_17971,N_16147);
nand U19001 (N_19001,N_17552,N_17719);
nand U19002 (N_19002,N_16139,N_17697);
xnor U19003 (N_19003,N_16070,N_16151);
nand U19004 (N_19004,N_16780,N_16488);
nand U19005 (N_19005,N_17324,N_16796);
xor U19006 (N_19006,N_16210,N_17997);
or U19007 (N_19007,N_17375,N_17598);
xnor U19008 (N_19008,N_17512,N_17853);
xor U19009 (N_19009,N_17650,N_16115);
nand U19010 (N_19010,N_17531,N_16355);
nor U19011 (N_19011,N_17509,N_16863);
nand U19012 (N_19012,N_17965,N_16603);
or U19013 (N_19013,N_16992,N_17495);
nand U19014 (N_19014,N_16392,N_17308);
or U19015 (N_19015,N_16417,N_17029);
nor U19016 (N_19016,N_16281,N_17544);
or U19017 (N_19017,N_16896,N_17460);
and U19018 (N_19018,N_16501,N_16638);
xnor U19019 (N_19019,N_17764,N_17035);
and U19020 (N_19020,N_17916,N_16332);
and U19021 (N_19021,N_16682,N_16915);
or U19022 (N_19022,N_17184,N_17892);
xnor U19023 (N_19023,N_16487,N_17046);
or U19024 (N_19024,N_17305,N_16835);
or U19025 (N_19025,N_17715,N_17744);
and U19026 (N_19026,N_16664,N_17318);
and U19027 (N_19027,N_16182,N_16837);
or U19028 (N_19028,N_16018,N_16809);
nor U19029 (N_19029,N_17479,N_17818);
xnor U19030 (N_19030,N_16957,N_16165);
and U19031 (N_19031,N_17421,N_16113);
and U19032 (N_19032,N_16181,N_16845);
and U19033 (N_19033,N_17232,N_17308);
nand U19034 (N_19034,N_17824,N_16833);
and U19035 (N_19035,N_16584,N_16826);
nand U19036 (N_19036,N_17159,N_17308);
or U19037 (N_19037,N_16217,N_17375);
nand U19038 (N_19038,N_17450,N_16897);
nand U19039 (N_19039,N_16330,N_16679);
xor U19040 (N_19040,N_16250,N_17750);
nand U19041 (N_19041,N_17577,N_17249);
xnor U19042 (N_19042,N_16607,N_16663);
nor U19043 (N_19043,N_16635,N_16700);
nor U19044 (N_19044,N_17536,N_16208);
and U19045 (N_19045,N_16226,N_16317);
and U19046 (N_19046,N_17728,N_16561);
or U19047 (N_19047,N_17580,N_17116);
xor U19048 (N_19048,N_17256,N_17121);
xor U19049 (N_19049,N_17632,N_16216);
nor U19050 (N_19050,N_16255,N_16351);
and U19051 (N_19051,N_16526,N_16956);
nor U19052 (N_19052,N_16213,N_17924);
and U19053 (N_19053,N_17835,N_17571);
and U19054 (N_19054,N_17355,N_16700);
nor U19055 (N_19055,N_16327,N_16814);
xor U19056 (N_19056,N_17585,N_16882);
xor U19057 (N_19057,N_17864,N_17677);
or U19058 (N_19058,N_16902,N_16393);
nand U19059 (N_19059,N_17064,N_17992);
nand U19060 (N_19060,N_16267,N_16796);
nand U19061 (N_19061,N_17903,N_17060);
nand U19062 (N_19062,N_17800,N_16882);
and U19063 (N_19063,N_17896,N_16073);
or U19064 (N_19064,N_17841,N_16244);
nor U19065 (N_19065,N_16908,N_16920);
xnor U19066 (N_19066,N_16692,N_17652);
nor U19067 (N_19067,N_16684,N_17600);
nand U19068 (N_19068,N_17589,N_17539);
or U19069 (N_19069,N_16645,N_17700);
nand U19070 (N_19070,N_17114,N_17996);
and U19071 (N_19071,N_17540,N_17638);
xnor U19072 (N_19072,N_16805,N_17523);
and U19073 (N_19073,N_17880,N_17020);
or U19074 (N_19074,N_16424,N_17035);
xnor U19075 (N_19075,N_16992,N_17465);
or U19076 (N_19076,N_16422,N_16203);
xor U19077 (N_19077,N_16727,N_17368);
nor U19078 (N_19078,N_17084,N_16353);
xnor U19079 (N_19079,N_17899,N_17821);
nor U19080 (N_19080,N_16711,N_17237);
and U19081 (N_19081,N_17941,N_17733);
nor U19082 (N_19082,N_17949,N_17359);
nand U19083 (N_19083,N_17590,N_16613);
xor U19084 (N_19084,N_16935,N_17523);
and U19085 (N_19085,N_17097,N_17490);
nand U19086 (N_19086,N_17556,N_17045);
xor U19087 (N_19087,N_17542,N_16835);
or U19088 (N_19088,N_17743,N_17047);
nor U19089 (N_19089,N_16174,N_16810);
xnor U19090 (N_19090,N_17982,N_17844);
nor U19091 (N_19091,N_16415,N_16737);
xnor U19092 (N_19092,N_17754,N_16253);
or U19093 (N_19093,N_17413,N_17214);
or U19094 (N_19094,N_17712,N_16740);
or U19095 (N_19095,N_17208,N_16675);
and U19096 (N_19096,N_16595,N_17699);
or U19097 (N_19097,N_16127,N_16482);
or U19098 (N_19098,N_17254,N_17775);
or U19099 (N_19099,N_17170,N_17751);
nor U19100 (N_19100,N_16045,N_17340);
nor U19101 (N_19101,N_16496,N_17221);
and U19102 (N_19102,N_17818,N_16163);
and U19103 (N_19103,N_17430,N_17296);
nor U19104 (N_19104,N_17889,N_16928);
xnor U19105 (N_19105,N_17762,N_17492);
or U19106 (N_19106,N_16206,N_17913);
nor U19107 (N_19107,N_16830,N_17861);
or U19108 (N_19108,N_17932,N_17956);
nor U19109 (N_19109,N_17728,N_16106);
and U19110 (N_19110,N_16390,N_16479);
nand U19111 (N_19111,N_17238,N_16064);
nor U19112 (N_19112,N_16526,N_16183);
xor U19113 (N_19113,N_16111,N_17245);
nor U19114 (N_19114,N_16455,N_16966);
and U19115 (N_19115,N_17076,N_16736);
nand U19116 (N_19116,N_16103,N_17084);
nand U19117 (N_19117,N_16927,N_16395);
nand U19118 (N_19118,N_16493,N_16659);
and U19119 (N_19119,N_17319,N_16232);
or U19120 (N_19120,N_16802,N_17721);
and U19121 (N_19121,N_17857,N_16874);
and U19122 (N_19122,N_16820,N_16225);
nand U19123 (N_19123,N_17024,N_16939);
or U19124 (N_19124,N_16246,N_16701);
nor U19125 (N_19125,N_16998,N_16240);
or U19126 (N_19126,N_17929,N_16592);
xnor U19127 (N_19127,N_17872,N_17816);
nor U19128 (N_19128,N_17938,N_16301);
nor U19129 (N_19129,N_17780,N_16372);
xnor U19130 (N_19130,N_17375,N_17086);
or U19131 (N_19131,N_17506,N_17233);
and U19132 (N_19132,N_16155,N_16428);
and U19133 (N_19133,N_17377,N_17237);
or U19134 (N_19134,N_17627,N_16426);
nand U19135 (N_19135,N_16706,N_17050);
xor U19136 (N_19136,N_16066,N_16959);
nor U19137 (N_19137,N_16383,N_17940);
xnor U19138 (N_19138,N_17840,N_17311);
or U19139 (N_19139,N_16968,N_16607);
nand U19140 (N_19140,N_17415,N_17194);
nand U19141 (N_19141,N_17146,N_17532);
nand U19142 (N_19142,N_16415,N_16768);
and U19143 (N_19143,N_16974,N_17649);
or U19144 (N_19144,N_17805,N_17072);
xnor U19145 (N_19145,N_16188,N_16657);
or U19146 (N_19146,N_16750,N_17378);
and U19147 (N_19147,N_16975,N_16595);
nand U19148 (N_19148,N_17877,N_16979);
nor U19149 (N_19149,N_17789,N_17321);
nor U19150 (N_19150,N_16327,N_17776);
nor U19151 (N_19151,N_16496,N_17190);
nor U19152 (N_19152,N_17278,N_16860);
xnor U19153 (N_19153,N_16133,N_16942);
nor U19154 (N_19154,N_17663,N_16124);
nor U19155 (N_19155,N_16320,N_17909);
nand U19156 (N_19156,N_17917,N_17121);
nand U19157 (N_19157,N_16150,N_16126);
nand U19158 (N_19158,N_16684,N_17766);
xnor U19159 (N_19159,N_16743,N_16559);
nand U19160 (N_19160,N_17632,N_16227);
xor U19161 (N_19161,N_16612,N_16433);
nand U19162 (N_19162,N_16636,N_16234);
nand U19163 (N_19163,N_17128,N_16503);
and U19164 (N_19164,N_17771,N_16023);
or U19165 (N_19165,N_17737,N_16658);
or U19166 (N_19166,N_16549,N_16618);
xor U19167 (N_19167,N_17430,N_16341);
nand U19168 (N_19168,N_17632,N_17093);
nor U19169 (N_19169,N_16081,N_17287);
or U19170 (N_19170,N_16486,N_16318);
nand U19171 (N_19171,N_17118,N_17676);
nor U19172 (N_19172,N_17168,N_17740);
nand U19173 (N_19173,N_16432,N_17487);
nand U19174 (N_19174,N_16068,N_17308);
xnor U19175 (N_19175,N_16605,N_16304);
nand U19176 (N_19176,N_17314,N_16837);
and U19177 (N_19177,N_16292,N_17755);
nand U19178 (N_19178,N_17588,N_16153);
nor U19179 (N_19179,N_16490,N_16751);
xor U19180 (N_19180,N_17232,N_16426);
nand U19181 (N_19181,N_16440,N_17516);
and U19182 (N_19182,N_16611,N_16656);
xor U19183 (N_19183,N_17461,N_16402);
and U19184 (N_19184,N_17381,N_16689);
nand U19185 (N_19185,N_16614,N_17067);
xor U19186 (N_19186,N_16802,N_17575);
nor U19187 (N_19187,N_17600,N_17203);
xor U19188 (N_19188,N_16225,N_17872);
nand U19189 (N_19189,N_16453,N_17711);
or U19190 (N_19190,N_17641,N_16937);
or U19191 (N_19191,N_17217,N_16540);
and U19192 (N_19192,N_16143,N_16441);
or U19193 (N_19193,N_17363,N_17075);
nor U19194 (N_19194,N_17336,N_16654);
nand U19195 (N_19195,N_17875,N_17650);
xor U19196 (N_19196,N_17385,N_17343);
or U19197 (N_19197,N_17171,N_17000);
nand U19198 (N_19198,N_16281,N_16060);
nor U19199 (N_19199,N_17002,N_17539);
nand U19200 (N_19200,N_16993,N_17141);
and U19201 (N_19201,N_16000,N_16280);
nor U19202 (N_19202,N_16340,N_16387);
and U19203 (N_19203,N_16434,N_17460);
nand U19204 (N_19204,N_17531,N_16333);
and U19205 (N_19205,N_17080,N_17993);
nand U19206 (N_19206,N_16539,N_16197);
nand U19207 (N_19207,N_16314,N_16034);
nand U19208 (N_19208,N_16270,N_17432);
and U19209 (N_19209,N_17842,N_16955);
and U19210 (N_19210,N_16813,N_17588);
and U19211 (N_19211,N_17423,N_17837);
or U19212 (N_19212,N_16658,N_17421);
nor U19213 (N_19213,N_17997,N_17179);
nor U19214 (N_19214,N_16895,N_17909);
xor U19215 (N_19215,N_17721,N_17429);
or U19216 (N_19216,N_17872,N_16141);
and U19217 (N_19217,N_16181,N_17318);
nor U19218 (N_19218,N_16174,N_17489);
nand U19219 (N_19219,N_16916,N_17992);
nand U19220 (N_19220,N_17095,N_17248);
nand U19221 (N_19221,N_17472,N_16109);
nand U19222 (N_19222,N_16798,N_17952);
and U19223 (N_19223,N_17409,N_17069);
nor U19224 (N_19224,N_17286,N_17566);
and U19225 (N_19225,N_17057,N_17810);
and U19226 (N_19226,N_16899,N_16313);
nor U19227 (N_19227,N_16478,N_17266);
nor U19228 (N_19228,N_16796,N_16134);
xor U19229 (N_19229,N_16163,N_17325);
and U19230 (N_19230,N_17139,N_17176);
nand U19231 (N_19231,N_17627,N_16145);
xnor U19232 (N_19232,N_16959,N_17716);
and U19233 (N_19233,N_16293,N_17777);
xnor U19234 (N_19234,N_16566,N_17267);
or U19235 (N_19235,N_16032,N_17630);
or U19236 (N_19236,N_16988,N_17067);
and U19237 (N_19237,N_16547,N_16903);
and U19238 (N_19238,N_16898,N_17804);
or U19239 (N_19239,N_16836,N_17704);
nor U19240 (N_19240,N_16496,N_17747);
nor U19241 (N_19241,N_16360,N_16130);
xor U19242 (N_19242,N_17912,N_16190);
and U19243 (N_19243,N_17446,N_17288);
and U19244 (N_19244,N_16099,N_17247);
nand U19245 (N_19245,N_16338,N_16439);
and U19246 (N_19246,N_17836,N_16447);
and U19247 (N_19247,N_16160,N_16206);
and U19248 (N_19248,N_17404,N_16526);
xnor U19249 (N_19249,N_16234,N_17401);
and U19250 (N_19250,N_16059,N_17806);
xor U19251 (N_19251,N_16884,N_16773);
and U19252 (N_19252,N_16864,N_17715);
nor U19253 (N_19253,N_16593,N_17609);
nor U19254 (N_19254,N_17543,N_16967);
xor U19255 (N_19255,N_16621,N_17363);
and U19256 (N_19256,N_17859,N_16965);
nand U19257 (N_19257,N_17626,N_17385);
or U19258 (N_19258,N_17239,N_16670);
nor U19259 (N_19259,N_16102,N_17051);
nor U19260 (N_19260,N_16735,N_16750);
nor U19261 (N_19261,N_16509,N_16521);
nor U19262 (N_19262,N_16336,N_16575);
nor U19263 (N_19263,N_17447,N_16034);
nor U19264 (N_19264,N_16276,N_17330);
xor U19265 (N_19265,N_16032,N_17297);
nand U19266 (N_19266,N_17154,N_17033);
nor U19267 (N_19267,N_17931,N_16998);
nor U19268 (N_19268,N_17808,N_17114);
xor U19269 (N_19269,N_16330,N_16529);
nand U19270 (N_19270,N_17456,N_16016);
or U19271 (N_19271,N_17216,N_17757);
xnor U19272 (N_19272,N_17022,N_16105);
xnor U19273 (N_19273,N_17009,N_16611);
xnor U19274 (N_19274,N_16903,N_16105);
nor U19275 (N_19275,N_16986,N_16011);
nor U19276 (N_19276,N_16154,N_17553);
nand U19277 (N_19277,N_17042,N_16474);
and U19278 (N_19278,N_17139,N_17705);
nand U19279 (N_19279,N_16195,N_17456);
nand U19280 (N_19280,N_16712,N_16375);
or U19281 (N_19281,N_16730,N_16343);
nand U19282 (N_19282,N_16933,N_16673);
xnor U19283 (N_19283,N_16383,N_16838);
nor U19284 (N_19284,N_17720,N_16842);
nand U19285 (N_19285,N_16394,N_16179);
nand U19286 (N_19286,N_16275,N_17827);
nor U19287 (N_19287,N_16480,N_17855);
xnor U19288 (N_19288,N_17354,N_17043);
or U19289 (N_19289,N_16285,N_17287);
xnor U19290 (N_19290,N_16423,N_17528);
and U19291 (N_19291,N_17861,N_17747);
xor U19292 (N_19292,N_16593,N_17885);
nand U19293 (N_19293,N_16593,N_17480);
xnor U19294 (N_19294,N_16346,N_16136);
and U19295 (N_19295,N_17214,N_17500);
and U19296 (N_19296,N_17820,N_17258);
xor U19297 (N_19297,N_17172,N_17724);
or U19298 (N_19298,N_17760,N_16723);
xor U19299 (N_19299,N_16883,N_16905);
or U19300 (N_19300,N_16581,N_16971);
or U19301 (N_19301,N_17400,N_16336);
nor U19302 (N_19302,N_16782,N_17388);
nand U19303 (N_19303,N_16930,N_16581);
xor U19304 (N_19304,N_17396,N_17638);
nor U19305 (N_19305,N_17322,N_17545);
and U19306 (N_19306,N_16711,N_16761);
or U19307 (N_19307,N_17466,N_16342);
or U19308 (N_19308,N_16595,N_17536);
and U19309 (N_19309,N_17868,N_17665);
nand U19310 (N_19310,N_17683,N_17154);
and U19311 (N_19311,N_16918,N_17328);
and U19312 (N_19312,N_17312,N_16941);
nor U19313 (N_19313,N_17350,N_16120);
and U19314 (N_19314,N_17925,N_17339);
nor U19315 (N_19315,N_16328,N_16018);
or U19316 (N_19316,N_16656,N_17359);
and U19317 (N_19317,N_17383,N_16968);
nor U19318 (N_19318,N_17163,N_16014);
or U19319 (N_19319,N_17561,N_16565);
nor U19320 (N_19320,N_16487,N_17423);
and U19321 (N_19321,N_16986,N_17696);
xnor U19322 (N_19322,N_16571,N_16030);
nand U19323 (N_19323,N_17923,N_16921);
and U19324 (N_19324,N_17443,N_17587);
nor U19325 (N_19325,N_16851,N_16052);
nor U19326 (N_19326,N_17744,N_17060);
xnor U19327 (N_19327,N_16178,N_17884);
xnor U19328 (N_19328,N_16435,N_16278);
or U19329 (N_19329,N_16977,N_17869);
nor U19330 (N_19330,N_16575,N_17062);
nor U19331 (N_19331,N_16644,N_16864);
and U19332 (N_19332,N_16999,N_17356);
xnor U19333 (N_19333,N_17731,N_17272);
xor U19334 (N_19334,N_16374,N_17205);
nand U19335 (N_19335,N_17166,N_16138);
nand U19336 (N_19336,N_16505,N_17240);
and U19337 (N_19337,N_16405,N_17223);
nand U19338 (N_19338,N_16048,N_17578);
nor U19339 (N_19339,N_17593,N_17843);
nand U19340 (N_19340,N_17279,N_17998);
and U19341 (N_19341,N_17589,N_17107);
or U19342 (N_19342,N_17990,N_16753);
nand U19343 (N_19343,N_16371,N_17971);
or U19344 (N_19344,N_17727,N_17626);
and U19345 (N_19345,N_16969,N_16038);
xor U19346 (N_19346,N_17842,N_17084);
and U19347 (N_19347,N_16002,N_17370);
and U19348 (N_19348,N_16888,N_16454);
or U19349 (N_19349,N_17941,N_17058);
and U19350 (N_19350,N_17652,N_17960);
or U19351 (N_19351,N_17023,N_16978);
and U19352 (N_19352,N_16666,N_16780);
nand U19353 (N_19353,N_17659,N_17034);
and U19354 (N_19354,N_17692,N_17169);
and U19355 (N_19355,N_17429,N_17897);
xnor U19356 (N_19356,N_17028,N_17836);
xor U19357 (N_19357,N_17434,N_16628);
nand U19358 (N_19358,N_16792,N_16923);
nand U19359 (N_19359,N_17826,N_16047);
and U19360 (N_19360,N_16279,N_16076);
xor U19361 (N_19361,N_17771,N_17076);
nor U19362 (N_19362,N_17377,N_17279);
xnor U19363 (N_19363,N_17472,N_17756);
nand U19364 (N_19364,N_16957,N_16585);
nor U19365 (N_19365,N_16870,N_17945);
xnor U19366 (N_19366,N_17104,N_16677);
nor U19367 (N_19367,N_17624,N_17059);
xnor U19368 (N_19368,N_16441,N_16977);
xnor U19369 (N_19369,N_17859,N_16743);
xor U19370 (N_19370,N_17305,N_17375);
and U19371 (N_19371,N_17610,N_17341);
nor U19372 (N_19372,N_16339,N_17698);
nand U19373 (N_19373,N_17857,N_17279);
xnor U19374 (N_19374,N_17848,N_17672);
or U19375 (N_19375,N_16298,N_16055);
and U19376 (N_19376,N_17767,N_16072);
or U19377 (N_19377,N_16513,N_17513);
nor U19378 (N_19378,N_16331,N_17435);
or U19379 (N_19379,N_16380,N_17454);
nor U19380 (N_19380,N_17296,N_16404);
nor U19381 (N_19381,N_17955,N_17240);
or U19382 (N_19382,N_17665,N_17842);
nand U19383 (N_19383,N_16964,N_17269);
and U19384 (N_19384,N_17262,N_16025);
xnor U19385 (N_19385,N_17490,N_16664);
xor U19386 (N_19386,N_17284,N_16588);
nand U19387 (N_19387,N_16270,N_17157);
or U19388 (N_19388,N_17756,N_16811);
xor U19389 (N_19389,N_16578,N_16160);
nor U19390 (N_19390,N_16821,N_16885);
and U19391 (N_19391,N_17831,N_16253);
xnor U19392 (N_19392,N_16428,N_16378);
nand U19393 (N_19393,N_17743,N_16898);
xnor U19394 (N_19394,N_17028,N_17623);
nor U19395 (N_19395,N_16101,N_17871);
or U19396 (N_19396,N_17568,N_16747);
and U19397 (N_19397,N_17364,N_16553);
xnor U19398 (N_19398,N_16507,N_17432);
xnor U19399 (N_19399,N_17292,N_16527);
xnor U19400 (N_19400,N_17350,N_17985);
xor U19401 (N_19401,N_16387,N_16483);
nor U19402 (N_19402,N_16605,N_17682);
and U19403 (N_19403,N_17674,N_17910);
or U19404 (N_19404,N_17386,N_17581);
or U19405 (N_19405,N_16014,N_17028);
nand U19406 (N_19406,N_16564,N_17701);
nand U19407 (N_19407,N_17688,N_16046);
and U19408 (N_19408,N_17696,N_16380);
nand U19409 (N_19409,N_16354,N_17377);
nand U19410 (N_19410,N_17330,N_17502);
or U19411 (N_19411,N_17215,N_17906);
nand U19412 (N_19412,N_17526,N_17964);
or U19413 (N_19413,N_17361,N_17659);
or U19414 (N_19414,N_17506,N_17630);
nor U19415 (N_19415,N_16461,N_17087);
or U19416 (N_19416,N_16503,N_17217);
and U19417 (N_19417,N_16313,N_16463);
or U19418 (N_19418,N_17866,N_16551);
xnor U19419 (N_19419,N_16231,N_17639);
nor U19420 (N_19420,N_16769,N_16212);
or U19421 (N_19421,N_17610,N_16289);
nor U19422 (N_19422,N_17711,N_17008);
xnor U19423 (N_19423,N_17945,N_16287);
and U19424 (N_19424,N_16595,N_17288);
or U19425 (N_19425,N_16040,N_16892);
nand U19426 (N_19426,N_17356,N_17133);
nand U19427 (N_19427,N_16751,N_16505);
nand U19428 (N_19428,N_16172,N_17255);
and U19429 (N_19429,N_17014,N_17551);
nor U19430 (N_19430,N_17365,N_16151);
and U19431 (N_19431,N_16962,N_17335);
or U19432 (N_19432,N_17850,N_16660);
nand U19433 (N_19433,N_17733,N_17845);
nor U19434 (N_19434,N_17667,N_16375);
and U19435 (N_19435,N_17956,N_17553);
and U19436 (N_19436,N_16962,N_17716);
nor U19437 (N_19437,N_16990,N_16614);
nand U19438 (N_19438,N_16671,N_16094);
nand U19439 (N_19439,N_17569,N_16080);
and U19440 (N_19440,N_16509,N_17824);
or U19441 (N_19441,N_16751,N_17337);
and U19442 (N_19442,N_16070,N_16389);
or U19443 (N_19443,N_17903,N_16597);
and U19444 (N_19444,N_16061,N_17686);
nand U19445 (N_19445,N_16946,N_17355);
and U19446 (N_19446,N_16160,N_17110);
nand U19447 (N_19447,N_17619,N_16516);
nor U19448 (N_19448,N_16832,N_16530);
xnor U19449 (N_19449,N_17394,N_17686);
nor U19450 (N_19450,N_17427,N_17084);
nand U19451 (N_19451,N_17977,N_17257);
or U19452 (N_19452,N_17238,N_17332);
nor U19453 (N_19453,N_17990,N_16302);
or U19454 (N_19454,N_17592,N_16752);
nand U19455 (N_19455,N_17851,N_17550);
nand U19456 (N_19456,N_17447,N_16655);
xnor U19457 (N_19457,N_16975,N_17959);
and U19458 (N_19458,N_16847,N_17641);
xnor U19459 (N_19459,N_17213,N_16884);
and U19460 (N_19460,N_17954,N_16631);
and U19461 (N_19461,N_16833,N_16522);
or U19462 (N_19462,N_16627,N_17460);
xor U19463 (N_19463,N_16425,N_17848);
and U19464 (N_19464,N_16816,N_17841);
or U19465 (N_19465,N_16675,N_16113);
or U19466 (N_19466,N_16964,N_17699);
or U19467 (N_19467,N_17339,N_17049);
nor U19468 (N_19468,N_17195,N_17567);
or U19469 (N_19469,N_16092,N_16051);
nor U19470 (N_19470,N_17837,N_17343);
xor U19471 (N_19471,N_17737,N_17541);
nor U19472 (N_19472,N_17855,N_17093);
nor U19473 (N_19473,N_16158,N_16310);
or U19474 (N_19474,N_17306,N_16884);
nand U19475 (N_19475,N_17276,N_17624);
or U19476 (N_19476,N_17506,N_16454);
or U19477 (N_19477,N_16842,N_16203);
nor U19478 (N_19478,N_16353,N_17373);
xor U19479 (N_19479,N_17289,N_17602);
xor U19480 (N_19480,N_17063,N_17931);
or U19481 (N_19481,N_16992,N_17751);
and U19482 (N_19482,N_16026,N_17388);
xnor U19483 (N_19483,N_17415,N_17012);
nor U19484 (N_19484,N_16673,N_16725);
xnor U19485 (N_19485,N_16792,N_17633);
nor U19486 (N_19486,N_17722,N_17898);
and U19487 (N_19487,N_16794,N_16399);
nor U19488 (N_19488,N_17103,N_17670);
and U19489 (N_19489,N_17470,N_17436);
or U19490 (N_19490,N_16236,N_16746);
nor U19491 (N_19491,N_17469,N_16265);
and U19492 (N_19492,N_16865,N_17729);
and U19493 (N_19493,N_17531,N_17280);
or U19494 (N_19494,N_17338,N_16031);
xor U19495 (N_19495,N_17527,N_17052);
and U19496 (N_19496,N_16687,N_17493);
nor U19497 (N_19497,N_16050,N_17119);
nor U19498 (N_19498,N_17372,N_17996);
nor U19499 (N_19499,N_17184,N_16153);
nor U19500 (N_19500,N_16905,N_17314);
nor U19501 (N_19501,N_16911,N_16488);
nor U19502 (N_19502,N_16184,N_16112);
and U19503 (N_19503,N_16076,N_17420);
nand U19504 (N_19504,N_17489,N_17728);
nand U19505 (N_19505,N_17458,N_17273);
and U19506 (N_19506,N_17151,N_16455);
xnor U19507 (N_19507,N_16751,N_17262);
nor U19508 (N_19508,N_17046,N_17340);
or U19509 (N_19509,N_16827,N_17937);
or U19510 (N_19510,N_17315,N_16854);
nor U19511 (N_19511,N_17625,N_17642);
nand U19512 (N_19512,N_16198,N_16837);
and U19513 (N_19513,N_16701,N_17397);
or U19514 (N_19514,N_16830,N_17593);
nand U19515 (N_19515,N_16217,N_16789);
and U19516 (N_19516,N_17908,N_16132);
nor U19517 (N_19517,N_16385,N_17298);
nand U19518 (N_19518,N_17515,N_17455);
or U19519 (N_19519,N_16447,N_16155);
xnor U19520 (N_19520,N_17409,N_17860);
nor U19521 (N_19521,N_16095,N_17833);
nor U19522 (N_19522,N_17426,N_16233);
xnor U19523 (N_19523,N_17822,N_16822);
and U19524 (N_19524,N_17471,N_16445);
nor U19525 (N_19525,N_17423,N_16900);
or U19526 (N_19526,N_16488,N_17143);
xnor U19527 (N_19527,N_16408,N_16452);
or U19528 (N_19528,N_16879,N_17294);
nand U19529 (N_19529,N_17941,N_16481);
or U19530 (N_19530,N_16779,N_17516);
and U19531 (N_19531,N_16348,N_17896);
nand U19532 (N_19532,N_17328,N_16016);
or U19533 (N_19533,N_17554,N_16522);
and U19534 (N_19534,N_16677,N_17496);
nand U19535 (N_19535,N_17436,N_17685);
nor U19536 (N_19536,N_17948,N_17834);
and U19537 (N_19537,N_16493,N_17157);
xor U19538 (N_19538,N_17382,N_17558);
and U19539 (N_19539,N_16125,N_16438);
and U19540 (N_19540,N_16219,N_16169);
and U19541 (N_19541,N_16904,N_16498);
nand U19542 (N_19542,N_17515,N_16282);
xor U19543 (N_19543,N_17298,N_17017);
nor U19544 (N_19544,N_16080,N_17059);
or U19545 (N_19545,N_17689,N_16358);
xnor U19546 (N_19546,N_17152,N_16368);
nand U19547 (N_19547,N_17133,N_17558);
or U19548 (N_19548,N_17424,N_17515);
nand U19549 (N_19549,N_16636,N_16637);
and U19550 (N_19550,N_17636,N_16697);
and U19551 (N_19551,N_16917,N_17136);
or U19552 (N_19552,N_17310,N_16532);
or U19553 (N_19553,N_17225,N_17105);
nor U19554 (N_19554,N_16001,N_17064);
and U19555 (N_19555,N_16302,N_17849);
nand U19556 (N_19556,N_16217,N_16015);
xor U19557 (N_19557,N_16267,N_17613);
nor U19558 (N_19558,N_17211,N_17109);
xnor U19559 (N_19559,N_17982,N_16565);
nand U19560 (N_19560,N_17024,N_16607);
nor U19561 (N_19561,N_16635,N_16014);
or U19562 (N_19562,N_16470,N_17235);
or U19563 (N_19563,N_17826,N_17853);
nor U19564 (N_19564,N_17692,N_16289);
or U19565 (N_19565,N_16252,N_16905);
xnor U19566 (N_19566,N_17135,N_16769);
or U19567 (N_19567,N_16670,N_17045);
nand U19568 (N_19568,N_16282,N_17699);
xor U19569 (N_19569,N_16255,N_17906);
or U19570 (N_19570,N_16207,N_16431);
xor U19571 (N_19571,N_16096,N_16753);
nor U19572 (N_19572,N_17494,N_16784);
or U19573 (N_19573,N_16801,N_16900);
xnor U19574 (N_19574,N_17439,N_16712);
and U19575 (N_19575,N_17294,N_16934);
or U19576 (N_19576,N_17766,N_17801);
nand U19577 (N_19577,N_17348,N_17259);
nor U19578 (N_19578,N_16117,N_17103);
or U19579 (N_19579,N_17311,N_17783);
nor U19580 (N_19580,N_17438,N_17181);
nand U19581 (N_19581,N_16337,N_16049);
or U19582 (N_19582,N_16749,N_16065);
nand U19583 (N_19583,N_17370,N_16251);
xnor U19584 (N_19584,N_16120,N_16783);
and U19585 (N_19585,N_17809,N_17250);
or U19586 (N_19586,N_16395,N_16449);
nor U19587 (N_19587,N_17998,N_17934);
nor U19588 (N_19588,N_16513,N_17679);
or U19589 (N_19589,N_17536,N_16019);
and U19590 (N_19590,N_16479,N_17668);
xnor U19591 (N_19591,N_16706,N_16152);
nand U19592 (N_19592,N_17548,N_17026);
xnor U19593 (N_19593,N_16126,N_17627);
and U19594 (N_19594,N_17211,N_17975);
xor U19595 (N_19595,N_16532,N_16117);
nand U19596 (N_19596,N_17389,N_17406);
xnor U19597 (N_19597,N_16242,N_17872);
xnor U19598 (N_19598,N_16438,N_17593);
nor U19599 (N_19599,N_17654,N_17976);
nor U19600 (N_19600,N_16295,N_16809);
or U19601 (N_19601,N_16656,N_16252);
or U19602 (N_19602,N_17912,N_16787);
xnor U19603 (N_19603,N_16410,N_17141);
or U19604 (N_19604,N_16467,N_16452);
and U19605 (N_19605,N_17292,N_16597);
or U19606 (N_19606,N_17453,N_17815);
or U19607 (N_19607,N_16106,N_17381);
and U19608 (N_19608,N_17371,N_16097);
or U19609 (N_19609,N_16012,N_17273);
or U19610 (N_19610,N_16046,N_17190);
or U19611 (N_19611,N_16280,N_16695);
nor U19612 (N_19612,N_16838,N_16049);
nor U19613 (N_19613,N_17148,N_16442);
nor U19614 (N_19614,N_16145,N_16538);
nor U19615 (N_19615,N_16208,N_17532);
and U19616 (N_19616,N_16525,N_17815);
and U19617 (N_19617,N_17300,N_16304);
nand U19618 (N_19618,N_16927,N_17792);
nand U19619 (N_19619,N_16994,N_17839);
and U19620 (N_19620,N_17127,N_17372);
xor U19621 (N_19621,N_16281,N_17551);
xnor U19622 (N_19622,N_16905,N_16668);
xnor U19623 (N_19623,N_17018,N_16733);
nand U19624 (N_19624,N_17755,N_16110);
xnor U19625 (N_19625,N_17904,N_16421);
xor U19626 (N_19626,N_17796,N_17919);
and U19627 (N_19627,N_17215,N_16514);
or U19628 (N_19628,N_16095,N_16777);
xor U19629 (N_19629,N_16890,N_16156);
nor U19630 (N_19630,N_17478,N_17716);
xnor U19631 (N_19631,N_16614,N_17761);
xor U19632 (N_19632,N_16653,N_17598);
and U19633 (N_19633,N_16341,N_17992);
xor U19634 (N_19634,N_16359,N_17051);
or U19635 (N_19635,N_17042,N_16131);
nor U19636 (N_19636,N_16321,N_17166);
nand U19637 (N_19637,N_17327,N_17997);
xor U19638 (N_19638,N_16959,N_17115);
or U19639 (N_19639,N_17796,N_17669);
or U19640 (N_19640,N_16082,N_17174);
xor U19641 (N_19641,N_16202,N_17862);
xnor U19642 (N_19642,N_16597,N_16900);
or U19643 (N_19643,N_16932,N_17567);
and U19644 (N_19644,N_17811,N_16872);
and U19645 (N_19645,N_16174,N_16250);
xnor U19646 (N_19646,N_17499,N_17994);
or U19647 (N_19647,N_16100,N_17641);
and U19648 (N_19648,N_17474,N_16122);
or U19649 (N_19649,N_17100,N_17429);
nand U19650 (N_19650,N_17402,N_16729);
or U19651 (N_19651,N_17949,N_17695);
and U19652 (N_19652,N_17684,N_16003);
and U19653 (N_19653,N_17753,N_16156);
nand U19654 (N_19654,N_17651,N_17205);
or U19655 (N_19655,N_17092,N_16972);
nor U19656 (N_19656,N_17284,N_16156);
xnor U19657 (N_19657,N_16059,N_16848);
and U19658 (N_19658,N_16634,N_17039);
nor U19659 (N_19659,N_16943,N_17272);
or U19660 (N_19660,N_16314,N_17310);
or U19661 (N_19661,N_17573,N_16756);
nand U19662 (N_19662,N_17232,N_16534);
nand U19663 (N_19663,N_16078,N_16984);
nand U19664 (N_19664,N_16932,N_16439);
and U19665 (N_19665,N_17776,N_16159);
or U19666 (N_19666,N_17581,N_16365);
and U19667 (N_19667,N_16704,N_17838);
nand U19668 (N_19668,N_16673,N_17493);
and U19669 (N_19669,N_16811,N_16304);
and U19670 (N_19670,N_17667,N_17346);
nand U19671 (N_19671,N_16210,N_16192);
nand U19672 (N_19672,N_17335,N_16396);
xnor U19673 (N_19673,N_16202,N_16022);
nand U19674 (N_19674,N_16003,N_16566);
or U19675 (N_19675,N_17149,N_17398);
or U19676 (N_19676,N_16332,N_17619);
nand U19677 (N_19677,N_16565,N_17544);
nand U19678 (N_19678,N_16842,N_16775);
xnor U19679 (N_19679,N_17818,N_17601);
and U19680 (N_19680,N_17530,N_17086);
nand U19681 (N_19681,N_17677,N_17567);
and U19682 (N_19682,N_16857,N_17572);
nor U19683 (N_19683,N_16013,N_17763);
nand U19684 (N_19684,N_17349,N_17667);
nor U19685 (N_19685,N_16632,N_17257);
xnor U19686 (N_19686,N_17314,N_17133);
nor U19687 (N_19687,N_17190,N_16644);
or U19688 (N_19688,N_16116,N_17633);
or U19689 (N_19689,N_17649,N_16876);
nor U19690 (N_19690,N_17399,N_17453);
nor U19691 (N_19691,N_17904,N_16854);
nand U19692 (N_19692,N_17461,N_17268);
nand U19693 (N_19693,N_16574,N_16778);
nand U19694 (N_19694,N_16741,N_16941);
nand U19695 (N_19695,N_16288,N_16115);
xnor U19696 (N_19696,N_16304,N_16734);
nand U19697 (N_19697,N_16346,N_16553);
nand U19698 (N_19698,N_16715,N_17664);
and U19699 (N_19699,N_17168,N_16945);
nor U19700 (N_19700,N_17602,N_17078);
xor U19701 (N_19701,N_16699,N_16812);
xnor U19702 (N_19702,N_17468,N_16791);
nor U19703 (N_19703,N_16720,N_17876);
or U19704 (N_19704,N_16877,N_17961);
nand U19705 (N_19705,N_17986,N_17119);
nand U19706 (N_19706,N_16663,N_16045);
xnor U19707 (N_19707,N_17678,N_17347);
nand U19708 (N_19708,N_17595,N_16886);
xnor U19709 (N_19709,N_17386,N_16498);
nand U19710 (N_19710,N_16645,N_16713);
nor U19711 (N_19711,N_17761,N_16135);
xnor U19712 (N_19712,N_17999,N_16629);
xnor U19713 (N_19713,N_16687,N_17483);
nand U19714 (N_19714,N_17078,N_17601);
or U19715 (N_19715,N_16420,N_17673);
or U19716 (N_19716,N_17644,N_17756);
and U19717 (N_19717,N_16870,N_16221);
nand U19718 (N_19718,N_16552,N_16178);
and U19719 (N_19719,N_16355,N_17172);
xor U19720 (N_19720,N_16350,N_16113);
xnor U19721 (N_19721,N_17184,N_17147);
nor U19722 (N_19722,N_17951,N_16710);
nand U19723 (N_19723,N_16959,N_16530);
nor U19724 (N_19724,N_16371,N_17756);
nand U19725 (N_19725,N_16830,N_17036);
nor U19726 (N_19726,N_17024,N_17773);
or U19727 (N_19727,N_17781,N_16777);
nor U19728 (N_19728,N_17921,N_17999);
or U19729 (N_19729,N_17937,N_17972);
nand U19730 (N_19730,N_16838,N_16845);
nand U19731 (N_19731,N_17631,N_17330);
nand U19732 (N_19732,N_16662,N_17338);
xor U19733 (N_19733,N_17255,N_16361);
nand U19734 (N_19734,N_16597,N_16573);
or U19735 (N_19735,N_17112,N_17030);
and U19736 (N_19736,N_16458,N_17889);
and U19737 (N_19737,N_17128,N_16694);
nor U19738 (N_19738,N_16598,N_17119);
or U19739 (N_19739,N_16881,N_17252);
xor U19740 (N_19740,N_17032,N_16978);
and U19741 (N_19741,N_17471,N_16072);
and U19742 (N_19742,N_16216,N_17738);
nor U19743 (N_19743,N_16917,N_17392);
nor U19744 (N_19744,N_16643,N_16481);
nand U19745 (N_19745,N_17186,N_17557);
xor U19746 (N_19746,N_16181,N_17521);
nor U19747 (N_19747,N_16967,N_17876);
nor U19748 (N_19748,N_16713,N_16962);
xnor U19749 (N_19749,N_17965,N_17682);
nand U19750 (N_19750,N_16353,N_16248);
xnor U19751 (N_19751,N_17566,N_17180);
and U19752 (N_19752,N_17489,N_17353);
or U19753 (N_19753,N_17254,N_16652);
xor U19754 (N_19754,N_17373,N_17238);
nand U19755 (N_19755,N_17024,N_17419);
and U19756 (N_19756,N_17734,N_17800);
nor U19757 (N_19757,N_16600,N_17966);
or U19758 (N_19758,N_16890,N_17327);
and U19759 (N_19759,N_16149,N_16461);
or U19760 (N_19760,N_16059,N_16945);
and U19761 (N_19761,N_16172,N_16883);
or U19762 (N_19762,N_16758,N_16754);
nor U19763 (N_19763,N_16217,N_17721);
nor U19764 (N_19764,N_16195,N_16510);
nor U19765 (N_19765,N_16404,N_16470);
nand U19766 (N_19766,N_17835,N_17775);
xnor U19767 (N_19767,N_17273,N_16107);
or U19768 (N_19768,N_17039,N_17116);
or U19769 (N_19769,N_16102,N_17707);
xnor U19770 (N_19770,N_17673,N_17923);
nand U19771 (N_19771,N_16692,N_17204);
xor U19772 (N_19772,N_17617,N_17538);
xnor U19773 (N_19773,N_17658,N_17478);
nor U19774 (N_19774,N_16687,N_16355);
or U19775 (N_19775,N_17834,N_17464);
nand U19776 (N_19776,N_17395,N_16457);
nor U19777 (N_19777,N_17980,N_16620);
or U19778 (N_19778,N_16540,N_17024);
xnor U19779 (N_19779,N_16993,N_16781);
and U19780 (N_19780,N_16406,N_16997);
nor U19781 (N_19781,N_16525,N_17583);
nor U19782 (N_19782,N_17797,N_16452);
nand U19783 (N_19783,N_16059,N_17024);
nor U19784 (N_19784,N_16118,N_17396);
nor U19785 (N_19785,N_17770,N_17311);
xnor U19786 (N_19786,N_16473,N_17422);
xnor U19787 (N_19787,N_16111,N_16583);
and U19788 (N_19788,N_16422,N_16443);
nand U19789 (N_19789,N_16376,N_16542);
or U19790 (N_19790,N_17594,N_17849);
xor U19791 (N_19791,N_17927,N_17772);
nor U19792 (N_19792,N_17037,N_17365);
and U19793 (N_19793,N_16971,N_17162);
xor U19794 (N_19794,N_16080,N_17557);
and U19795 (N_19795,N_16335,N_17339);
or U19796 (N_19796,N_17021,N_17898);
nand U19797 (N_19797,N_16038,N_17953);
or U19798 (N_19798,N_16551,N_17216);
nor U19799 (N_19799,N_16490,N_17021);
and U19800 (N_19800,N_17645,N_17474);
or U19801 (N_19801,N_17874,N_17484);
xnor U19802 (N_19802,N_17244,N_16268);
xnor U19803 (N_19803,N_17466,N_16595);
or U19804 (N_19804,N_16450,N_16473);
or U19805 (N_19805,N_17118,N_17033);
nor U19806 (N_19806,N_17201,N_17610);
nor U19807 (N_19807,N_17070,N_16813);
xnor U19808 (N_19808,N_17570,N_17694);
nand U19809 (N_19809,N_16962,N_16790);
and U19810 (N_19810,N_17673,N_16152);
nor U19811 (N_19811,N_17418,N_16400);
xnor U19812 (N_19812,N_17872,N_16979);
nor U19813 (N_19813,N_16203,N_16258);
or U19814 (N_19814,N_17683,N_16819);
nand U19815 (N_19815,N_17089,N_17164);
nor U19816 (N_19816,N_16470,N_17646);
or U19817 (N_19817,N_16813,N_17323);
nor U19818 (N_19818,N_17942,N_17650);
or U19819 (N_19819,N_16646,N_16582);
or U19820 (N_19820,N_17849,N_17707);
nand U19821 (N_19821,N_17802,N_16937);
xnor U19822 (N_19822,N_16621,N_16323);
nand U19823 (N_19823,N_16233,N_16613);
or U19824 (N_19824,N_16719,N_17416);
nor U19825 (N_19825,N_16431,N_17450);
and U19826 (N_19826,N_16861,N_17290);
nor U19827 (N_19827,N_17667,N_17208);
nor U19828 (N_19828,N_16618,N_16277);
nand U19829 (N_19829,N_17569,N_17637);
or U19830 (N_19830,N_17274,N_16664);
or U19831 (N_19831,N_17482,N_16541);
nor U19832 (N_19832,N_17948,N_16197);
and U19833 (N_19833,N_17685,N_16542);
and U19834 (N_19834,N_16681,N_16345);
or U19835 (N_19835,N_17596,N_17095);
nor U19836 (N_19836,N_17636,N_17984);
nor U19837 (N_19837,N_16621,N_16225);
or U19838 (N_19838,N_16433,N_16078);
xnor U19839 (N_19839,N_17219,N_17305);
nor U19840 (N_19840,N_17613,N_17182);
nand U19841 (N_19841,N_17086,N_17642);
xnor U19842 (N_19842,N_17847,N_17088);
nand U19843 (N_19843,N_17023,N_17163);
and U19844 (N_19844,N_17676,N_16299);
nor U19845 (N_19845,N_17129,N_17110);
or U19846 (N_19846,N_16993,N_16367);
or U19847 (N_19847,N_16618,N_16367);
or U19848 (N_19848,N_17879,N_17226);
nor U19849 (N_19849,N_16920,N_16310);
or U19850 (N_19850,N_16820,N_16855);
or U19851 (N_19851,N_17170,N_17252);
xnor U19852 (N_19852,N_16256,N_16452);
nor U19853 (N_19853,N_17089,N_16877);
and U19854 (N_19854,N_17962,N_16839);
and U19855 (N_19855,N_17892,N_16053);
nand U19856 (N_19856,N_17790,N_16961);
or U19857 (N_19857,N_16256,N_17086);
and U19858 (N_19858,N_17466,N_16080);
nand U19859 (N_19859,N_17971,N_17098);
xnor U19860 (N_19860,N_17510,N_16356);
or U19861 (N_19861,N_17027,N_16970);
nand U19862 (N_19862,N_17815,N_16881);
xor U19863 (N_19863,N_16492,N_16928);
xor U19864 (N_19864,N_17079,N_16617);
nor U19865 (N_19865,N_16294,N_17991);
and U19866 (N_19866,N_17980,N_16889);
or U19867 (N_19867,N_17219,N_17978);
and U19868 (N_19868,N_17097,N_17008);
xor U19869 (N_19869,N_16400,N_17933);
or U19870 (N_19870,N_17330,N_16678);
nor U19871 (N_19871,N_17576,N_16236);
nor U19872 (N_19872,N_16911,N_17646);
or U19873 (N_19873,N_16935,N_17744);
or U19874 (N_19874,N_16925,N_17558);
and U19875 (N_19875,N_17050,N_16036);
nand U19876 (N_19876,N_16448,N_16624);
nand U19877 (N_19877,N_17538,N_16154);
and U19878 (N_19878,N_17452,N_17541);
nand U19879 (N_19879,N_16296,N_16662);
nor U19880 (N_19880,N_17318,N_17494);
nand U19881 (N_19881,N_17428,N_16899);
nand U19882 (N_19882,N_17618,N_17643);
or U19883 (N_19883,N_17760,N_16145);
and U19884 (N_19884,N_17627,N_16835);
nand U19885 (N_19885,N_16264,N_16203);
or U19886 (N_19886,N_17179,N_17565);
xnor U19887 (N_19887,N_16306,N_16597);
and U19888 (N_19888,N_17661,N_16641);
and U19889 (N_19889,N_17193,N_16271);
or U19890 (N_19890,N_16630,N_17380);
nand U19891 (N_19891,N_16441,N_17100);
and U19892 (N_19892,N_16650,N_16067);
or U19893 (N_19893,N_17197,N_17451);
and U19894 (N_19894,N_16641,N_17308);
nand U19895 (N_19895,N_17339,N_16118);
or U19896 (N_19896,N_17824,N_17672);
xor U19897 (N_19897,N_17468,N_16758);
nor U19898 (N_19898,N_17751,N_17854);
or U19899 (N_19899,N_16149,N_16765);
or U19900 (N_19900,N_17743,N_16248);
xnor U19901 (N_19901,N_17078,N_17503);
xor U19902 (N_19902,N_17788,N_17914);
or U19903 (N_19903,N_16482,N_17515);
or U19904 (N_19904,N_16520,N_17754);
or U19905 (N_19905,N_17147,N_17926);
and U19906 (N_19906,N_16156,N_16107);
nand U19907 (N_19907,N_16180,N_16271);
nand U19908 (N_19908,N_16095,N_17659);
nor U19909 (N_19909,N_17947,N_17090);
xor U19910 (N_19910,N_16881,N_16304);
nor U19911 (N_19911,N_17904,N_17259);
xnor U19912 (N_19912,N_17971,N_17225);
or U19913 (N_19913,N_17125,N_17025);
nor U19914 (N_19914,N_16096,N_16396);
or U19915 (N_19915,N_16704,N_16180);
or U19916 (N_19916,N_16575,N_16686);
and U19917 (N_19917,N_16403,N_16502);
xor U19918 (N_19918,N_16157,N_16203);
nor U19919 (N_19919,N_16433,N_16482);
and U19920 (N_19920,N_17199,N_16159);
or U19921 (N_19921,N_17575,N_17078);
and U19922 (N_19922,N_16797,N_17027);
nor U19923 (N_19923,N_16738,N_17796);
xor U19924 (N_19924,N_17031,N_17552);
xnor U19925 (N_19925,N_17405,N_17682);
and U19926 (N_19926,N_17927,N_17890);
and U19927 (N_19927,N_16730,N_17583);
nor U19928 (N_19928,N_16384,N_16489);
nand U19929 (N_19929,N_16792,N_17172);
nor U19930 (N_19930,N_17833,N_16448);
nand U19931 (N_19931,N_17501,N_16914);
nor U19932 (N_19932,N_17909,N_16828);
xor U19933 (N_19933,N_16709,N_17616);
nand U19934 (N_19934,N_16877,N_16505);
xor U19935 (N_19935,N_17450,N_16202);
and U19936 (N_19936,N_17310,N_17181);
xor U19937 (N_19937,N_16913,N_16364);
nand U19938 (N_19938,N_17859,N_16586);
or U19939 (N_19939,N_16964,N_17087);
nor U19940 (N_19940,N_17856,N_17377);
xor U19941 (N_19941,N_17094,N_17864);
nor U19942 (N_19942,N_17268,N_17336);
xnor U19943 (N_19943,N_16944,N_16566);
and U19944 (N_19944,N_16710,N_17811);
nand U19945 (N_19945,N_16831,N_17365);
and U19946 (N_19946,N_17105,N_17929);
and U19947 (N_19947,N_17537,N_16521);
nand U19948 (N_19948,N_16512,N_17486);
and U19949 (N_19949,N_17550,N_16670);
and U19950 (N_19950,N_17661,N_17105);
xor U19951 (N_19951,N_17846,N_17354);
nor U19952 (N_19952,N_17209,N_16337);
or U19953 (N_19953,N_17692,N_16477);
or U19954 (N_19954,N_16528,N_17279);
or U19955 (N_19955,N_17415,N_17106);
or U19956 (N_19956,N_16999,N_17099);
nor U19957 (N_19957,N_17637,N_16840);
or U19958 (N_19958,N_16123,N_16391);
xnor U19959 (N_19959,N_17726,N_17977);
xnor U19960 (N_19960,N_17340,N_16292);
nand U19961 (N_19961,N_16350,N_17173);
or U19962 (N_19962,N_17957,N_16198);
xor U19963 (N_19963,N_17267,N_16667);
xnor U19964 (N_19964,N_17722,N_17158);
and U19965 (N_19965,N_17711,N_16073);
or U19966 (N_19966,N_16888,N_16151);
xor U19967 (N_19967,N_17370,N_16394);
nand U19968 (N_19968,N_16684,N_17220);
nor U19969 (N_19969,N_17616,N_16839);
or U19970 (N_19970,N_16380,N_16997);
nand U19971 (N_19971,N_17114,N_17801);
nand U19972 (N_19972,N_17095,N_17075);
nor U19973 (N_19973,N_17065,N_17547);
nand U19974 (N_19974,N_17726,N_16132);
or U19975 (N_19975,N_16032,N_17956);
nor U19976 (N_19976,N_17994,N_16432);
xor U19977 (N_19977,N_17683,N_17306);
and U19978 (N_19978,N_17224,N_17871);
and U19979 (N_19979,N_16725,N_17795);
xnor U19980 (N_19980,N_16635,N_17950);
or U19981 (N_19981,N_17582,N_17212);
nor U19982 (N_19982,N_16964,N_17355);
nor U19983 (N_19983,N_17789,N_16838);
or U19984 (N_19984,N_17567,N_16730);
nor U19985 (N_19985,N_17662,N_16928);
or U19986 (N_19986,N_17734,N_16076);
nor U19987 (N_19987,N_17947,N_17876);
nor U19988 (N_19988,N_16909,N_16853);
nand U19989 (N_19989,N_17345,N_16611);
or U19990 (N_19990,N_16755,N_17785);
and U19991 (N_19991,N_16419,N_17211);
xor U19992 (N_19992,N_17697,N_16676);
or U19993 (N_19993,N_17590,N_16671);
or U19994 (N_19994,N_16307,N_16607);
xor U19995 (N_19995,N_16237,N_17066);
xor U19996 (N_19996,N_16024,N_17895);
or U19997 (N_19997,N_16153,N_17083);
nand U19998 (N_19998,N_16308,N_16624);
xnor U19999 (N_19999,N_16736,N_16616);
xor U20000 (N_20000,N_19293,N_18546);
nand U20001 (N_20001,N_18919,N_19927);
xnor U20002 (N_20002,N_18849,N_19942);
nand U20003 (N_20003,N_18569,N_18840);
or U20004 (N_20004,N_19678,N_18627);
and U20005 (N_20005,N_19684,N_18054);
nand U20006 (N_20006,N_18322,N_19598);
or U20007 (N_20007,N_18685,N_18346);
and U20008 (N_20008,N_18571,N_18532);
nor U20009 (N_20009,N_19994,N_19680);
and U20010 (N_20010,N_18999,N_19246);
nor U20011 (N_20011,N_19581,N_19758);
nand U20012 (N_20012,N_19075,N_19998);
and U20013 (N_20013,N_19802,N_18312);
and U20014 (N_20014,N_18468,N_19688);
nand U20015 (N_20015,N_18835,N_19773);
nor U20016 (N_20016,N_18824,N_19567);
nand U20017 (N_20017,N_19182,N_18146);
nor U20018 (N_20018,N_19560,N_19670);
xnor U20019 (N_20019,N_18708,N_19760);
and U20020 (N_20020,N_19025,N_19762);
nand U20021 (N_20021,N_18517,N_19558);
nand U20022 (N_20022,N_19769,N_19072);
xor U20023 (N_20023,N_18389,N_19894);
nor U20024 (N_20024,N_19779,N_18747);
or U20025 (N_20025,N_18308,N_19727);
or U20026 (N_20026,N_18189,N_18327);
and U20027 (N_20027,N_19631,N_18917);
and U20028 (N_20028,N_19857,N_18429);
nor U20029 (N_20029,N_19124,N_18832);
nor U20030 (N_20030,N_19549,N_19990);
and U20031 (N_20031,N_19322,N_19430);
nor U20032 (N_20032,N_18823,N_19064);
xor U20033 (N_20033,N_18127,N_18606);
nor U20034 (N_20034,N_18581,N_18080);
nor U20035 (N_20035,N_19589,N_18420);
or U20036 (N_20036,N_19432,N_19556);
and U20037 (N_20037,N_19867,N_19939);
or U20038 (N_20038,N_19775,N_19256);
xnor U20039 (N_20039,N_18197,N_19418);
and U20040 (N_20040,N_18720,N_18195);
nand U20041 (N_20041,N_19685,N_18169);
and U20042 (N_20042,N_18699,N_18210);
nand U20043 (N_20043,N_18001,N_19711);
or U20044 (N_20044,N_19066,N_18249);
nor U20045 (N_20045,N_19453,N_19481);
nor U20046 (N_20046,N_18303,N_18209);
and U20047 (N_20047,N_18120,N_18461);
nand U20048 (N_20048,N_18180,N_18175);
nand U20049 (N_20049,N_19340,N_19706);
nor U20050 (N_20050,N_18889,N_19753);
nor U20051 (N_20051,N_18271,N_18930);
or U20052 (N_20052,N_19111,N_19972);
and U20053 (N_20053,N_19341,N_18914);
and U20054 (N_20054,N_19180,N_19236);
xor U20055 (N_20055,N_19726,N_19023);
xnor U20056 (N_20056,N_18050,N_18217);
nand U20057 (N_20057,N_18753,N_19737);
and U20058 (N_20058,N_18070,N_18359);
nor U20059 (N_20059,N_19744,N_18423);
xor U20060 (N_20060,N_19539,N_19468);
xnor U20061 (N_20061,N_19980,N_18960);
nor U20062 (N_20062,N_19687,N_19291);
nand U20063 (N_20063,N_19877,N_19208);
xor U20064 (N_20064,N_18990,N_18037);
and U20065 (N_20065,N_19082,N_19100);
nand U20066 (N_20066,N_19911,N_18785);
or U20067 (N_20067,N_19078,N_19168);
or U20068 (N_20068,N_19908,N_19020);
or U20069 (N_20069,N_19081,N_18230);
nor U20070 (N_20070,N_18506,N_19067);
nand U20071 (N_20071,N_18640,N_19542);
or U20072 (N_20072,N_18036,N_18148);
nor U20073 (N_20073,N_18595,N_18692);
or U20074 (N_20074,N_18323,N_18582);
xnor U20075 (N_20075,N_18167,N_19467);
and U20076 (N_20076,N_18847,N_19752);
and U20077 (N_20077,N_18244,N_18969);
and U20078 (N_20078,N_18728,N_18207);
xnor U20079 (N_20079,N_19610,N_19056);
or U20080 (N_20080,N_19105,N_18259);
nor U20081 (N_20081,N_19130,N_18289);
and U20082 (N_20082,N_18239,N_18181);
nand U20083 (N_20083,N_18915,N_18446);
xnor U20084 (N_20084,N_18187,N_19645);
or U20085 (N_20085,N_19926,N_19283);
or U20086 (N_20086,N_19826,N_19335);
and U20087 (N_20087,N_19673,N_18311);
or U20088 (N_20088,N_18428,N_19561);
nor U20089 (N_20089,N_18220,N_18851);
or U20090 (N_20090,N_19698,N_18669);
and U20091 (N_20091,N_19320,N_18119);
or U20092 (N_20092,N_19859,N_18283);
and U20093 (N_20093,N_18171,N_19931);
nand U20094 (N_20094,N_18503,N_18224);
nand U20095 (N_20095,N_18857,N_18122);
nand U20096 (N_20096,N_18719,N_19494);
xnor U20097 (N_20097,N_18584,N_18600);
xnor U20098 (N_20098,N_18649,N_19250);
nor U20099 (N_20099,N_19169,N_19951);
and U20100 (N_20100,N_19203,N_18853);
nand U20101 (N_20101,N_19328,N_18592);
nand U20102 (N_20102,N_19640,N_19805);
nand U20103 (N_20103,N_19748,N_18309);
xnor U20104 (N_20104,N_18299,N_18878);
xor U20105 (N_20105,N_18086,N_18547);
nor U20106 (N_20106,N_18644,N_19351);
or U20107 (N_20107,N_18011,N_19646);
xor U20108 (N_20108,N_19836,N_19407);
or U20109 (N_20109,N_19162,N_19772);
nor U20110 (N_20110,N_19833,N_18602);
xor U20111 (N_20111,N_19403,N_18085);
and U20112 (N_20112,N_19152,N_18399);
nand U20113 (N_20113,N_19574,N_18083);
and U20114 (N_20114,N_18324,N_18464);
nand U20115 (N_20115,N_18158,N_19912);
xnor U20116 (N_20116,N_19932,N_19683);
nand U20117 (N_20117,N_18129,N_19822);
nand U20118 (N_20118,N_18727,N_19039);
nor U20119 (N_20119,N_18937,N_18409);
nor U20120 (N_20120,N_19551,N_18372);
and U20121 (N_20121,N_18163,N_19317);
nor U20122 (N_20122,N_18069,N_18347);
and U20123 (N_20123,N_19720,N_18485);
nand U20124 (N_20124,N_19140,N_19393);
and U20125 (N_20125,N_18936,N_19557);
nand U20126 (N_20126,N_18358,N_18174);
nor U20127 (N_20127,N_18901,N_18340);
nor U20128 (N_20128,N_18710,N_18918);
nand U20129 (N_20129,N_18132,N_19389);
nor U20130 (N_20130,N_18574,N_18599);
nor U20131 (N_20131,N_18381,N_18457);
xnor U20132 (N_20132,N_19710,N_19435);
or U20133 (N_20133,N_18537,N_18084);
xor U20134 (N_20134,N_18670,N_19968);
or U20135 (N_20135,N_18360,N_19623);
nor U20136 (N_20136,N_19840,N_18596);
or U20137 (N_20137,N_18892,N_18183);
nor U20138 (N_20138,N_19944,N_19212);
and U20139 (N_20139,N_18248,N_18388);
or U20140 (N_20140,N_18726,N_19599);
and U20141 (N_20141,N_18612,N_19423);
and U20142 (N_20142,N_19337,N_19218);
xnor U20143 (N_20143,N_18135,N_19537);
xor U20144 (N_20144,N_18405,N_18236);
xor U20145 (N_20145,N_19902,N_18293);
nor U20146 (N_20146,N_19545,N_18425);
nand U20147 (N_20147,N_18868,N_18958);
or U20148 (N_20148,N_19451,N_18711);
xor U20149 (N_20149,N_19641,N_19483);
nor U20150 (N_20150,N_18630,N_19178);
nor U20151 (N_20151,N_18752,N_18281);
nand U20152 (N_20152,N_18385,N_19681);
and U20153 (N_20153,N_19277,N_19976);
and U20154 (N_20154,N_18294,N_19366);
and U20155 (N_20155,N_19898,N_18679);
or U20156 (N_20156,N_19864,N_18774);
or U20157 (N_20157,N_19500,N_19047);
and U20158 (N_20158,N_18557,N_18314);
nand U20159 (N_20159,N_18900,N_18106);
or U20160 (N_20160,N_19866,N_19970);
nand U20161 (N_20161,N_19149,N_18343);
nand U20162 (N_20162,N_19353,N_18512);
and U20163 (N_20163,N_19440,N_18306);
xor U20164 (N_20164,N_19632,N_18020);
or U20165 (N_20165,N_19264,N_18071);
nand U20166 (N_20166,N_19831,N_19402);
or U20167 (N_20167,N_18952,N_19835);
and U20168 (N_20168,N_19127,N_18641);
or U20169 (N_20169,N_19458,N_18583);
and U20170 (N_20170,N_18540,N_19071);
nor U20171 (N_20171,N_18435,N_19445);
or U20172 (N_20172,N_18904,N_19904);
or U20173 (N_20173,N_18304,N_18921);
or U20174 (N_20174,N_19181,N_19801);
or U20175 (N_20175,N_18130,N_19583);
nor U20176 (N_20176,N_18784,N_18791);
or U20177 (N_20177,N_18162,N_19425);
nor U20178 (N_20178,N_19281,N_19906);
and U20179 (N_20179,N_19997,N_18707);
nand U20180 (N_20180,N_18643,N_18749);
or U20181 (N_20181,N_18103,N_19154);
nand U20182 (N_20182,N_18782,N_18221);
or U20183 (N_20183,N_19136,N_18615);
nand U20184 (N_20184,N_19333,N_19210);
nand U20185 (N_20185,N_18943,N_18780);
and U20186 (N_20186,N_19360,N_18042);
or U20187 (N_20187,N_19702,N_18535);
nand U20188 (N_20188,N_18855,N_18695);
nand U20189 (N_20189,N_19068,N_19963);
xnor U20190 (N_20190,N_18396,N_19249);
nor U20191 (N_20191,N_19234,N_19095);
nand U20192 (N_20192,N_18959,N_19295);
and U20193 (N_20193,N_18502,N_19666);
nand U20194 (N_20194,N_19480,N_19695);
and U20195 (N_20195,N_19883,N_19579);
xnor U20196 (N_20196,N_19416,N_18745);
nor U20197 (N_20197,N_19251,N_18949);
nor U20198 (N_20198,N_19575,N_18687);
nor U20199 (N_20199,N_19848,N_19896);
and U20200 (N_20200,N_18625,N_18539);
nor U20201 (N_20201,N_19312,N_18718);
nor U20202 (N_20202,N_18704,N_19895);
nor U20203 (N_20203,N_19431,N_18763);
or U20204 (N_20204,N_18934,N_18986);
xnor U20205 (N_20205,N_19934,N_18770);
nor U20206 (N_20206,N_19400,N_19396);
xnor U20207 (N_20207,N_18160,N_19187);
and U20208 (N_20208,N_18508,N_19648);
or U20209 (N_20209,N_19446,N_18626);
and U20210 (N_20210,N_18184,N_19070);
nor U20211 (N_20211,N_18672,N_19390);
xor U20212 (N_20212,N_19099,N_19655);
and U20213 (N_20213,N_19290,N_18074);
nand U20214 (N_20214,N_19030,N_18144);
nand U20215 (N_20215,N_19365,N_19049);
nor U20216 (N_20216,N_19671,N_19215);
or U20217 (N_20217,N_19343,N_19043);
or U20218 (N_20218,N_18864,N_18920);
xor U20219 (N_20219,N_19986,N_19201);
nand U20220 (N_20220,N_18484,N_18497);
and U20221 (N_20221,N_18676,N_19224);
nor U20222 (N_20222,N_19311,N_19767);
and U20223 (N_20223,N_19868,N_19816);
or U20224 (N_20224,N_19382,N_19026);
or U20225 (N_20225,N_18737,N_18262);
or U20226 (N_20226,N_19113,N_18393);
nand U20227 (N_20227,N_19268,N_18362);
nor U20228 (N_20228,N_19958,N_19634);
nand U20229 (N_20229,N_18964,N_19091);
nor U20230 (N_20230,N_19288,N_19624);
xor U20231 (N_20231,N_19447,N_19792);
xnor U20232 (N_20232,N_18471,N_19949);
and U20233 (N_20233,N_18452,N_19809);
xnor U20234 (N_20234,N_18227,N_19263);
xnor U20235 (N_20235,N_19073,N_19369);
nand U20236 (N_20236,N_19090,N_18049);
xor U20237 (N_20237,N_19576,N_19886);
or U20238 (N_20238,N_18716,N_19144);
nor U20239 (N_20239,N_18002,N_18081);
nor U20240 (N_20240,N_18177,N_18783);
nand U20241 (N_20241,N_18666,N_19229);
nor U20242 (N_20242,N_19392,N_18712);
nor U20243 (N_20243,N_19231,N_18993);
xor U20244 (N_20244,N_19935,N_19057);
and U20245 (N_20245,N_19338,N_18430);
xnor U20246 (N_20246,N_18799,N_18825);
nor U20247 (N_20247,N_18056,N_19409);
or U20248 (N_20248,N_19945,N_19652);
or U20249 (N_20249,N_19804,N_19987);
nand U20250 (N_20250,N_18565,N_19692);
xor U20251 (N_20251,N_19928,N_19289);
nor U20252 (N_20252,N_19045,N_19088);
and U20253 (N_20253,N_18809,N_18156);
nor U20254 (N_20254,N_19035,N_19241);
and U20255 (N_20255,N_18821,N_19862);
nand U20256 (N_20256,N_18524,N_19044);
and U20257 (N_20257,N_18141,N_19190);
nand U20258 (N_20258,N_18639,N_18820);
and U20259 (N_20259,N_18058,N_19490);
or U20260 (N_20260,N_19211,N_18664);
or U20261 (N_20261,N_19741,N_18881);
and U20262 (N_20262,N_19243,N_18651);
nand U20263 (N_20263,N_18637,N_19391);
nand U20264 (N_20264,N_19721,N_19514);
and U20265 (N_20265,N_19342,N_19011);
and U20266 (N_20266,N_18115,N_18223);
nor U20267 (N_20267,N_19093,N_18948);
nand U20268 (N_20268,N_19756,N_19461);
nand U20269 (N_20269,N_19334,N_19098);
nand U20270 (N_20270,N_18498,N_18678);
or U20271 (N_20271,N_19959,N_18590);
or U20272 (N_20272,N_18991,N_18538);
and U20273 (N_20273,N_19206,N_18761);
xnor U20274 (N_20274,N_18872,N_19327);
nor U20275 (N_20275,N_19660,N_19584);
or U20276 (N_20276,N_18449,N_19000);
or U20277 (N_20277,N_18586,N_18269);
xnor U20278 (N_20278,N_18732,N_18758);
xor U20279 (N_20279,N_18336,N_19853);
and U20280 (N_20280,N_18795,N_18977);
or U20281 (N_20281,N_18234,N_19903);
and U20282 (N_20282,N_18767,N_19257);
or U20283 (N_20283,N_18033,N_18505);
and U20284 (N_20284,N_19719,N_18124);
xor U20285 (N_20285,N_19530,N_19807);
xnor U20286 (N_20286,N_19374,N_19621);
nand U20287 (N_20287,N_19601,N_18924);
xor U20288 (N_20288,N_19475,N_19725);
xnor U20289 (N_20289,N_18113,N_19981);
and U20290 (N_20290,N_18355,N_18885);
or U20291 (N_20291,N_18973,N_18241);
and U20292 (N_20292,N_19254,N_18076);
xnor U20293 (N_20293,N_19937,N_18316);
xor U20294 (N_20294,N_19298,N_18077);
or U20295 (N_20295,N_18700,N_19485);
xnor U20296 (N_20296,N_18196,N_19259);
xnor U20297 (N_20297,N_18317,N_19129);
and U20298 (N_20298,N_18198,N_19300);
nor U20299 (N_20299,N_18302,N_18380);
or U20300 (N_20300,N_18989,N_19377);
nor U20301 (N_20301,N_18650,N_18418);
nor U20302 (N_20302,N_19993,N_19543);
and U20303 (N_20303,N_18486,N_18140);
nor U20304 (N_20304,N_18490,N_18812);
and U20305 (N_20305,N_19803,N_18378);
or U20306 (N_20306,N_18671,N_19768);
nand U20307 (N_20307,N_19754,N_18143);
or U20308 (N_20308,N_18007,N_18473);
and U20309 (N_20309,N_18255,N_18391);
nor U20310 (N_20310,N_19414,N_19618);
xor U20311 (N_20311,N_19214,N_19386);
or U20312 (N_20312,N_19996,N_18172);
or U20313 (N_20313,N_19008,N_18897);
nand U20314 (N_20314,N_19107,N_19914);
nand U20315 (N_20315,N_19294,N_19370);
nor U20316 (N_20316,N_19110,N_18604);
or U20317 (N_20317,N_19448,N_18291);
or U20318 (N_20318,N_18724,N_19844);
or U20319 (N_20319,N_18845,N_18587);
or U20320 (N_20320,N_19787,N_19131);
xnor U20321 (N_20321,N_18520,N_19971);
nand U20322 (N_20322,N_19395,N_18890);
or U20323 (N_20323,N_18110,N_19006);
and U20324 (N_20324,N_19689,N_18815);
nand U20325 (N_20325,N_18088,N_19122);
and U20326 (N_20326,N_19843,N_19094);
nand U20327 (N_20327,N_19955,N_19983);
xnor U20328 (N_20328,N_18191,N_18290);
nand U20329 (N_20329,N_18658,N_18102);
nor U20330 (N_20330,N_19650,N_19001);
nor U20331 (N_20331,N_18739,N_19845);
nor U20332 (N_20332,N_19554,N_19097);
xnor U20333 (N_20333,N_18798,N_19329);
nor U20334 (N_20334,N_18364,N_19399);
xnor U20335 (N_20335,N_18017,N_18746);
or U20336 (N_20336,N_18038,N_18453);
xor U20337 (N_20337,N_18242,N_18427);
and U20338 (N_20338,N_19513,N_19946);
and U20339 (N_20339,N_19145,N_18014);
or U20340 (N_20340,N_19040,N_18376);
or U20341 (N_20341,N_18764,N_19989);
xor U20342 (N_20342,N_18475,N_18178);
xor U20343 (N_20343,N_18865,N_18318);
xor U20344 (N_20344,N_19137,N_19882);
nand U20345 (N_20345,N_18591,N_18722);
xor U20346 (N_20346,N_19018,N_19273);
xor U20347 (N_20347,N_18480,N_19498);
xor U20348 (N_20348,N_19383,N_19552);
nand U20349 (N_20349,N_19315,N_19757);
nand U20350 (N_20350,N_18802,N_19367);
or U20351 (N_20351,N_19879,N_18603);
or U20352 (N_20352,N_19235,N_18394);
nand U20353 (N_20353,N_19087,N_19260);
nor U20354 (N_20354,N_19270,N_18775);
nand U20355 (N_20355,N_18450,N_19454);
or U20356 (N_20356,N_19482,N_18168);
or U20357 (N_20357,N_19510,N_19196);
nor U20358 (N_20358,N_19069,N_18375);
and U20359 (N_20359,N_18947,N_19881);
nor U20360 (N_20360,N_19507,N_19967);
nand U20361 (N_20361,N_19774,N_18597);
xnor U20362 (N_20362,N_19724,N_19707);
nand U20363 (N_20363,N_19755,N_19799);
or U20364 (N_20364,N_18663,N_19776);
nor U20365 (N_20365,N_19922,N_18944);
xor U20366 (N_20366,N_18622,N_18448);
or U20367 (N_20367,N_18406,N_18212);
and U20368 (N_20368,N_18577,N_18580);
or U20369 (N_20369,N_19887,N_19873);
nor U20370 (N_20370,N_18624,N_18267);
or U20371 (N_20371,N_18877,N_18706);
nor U20372 (N_20372,N_19874,N_19905);
xor U20373 (N_20373,N_19427,N_19207);
or U20374 (N_20374,N_18957,N_18190);
nor U20375 (N_20375,N_18206,N_18933);
nand U20376 (N_20376,N_19258,N_18982);
and U20377 (N_20377,N_18981,N_19139);
or U20378 (N_20378,N_19723,N_18431);
nand U20379 (N_20379,N_19420,N_18811);
or U20380 (N_20380,N_19248,N_19920);
nand U20381 (N_20381,N_18186,N_19718);
xnor U20382 (N_20382,N_18558,N_18608);
and U20383 (N_20383,N_19825,N_19793);
nand U20384 (N_20384,N_19021,N_19999);
xor U20385 (N_20385,N_19488,N_18810);
xnor U20386 (N_20386,N_18536,N_18713);
xnor U20387 (N_20387,N_19349,N_18564);
and U20388 (N_20388,N_19104,N_18776);
or U20389 (N_20389,N_19385,N_18866);
xor U20390 (N_20390,N_19063,N_18734);
nor U20391 (N_20391,N_18252,N_19603);
nor U20392 (N_20392,N_18545,N_18032);
and U20393 (N_20393,N_19036,N_19703);
and U20394 (N_20394,N_18500,N_18023);
nand U20395 (N_20395,N_18805,N_18585);
nor U20396 (N_20396,N_18170,N_18852);
and U20397 (N_20397,N_18413,N_19850);
xor U20398 (N_20398,N_18016,N_19166);
nor U20399 (N_20399,N_18467,N_18554);
xor U20400 (N_20400,N_19153,N_18751);
nand U20401 (N_20401,N_18407,N_19496);
xnor U20402 (N_20402,N_19050,N_19279);
nand U20403 (N_20403,N_19694,N_18688);
nor U20404 (N_20404,N_18109,N_19643);
xor U20405 (N_20405,N_19160,N_18908);
xor U20406 (N_20406,N_18082,N_18041);
xnor U20407 (N_20407,N_19974,N_19619);
nor U20408 (N_20408,N_19272,N_19607);
xnor U20409 (N_20409,N_19841,N_18909);
and U20410 (N_20410,N_19463,N_18647);
or U20411 (N_20411,N_18287,N_18436);
nand U20412 (N_20412,N_19125,N_18131);
nor U20413 (N_20413,N_18522,N_19204);
xor U20414 (N_20414,N_19456,N_19376);
xnor U20415 (N_20415,N_19265,N_19674);
and U20416 (N_20416,N_19676,N_19037);
and U20417 (N_20417,N_18528,N_19795);
nor U20418 (N_20418,N_19714,N_19318);
nor U20419 (N_20419,N_19661,N_19875);
xor U20420 (N_20420,N_18594,N_19076);
or U20421 (N_20421,N_19146,N_18326);
and U20422 (N_20422,N_19261,N_18395);
nor U20423 (N_20423,N_19740,N_18208);
or U20424 (N_20424,N_19709,N_19956);
nor U20425 (N_20425,N_19770,N_19854);
nor U20426 (N_20426,N_19665,N_18321);
or U20427 (N_20427,N_18319,N_19474);
nor U20428 (N_20428,N_19637,N_18310);
nor U20429 (N_20429,N_18863,N_18035);
or U20430 (N_20430,N_18862,N_18465);
or U20431 (N_20431,N_19192,N_18705);
nand U20432 (N_20432,N_19228,N_19915);
and U20433 (N_20433,N_19116,N_18185);
nand U20434 (N_20434,N_19789,N_18495);
nor U20435 (N_20435,N_19749,N_18344);
nor U20436 (N_20436,N_18066,N_19222);
and U20437 (N_20437,N_19114,N_18850);
and U20438 (N_20438,N_18839,N_18786);
or U20439 (N_20439,N_19988,N_19041);
or U20440 (N_20440,N_18416,N_18955);
and U20441 (N_20441,N_18356,N_18368);
and U20442 (N_20442,N_19005,N_18985);
or U20443 (N_20443,N_18556,N_19910);
xor U20444 (N_20444,N_19553,N_18510);
nand U20445 (N_20445,N_19642,N_18563);
and U20446 (N_20446,N_19083,N_18087);
nor U20447 (N_20447,N_19991,N_18962);
or U20448 (N_20448,N_18442,N_19628);
and U20449 (N_20449,N_19582,N_19060);
nor U20450 (N_20450,N_19715,N_19232);
or U20451 (N_20451,N_19960,N_19829);
xor U20452 (N_20452,N_18126,N_18149);
nand U20453 (N_20453,N_19388,N_19185);
or U20454 (N_20454,N_18794,N_19616);
nand U20455 (N_20455,N_18633,N_19027);
nor U20456 (N_20456,N_19278,N_18731);
or U20457 (N_20457,N_19171,N_19531);
nor U20458 (N_20458,N_18527,N_18494);
xor U20459 (N_20459,N_19230,N_18741);
nand U20460 (N_20460,N_19449,N_18004);
and U20461 (N_20461,N_18634,N_18218);
or U20462 (N_20462,N_19119,N_18329);
xnor U20463 (N_20463,N_19512,N_19470);
nand U20464 (N_20464,N_18463,N_18523);
and U20465 (N_20465,N_18137,N_19526);
nand U20466 (N_20466,N_18501,N_19763);
nand U20467 (N_20467,N_18292,N_18027);
or U20468 (N_20468,N_18157,N_18736);
and U20469 (N_20469,N_19085,N_18531);
and U20470 (N_20470,N_18469,N_19699);
or U20471 (N_20471,N_19953,N_19310);
and U20472 (N_20472,N_18243,N_19301);
or U20473 (N_20473,N_19032,N_19269);
xor U20474 (N_20474,N_18907,N_19141);
xnor U20475 (N_20475,N_19319,N_18974);
nor U20476 (N_20476,N_19364,N_18946);
and U20477 (N_20477,N_19436,N_18929);
or U20478 (N_20478,N_19062,N_19471);
xor U20479 (N_20479,N_18858,N_18279);
nand U20480 (N_20480,N_19533,N_19863);
nand U20481 (N_20481,N_19856,N_18458);
nor U20482 (N_20482,N_19849,N_19499);
and U20483 (N_20483,N_18213,N_18827);
or U20484 (N_20484,N_18661,N_19569);
xnor U20485 (N_20485,N_19159,N_18108);
or U20486 (N_20486,N_18397,N_19653);
and U20487 (N_20487,N_19079,N_18880);
and U20488 (N_20488,N_18579,N_18911);
or U20489 (N_20489,N_19356,N_18682);
nand U20490 (N_20490,N_19964,N_19452);
or U20491 (N_20491,N_18348,N_18338);
and U20492 (N_20492,N_19084,N_18193);
xnor U20493 (N_20493,N_19693,N_19275);
or U20494 (N_20494,N_19817,N_19484);
nand U20495 (N_20495,N_18951,N_19151);
and U20496 (N_20496,N_19913,N_19712);
nor U20497 (N_20497,N_18462,N_18601);
and U20498 (N_20498,N_18489,N_19143);
nor U20499 (N_20499,N_18118,N_19780);
nand U20500 (N_20500,N_19823,N_18575);
or U20501 (N_20501,N_19307,N_18927);
nor U20502 (N_20502,N_19878,N_19975);
nand U20503 (N_20503,N_18142,N_18572);
or U20504 (N_20504,N_18100,N_19924);
xnor U20505 (N_20505,N_18961,N_18470);
xnor U20506 (N_20506,N_19532,N_18836);
or U20507 (N_20507,N_19292,N_18367);
nand U20508 (N_20508,N_19359,N_19834);
and U20509 (N_20509,N_18040,N_19200);
nor U20510 (N_20510,N_19751,N_18683);
or U20511 (N_20511,N_19003,N_19861);
xnor U20512 (N_20512,N_19808,N_18226);
nor U20513 (N_20513,N_18478,N_18806);
xor U20514 (N_20514,N_19033,N_18440);
nand U20515 (N_20515,N_18529,N_18605);
or U20516 (N_20516,N_19839,N_18147);
or U20517 (N_20517,N_18942,N_19013);
nand U20518 (N_20518,N_18978,N_19516);
or U20519 (N_20519,N_18804,N_19790);
nor U20520 (N_20520,N_19778,N_18097);
or U20521 (N_20521,N_19851,N_18668);
or U20522 (N_20522,N_18025,N_18298);
xor U20523 (N_20523,N_19788,N_19900);
or U20524 (N_20524,N_19966,N_18987);
nor U20525 (N_20525,N_18648,N_19613);
or U20526 (N_20526,N_18816,N_19798);
nor U20527 (N_20527,N_18834,N_19509);
or U20528 (N_20528,N_18151,N_19074);
nor U20529 (N_20529,N_18972,N_19677);
nor U20530 (N_20530,N_18021,N_19372);
and U20531 (N_20531,N_18288,N_18089);
nand U20532 (N_20532,N_19106,N_19493);
xor U20533 (N_20533,N_18095,N_19424);
nand U20534 (N_20534,N_19739,N_19308);
xnor U20535 (N_20535,N_18060,N_18525);
nor U20536 (N_20536,N_18988,N_18472);
nand U20537 (N_20537,N_19810,N_18112);
xnor U20538 (N_20538,N_19501,N_18689);
nor U20539 (N_20539,N_19186,N_18459);
nor U20540 (N_20540,N_18725,N_19523);
nand U20541 (N_20541,N_19252,N_19586);
xnor U20542 (N_20542,N_19157,N_19781);
and U20543 (N_20543,N_18616,N_18159);
xnor U20544 (N_20544,N_18349,N_19477);
xor U20545 (N_20545,N_19750,N_18246);
or U20546 (N_20546,N_19686,N_18859);
xor U20547 (N_20547,N_19002,N_19890);
nor U20548 (N_20548,N_18211,N_18128);
nor U20549 (N_20549,N_18256,N_18010);
xnor U20550 (N_20550,N_18559,N_18701);
and U20551 (N_20551,N_18039,N_18153);
nor U20552 (N_20552,N_18928,N_19237);
or U20553 (N_20553,N_18231,N_18526);
and U20554 (N_20554,N_19590,N_18477);
or U20555 (N_20555,N_18415,N_18005);
xor U20556 (N_20556,N_19042,N_18410);
and U20557 (N_20557,N_18980,N_19528);
and U20558 (N_20558,N_18869,N_18922);
xnor U20559 (N_20559,N_19135,N_19491);
xnor U20560 (N_20560,N_19568,N_18125);
and U20561 (N_20561,N_18411,N_19538);
and U20562 (N_20562,N_19664,N_19722);
or U20563 (N_20563,N_19544,N_18345);
and U20564 (N_20564,N_19227,N_19012);
nand U20565 (N_20565,N_18164,N_19705);
or U20566 (N_20566,N_18619,N_18046);
nor U20567 (N_20567,N_18521,N_18693);
nor U20568 (N_20568,N_19620,N_19358);
or U20569 (N_20569,N_19995,N_19521);
nand U20570 (N_20570,N_18398,N_19242);
nor U20571 (N_20571,N_18801,N_18673);
nand U20572 (N_20572,N_18511,N_19195);
and U20573 (N_20573,N_19173,N_18533);
or U20574 (N_20574,N_18382,N_18332);
and U20575 (N_20575,N_18754,N_18412);
nor U20576 (N_20576,N_18134,N_19546);
nor U20577 (N_20577,N_19785,N_18618);
and U20578 (N_20578,N_18337,N_18883);
xnor U20579 (N_20579,N_19492,N_18092);
nor U20580 (N_20580,N_18796,N_19148);
nand U20581 (N_20581,N_18059,N_18570);
nor U20582 (N_20582,N_19865,N_19917);
and U20583 (N_20583,N_19410,N_18874);
or U20584 (N_20584,N_18534,N_19240);
and U20585 (N_20585,N_18609,N_19010);
or U20586 (N_20586,N_18012,N_18297);
nor U20587 (N_20587,N_18513,N_19742);
or U20588 (N_20588,N_18610,N_19747);
and U20589 (N_20589,N_18576,N_19175);
nand U20590 (N_20590,N_18204,N_19165);
nor U20591 (N_20591,N_19548,N_19614);
xnor U20592 (N_20592,N_19884,N_19682);
nor U20593 (N_20593,N_19120,N_19907);
and U20594 (N_20594,N_19784,N_19197);
nor U20595 (N_20595,N_18873,N_18814);
xor U20596 (N_20596,N_19746,N_18325);
nand U20597 (N_20597,N_18551,N_18179);
and U20598 (N_20598,N_18560,N_19961);
and U20599 (N_20599,N_19690,N_18656);
xnor U20600 (N_20600,N_18222,N_18923);
nor U20601 (N_20601,N_18028,N_19332);
xor U20602 (N_20602,N_19638,N_19824);
or U20603 (N_20603,N_18067,N_19771);
or U20604 (N_20604,N_18925,N_19639);
nand U20605 (N_20605,N_18333,N_19654);
or U20606 (N_20606,N_18898,N_18053);
nand U20607 (N_20607,N_18034,N_18765);
or U20608 (N_20608,N_18833,N_18263);
xnor U20609 (N_20609,N_18762,N_19324);
nor U20610 (N_20610,N_19858,N_19936);
and U20611 (N_20611,N_19901,N_19571);
or U20612 (N_20612,N_19437,N_19667);
and U20613 (N_20613,N_19591,N_19193);
and U20614 (N_20614,N_18432,N_18894);
or U20615 (N_20615,N_19022,N_18098);
or U20616 (N_20616,N_18516,N_18386);
nand U20617 (N_20617,N_18975,N_18514);
or U20618 (N_20618,N_18300,N_18940);
nor U20619 (N_20619,N_19818,N_19644);
or U20620 (N_20620,N_18738,N_19465);
and U20621 (N_20621,N_19592,N_19600);
xnor U20622 (N_20622,N_18939,N_18264);
nand U20623 (N_20623,N_19053,N_19016);
and U20624 (N_20624,N_19126,N_19347);
nand U20625 (N_20625,N_19604,N_18339);
nor U20626 (N_20626,N_19271,N_19508);
and U20627 (N_20627,N_19109,N_18225);
xnor U20628 (N_20628,N_19502,N_18492);
xnor U20629 (N_20629,N_18421,N_19947);
nor U20630 (N_20630,N_18519,N_18133);
nor U20631 (N_20631,N_18090,N_19102);
or U20632 (N_20632,N_18994,N_18910);
nor U20633 (N_20633,N_18201,N_18445);
and U20634 (N_20634,N_19622,N_19302);
and U20635 (N_20635,N_19679,N_19938);
or U20636 (N_20636,N_18383,N_18968);
and U20637 (N_20637,N_19668,N_19701);
nand U20638 (N_20638,N_19363,N_19814);
or U20639 (N_20639,N_19657,N_19314);
xnor U20640 (N_20640,N_19287,N_19594);
nor U20641 (N_20641,N_19054,N_19034);
nor U20642 (N_20642,N_18315,N_19096);
xor U20643 (N_20643,N_19478,N_18677);
xnor U20644 (N_20644,N_19891,N_18205);
nor U20645 (N_20645,N_19061,N_19077);
nand U20646 (N_20646,N_18048,N_19128);
xnor U20647 (N_20647,N_19239,N_18848);
xor U20648 (N_20648,N_19606,N_18476);
xor U20649 (N_20649,N_19009,N_18632);
nand U20650 (N_20650,N_18414,N_18694);
nor U20651 (N_20651,N_19244,N_19163);
xor U20652 (N_20652,N_19738,N_19408);
xnor U20653 (N_20653,N_19696,N_19524);
nor U20654 (N_20654,N_18926,N_19172);
or U20655 (N_20655,N_18846,N_18653);
or U20656 (N_20656,N_19943,N_19626);
xnor U20657 (N_20657,N_18790,N_18899);
nand U20658 (N_20658,N_18655,N_18334);
nor U20659 (N_20659,N_19717,N_19361);
and U20660 (N_20660,N_18646,N_18176);
nor U20661 (N_20661,N_18976,N_18003);
nor U20662 (N_20662,N_18121,N_19649);
nor U20663 (N_20663,N_19220,N_18203);
xor U20664 (N_20664,N_18882,N_18078);
nor U20665 (N_20665,N_19419,N_19303);
or U20666 (N_20666,N_19017,N_19304);
nand U20667 (N_20667,N_19728,N_19183);
xnor U20668 (N_20668,N_19373,N_18759);
or U20669 (N_20669,N_19323,N_19765);
or U20670 (N_20670,N_19984,N_18766);
and U20671 (N_20671,N_18296,N_18301);
xor U20672 (N_20672,N_19147,N_19734);
or U20673 (N_20673,N_19578,N_18285);
xor U20674 (N_20674,N_19038,N_19103);
and U20675 (N_20675,N_19014,N_19176);
nor U20676 (N_20676,N_19326,N_19566);
nor U20677 (N_20677,N_19401,N_19791);
nand U20678 (N_20678,N_18441,N_19344);
or U20679 (N_20679,N_18748,N_18567);
nand U20680 (N_20680,N_19150,N_19205);
or U20681 (N_20681,N_19517,N_18366);
or U20682 (N_20682,N_19957,N_19443);
nor U20683 (N_20683,N_19306,N_19226);
nor U20684 (N_20684,N_18474,N_19617);
xnor U20685 (N_20685,N_19284,N_18886);
nand U20686 (N_20686,N_19469,N_18636);
nor U20687 (N_20687,N_18553,N_18589);
or U20688 (N_20688,N_19933,N_19439);
or U20689 (N_20689,N_18379,N_19417);
nor U20690 (N_20690,N_18305,N_18854);
xor U20691 (N_20691,N_18276,N_18703);
xor U20692 (N_20692,N_19142,N_19080);
and U20693 (N_20693,N_18844,N_18654);
and U20694 (N_20694,N_18837,N_18258);
or U20695 (N_20695,N_19609,N_18328);
xnor U20696 (N_20696,N_19588,N_18965);
or U20697 (N_20697,N_19506,N_19167);
nand U20698 (N_20698,N_18447,N_18051);
and U20699 (N_20699,N_18771,N_19585);
and U20700 (N_20700,N_18818,N_18891);
or U20701 (N_20701,N_18635,N_19380);
nand U20702 (N_20702,N_19659,N_19486);
xnor U20703 (N_20703,N_19379,N_18876);
and U20704 (N_20704,N_18335,N_18247);
nor U20705 (N_20705,N_19309,N_18214);
and U20706 (N_20706,N_18352,N_19274);
and U20707 (N_20707,N_19371,N_18902);
or U20708 (N_20708,N_19745,N_19615);
xnor U20709 (N_20709,N_18750,N_18778);
xor U20710 (N_20710,N_18686,N_18434);
nand U20711 (N_20711,N_18642,N_18697);
nor U20712 (N_20712,N_19133,N_18568);
xnor U20713 (N_20713,N_18482,N_19476);
xnor U20714 (N_20714,N_19716,N_18884);
or U20715 (N_20715,N_18896,N_19794);
nor U20716 (N_20716,N_18681,N_18542);
or U20717 (N_20717,N_19838,N_19426);
xnor U20718 (N_20718,N_18013,N_19194);
xnor U20719 (N_20719,N_18354,N_18721);
or U20720 (N_20720,N_18064,N_18807);
nor U20721 (N_20721,N_18995,N_19155);
and U20722 (N_20722,N_19837,N_18548);
nand U20723 (N_20723,N_18274,N_19527);
nand U20724 (N_20724,N_19497,N_18072);
nand U20725 (N_20725,N_19669,N_19352);
xnor U20726 (N_20726,N_19065,N_18970);
and U20727 (N_20727,N_19375,N_18992);
and U20728 (N_20728,N_18789,N_19520);
nor U20729 (N_20729,N_18645,N_18887);
nand U20730 (N_20730,N_19164,N_18044);
nand U20731 (N_20731,N_19348,N_19422);
xnor U20732 (N_20732,N_19355,N_19732);
or U20733 (N_20733,N_19473,N_19028);
and U20734 (N_20734,N_18026,N_18006);
and U20735 (N_20735,N_19108,N_19729);
nand U20736 (N_20736,N_18116,N_18861);
nor U20737 (N_20737,N_18998,N_19134);
or U20738 (N_20738,N_18530,N_19209);
xor U20739 (N_20739,N_18509,N_18623);
xnor U20740 (N_20740,N_19534,N_18245);
or U20741 (N_20741,N_19313,N_19821);
and U20742 (N_20742,N_19339,N_19736);
xnor U20743 (N_20743,N_19255,N_18192);
nor U20744 (N_20744,N_18667,N_19441);
nand U20745 (N_20745,N_18253,N_19297);
and U20746 (N_20746,N_19608,N_18400);
or U20747 (N_20747,N_19202,N_18188);
and U20748 (N_20748,N_19029,N_18662);
xor U20749 (N_20749,N_18709,N_19731);
nor U20750 (N_20750,N_18377,N_19885);
or U20751 (N_20751,N_18307,N_19428);
xnor U20752 (N_20752,N_19813,N_19547);
nor U20753 (N_20753,N_19782,N_18240);
nor U20754 (N_20754,N_18229,N_19525);
nor U20755 (N_20755,N_19253,N_18690);
xor U20756 (N_20756,N_19979,N_19223);
nand U20757 (N_20757,N_19730,N_19572);
and U20758 (N_20758,N_19559,N_19871);
xnor U20759 (N_20759,N_19398,N_18275);
and U20760 (N_20760,N_19046,N_19899);
and U20761 (N_20761,N_19123,N_18165);
xnor U20762 (N_20762,N_18613,N_18075);
or U20763 (N_20763,N_19602,N_18284);
or U20764 (N_20764,N_18491,N_18757);
xnor U20765 (N_20765,N_18117,N_18755);
nand U20766 (N_20766,N_18963,N_18588);
nor U20767 (N_20767,N_18093,N_18504);
nor U20768 (N_20768,N_19384,N_18652);
nor U20769 (N_20769,N_19286,N_19565);
nand U20770 (N_20770,N_18938,N_19170);
xor U20771 (N_20771,N_18330,N_18691);
or U20772 (N_20772,N_19555,N_18518);
and U20773 (N_20773,N_19962,N_19438);
and U20774 (N_20774,N_19245,N_18826);
nand U20775 (N_20775,N_18365,N_18931);
xor U20776 (N_20776,N_18561,N_18723);
nand U20777 (N_20777,N_18715,N_18628);
xnor U20778 (N_20778,N_18956,N_19733);
or U20779 (N_20779,N_18830,N_19345);
nor U20780 (N_20780,N_18932,N_18219);
xnor U20781 (N_20781,N_18696,N_18543);
and U20782 (N_20782,N_19536,N_18842);
nand U20783 (N_20783,N_18598,N_19444);
or U20784 (N_20784,N_18200,N_18841);
and U20785 (N_20785,N_19121,N_19743);
or U20786 (N_20786,N_19605,N_19828);
nor U20787 (N_20787,N_19412,N_18353);
nor U20788 (N_20788,N_19704,N_19580);
xnor U20789 (N_20789,N_18426,N_18111);
nand U20790 (N_20790,N_19238,N_18496);
nor U20791 (N_20791,N_18867,N_19198);
nand U20792 (N_20792,N_18544,N_18903);
or U20793 (N_20793,N_18363,N_18065);
or U20794 (N_20794,N_19378,N_18373);
nor U20795 (N_20795,N_18698,N_19019);
or U20796 (N_20796,N_18000,N_18680);
and U20797 (N_20797,N_19522,N_19296);
xor U20798 (N_20798,N_19855,N_18843);
or U20799 (N_20799,N_18787,N_18760);
nand U20800 (N_20800,N_18674,N_18813);
or U20801 (N_20801,N_18443,N_19672);
and U20802 (N_20802,N_19413,N_19897);
or U20803 (N_20803,N_18954,N_18714);
or U20804 (N_20804,N_19460,N_19691);
and U20805 (N_20805,N_19495,N_19161);
nor U20806 (N_20806,N_18417,N_18549);
nor U20807 (N_20807,N_18350,N_19515);
xnor U20808 (N_20808,N_19503,N_19766);
and U20809 (N_20809,N_19827,N_18277);
nor U20810 (N_20810,N_18913,N_18152);
xor U20811 (N_20811,N_19368,N_19421);
nand U20812 (N_20812,N_18107,N_18073);
and U20813 (N_20813,N_19954,N_19633);
xor U20814 (N_20814,N_19504,N_19573);
xnor U20815 (N_20815,N_19267,N_19662);
nand U20816 (N_20816,N_19411,N_19112);
and U20817 (N_20817,N_18660,N_19132);
nor U20818 (N_20818,N_18779,N_18392);
xnor U20819 (N_20819,N_18487,N_18320);
or U20820 (N_20820,N_18870,N_18768);
nand U20821 (N_20821,N_18451,N_18295);
and U20822 (N_20822,N_19978,N_18150);
and U20823 (N_20823,N_19299,N_18215);
nand U20824 (N_20824,N_19479,N_19221);
or U20825 (N_20825,N_18800,N_18797);
nor U20826 (N_20826,N_19832,N_18657);
xnor U20827 (N_20827,N_19464,N_19052);
or U20828 (N_20828,N_19199,N_18659);
xor U20829 (N_20829,N_19806,N_18507);
nor U20830 (N_20830,N_18979,N_19629);
or U20831 (N_20831,N_18270,N_18370);
nand U20832 (N_20832,N_18031,N_19597);
nor U20833 (N_20833,N_19225,N_18593);
and U20834 (N_20834,N_19948,N_19697);
or U20835 (N_20835,N_18555,N_18384);
xor U20836 (N_20836,N_19647,N_18479);
or U20837 (N_20837,N_18166,N_19394);
or U20838 (N_20838,N_18945,N_18675);
or U20839 (N_20839,N_18401,N_18404);
nand U20840 (N_20840,N_19179,N_19952);
nor U20841 (N_20841,N_18455,N_18139);
nor U20842 (N_20842,N_19876,N_18438);
nand U20843 (N_20843,N_19541,N_18237);
nand U20844 (N_20844,N_18052,N_19812);
or U20845 (N_20845,N_18793,N_19982);
xnor U20846 (N_20846,N_18792,N_18265);
and U20847 (N_20847,N_18062,N_18733);
xnor U20848 (N_20848,N_19219,N_18456);
and U20849 (N_20849,N_18744,N_18483);
nand U20850 (N_20850,N_19842,N_19819);
nor U20851 (N_20851,N_19611,N_18390);
nor U20852 (N_20852,N_19761,N_19596);
and U20853 (N_20853,N_18068,N_19184);
xor U20854 (N_20854,N_18433,N_18374);
nand U20855 (N_20855,N_19462,N_18953);
nor U20856 (N_20856,N_19051,N_18772);
or U20857 (N_20857,N_19992,N_19909);
xor U20858 (N_20858,N_19636,N_19651);
nand U20859 (N_20859,N_18402,N_19570);
nor U20860 (N_20860,N_19918,N_19055);
xnor U20861 (N_20861,N_19233,N_19973);
or U20862 (N_20862,N_19285,N_18261);
and U20863 (N_20863,N_19321,N_19929);
nand U20864 (N_20864,N_19158,N_19007);
xnor U20865 (N_20865,N_18460,N_18341);
nor U20866 (N_20866,N_19450,N_18268);
xnor U20867 (N_20867,N_19846,N_18424);
xnor U20868 (N_20868,N_18235,N_18871);
xor U20869 (N_20869,N_18971,N_18238);
xor U20870 (N_20870,N_18966,N_18055);
or U20871 (N_20871,N_19919,N_18342);
or U20872 (N_20872,N_19434,N_19247);
xnor U20873 (N_20873,N_19612,N_19675);
or U20874 (N_20874,N_19466,N_18828);
or U20875 (N_20875,N_18101,N_19189);
nand U20876 (N_20876,N_19535,N_19015);
nor U20877 (N_20877,N_19735,N_18260);
nand U20878 (N_20878,N_18756,N_18361);
nand U20879 (N_20879,N_19764,N_19860);
and U20880 (N_20880,N_19985,N_18829);
nor U20881 (N_20881,N_19048,N_18202);
nand U20882 (N_20882,N_19511,N_19872);
or U20883 (N_20883,N_18357,N_18047);
or U20884 (N_20884,N_19156,N_18573);
or U20885 (N_20885,N_19101,N_19869);
xnor U20886 (N_20886,N_19505,N_18114);
nand U20887 (N_20887,N_18282,N_18094);
and U20888 (N_20888,N_19086,N_18803);
or U20889 (N_20889,N_18838,N_19893);
nor U20890 (N_20890,N_19783,N_19870);
xor U20891 (N_20891,N_19397,N_19031);
xor U20892 (N_20892,N_19174,N_18286);
or U20893 (N_20893,N_19406,N_18105);
xor U20894 (N_20894,N_18856,N_19852);
nor U20895 (N_20895,N_18437,N_19940);
nor U20896 (N_20896,N_18631,N_18280);
nand U20897 (N_20897,N_18562,N_19276);
nand U20898 (N_20898,N_18822,N_18481);
xor U20899 (N_20899,N_19089,N_19663);
nor U20900 (N_20900,N_18009,N_19433);
and U20901 (N_20901,N_18018,N_18123);
and U20902 (N_20902,N_18233,N_19429);
xnor U20903 (N_20903,N_19529,N_19004);
nor U20904 (N_20904,N_18629,N_18228);
nor U20905 (N_20905,N_19889,N_18387);
nand U20906 (N_20906,N_18272,N_19092);
xnor U20907 (N_20907,N_19811,N_18019);
nor U20908 (N_20908,N_19950,N_19563);
and U20909 (N_20909,N_18740,N_18096);
and U20910 (N_20910,N_18422,N_18620);
nand U20911 (N_20911,N_19442,N_19217);
and U20912 (N_20912,N_18566,N_18743);
xor U20913 (N_20913,N_18541,N_19331);
or U20914 (N_20914,N_18232,N_19350);
nand U20915 (N_20915,N_19115,N_18403);
nand U20916 (N_20916,N_18621,N_19593);
xor U20917 (N_20917,N_18607,N_19024);
or U20918 (N_20918,N_18781,N_18154);
and U20919 (N_20919,N_18614,N_19550);
or U20920 (N_20920,N_19387,N_18194);
nor U20921 (N_20921,N_18735,N_19923);
nor U20922 (N_20922,N_19630,N_19305);
or U20923 (N_20923,N_18684,N_18893);
or U20924 (N_20924,N_18371,N_19658);
nand U20925 (N_20925,N_18773,N_18199);
or U20926 (N_20926,N_18063,N_19191);
or U20927 (N_20927,N_19916,N_19800);
or U20928 (N_20928,N_18408,N_19354);
nand U20929 (N_20929,N_19777,N_18996);
nand U20930 (N_20930,N_19519,N_19830);
xnor U20931 (N_20931,N_19188,N_19404);
nor U20932 (N_20932,N_18015,N_18912);
and U20933 (N_20933,N_19713,N_18831);
xor U20934 (N_20934,N_18499,N_18266);
xor U20935 (N_20935,N_18173,N_18967);
and U20936 (N_20936,N_18254,N_18906);
or U20937 (N_20937,N_18030,N_19455);
or U20938 (N_20938,N_19262,N_18155);
and U20939 (N_20939,N_18466,N_18860);
nand U20940 (N_20940,N_19930,N_19977);
nand U20941 (N_20941,N_18488,N_19815);
nor U20942 (N_20942,N_19489,N_18769);
nand U20943 (N_20943,N_18043,N_18313);
and U20944 (N_20944,N_18515,N_18493);
xnor U20945 (N_20945,N_19059,N_18250);
nor U20946 (N_20946,N_18099,N_19796);
or U20947 (N_20947,N_18950,N_19700);
and U20948 (N_20948,N_18251,N_18351);
and U20949 (N_20949,N_18941,N_18444);
or U20950 (N_20950,N_19058,N_19625);
xnor U20951 (N_20951,N_19316,N_19708);
or U20952 (N_20952,N_18983,N_18419);
nand U20953 (N_20953,N_18717,N_18879);
nor U20954 (N_20954,N_18742,N_18278);
nand U20955 (N_20955,N_18788,N_19118);
xnor U20956 (N_20956,N_19656,N_18817);
or U20957 (N_20957,N_19925,N_18331);
xor U20958 (N_20958,N_19266,N_18024);
or U20959 (N_20959,N_18984,N_18550);
and U20960 (N_20960,N_18182,N_19138);
and U20961 (N_20961,N_18730,N_19786);
and U20962 (N_20962,N_19820,N_19564);
and U20963 (N_20963,N_19459,N_19457);
nor U20964 (N_20964,N_18777,N_19177);
or U20965 (N_20965,N_18136,N_18145);
xnor U20966 (N_20966,N_18216,N_19577);
and U20967 (N_20967,N_18875,N_18061);
or U20968 (N_20968,N_19892,N_19847);
nor U20969 (N_20969,N_18104,N_19635);
xor U20970 (N_20970,N_19562,N_18916);
nand U20971 (N_20971,N_19921,N_18008);
nand U20972 (N_20972,N_19362,N_18997);
and U20973 (N_20973,N_18895,N_19627);
nand U20974 (N_20974,N_19117,N_18091);
or U20975 (N_20975,N_18888,N_19472);
and U20976 (N_20976,N_19941,N_19282);
xor U20977 (N_20977,N_18638,N_18257);
xor U20978 (N_20978,N_19880,N_18578);
nand U20979 (N_20979,N_18369,N_19888);
xor U20980 (N_20980,N_18729,N_18029);
xor U20981 (N_20981,N_19280,N_19381);
nor U20982 (N_20982,N_18161,N_18022);
and U20983 (N_20983,N_19346,N_19587);
and U20984 (N_20984,N_19405,N_18045);
nor U20985 (N_20985,N_19325,N_18808);
nand U20986 (N_20986,N_19216,N_18617);
xnor U20987 (N_20987,N_19487,N_18439);
and U20988 (N_20988,N_18138,N_19797);
or U20989 (N_20989,N_18905,N_19213);
and U20990 (N_20990,N_18454,N_18552);
nand U20991 (N_20991,N_18935,N_19595);
xnor U20992 (N_20992,N_18665,N_19540);
and U20993 (N_20993,N_19965,N_18611);
or U20994 (N_20994,N_18079,N_18057);
nor U20995 (N_20995,N_19518,N_19330);
nand U20996 (N_20996,N_19357,N_19759);
xor U20997 (N_20997,N_19336,N_18273);
xnor U20998 (N_20998,N_18702,N_18819);
nor U20999 (N_20999,N_19415,N_19969);
xnor U21000 (N_21000,N_19705,N_19234);
nand U21001 (N_21001,N_18514,N_18447);
nor U21002 (N_21002,N_19882,N_18896);
xor U21003 (N_21003,N_18374,N_19471);
nand U21004 (N_21004,N_18278,N_19780);
nand U21005 (N_21005,N_18196,N_18833);
xnor U21006 (N_21006,N_18786,N_18764);
and U21007 (N_21007,N_18915,N_18975);
nand U21008 (N_21008,N_19128,N_18130);
nor U21009 (N_21009,N_19145,N_19938);
nor U21010 (N_21010,N_19649,N_19858);
nor U21011 (N_21011,N_18062,N_18510);
nand U21012 (N_21012,N_19492,N_18004);
xor U21013 (N_21013,N_19712,N_18862);
nand U21014 (N_21014,N_18913,N_18127);
nor U21015 (N_21015,N_18762,N_19264);
xnor U21016 (N_21016,N_19947,N_19341);
nand U21017 (N_21017,N_19142,N_18681);
xor U21018 (N_21018,N_19263,N_18935);
and U21019 (N_21019,N_18408,N_19072);
nand U21020 (N_21020,N_18507,N_18397);
or U21021 (N_21021,N_18883,N_19575);
and U21022 (N_21022,N_19420,N_19270);
or U21023 (N_21023,N_19585,N_18107);
or U21024 (N_21024,N_18185,N_18378);
nand U21025 (N_21025,N_18676,N_18040);
xor U21026 (N_21026,N_18873,N_19476);
nand U21027 (N_21027,N_18463,N_18534);
and U21028 (N_21028,N_18213,N_19162);
xor U21029 (N_21029,N_19644,N_18680);
nor U21030 (N_21030,N_19073,N_19679);
or U21031 (N_21031,N_18247,N_18415);
and U21032 (N_21032,N_18952,N_19805);
nor U21033 (N_21033,N_19050,N_19338);
and U21034 (N_21034,N_19640,N_19151);
xnor U21035 (N_21035,N_18093,N_19222);
xnor U21036 (N_21036,N_19743,N_19501);
and U21037 (N_21037,N_18935,N_19161);
xnor U21038 (N_21038,N_19130,N_19411);
and U21039 (N_21039,N_19832,N_18454);
xor U21040 (N_21040,N_19331,N_18839);
xor U21041 (N_21041,N_18011,N_18351);
xnor U21042 (N_21042,N_19959,N_19700);
and U21043 (N_21043,N_18233,N_19741);
nand U21044 (N_21044,N_19335,N_19324);
xor U21045 (N_21045,N_18770,N_19617);
nor U21046 (N_21046,N_18567,N_18899);
nor U21047 (N_21047,N_18753,N_18270);
and U21048 (N_21048,N_18340,N_19875);
nor U21049 (N_21049,N_19795,N_19844);
nor U21050 (N_21050,N_19479,N_18622);
nor U21051 (N_21051,N_18061,N_19398);
nand U21052 (N_21052,N_18127,N_19868);
or U21053 (N_21053,N_19798,N_19355);
nand U21054 (N_21054,N_19822,N_19163);
and U21055 (N_21055,N_19866,N_19094);
or U21056 (N_21056,N_18492,N_19472);
nand U21057 (N_21057,N_19336,N_19823);
nor U21058 (N_21058,N_18736,N_18240);
or U21059 (N_21059,N_19511,N_19634);
or U21060 (N_21060,N_19416,N_18327);
nor U21061 (N_21061,N_19164,N_18511);
nor U21062 (N_21062,N_19235,N_18300);
nor U21063 (N_21063,N_19529,N_18501);
and U21064 (N_21064,N_19581,N_19781);
nor U21065 (N_21065,N_19629,N_18595);
nor U21066 (N_21066,N_19041,N_19464);
or U21067 (N_21067,N_18230,N_19487);
and U21068 (N_21068,N_18395,N_18010);
and U21069 (N_21069,N_19546,N_18734);
nand U21070 (N_21070,N_18767,N_19292);
nand U21071 (N_21071,N_18097,N_19821);
and U21072 (N_21072,N_18009,N_18809);
nand U21073 (N_21073,N_19320,N_19726);
and U21074 (N_21074,N_18057,N_18017);
nor U21075 (N_21075,N_19224,N_19838);
xnor U21076 (N_21076,N_18952,N_19628);
or U21077 (N_21077,N_19143,N_19523);
or U21078 (N_21078,N_19652,N_18723);
nand U21079 (N_21079,N_18949,N_19180);
or U21080 (N_21080,N_18237,N_18022);
or U21081 (N_21081,N_19411,N_18885);
and U21082 (N_21082,N_19240,N_19378);
nand U21083 (N_21083,N_19478,N_19212);
or U21084 (N_21084,N_18646,N_19410);
xor U21085 (N_21085,N_18579,N_18275);
nand U21086 (N_21086,N_18615,N_19771);
xnor U21087 (N_21087,N_18834,N_19117);
nand U21088 (N_21088,N_19440,N_18912);
and U21089 (N_21089,N_19386,N_18426);
nor U21090 (N_21090,N_18080,N_18663);
and U21091 (N_21091,N_19717,N_18756);
or U21092 (N_21092,N_18729,N_18534);
xor U21093 (N_21093,N_19090,N_19789);
and U21094 (N_21094,N_19257,N_18368);
xnor U21095 (N_21095,N_19756,N_18562);
nor U21096 (N_21096,N_18281,N_19680);
nor U21097 (N_21097,N_18555,N_19235);
and U21098 (N_21098,N_19232,N_18599);
nand U21099 (N_21099,N_19881,N_19149);
or U21100 (N_21100,N_19718,N_18876);
or U21101 (N_21101,N_19056,N_18116);
or U21102 (N_21102,N_18549,N_19717);
and U21103 (N_21103,N_19584,N_19810);
nand U21104 (N_21104,N_18231,N_18303);
or U21105 (N_21105,N_19982,N_19623);
nor U21106 (N_21106,N_19895,N_19299);
nand U21107 (N_21107,N_18692,N_19343);
nand U21108 (N_21108,N_18109,N_19505);
or U21109 (N_21109,N_18461,N_18879);
and U21110 (N_21110,N_18798,N_19321);
nor U21111 (N_21111,N_19487,N_18093);
or U21112 (N_21112,N_18140,N_18854);
or U21113 (N_21113,N_19786,N_18441);
xor U21114 (N_21114,N_19320,N_19785);
xnor U21115 (N_21115,N_18733,N_18875);
and U21116 (N_21116,N_19867,N_19037);
nor U21117 (N_21117,N_18737,N_19004);
and U21118 (N_21118,N_19572,N_18915);
xnor U21119 (N_21119,N_19833,N_18006);
xnor U21120 (N_21120,N_18367,N_19619);
nor U21121 (N_21121,N_18668,N_18650);
xor U21122 (N_21122,N_18320,N_19624);
nand U21123 (N_21123,N_19871,N_19312);
xnor U21124 (N_21124,N_19258,N_19744);
nand U21125 (N_21125,N_19780,N_19226);
nor U21126 (N_21126,N_18953,N_19185);
nand U21127 (N_21127,N_19408,N_19178);
and U21128 (N_21128,N_19474,N_18307);
and U21129 (N_21129,N_18386,N_18204);
nand U21130 (N_21130,N_19282,N_19951);
nand U21131 (N_21131,N_18274,N_19526);
nor U21132 (N_21132,N_18491,N_18060);
and U21133 (N_21133,N_19224,N_19969);
nand U21134 (N_21134,N_19513,N_18897);
or U21135 (N_21135,N_19960,N_19010);
nor U21136 (N_21136,N_18602,N_19697);
or U21137 (N_21137,N_19726,N_19851);
or U21138 (N_21138,N_18636,N_18275);
nand U21139 (N_21139,N_18934,N_18591);
xnor U21140 (N_21140,N_19858,N_19747);
and U21141 (N_21141,N_19898,N_18113);
nor U21142 (N_21142,N_19111,N_19795);
nand U21143 (N_21143,N_18565,N_18979);
nand U21144 (N_21144,N_19834,N_19100);
nor U21145 (N_21145,N_19602,N_19238);
nor U21146 (N_21146,N_18752,N_18520);
and U21147 (N_21147,N_18038,N_19244);
or U21148 (N_21148,N_18898,N_18567);
nor U21149 (N_21149,N_18747,N_18540);
xor U21150 (N_21150,N_19184,N_19003);
xor U21151 (N_21151,N_18446,N_19438);
nand U21152 (N_21152,N_19098,N_19391);
nand U21153 (N_21153,N_18186,N_18590);
xor U21154 (N_21154,N_19048,N_18170);
xor U21155 (N_21155,N_18993,N_18923);
xor U21156 (N_21156,N_18855,N_18361);
and U21157 (N_21157,N_18635,N_18574);
xnor U21158 (N_21158,N_18654,N_19410);
and U21159 (N_21159,N_18671,N_18730);
nand U21160 (N_21160,N_19853,N_19499);
or U21161 (N_21161,N_18343,N_18464);
and U21162 (N_21162,N_19187,N_19018);
and U21163 (N_21163,N_19334,N_18822);
nand U21164 (N_21164,N_19313,N_18745);
or U21165 (N_21165,N_19387,N_19189);
xnor U21166 (N_21166,N_18440,N_18893);
nand U21167 (N_21167,N_18034,N_19434);
or U21168 (N_21168,N_18042,N_18949);
nor U21169 (N_21169,N_18151,N_18362);
nand U21170 (N_21170,N_19686,N_19159);
nand U21171 (N_21171,N_18109,N_19456);
nand U21172 (N_21172,N_19887,N_19127);
and U21173 (N_21173,N_18587,N_18016);
nor U21174 (N_21174,N_18478,N_18702);
nand U21175 (N_21175,N_18977,N_18663);
xor U21176 (N_21176,N_18604,N_18037);
nor U21177 (N_21177,N_18468,N_18496);
or U21178 (N_21178,N_18336,N_18068);
nor U21179 (N_21179,N_18814,N_19416);
nor U21180 (N_21180,N_19537,N_18795);
nand U21181 (N_21181,N_19261,N_18971);
nor U21182 (N_21182,N_18674,N_18138);
xnor U21183 (N_21183,N_18082,N_19242);
or U21184 (N_21184,N_18688,N_18008);
or U21185 (N_21185,N_19868,N_18520);
or U21186 (N_21186,N_19178,N_18746);
nor U21187 (N_21187,N_19666,N_19669);
nor U21188 (N_21188,N_18701,N_18232);
or U21189 (N_21189,N_19424,N_19022);
nand U21190 (N_21190,N_19390,N_18199);
and U21191 (N_21191,N_19132,N_18716);
nand U21192 (N_21192,N_18058,N_19227);
or U21193 (N_21193,N_19645,N_18125);
and U21194 (N_21194,N_19522,N_19690);
nor U21195 (N_21195,N_18591,N_18869);
or U21196 (N_21196,N_19126,N_19747);
nand U21197 (N_21197,N_19409,N_19765);
nand U21198 (N_21198,N_18067,N_19652);
and U21199 (N_21199,N_19118,N_18298);
and U21200 (N_21200,N_18894,N_18723);
xnor U21201 (N_21201,N_19914,N_18748);
nand U21202 (N_21202,N_18592,N_19381);
or U21203 (N_21203,N_18736,N_18020);
nor U21204 (N_21204,N_18060,N_19794);
xor U21205 (N_21205,N_19346,N_19463);
nor U21206 (N_21206,N_19778,N_19254);
or U21207 (N_21207,N_19599,N_18183);
or U21208 (N_21208,N_18102,N_18089);
xor U21209 (N_21209,N_19961,N_19628);
xnor U21210 (N_21210,N_19185,N_18652);
xnor U21211 (N_21211,N_18073,N_19414);
nand U21212 (N_21212,N_18307,N_18737);
and U21213 (N_21213,N_19868,N_18374);
or U21214 (N_21214,N_18694,N_18472);
xnor U21215 (N_21215,N_19686,N_19299);
xnor U21216 (N_21216,N_19943,N_18976);
xnor U21217 (N_21217,N_19038,N_19759);
nand U21218 (N_21218,N_18125,N_18820);
nand U21219 (N_21219,N_19430,N_19298);
nor U21220 (N_21220,N_18415,N_18131);
nor U21221 (N_21221,N_18164,N_18674);
nor U21222 (N_21222,N_18532,N_19272);
nor U21223 (N_21223,N_18602,N_18740);
or U21224 (N_21224,N_19192,N_19475);
nand U21225 (N_21225,N_18101,N_18701);
xor U21226 (N_21226,N_18041,N_19630);
xnor U21227 (N_21227,N_18641,N_19111);
xnor U21228 (N_21228,N_19336,N_18367);
nand U21229 (N_21229,N_19356,N_19720);
or U21230 (N_21230,N_18312,N_18616);
and U21231 (N_21231,N_19631,N_18975);
nand U21232 (N_21232,N_19008,N_19131);
xnor U21233 (N_21233,N_19252,N_18388);
xor U21234 (N_21234,N_18349,N_18619);
nand U21235 (N_21235,N_18823,N_19794);
nor U21236 (N_21236,N_18995,N_18530);
nand U21237 (N_21237,N_19526,N_19428);
xnor U21238 (N_21238,N_18812,N_18408);
nand U21239 (N_21239,N_19693,N_19333);
nand U21240 (N_21240,N_19704,N_18921);
nand U21241 (N_21241,N_19061,N_19188);
xnor U21242 (N_21242,N_18605,N_18862);
xor U21243 (N_21243,N_19194,N_19580);
nor U21244 (N_21244,N_19183,N_19020);
or U21245 (N_21245,N_18098,N_19392);
and U21246 (N_21246,N_18843,N_18554);
nor U21247 (N_21247,N_18547,N_19572);
nor U21248 (N_21248,N_19613,N_19923);
and U21249 (N_21249,N_19773,N_19802);
and U21250 (N_21250,N_19533,N_19555);
and U21251 (N_21251,N_19946,N_18704);
and U21252 (N_21252,N_18861,N_19626);
and U21253 (N_21253,N_18140,N_18402);
xnor U21254 (N_21254,N_18051,N_18060);
nand U21255 (N_21255,N_19705,N_19573);
xor U21256 (N_21256,N_19628,N_18763);
and U21257 (N_21257,N_19146,N_19439);
nor U21258 (N_21258,N_19232,N_18019);
xnor U21259 (N_21259,N_19744,N_18796);
xnor U21260 (N_21260,N_19959,N_18914);
and U21261 (N_21261,N_19286,N_18222);
nand U21262 (N_21262,N_19640,N_19446);
nand U21263 (N_21263,N_19826,N_18618);
nor U21264 (N_21264,N_19565,N_19757);
nor U21265 (N_21265,N_19079,N_19307);
xnor U21266 (N_21266,N_18576,N_19264);
nand U21267 (N_21267,N_18188,N_19300);
or U21268 (N_21268,N_19223,N_19750);
xor U21269 (N_21269,N_18826,N_19906);
or U21270 (N_21270,N_18203,N_18542);
or U21271 (N_21271,N_18840,N_19009);
xnor U21272 (N_21272,N_19754,N_19912);
nor U21273 (N_21273,N_19113,N_19120);
or U21274 (N_21274,N_19083,N_18802);
and U21275 (N_21275,N_19927,N_19196);
or U21276 (N_21276,N_18695,N_18622);
xor U21277 (N_21277,N_18291,N_18703);
xor U21278 (N_21278,N_18890,N_18364);
and U21279 (N_21279,N_18229,N_18240);
or U21280 (N_21280,N_19381,N_19188);
nor U21281 (N_21281,N_19637,N_19697);
nand U21282 (N_21282,N_18723,N_19046);
or U21283 (N_21283,N_19536,N_18734);
xnor U21284 (N_21284,N_18626,N_19125);
nand U21285 (N_21285,N_19830,N_19441);
or U21286 (N_21286,N_18323,N_19994);
xnor U21287 (N_21287,N_19171,N_18356);
or U21288 (N_21288,N_19577,N_19465);
xor U21289 (N_21289,N_18093,N_18850);
nand U21290 (N_21290,N_18774,N_19768);
nor U21291 (N_21291,N_19766,N_19121);
nand U21292 (N_21292,N_19635,N_18849);
nor U21293 (N_21293,N_19141,N_19624);
xor U21294 (N_21294,N_19013,N_18242);
nand U21295 (N_21295,N_18902,N_19268);
nor U21296 (N_21296,N_18301,N_18516);
and U21297 (N_21297,N_18690,N_19218);
nand U21298 (N_21298,N_18496,N_18401);
or U21299 (N_21299,N_19269,N_19141);
nor U21300 (N_21300,N_18410,N_18452);
or U21301 (N_21301,N_18600,N_18371);
or U21302 (N_21302,N_18122,N_19089);
and U21303 (N_21303,N_18405,N_18452);
or U21304 (N_21304,N_18361,N_18992);
or U21305 (N_21305,N_19228,N_19490);
nor U21306 (N_21306,N_19262,N_18784);
and U21307 (N_21307,N_19726,N_19799);
or U21308 (N_21308,N_18049,N_18853);
nor U21309 (N_21309,N_19042,N_19471);
and U21310 (N_21310,N_19252,N_18517);
xnor U21311 (N_21311,N_18388,N_19101);
or U21312 (N_21312,N_18636,N_19083);
nor U21313 (N_21313,N_18804,N_18947);
xor U21314 (N_21314,N_18602,N_19053);
and U21315 (N_21315,N_19551,N_19854);
nor U21316 (N_21316,N_18504,N_18770);
xnor U21317 (N_21317,N_19142,N_19622);
or U21318 (N_21318,N_18699,N_18528);
nand U21319 (N_21319,N_19158,N_18032);
nand U21320 (N_21320,N_18079,N_19280);
xor U21321 (N_21321,N_19808,N_18860);
nand U21322 (N_21322,N_19468,N_19978);
nand U21323 (N_21323,N_18118,N_19174);
xnor U21324 (N_21324,N_18137,N_19177);
nand U21325 (N_21325,N_18527,N_19491);
xor U21326 (N_21326,N_18116,N_19410);
nor U21327 (N_21327,N_18534,N_18787);
xnor U21328 (N_21328,N_19153,N_18524);
xor U21329 (N_21329,N_19312,N_18871);
nor U21330 (N_21330,N_18847,N_18249);
and U21331 (N_21331,N_19931,N_18068);
xor U21332 (N_21332,N_18994,N_19560);
and U21333 (N_21333,N_18199,N_18072);
nor U21334 (N_21334,N_19555,N_18913);
nand U21335 (N_21335,N_19620,N_19294);
nor U21336 (N_21336,N_18201,N_18845);
nand U21337 (N_21337,N_18460,N_19196);
nand U21338 (N_21338,N_18923,N_18381);
xnor U21339 (N_21339,N_19130,N_18911);
or U21340 (N_21340,N_19383,N_19999);
xnor U21341 (N_21341,N_19861,N_19169);
nor U21342 (N_21342,N_19926,N_19079);
nand U21343 (N_21343,N_19292,N_18620);
nor U21344 (N_21344,N_19667,N_19675);
nand U21345 (N_21345,N_19666,N_18079);
and U21346 (N_21346,N_19892,N_18621);
nand U21347 (N_21347,N_18002,N_18543);
nor U21348 (N_21348,N_19346,N_18200);
nor U21349 (N_21349,N_18953,N_18295);
nand U21350 (N_21350,N_18271,N_18686);
nor U21351 (N_21351,N_19042,N_18669);
nor U21352 (N_21352,N_19880,N_19477);
xnor U21353 (N_21353,N_19329,N_18719);
nor U21354 (N_21354,N_18343,N_19091);
nand U21355 (N_21355,N_18625,N_19577);
and U21356 (N_21356,N_18228,N_19548);
nor U21357 (N_21357,N_18970,N_19161);
xnor U21358 (N_21358,N_18801,N_18489);
or U21359 (N_21359,N_19163,N_18353);
xnor U21360 (N_21360,N_18751,N_18625);
xor U21361 (N_21361,N_18251,N_18533);
xor U21362 (N_21362,N_18508,N_18019);
nor U21363 (N_21363,N_18152,N_19055);
nand U21364 (N_21364,N_18514,N_18661);
and U21365 (N_21365,N_18002,N_18256);
nor U21366 (N_21366,N_18252,N_19562);
nand U21367 (N_21367,N_18369,N_18278);
or U21368 (N_21368,N_19276,N_19671);
nor U21369 (N_21369,N_18317,N_19955);
xor U21370 (N_21370,N_18270,N_19131);
and U21371 (N_21371,N_18491,N_18298);
nand U21372 (N_21372,N_19445,N_19254);
xor U21373 (N_21373,N_19174,N_19588);
and U21374 (N_21374,N_18285,N_18111);
nor U21375 (N_21375,N_18169,N_19373);
and U21376 (N_21376,N_19005,N_19890);
and U21377 (N_21377,N_18377,N_18886);
nand U21378 (N_21378,N_18163,N_19683);
nand U21379 (N_21379,N_18669,N_19916);
nand U21380 (N_21380,N_19864,N_19124);
nor U21381 (N_21381,N_19042,N_18808);
and U21382 (N_21382,N_19007,N_18235);
nand U21383 (N_21383,N_19691,N_18324);
nand U21384 (N_21384,N_18776,N_18707);
or U21385 (N_21385,N_18510,N_19575);
and U21386 (N_21386,N_19772,N_19602);
and U21387 (N_21387,N_19655,N_18866);
xor U21388 (N_21388,N_18458,N_19884);
or U21389 (N_21389,N_18551,N_19918);
nand U21390 (N_21390,N_18935,N_18035);
nand U21391 (N_21391,N_19420,N_19496);
nor U21392 (N_21392,N_19795,N_19381);
nor U21393 (N_21393,N_18256,N_19881);
xnor U21394 (N_21394,N_19411,N_18637);
nand U21395 (N_21395,N_18493,N_18340);
and U21396 (N_21396,N_19502,N_18571);
nor U21397 (N_21397,N_19288,N_18215);
nand U21398 (N_21398,N_19696,N_18522);
nand U21399 (N_21399,N_18867,N_18534);
or U21400 (N_21400,N_19532,N_18589);
and U21401 (N_21401,N_18215,N_19717);
and U21402 (N_21402,N_19838,N_18850);
nand U21403 (N_21403,N_19219,N_19856);
or U21404 (N_21404,N_18755,N_19457);
nand U21405 (N_21405,N_19705,N_19620);
nor U21406 (N_21406,N_19357,N_18467);
nand U21407 (N_21407,N_18397,N_18503);
or U21408 (N_21408,N_19623,N_18125);
xor U21409 (N_21409,N_18307,N_18842);
nand U21410 (N_21410,N_19312,N_18939);
or U21411 (N_21411,N_19861,N_18319);
and U21412 (N_21412,N_19995,N_18615);
and U21413 (N_21413,N_18312,N_18339);
and U21414 (N_21414,N_19584,N_18595);
or U21415 (N_21415,N_19994,N_19539);
or U21416 (N_21416,N_19563,N_19821);
and U21417 (N_21417,N_18878,N_19294);
nor U21418 (N_21418,N_19910,N_18127);
and U21419 (N_21419,N_19333,N_19689);
nand U21420 (N_21420,N_18328,N_19433);
nor U21421 (N_21421,N_19415,N_19978);
and U21422 (N_21422,N_18023,N_19115);
or U21423 (N_21423,N_18867,N_19070);
nand U21424 (N_21424,N_19668,N_18001);
xnor U21425 (N_21425,N_19324,N_18285);
or U21426 (N_21426,N_18483,N_18794);
and U21427 (N_21427,N_18113,N_19083);
or U21428 (N_21428,N_18774,N_18533);
and U21429 (N_21429,N_18360,N_19497);
nor U21430 (N_21430,N_18940,N_18470);
xnor U21431 (N_21431,N_19566,N_19951);
or U21432 (N_21432,N_19525,N_18060);
and U21433 (N_21433,N_19734,N_19421);
nand U21434 (N_21434,N_19272,N_19714);
and U21435 (N_21435,N_18794,N_18247);
xnor U21436 (N_21436,N_18141,N_18810);
and U21437 (N_21437,N_18558,N_19810);
nor U21438 (N_21438,N_19771,N_18062);
nand U21439 (N_21439,N_19412,N_18427);
nand U21440 (N_21440,N_19492,N_18291);
and U21441 (N_21441,N_18860,N_19290);
xor U21442 (N_21442,N_19480,N_19264);
or U21443 (N_21443,N_19081,N_18739);
xor U21444 (N_21444,N_19237,N_19160);
and U21445 (N_21445,N_18328,N_18863);
nor U21446 (N_21446,N_18209,N_19510);
nand U21447 (N_21447,N_18850,N_18514);
or U21448 (N_21448,N_18739,N_18220);
nor U21449 (N_21449,N_18413,N_19361);
nand U21450 (N_21450,N_18100,N_18817);
or U21451 (N_21451,N_19012,N_19649);
nor U21452 (N_21452,N_19857,N_19176);
nand U21453 (N_21453,N_18169,N_19126);
nand U21454 (N_21454,N_18722,N_18346);
or U21455 (N_21455,N_19720,N_19976);
nand U21456 (N_21456,N_19179,N_19182);
nand U21457 (N_21457,N_19528,N_19082);
nor U21458 (N_21458,N_19441,N_18946);
or U21459 (N_21459,N_19525,N_18848);
or U21460 (N_21460,N_19589,N_18045);
and U21461 (N_21461,N_18486,N_19346);
xnor U21462 (N_21462,N_18468,N_19528);
and U21463 (N_21463,N_18928,N_19396);
and U21464 (N_21464,N_19250,N_19781);
nand U21465 (N_21465,N_19639,N_18359);
xor U21466 (N_21466,N_18999,N_19112);
xor U21467 (N_21467,N_18018,N_19373);
xor U21468 (N_21468,N_18667,N_18165);
xnor U21469 (N_21469,N_19270,N_19319);
xnor U21470 (N_21470,N_18078,N_19887);
or U21471 (N_21471,N_18086,N_18535);
and U21472 (N_21472,N_19226,N_18976);
and U21473 (N_21473,N_18420,N_18879);
nor U21474 (N_21474,N_18863,N_19253);
nand U21475 (N_21475,N_19431,N_19271);
nor U21476 (N_21476,N_19214,N_19796);
and U21477 (N_21477,N_18926,N_19471);
and U21478 (N_21478,N_19249,N_19984);
or U21479 (N_21479,N_18125,N_18976);
nor U21480 (N_21480,N_18988,N_18462);
nor U21481 (N_21481,N_19989,N_18398);
or U21482 (N_21482,N_19386,N_19747);
or U21483 (N_21483,N_19280,N_18587);
nand U21484 (N_21484,N_19409,N_19256);
and U21485 (N_21485,N_19036,N_18660);
nand U21486 (N_21486,N_18631,N_19679);
xnor U21487 (N_21487,N_19236,N_19257);
and U21488 (N_21488,N_19990,N_18325);
and U21489 (N_21489,N_18521,N_18216);
and U21490 (N_21490,N_18398,N_19403);
nor U21491 (N_21491,N_19822,N_19678);
or U21492 (N_21492,N_18712,N_19895);
nor U21493 (N_21493,N_19180,N_18647);
xnor U21494 (N_21494,N_19054,N_19720);
nor U21495 (N_21495,N_18908,N_19062);
and U21496 (N_21496,N_19877,N_19248);
and U21497 (N_21497,N_18719,N_18744);
xor U21498 (N_21498,N_19584,N_18137);
or U21499 (N_21499,N_19686,N_19688);
nand U21500 (N_21500,N_19391,N_18861);
or U21501 (N_21501,N_18800,N_18902);
or U21502 (N_21502,N_18073,N_18019);
and U21503 (N_21503,N_19715,N_19348);
nand U21504 (N_21504,N_19802,N_19430);
and U21505 (N_21505,N_19502,N_19932);
and U21506 (N_21506,N_18874,N_18868);
nor U21507 (N_21507,N_18065,N_19149);
and U21508 (N_21508,N_19968,N_18241);
and U21509 (N_21509,N_19803,N_19974);
xor U21510 (N_21510,N_19255,N_19454);
xor U21511 (N_21511,N_19147,N_18196);
nand U21512 (N_21512,N_19664,N_19226);
nand U21513 (N_21513,N_18533,N_19341);
and U21514 (N_21514,N_18322,N_19596);
xor U21515 (N_21515,N_18973,N_18536);
nand U21516 (N_21516,N_19519,N_19191);
xnor U21517 (N_21517,N_18091,N_18285);
or U21518 (N_21518,N_19207,N_19888);
or U21519 (N_21519,N_18057,N_19242);
xnor U21520 (N_21520,N_19921,N_19542);
or U21521 (N_21521,N_19004,N_19864);
nor U21522 (N_21522,N_18196,N_18975);
xor U21523 (N_21523,N_19155,N_19310);
and U21524 (N_21524,N_18957,N_19556);
nor U21525 (N_21525,N_19623,N_18019);
or U21526 (N_21526,N_18080,N_19553);
xnor U21527 (N_21527,N_18084,N_18163);
and U21528 (N_21528,N_19544,N_18167);
xnor U21529 (N_21529,N_19468,N_18102);
nand U21530 (N_21530,N_18378,N_19416);
nor U21531 (N_21531,N_18071,N_18284);
or U21532 (N_21532,N_19863,N_19133);
nor U21533 (N_21533,N_18353,N_19313);
and U21534 (N_21534,N_19042,N_18468);
nor U21535 (N_21535,N_18589,N_18874);
or U21536 (N_21536,N_19172,N_18024);
xor U21537 (N_21537,N_18034,N_19806);
nor U21538 (N_21538,N_19906,N_19347);
nand U21539 (N_21539,N_18752,N_19422);
and U21540 (N_21540,N_18606,N_18800);
nand U21541 (N_21541,N_18535,N_18574);
and U21542 (N_21542,N_19427,N_19470);
nand U21543 (N_21543,N_18972,N_19440);
and U21544 (N_21544,N_18957,N_19922);
nand U21545 (N_21545,N_19342,N_18674);
nand U21546 (N_21546,N_18509,N_18222);
or U21547 (N_21547,N_19772,N_19578);
nand U21548 (N_21548,N_19967,N_19021);
and U21549 (N_21549,N_19234,N_18291);
nand U21550 (N_21550,N_19501,N_18708);
xor U21551 (N_21551,N_19209,N_19191);
and U21552 (N_21552,N_18177,N_19779);
nor U21553 (N_21553,N_18682,N_19916);
nand U21554 (N_21554,N_18253,N_19579);
xor U21555 (N_21555,N_19969,N_19328);
nor U21556 (N_21556,N_18988,N_18297);
nand U21557 (N_21557,N_19165,N_19603);
or U21558 (N_21558,N_19374,N_18647);
nand U21559 (N_21559,N_19681,N_19716);
or U21560 (N_21560,N_19276,N_18574);
xnor U21561 (N_21561,N_18891,N_19244);
and U21562 (N_21562,N_19465,N_19914);
and U21563 (N_21563,N_19837,N_18630);
or U21564 (N_21564,N_19533,N_19460);
nor U21565 (N_21565,N_19446,N_19531);
xor U21566 (N_21566,N_19240,N_18876);
and U21567 (N_21567,N_18933,N_19341);
and U21568 (N_21568,N_19248,N_18531);
xnor U21569 (N_21569,N_19166,N_19034);
nor U21570 (N_21570,N_18435,N_18348);
and U21571 (N_21571,N_19398,N_18749);
nand U21572 (N_21572,N_19567,N_18459);
nand U21573 (N_21573,N_18556,N_19700);
and U21574 (N_21574,N_19371,N_19464);
xnor U21575 (N_21575,N_18907,N_18709);
or U21576 (N_21576,N_19847,N_18432);
and U21577 (N_21577,N_18015,N_18274);
nor U21578 (N_21578,N_19779,N_18984);
and U21579 (N_21579,N_18557,N_18780);
nand U21580 (N_21580,N_19433,N_19256);
nand U21581 (N_21581,N_19558,N_18141);
nor U21582 (N_21582,N_19218,N_19481);
and U21583 (N_21583,N_18317,N_18422);
nor U21584 (N_21584,N_18025,N_18468);
nand U21585 (N_21585,N_19516,N_18225);
or U21586 (N_21586,N_19062,N_18451);
nand U21587 (N_21587,N_18123,N_18290);
xnor U21588 (N_21588,N_18076,N_18246);
or U21589 (N_21589,N_19814,N_18032);
nand U21590 (N_21590,N_19956,N_19804);
and U21591 (N_21591,N_19570,N_19748);
xor U21592 (N_21592,N_18615,N_19202);
or U21593 (N_21593,N_19972,N_18438);
and U21594 (N_21594,N_18440,N_19990);
nand U21595 (N_21595,N_18305,N_18734);
nand U21596 (N_21596,N_19527,N_19491);
or U21597 (N_21597,N_18417,N_19707);
nand U21598 (N_21598,N_18026,N_18942);
nor U21599 (N_21599,N_18167,N_18348);
or U21600 (N_21600,N_18810,N_18535);
nor U21601 (N_21601,N_18171,N_19612);
xnor U21602 (N_21602,N_19386,N_18863);
nand U21603 (N_21603,N_19962,N_19911);
nand U21604 (N_21604,N_19477,N_18041);
nand U21605 (N_21605,N_19094,N_19367);
and U21606 (N_21606,N_18291,N_19348);
or U21607 (N_21607,N_19497,N_18273);
or U21608 (N_21608,N_18628,N_19092);
nand U21609 (N_21609,N_19887,N_19334);
nor U21610 (N_21610,N_19311,N_19274);
and U21611 (N_21611,N_19344,N_19732);
or U21612 (N_21612,N_19338,N_19738);
nor U21613 (N_21613,N_18848,N_19533);
and U21614 (N_21614,N_18619,N_18726);
nor U21615 (N_21615,N_18092,N_18579);
and U21616 (N_21616,N_19897,N_19524);
nand U21617 (N_21617,N_18303,N_18623);
nand U21618 (N_21618,N_18775,N_19619);
nand U21619 (N_21619,N_18557,N_19146);
and U21620 (N_21620,N_18492,N_18923);
or U21621 (N_21621,N_19749,N_19157);
and U21622 (N_21622,N_18374,N_18577);
and U21623 (N_21623,N_18031,N_19582);
xor U21624 (N_21624,N_19223,N_18614);
nand U21625 (N_21625,N_19726,N_18799);
and U21626 (N_21626,N_19157,N_18053);
xor U21627 (N_21627,N_18670,N_19240);
and U21628 (N_21628,N_18018,N_19908);
or U21629 (N_21629,N_18406,N_19022);
nor U21630 (N_21630,N_19365,N_19819);
or U21631 (N_21631,N_18701,N_19240);
or U21632 (N_21632,N_18985,N_18441);
or U21633 (N_21633,N_18805,N_18692);
xor U21634 (N_21634,N_19528,N_19742);
and U21635 (N_21635,N_19253,N_18014);
nand U21636 (N_21636,N_18101,N_18999);
nand U21637 (N_21637,N_18693,N_18244);
nand U21638 (N_21638,N_19571,N_19658);
nor U21639 (N_21639,N_18189,N_19989);
nand U21640 (N_21640,N_19049,N_19460);
nand U21641 (N_21641,N_18443,N_18706);
nor U21642 (N_21642,N_19493,N_19074);
nor U21643 (N_21643,N_18872,N_19310);
nand U21644 (N_21644,N_18914,N_18864);
and U21645 (N_21645,N_19856,N_18456);
xor U21646 (N_21646,N_19065,N_18126);
nor U21647 (N_21647,N_19068,N_19409);
nand U21648 (N_21648,N_18087,N_19511);
nand U21649 (N_21649,N_19050,N_19277);
or U21650 (N_21650,N_19014,N_19845);
nand U21651 (N_21651,N_18379,N_19476);
and U21652 (N_21652,N_18598,N_18981);
xnor U21653 (N_21653,N_19528,N_18907);
or U21654 (N_21654,N_18048,N_19953);
and U21655 (N_21655,N_18714,N_18420);
nand U21656 (N_21656,N_19344,N_19304);
xnor U21657 (N_21657,N_18287,N_18816);
nand U21658 (N_21658,N_19860,N_18271);
nand U21659 (N_21659,N_19568,N_19279);
nor U21660 (N_21660,N_18739,N_19364);
or U21661 (N_21661,N_19948,N_18472);
nand U21662 (N_21662,N_19859,N_19601);
nor U21663 (N_21663,N_18775,N_19238);
nand U21664 (N_21664,N_19581,N_19200);
xnor U21665 (N_21665,N_18440,N_18650);
xor U21666 (N_21666,N_19250,N_19956);
xor U21667 (N_21667,N_18934,N_18232);
nand U21668 (N_21668,N_19852,N_18361);
or U21669 (N_21669,N_19458,N_19079);
xnor U21670 (N_21670,N_19636,N_19298);
nor U21671 (N_21671,N_18178,N_18699);
nor U21672 (N_21672,N_18284,N_19039);
nand U21673 (N_21673,N_18464,N_19452);
or U21674 (N_21674,N_19271,N_19679);
and U21675 (N_21675,N_19784,N_18006);
or U21676 (N_21676,N_19174,N_19008);
xnor U21677 (N_21677,N_18714,N_19621);
nor U21678 (N_21678,N_18842,N_19295);
and U21679 (N_21679,N_18878,N_19242);
xnor U21680 (N_21680,N_19726,N_19903);
or U21681 (N_21681,N_19150,N_18848);
and U21682 (N_21682,N_18735,N_19152);
and U21683 (N_21683,N_19327,N_19634);
and U21684 (N_21684,N_19338,N_18085);
and U21685 (N_21685,N_19657,N_19589);
nand U21686 (N_21686,N_19478,N_19835);
or U21687 (N_21687,N_18749,N_18041);
nor U21688 (N_21688,N_18676,N_19641);
nor U21689 (N_21689,N_19158,N_19708);
or U21690 (N_21690,N_18488,N_19034);
nand U21691 (N_21691,N_19489,N_18374);
xor U21692 (N_21692,N_18240,N_18571);
or U21693 (N_21693,N_19164,N_19220);
nand U21694 (N_21694,N_19034,N_19057);
and U21695 (N_21695,N_19595,N_19252);
or U21696 (N_21696,N_19042,N_18185);
and U21697 (N_21697,N_18706,N_19686);
nor U21698 (N_21698,N_19247,N_18903);
nand U21699 (N_21699,N_19198,N_19657);
or U21700 (N_21700,N_18350,N_18617);
nor U21701 (N_21701,N_18800,N_18765);
nor U21702 (N_21702,N_18733,N_19066);
and U21703 (N_21703,N_18962,N_18807);
and U21704 (N_21704,N_19695,N_18826);
nor U21705 (N_21705,N_19574,N_19572);
nor U21706 (N_21706,N_19336,N_18984);
nor U21707 (N_21707,N_19702,N_18358);
nand U21708 (N_21708,N_18686,N_18136);
nor U21709 (N_21709,N_18167,N_18652);
or U21710 (N_21710,N_19678,N_18612);
nand U21711 (N_21711,N_19775,N_18429);
or U21712 (N_21712,N_18881,N_19270);
and U21713 (N_21713,N_19601,N_19974);
and U21714 (N_21714,N_18320,N_19080);
or U21715 (N_21715,N_18851,N_19086);
or U21716 (N_21716,N_19549,N_19519);
nor U21717 (N_21717,N_19515,N_18362);
and U21718 (N_21718,N_19213,N_18789);
or U21719 (N_21719,N_19889,N_19856);
and U21720 (N_21720,N_18765,N_18100);
nand U21721 (N_21721,N_18908,N_19340);
xor U21722 (N_21722,N_19751,N_18644);
xor U21723 (N_21723,N_19573,N_18355);
and U21724 (N_21724,N_18556,N_19638);
or U21725 (N_21725,N_19661,N_19611);
xor U21726 (N_21726,N_18029,N_18429);
nand U21727 (N_21727,N_18267,N_18378);
xnor U21728 (N_21728,N_19608,N_19241);
and U21729 (N_21729,N_19770,N_18744);
and U21730 (N_21730,N_18972,N_19522);
and U21731 (N_21731,N_18861,N_19364);
xor U21732 (N_21732,N_18065,N_18367);
and U21733 (N_21733,N_18288,N_18989);
and U21734 (N_21734,N_19081,N_18898);
nand U21735 (N_21735,N_18943,N_18540);
nor U21736 (N_21736,N_19940,N_18110);
xnor U21737 (N_21737,N_19809,N_19520);
or U21738 (N_21738,N_18166,N_18670);
or U21739 (N_21739,N_19551,N_19511);
nand U21740 (N_21740,N_18906,N_19604);
or U21741 (N_21741,N_19123,N_19637);
nor U21742 (N_21742,N_18399,N_19714);
nand U21743 (N_21743,N_19581,N_19751);
and U21744 (N_21744,N_19298,N_19141);
xnor U21745 (N_21745,N_18136,N_19982);
nor U21746 (N_21746,N_18615,N_19188);
nand U21747 (N_21747,N_19048,N_19761);
or U21748 (N_21748,N_19817,N_19353);
xnor U21749 (N_21749,N_19313,N_19938);
and U21750 (N_21750,N_18473,N_18247);
nand U21751 (N_21751,N_18647,N_19526);
nor U21752 (N_21752,N_19183,N_18219);
xor U21753 (N_21753,N_19008,N_19223);
and U21754 (N_21754,N_18930,N_19958);
or U21755 (N_21755,N_19730,N_19335);
nand U21756 (N_21756,N_19032,N_18886);
nand U21757 (N_21757,N_18841,N_19612);
nand U21758 (N_21758,N_18557,N_19413);
nand U21759 (N_21759,N_18597,N_19898);
nor U21760 (N_21760,N_18066,N_18609);
nand U21761 (N_21761,N_18214,N_18742);
or U21762 (N_21762,N_19897,N_19703);
nand U21763 (N_21763,N_19644,N_19077);
xnor U21764 (N_21764,N_19481,N_18578);
or U21765 (N_21765,N_19061,N_18340);
nor U21766 (N_21766,N_18400,N_19257);
and U21767 (N_21767,N_18593,N_19806);
xor U21768 (N_21768,N_18336,N_18938);
xor U21769 (N_21769,N_18300,N_19992);
nor U21770 (N_21770,N_19198,N_18231);
or U21771 (N_21771,N_18954,N_19260);
or U21772 (N_21772,N_19675,N_19272);
or U21773 (N_21773,N_19192,N_18666);
nand U21774 (N_21774,N_18116,N_18564);
or U21775 (N_21775,N_18970,N_19426);
nand U21776 (N_21776,N_19318,N_18364);
nor U21777 (N_21777,N_19658,N_18227);
or U21778 (N_21778,N_18689,N_18796);
and U21779 (N_21779,N_19707,N_18467);
nand U21780 (N_21780,N_18886,N_18726);
nor U21781 (N_21781,N_18285,N_19555);
or U21782 (N_21782,N_19539,N_19326);
nand U21783 (N_21783,N_18220,N_18271);
xor U21784 (N_21784,N_18722,N_19718);
nor U21785 (N_21785,N_19128,N_18872);
and U21786 (N_21786,N_19690,N_19921);
xor U21787 (N_21787,N_18896,N_19511);
nor U21788 (N_21788,N_19886,N_18710);
and U21789 (N_21789,N_18798,N_19769);
and U21790 (N_21790,N_18497,N_18479);
xnor U21791 (N_21791,N_18979,N_19653);
xor U21792 (N_21792,N_18383,N_18612);
nand U21793 (N_21793,N_18217,N_18013);
and U21794 (N_21794,N_19909,N_18832);
nor U21795 (N_21795,N_19067,N_18565);
xor U21796 (N_21796,N_19152,N_18918);
nor U21797 (N_21797,N_18626,N_18756);
and U21798 (N_21798,N_18055,N_18612);
xor U21799 (N_21799,N_19784,N_18605);
and U21800 (N_21800,N_18766,N_18854);
xnor U21801 (N_21801,N_19982,N_18221);
nand U21802 (N_21802,N_19486,N_19048);
xor U21803 (N_21803,N_19568,N_19096);
and U21804 (N_21804,N_19820,N_19921);
and U21805 (N_21805,N_19930,N_19616);
nor U21806 (N_21806,N_19862,N_19186);
xor U21807 (N_21807,N_19784,N_19334);
xor U21808 (N_21808,N_19828,N_18071);
or U21809 (N_21809,N_18113,N_18945);
nor U21810 (N_21810,N_19478,N_18363);
or U21811 (N_21811,N_18570,N_19795);
or U21812 (N_21812,N_19473,N_18659);
or U21813 (N_21813,N_18700,N_19409);
or U21814 (N_21814,N_18042,N_19907);
nand U21815 (N_21815,N_19366,N_18733);
xor U21816 (N_21816,N_19625,N_18169);
and U21817 (N_21817,N_19463,N_19110);
xor U21818 (N_21818,N_19738,N_18694);
nand U21819 (N_21819,N_18959,N_19729);
and U21820 (N_21820,N_19857,N_18929);
nand U21821 (N_21821,N_19417,N_19050);
nor U21822 (N_21822,N_18300,N_18401);
nor U21823 (N_21823,N_18944,N_19540);
and U21824 (N_21824,N_19185,N_19283);
nor U21825 (N_21825,N_19765,N_19246);
nand U21826 (N_21826,N_19542,N_18496);
nor U21827 (N_21827,N_19497,N_18313);
nand U21828 (N_21828,N_19489,N_19740);
and U21829 (N_21829,N_18530,N_19813);
or U21830 (N_21830,N_18304,N_18761);
nand U21831 (N_21831,N_19202,N_18441);
or U21832 (N_21832,N_19598,N_18477);
or U21833 (N_21833,N_19124,N_18003);
xor U21834 (N_21834,N_18197,N_18887);
nand U21835 (N_21835,N_18943,N_19192);
or U21836 (N_21836,N_18315,N_18842);
or U21837 (N_21837,N_18224,N_18644);
xnor U21838 (N_21838,N_18000,N_18914);
and U21839 (N_21839,N_19467,N_19057);
nand U21840 (N_21840,N_19806,N_18758);
nor U21841 (N_21841,N_19493,N_19618);
xor U21842 (N_21842,N_18637,N_19584);
and U21843 (N_21843,N_19290,N_19613);
and U21844 (N_21844,N_18319,N_19039);
xor U21845 (N_21845,N_19732,N_19508);
or U21846 (N_21846,N_18813,N_18761);
nor U21847 (N_21847,N_19107,N_19314);
nor U21848 (N_21848,N_18158,N_18570);
and U21849 (N_21849,N_18231,N_19145);
xor U21850 (N_21850,N_19378,N_19506);
or U21851 (N_21851,N_19834,N_18825);
nor U21852 (N_21852,N_19029,N_19714);
nand U21853 (N_21853,N_19302,N_19835);
and U21854 (N_21854,N_18783,N_18514);
and U21855 (N_21855,N_19478,N_19897);
nor U21856 (N_21856,N_19916,N_18679);
nand U21857 (N_21857,N_19845,N_18758);
nor U21858 (N_21858,N_18245,N_19495);
nand U21859 (N_21859,N_18077,N_19532);
nand U21860 (N_21860,N_18951,N_18696);
nand U21861 (N_21861,N_19276,N_19231);
nor U21862 (N_21862,N_19530,N_18641);
and U21863 (N_21863,N_18847,N_18425);
xor U21864 (N_21864,N_19655,N_19758);
nor U21865 (N_21865,N_19391,N_19419);
or U21866 (N_21866,N_19848,N_19273);
xor U21867 (N_21867,N_18034,N_18222);
or U21868 (N_21868,N_19135,N_19004);
and U21869 (N_21869,N_18481,N_18734);
nand U21870 (N_21870,N_18176,N_19283);
and U21871 (N_21871,N_18731,N_19262);
nand U21872 (N_21872,N_19422,N_19810);
and U21873 (N_21873,N_18687,N_18804);
nand U21874 (N_21874,N_18186,N_19425);
xnor U21875 (N_21875,N_19719,N_19672);
and U21876 (N_21876,N_18661,N_19730);
nand U21877 (N_21877,N_18399,N_18672);
and U21878 (N_21878,N_19483,N_19366);
nand U21879 (N_21879,N_18878,N_18178);
xnor U21880 (N_21880,N_18556,N_18704);
nor U21881 (N_21881,N_18050,N_19744);
xor U21882 (N_21882,N_18976,N_19481);
or U21883 (N_21883,N_19134,N_19487);
xnor U21884 (N_21884,N_18383,N_19956);
xor U21885 (N_21885,N_18786,N_18223);
xor U21886 (N_21886,N_19922,N_18598);
or U21887 (N_21887,N_18318,N_18975);
or U21888 (N_21888,N_18400,N_18746);
nor U21889 (N_21889,N_19114,N_19053);
and U21890 (N_21890,N_19445,N_18811);
nor U21891 (N_21891,N_19250,N_19316);
nor U21892 (N_21892,N_19483,N_19571);
and U21893 (N_21893,N_18793,N_19691);
nand U21894 (N_21894,N_19190,N_19681);
nand U21895 (N_21895,N_19218,N_19120);
and U21896 (N_21896,N_18960,N_19566);
or U21897 (N_21897,N_18950,N_18334);
or U21898 (N_21898,N_19153,N_18552);
nand U21899 (N_21899,N_18684,N_19281);
nand U21900 (N_21900,N_18786,N_18116);
or U21901 (N_21901,N_19917,N_18692);
xor U21902 (N_21902,N_19350,N_19299);
nand U21903 (N_21903,N_18323,N_19981);
or U21904 (N_21904,N_19500,N_18066);
nor U21905 (N_21905,N_18948,N_18013);
xnor U21906 (N_21906,N_18112,N_19469);
nand U21907 (N_21907,N_18981,N_19933);
or U21908 (N_21908,N_18988,N_18490);
nor U21909 (N_21909,N_18544,N_19033);
and U21910 (N_21910,N_19511,N_19807);
or U21911 (N_21911,N_19362,N_18667);
xnor U21912 (N_21912,N_19141,N_19341);
nor U21913 (N_21913,N_18707,N_19079);
xnor U21914 (N_21914,N_19802,N_19942);
xnor U21915 (N_21915,N_18065,N_19665);
and U21916 (N_21916,N_18284,N_18416);
nand U21917 (N_21917,N_18200,N_19249);
nand U21918 (N_21918,N_18378,N_19576);
nor U21919 (N_21919,N_18037,N_18418);
nand U21920 (N_21920,N_19284,N_18515);
and U21921 (N_21921,N_18663,N_19992);
xnor U21922 (N_21922,N_19578,N_18396);
and U21923 (N_21923,N_19637,N_18136);
and U21924 (N_21924,N_19785,N_19959);
and U21925 (N_21925,N_19681,N_19771);
nor U21926 (N_21926,N_19770,N_18666);
xor U21927 (N_21927,N_18955,N_19165);
nand U21928 (N_21928,N_19540,N_18821);
xor U21929 (N_21929,N_19207,N_19152);
nand U21930 (N_21930,N_18182,N_19381);
and U21931 (N_21931,N_18651,N_18376);
nor U21932 (N_21932,N_18513,N_19161);
and U21933 (N_21933,N_18070,N_18875);
and U21934 (N_21934,N_18473,N_18140);
xnor U21935 (N_21935,N_18305,N_18055);
or U21936 (N_21936,N_19978,N_18478);
or U21937 (N_21937,N_19394,N_19004);
or U21938 (N_21938,N_18246,N_18462);
nand U21939 (N_21939,N_18632,N_19005);
nor U21940 (N_21940,N_18043,N_19243);
or U21941 (N_21941,N_18550,N_19936);
xor U21942 (N_21942,N_18970,N_18362);
xor U21943 (N_21943,N_18968,N_19920);
or U21944 (N_21944,N_18387,N_19043);
nor U21945 (N_21945,N_19140,N_18737);
xor U21946 (N_21946,N_18324,N_18805);
nor U21947 (N_21947,N_18951,N_19088);
xor U21948 (N_21948,N_18011,N_18421);
and U21949 (N_21949,N_19726,N_19170);
and U21950 (N_21950,N_18088,N_18752);
or U21951 (N_21951,N_18546,N_18777);
nor U21952 (N_21952,N_18268,N_18472);
or U21953 (N_21953,N_19981,N_19587);
xnor U21954 (N_21954,N_18552,N_19691);
and U21955 (N_21955,N_18103,N_18716);
or U21956 (N_21956,N_19655,N_19793);
nand U21957 (N_21957,N_19235,N_18468);
nand U21958 (N_21958,N_19650,N_19109);
xnor U21959 (N_21959,N_18011,N_18417);
nand U21960 (N_21960,N_19161,N_18555);
and U21961 (N_21961,N_18985,N_18656);
xor U21962 (N_21962,N_18145,N_19323);
xor U21963 (N_21963,N_19385,N_19079);
nor U21964 (N_21964,N_18281,N_18227);
and U21965 (N_21965,N_18758,N_19610);
and U21966 (N_21966,N_18306,N_18578);
nand U21967 (N_21967,N_18433,N_18592);
nand U21968 (N_21968,N_19257,N_18670);
xnor U21969 (N_21969,N_19148,N_18476);
or U21970 (N_21970,N_19645,N_19186);
xor U21971 (N_21971,N_18570,N_18914);
xnor U21972 (N_21972,N_18065,N_19854);
and U21973 (N_21973,N_19329,N_18052);
nand U21974 (N_21974,N_19426,N_18449);
xnor U21975 (N_21975,N_18177,N_18219);
and U21976 (N_21976,N_18098,N_19100);
nor U21977 (N_21977,N_19254,N_18161);
and U21978 (N_21978,N_19427,N_18050);
or U21979 (N_21979,N_18530,N_18868);
nor U21980 (N_21980,N_18709,N_19755);
xnor U21981 (N_21981,N_18638,N_18547);
nor U21982 (N_21982,N_19754,N_19144);
and U21983 (N_21983,N_18905,N_19598);
or U21984 (N_21984,N_19650,N_18926);
or U21985 (N_21985,N_18620,N_18221);
nand U21986 (N_21986,N_19273,N_19994);
xnor U21987 (N_21987,N_19846,N_19144);
and U21988 (N_21988,N_19392,N_18762);
nand U21989 (N_21989,N_19382,N_18535);
and U21990 (N_21990,N_18654,N_19569);
nand U21991 (N_21991,N_18205,N_19418);
or U21992 (N_21992,N_19559,N_18282);
and U21993 (N_21993,N_18848,N_19754);
nor U21994 (N_21994,N_19094,N_19153);
xor U21995 (N_21995,N_19748,N_19481);
nand U21996 (N_21996,N_19167,N_19362);
and U21997 (N_21997,N_18024,N_18138);
xnor U21998 (N_21998,N_18806,N_19781);
or U21999 (N_21999,N_19209,N_18082);
xnor U22000 (N_22000,N_20979,N_20994);
nor U22001 (N_22001,N_20297,N_21370);
xor U22002 (N_22002,N_21132,N_20524);
or U22003 (N_22003,N_20447,N_20458);
nor U22004 (N_22004,N_20313,N_21025);
and U22005 (N_22005,N_21588,N_20263);
or U22006 (N_22006,N_20151,N_21937);
or U22007 (N_22007,N_21958,N_21286);
xnor U22008 (N_22008,N_20480,N_21854);
nand U22009 (N_22009,N_21753,N_20248);
and U22010 (N_22010,N_20354,N_21026);
xnor U22011 (N_22011,N_20476,N_20906);
nor U22012 (N_22012,N_20877,N_20680);
or U22013 (N_22013,N_21528,N_21624);
nor U22014 (N_22014,N_21084,N_21341);
nand U22015 (N_22015,N_21147,N_21758);
xnor U22016 (N_22016,N_20440,N_21351);
and U22017 (N_22017,N_21844,N_20580);
xor U22018 (N_22018,N_20791,N_21731);
xnor U22019 (N_22019,N_21041,N_21682);
or U22020 (N_22020,N_21740,N_21587);
or U22021 (N_22021,N_20742,N_21849);
or U22022 (N_22022,N_21651,N_21436);
nor U22023 (N_22023,N_20144,N_20006);
nor U22024 (N_22024,N_21563,N_21934);
nand U22025 (N_22025,N_21979,N_21853);
or U22026 (N_22026,N_21020,N_21851);
and U22027 (N_22027,N_21306,N_21035);
nor U22028 (N_22028,N_20556,N_20661);
and U22029 (N_22029,N_21835,N_21227);
and U22030 (N_22030,N_21989,N_20893);
nand U22031 (N_22031,N_21481,N_20783);
xnor U22032 (N_22032,N_21164,N_20504);
xnor U22033 (N_22033,N_20181,N_21745);
nor U22034 (N_22034,N_21580,N_20849);
nand U22035 (N_22035,N_20083,N_21906);
and U22036 (N_22036,N_20364,N_20891);
xnor U22037 (N_22037,N_20063,N_20406);
nand U22038 (N_22038,N_20434,N_21149);
xnor U22039 (N_22039,N_21640,N_21942);
or U22040 (N_22040,N_21022,N_21335);
nand U22041 (N_22041,N_20191,N_20179);
or U22042 (N_22042,N_20931,N_21644);
nand U22043 (N_22043,N_20190,N_21135);
xnor U22044 (N_22044,N_20127,N_20587);
xnor U22045 (N_22045,N_21977,N_20177);
and U22046 (N_22046,N_21599,N_21858);
xnor U22047 (N_22047,N_21703,N_21032);
nand U22048 (N_22048,N_20643,N_20465);
xnor U22049 (N_22049,N_20666,N_20638);
or U22050 (N_22050,N_20139,N_20096);
or U22051 (N_22051,N_20142,N_20820);
nand U22052 (N_22052,N_21260,N_20544);
xor U22053 (N_22053,N_21133,N_20763);
and U22054 (N_22054,N_20199,N_20284);
or U22055 (N_22055,N_20049,N_20419);
nand U22056 (N_22056,N_21261,N_21760);
nand U22057 (N_22057,N_21313,N_21500);
and U22058 (N_22058,N_21901,N_20082);
and U22059 (N_22059,N_20050,N_20795);
nand U22060 (N_22060,N_21179,N_20037);
nor U22061 (N_22061,N_20609,N_21560);
nand U22062 (N_22062,N_20414,N_21419);
and U22063 (N_22063,N_21607,N_20528);
nor U22064 (N_22064,N_21876,N_21982);
xor U22065 (N_22065,N_20123,N_20631);
or U22066 (N_22066,N_20099,N_21763);
nand U22067 (N_22067,N_21031,N_21669);
xnor U22068 (N_22068,N_20409,N_21966);
nor U22069 (N_22069,N_21173,N_21476);
or U22070 (N_22070,N_20101,N_21935);
xor U22071 (N_22071,N_20028,N_21023);
and U22072 (N_22072,N_20714,N_21027);
nor U22073 (N_22073,N_20615,N_20776);
and U22074 (N_22074,N_21093,N_21330);
nor U22075 (N_22075,N_20390,N_21076);
nand U22076 (N_22076,N_21533,N_21015);
nor U22077 (N_22077,N_21328,N_20016);
nand U22078 (N_22078,N_21984,N_21245);
nand U22079 (N_22079,N_20106,N_20278);
nor U22080 (N_22080,N_20721,N_20612);
and U22081 (N_22081,N_21929,N_20892);
or U22082 (N_22082,N_21034,N_21424);
nor U22083 (N_22083,N_20235,N_20244);
xor U22084 (N_22084,N_20208,N_20607);
nand U22085 (N_22085,N_20462,N_21111);
nand U22086 (N_22086,N_21878,N_21414);
and U22087 (N_22087,N_20232,N_20094);
nor U22088 (N_22088,N_21770,N_20936);
or U22089 (N_22089,N_21113,N_20922);
or U22090 (N_22090,N_21024,N_21812);
nor U22091 (N_22091,N_21267,N_20627);
nor U22092 (N_22092,N_21504,N_21470);
or U22093 (N_22093,N_20312,N_21983);
or U22094 (N_22094,N_20084,N_21761);
and U22095 (N_22095,N_20110,N_20300);
and U22096 (N_22096,N_21492,N_21114);
nand U22097 (N_22097,N_21038,N_20495);
nor U22098 (N_22098,N_21980,N_20808);
nand U22099 (N_22099,N_21943,N_20575);
nor U22100 (N_22100,N_20402,N_21695);
xnor U22101 (N_22101,N_21461,N_21386);
nand U22102 (N_22102,N_21143,N_20159);
xnor U22103 (N_22103,N_21350,N_20704);
xor U22104 (N_22104,N_20599,N_20441);
xor U22105 (N_22105,N_21839,N_20200);
xor U22106 (N_22106,N_21270,N_20145);
nand U22107 (N_22107,N_20549,N_21898);
or U22108 (N_22108,N_20424,N_20854);
or U22109 (N_22109,N_20886,N_21940);
nor U22110 (N_22110,N_20619,N_20956);
xor U22111 (N_22111,N_20362,N_21304);
xnor U22112 (N_22112,N_20233,N_20871);
and U22113 (N_22113,N_21180,N_20370);
or U22114 (N_22114,N_20448,N_20100);
xor U22115 (N_22115,N_20164,N_21401);
and U22116 (N_22116,N_20496,N_20209);
nor U22117 (N_22117,N_20740,N_21246);
xor U22118 (N_22118,N_20507,N_21442);
and U22119 (N_22119,N_20806,N_21207);
and U22120 (N_22120,N_21721,N_20058);
and U22121 (N_22121,N_20299,N_21961);
and U22122 (N_22122,N_20306,N_20111);
or U22123 (N_22123,N_20147,N_20366);
and U22124 (N_22124,N_21879,N_20463);
and U22125 (N_22125,N_20699,N_21790);
or U22126 (N_22126,N_20718,N_20966);
xnor U22127 (N_22127,N_21503,N_20819);
and U22128 (N_22128,N_20878,N_21441);
nor U22129 (N_22129,N_21948,N_20741);
nand U22130 (N_22130,N_20472,N_21774);
nor U22131 (N_22131,N_20780,N_20098);
nand U22132 (N_22132,N_20381,N_21360);
or U22133 (N_22133,N_20997,N_20959);
and U22134 (N_22134,N_20592,N_20771);
and U22135 (N_22135,N_21233,N_21719);
or U22136 (N_22136,N_20374,N_21174);
and U22137 (N_22137,N_20078,N_20621);
nand U22138 (N_22138,N_20501,N_21828);
xnor U22139 (N_22139,N_20657,N_20725);
xnor U22140 (N_22140,N_20843,N_20975);
or U22141 (N_22141,N_20952,N_21619);
or U22142 (N_22142,N_20969,N_20696);
nor U22143 (N_22143,N_21697,N_20750);
xor U22144 (N_22144,N_20829,N_21380);
or U22145 (N_22145,N_20076,N_20008);
or U22146 (N_22146,N_20392,N_21054);
nand U22147 (N_22147,N_21171,N_21403);
xnor U22148 (N_22148,N_21787,N_21616);
nand U22149 (N_22149,N_20971,N_21987);
xor U22150 (N_22150,N_21791,N_21850);
and U22151 (N_22151,N_20832,N_20389);
nor U22152 (N_22152,N_20505,N_20659);
nor U22153 (N_22153,N_21632,N_21316);
nor U22154 (N_22154,N_20681,N_21680);
or U22155 (N_22155,N_21674,N_21600);
xnor U22156 (N_22156,N_20155,N_20937);
nand U22157 (N_22157,N_20268,N_20410);
or U22158 (N_22158,N_20230,N_21230);
nor U22159 (N_22159,N_20394,N_20197);
and U22160 (N_22160,N_20017,N_21860);
nand U22161 (N_22161,N_21797,N_21451);
xor U22162 (N_22162,N_21488,N_20091);
xnor U22163 (N_22163,N_21271,N_20274);
nor U22164 (N_22164,N_20610,N_20396);
and U22165 (N_22165,N_20692,N_21101);
nand U22166 (N_22166,N_21275,N_20613);
and U22167 (N_22167,N_20803,N_20324);
nor U22168 (N_22168,N_20167,N_21310);
xnor U22169 (N_22169,N_21012,N_20921);
nor U22170 (N_22170,N_21389,N_20796);
nor U22171 (N_22171,N_21375,N_21910);
nand U22172 (N_22172,N_20563,N_21641);
and U22173 (N_22173,N_21709,N_20865);
or U22174 (N_22174,N_21257,N_20288);
nor U22175 (N_22175,N_21971,N_21900);
xnor U22176 (N_22176,N_21505,N_20557);
or U22177 (N_22177,N_20113,N_20383);
xor U22178 (N_22178,N_21339,N_20131);
nor U22179 (N_22179,N_20315,N_21816);
nand U22180 (N_22180,N_21094,N_21701);
or U22181 (N_22181,N_20298,N_20812);
nand U22182 (N_22182,N_21356,N_21265);
nand U22183 (N_22183,N_20015,N_20405);
xnor U22184 (N_22184,N_21725,N_21999);
nand U22185 (N_22185,N_20443,N_21516);
nor U22186 (N_22186,N_21540,N_20686);
xor U22187 (N_22187,N_20273,N_21371);
and U22188 (N_22188,N_21192,N_20941);
xor U22189 (N_22189,N_20851,N_21169);
xnor U22190 (N_22190,N_20107,N_20663);
and U22191 (N_22191,N_21362,N_20104);
nand U22192 (N_22192,N_21873,N_20719);
nand U22193 (N_22193,N_21303,N_21278);
nor U22194 (N_22194,N_21452,N_20207);
xnor U22195 (N_22195,N_20708,N_20259);
or U22196 (N_22196,N_21785,N_21355);
nor U22197 (N_22197,N_21444,N_21123);
xor U22198 (N_22198,N_21105,N_20514);
nor U22199 (N_22199,N_20030,N_21893);
or U22200 (N_22200,N_21450,N_21314);
nor U22201 (N_22201,N_21921,N_20327);
and U22202 (N_22202,N_20706,N_21733);
nand U22203 (N_22203,N_21391,N_20329);
nor U22204 (N_22204,N_20119,N_20055);
nand U22205 (N_22205,N_21794,N_21880);
nor U22206 (N_22206,N_20180,N_21583);
and U22207 (N_22207,N_20464,N_20021);
xnor U22208 (N_22208,N_20797,N_21796);
xor U22209 (N_22209,N_21678,N_20555);
or U22210 (N_22210,N_20925,N_20195);
or U22211 (N_22211,N_20067,N_21170);
xnor U22212 (N_22212,N_21119,N_21384);
nand U22213 (N_22213,N_20927,N_21933);
and U22214 (N_22214,N_21309,N_21736);
and U22215 (N_22215,N_20246,N_21626);
nand U22216 (N_22216,N_20988,N_21460);
nor U22217 (N_22217,N_20918,N_21274);
nand U22218 (N_22218,N_21962,N_20899);
nand U22219 (N_22219,N_20371,N_21550);
nor U22220 (N_22220,N_21675,N_20649);
nor U22221 (N_22221,N_20767,N_20031);
nand U22222 (N_22222,N_20368,N_21568);
nor U22223 (N_22223,N_20081,N_21046);
or U22224 (N_22224,N_21168,N_20814);
nand U22225 (N_22225,N_21637,N_21223);
nand U22226 (N_22226,N_21466,N_20048);
nor U22227 (N_22227,N_21575,N_21001);
xnor U22228 (N_22228,N_20545,N_20828);
nand U22229 (N_22229,N_20384,N_21923);
xnor U22230 (N_22230,N_20429,N_20069);
nor U22231 (N_22231,N_21479,N_20732);
nor U22232 (N_22232,N_21883,N_20001);
or U22233 (N_22233,N_20358,N_21807);
xnor U22234 (N_22234,N_20679,N_21527);
and U22235 (N_22235,N_20532,N_20539);
nand U22236 (N_22236,N_21200,N_20744);
nor U22237 (N_22237,N_21831,N_21726);
and U22238 (N_22238,N_20051,N_20056);
or U22239 (N_22239,N_20601,N_20574);
and U22240 (N_22240,N_21225,N_20225);
xnor U22241 (N_22241,N_20174,N_20748);
and U22242 (N_22242,N_21714,N_21617);
and U22243 (N_22243,N_21609,N_21432);
and U22244 (N_22244,N_21236,N_21250);
or U22245 (N_22245,N_20333,N_20729);
and U22246 (N_22246,N_20754,N_21213);
or U22247 (N_22247,N_20917,N_20606);
or U22248 (N_22248,N_21329,N_20880);
nor U22249 (N_22249,N_20827,N_20401);
or U22250 (N_22250,N_21231,N_21708);
nand U22251 (N_22251,N_20935,N_20249);
nand U22252 (N_22252,N_20261,N_21569);
and U22253 (N_22253,N_20597,N_20901);
or U22254 (N_22254,N_21478,N_21118);
nor U22255 (N_22255,N_21042,N_21829);
and U22256 (N_22256,N_21385,N_20702);
nand U22257 (N_22257,N_20137,N_21212);
nand U22258 (N_22258,N_20942,N_21894);
or U22259 (N_22259,N_20902,N_20486);
and U22260 (N_22260,N_21717,N_21885);
nor U22261 (N_22261,N_21218,N_21882);
and U22262 (N_22262,N_20487,N_20116);
nand U22263 (N_22263,N_21826,N_20385);
or U22264 (N_22264,N_21268,N_20134);
nand U22265 (N_22265,N_21743,N_20608);
or U22266 (N_22266,N_21066,N_21209);
nand U22267 (N_22267,N_21561,N_20430);
nand U22268 (N_22268,N_21017,N_20982);
xnor U22269 (N_22269,N_20962,N_21574);
and U22270 (N_22270,N_21083,N_21315);
xor U22271 (N_22271,N_21413,N_20426);
nand U22272 (N_22272,N_20290,N_20378);
xnor U22273 (N_22273,N_20347,N_21486);
or U22274 (N_22274,N_20240,N_20075);
nand U22275 (N_22275,N_20624,N_21198);
nand U22276 (N_22276,N_21160,N_20964);
nor U22277 (N_22277,N_20872,N_21348);
nand U22278 (N_22278,N_21764,N_21827);
and U22279 (N_22279,N_20816,N_21889);
or U22280 (N_22280,N_20662,N_21082);
nand U22281 (N_22281,N_20046,N_20227);
and U22282 (N_22282,N_20451,N_21166);
or U22283 (N_22283,N_20784,N_20432);
or U22284 (N_22284,N_20667,N_21875);
or U22285 (N_22285,N_21756,N_20913);
or U22286 (N_22286,N_21472,N_21021);
or U22287 (N_22287,N_20326,N_21802);
or U22288 (N_22288,N_21463,N_21089);
and U22289 (N_22289,N_20656,N_21102);
nor U22290 (N_22290,N_20171,N_21751);
xor U22291 (N_22291,N_21103,N_21454);
xor U22292 (N_22292,N_20033,N_21792);
nor U22293 (N_22293,N_20221,N_21959);
nor U22294 (N_22294,N_21992,N_20437);
xor U22295 (N_22295,N_21194,N_21811);
nand U22296 (N_22296,N_20277,N_20143);
xnor U22297 (N_22297,N_20639,N_21614);
nor U22298 (N_22298,N_20509,N_20452);
xnor U22299 (N_22299,N_21493,N_20963);
or U22300 (N_22300,N_21523,N_21221);
xnor U22301 (N_22301,N_20674,N_20090);
and U22302 (N_22302,N_21353,N_20325);
or U22303 (N_22303,N_21671,N_21543);
or U22304 (N_22304,N_21251,N_21960);
and U22305 (N_22305,N_20337,N_21117);
or U22306 (N_22306,N_20894,N_21446);
nand U22307 (N_22307,N_21566,N_20735);
xor U22308 (N_22308,N_20520,N_21418);
xor U22309 (N_22309,N_21810,N_20810);
or U22310 (N_22310,N_20086,N_20265);
nand U22311 (N_22311,N_21998,N_21468);
or U22312 (N_22312,N_20372,N_21145);
or U22313 (N_22313,N_20074,N_20883);
and U22314 (N_22314,N_20834,N_20547);
nand U22315 (N_22315,N_21321,N_21919);
xor U22316 (N_22316,N_21866,N_20045);
nor U22317 (N_22317,N_20237,N_21120);
nor U22318 (N_22318,N_21405,N_21646);
or U22319 (N_22319,N_21320,N_20204);
xor U22320 (N_22320,N_20126,N_20635);
nand U22321 (N_22321,N_21427,N_20940);
xor U22322 (N_22322,N_21228,N_20813);
nand U22323 (N_22323,N_20926,N_20904);
or U22324 (N_22324,N_20169,N_20178);
nor U22325 (N_22325,N_20512,N_21097);
xor U22326 (N_22326,N_21175,N_20752);
or U22327 (N_22327,N_20453,N_21429);
nand U22328 (N_22328,N_20998,N_20855);
nor U22329 (N_22329,N_20737,N_21475);
and U22330 (N_22330,N_20584,N_21287);
xor U22331 (N_22331,N_21045,N_20565);
nand U22332 (N_22332,N_21440,N_20972);
nor U22333 (N_22333,N_21474,N_20529);
and U22334 (N_22334,N_21975,N_21292);
nand U22335 (N_22335,N_21155,N_20160);
and U22336 (N_22336,N_21392,N_21673);
or U22337 (N_22337,N_21272,N_20822);
nor U22338 (N_22338,N_20567,N_21724);
or U22339 (N_22339,N_20889,N_20411);
xnor U22340 (N_22340,N_21229,N_21871);
and U22341 (N_22341,N_21577,N_20036);
xor U22342 (N_22342,N_20319,N_20720);
xnor U22343 (N_22343,N_20003,N_21300);
nand U22344 (N_22344,N_20571,N_20672);
or U22345 (N_22345,N_20590,N_21817);
and U22346 (N_22346,N_21480,N_21060);
nand U22347 (N_22347,N_21549,N_21555);
nor U22348 (N_22348,N_20576,N_20837);
nand U22349 (N_22349,N_20664,N_21859);
nor U22350 (N_22350,N_20749,N_20182);
nor U22351 (N_22351,N_21634,N_20218);
nand U22352 (N_22352,N_20054,N_21397);
nand U22353 (N_22353,N_20646,N_20782);
and U22354 (N_22354,N_21264,N_20882);
nand U22355 (N_22355,N_21576,N_21109);
xor U22356 (N_22356,N_21006,N_20488);
nand U22357 (N_22357,N_20561,N_20217);
nor U22358 (N_22358,N_21752,N_21704);
nor U22359 (N_22359,N_21242,N_20541);
or U22360 (N_22360,N_20665,N_21131);
nand U22361 (N_22361,N_20951,N_20043);
or U22362 (N_22362,N_20734,N_21165);
and U22363 (N_22363,N_21888,N_20196);
or U22364 (N_22364,N_21501,N_20421);
nor U22365 (N_22365,N_21459,N_21957);
and U22366 (N_22366,N_20617,N_21345);
nor U22367 (N_22367,N_21520,N_20356);
or U22368 (N_22368,N_21579,N_20467);
nor U22369 (N_22369,N_20009,N_21840);
nor U22370 (N_22370,N_20915,N_21650);
or U22371 (N_22371,N_21638,N_21630);
nand U22372 (N_22372,N_20953,N_20236);
nor U22373 (N_22373,N_21473,N_21902);
xor U22374 (N_22374,N_21772,N_21255);
nand U22375 (N_22375,N_20559,N_21605);
nand U22376 (N_22376,N_20459,N_21915);
and U22377 (N_22377,N_20811,N_20032);
nand U22378 (N_22378,N_21435,N_21047);
and U22379 (N_22379,N_20468,N_20436);
and U22380 (N_22380,N_20360,N_20778);
and U22381 (N_22381,N_21127,N_21620);
and U22382 (N_22382,N_21290,N_21707);
and U22383 (N_22383,N_21623,N_20690);
and U22384 (N_22384,N_21307,N_21532);
xnor U22385 (N_22385,N_20109,N_20577);
or U22386 (N_22386,N_20637,N_21057);
or U22387 (N_22387,N_20404,N_20391);
nor U22388 (N_22388,N_21542,N_20205);
xor U22389 (N_22389,N_20890,N_21603);
nand U22390 (N_22390,N_20794,N_21727);
xor U22391 (N_22391,N_20841,N_20731);
and U22392 (N_22392,N_21358,N_21841);
nor U22393 (N_22393,N_20546,N_21639);
nand U22394 (N_22394,N_21412,N_20117);
xor U22395 (N_22395,N_21586,N_20618);
and U22396 (N_22396,N_20628,N_21039);
xor U22397 (N_22397,N_20961,N_21720);
or U22398 (N_22398,N_21621,N_20336);
nor U22399 (N_22399,N_20641,N_20395);
xnor U22400 (N_22400,N_21154,N_21662);
or U22401 (N_22401,N_20620,N_21092);
and U22402 (N_22402,N_20438,N_21409);
nor U22403 (N_22403,N_21633,N_20747);
and U22404 (N_22404,N_21383,N_21676);
and U22405 (N_22405,N_21125,N_20755);
nand U22406 (N_22406,N_21730,N_20603);
xnor U22407 (N_22407,N_21053,N_20611);
and U22408 (N_22408,N_20586,N_20057);
and U22409 (N_22409,N_21837,N_21100);
xnor U22410 (N_22410,N_21106,N_20685);
nand U22411 (N_22411,N_20884,N_21498);
nor U22412 (N_22412,N_20760,N_21604);
nor U22413 (N_22413,N_20991,N_21453);
nand U22414 (N_22414,N_21202,N_21613);
and U22415 (N_22415,N_20152,N_21489);
xor U22416 (N_22416,N_21757,N_21947);
and U22417 (N_22417,N_21234,N_21030);
nor U22418 (N_22418,N_20651,N_20309);
nor U22419 (N_22419,N_20508,N_20616);
xnor U22420 (N_22420,N_21239,N_21417);
and U22421 (N_22421,N_20531,N_21711);
xor U22422 (N_22422,N_21028,N_21685);
and U22423 (N_22423,N_21477,N_20569);
or U22424 (N_22424,N_21819,N_20012);
and U22425 (N_22425,N_20594,N_20198);
nor U22426 (N_22426,N_21954,N_21856);
or U22427 (N_22427,N_20766,N_20289);
nand U22428 (N_22428,N_20490,N_20060);
nor U22429 (N_22429,N_20302,N_21014);
nand U22430 (N_22430,N_21136,N_21546);
xor U22431 (N_22431,N_21536,N_20984);
nand U22432 (N_22432,N_20713,N_21611);
or U22433 (N_22433,N_20976,N_21808);
and U22434 (N_22434,N_20990,N_21352);
nand U22435 (N_22435,N_21924,N_21618);
and U22436 (N_22436,N_21151,N_21996);
xor U22437 (N_22437,N_21464,N_20818);
xor U22438 (N_22438,N_21931,N_20642);
or U22439 (N_22439,N_20670,N_21467);
or U22440 (N_22440,N_21944,N_20138);
nand U22441 (N_22441,N_21273,N_20423);
xnor U22442 (N_22442,N_20562,N_21085);
nor U22443 (N_22443,N_21890,N_21129);
or U22444 (N_22444,N_21248,N_20420);
or U22445 (N_22445,N_21593,N_21897);
nor U22446 (N_22446,N_20064,N_21868);
and U22447 (N_22447,N_21184,N_20220);
nand U22448 (N_22448,N_20231,N_20156);
nand U22449 (N_22449,N_20772,N_20353);
nand U22450 (N_22450,N_20492,N_21696);
nand U22451 (N_22451,N_20296,N_21116);
and U22452 (N_22452,N_21469,N_21778);
xnor U22453 (N_22453,N_20916,N_21612);
nand U22454 (N_22454,N_20342,N_21997);
and U22455 (N_22455,N_21908,N_21657);
nor U22456 (N_22456,N_20867,N_21738);
xnor U22457 (N_22457,N_20470,N_21416);
nor U22458 (N_22458,N_20630,N_21318);
xnor U22459 (N_22459,N_20595,N_21359);
xor U22460 (N_22460,N_21050,N_21277);
nand U22461 (N_22461,N_20422,N_21055);
nand U22462 (N_22462,N_20632,N_21496);
xor U22463 (N_22463,N_20193,N_21596);
or U22464 (N_22464,N_20241,N_20777);
or U22465 (N_22465,N_20321,N_21535);
nand U22466 (N_22466,N_21573,N_21814);
nand U22467 (N_22467,N_21016,N_20591);
xnor U22468 (N_22468,N_21346,N_21508);
xnor U22469 (N_22469,N_21390,N_21506);
or U22470 (N_22470,N_21404,N_20516);
or U22471 (N_22471,N_21455,N_20482);
nor U22472 (N_22472,N_21216,N_21558);
or U22473 (N_22473,N_21767,N_20024);
nor U22474 (N_22474,N_20251,N_21056);
nor U22475 (N_22475,N_21728,N_21064);
or U22476 (N_22476,N_20558,N_20022);
and U22477 (N_22477,N_21559,N_20564);
or U22478 (N_22478,N_20427,N_20053);
nand U22479 (N_22479,N_21208,N_21693);
or U22480 (N_22480,N_20623,N_20910);
and U22481 (N_22481,N_20560,N_20187);
xnor U22482 (N_22482,N_21737,N_21421);
and U22483 (N_22483,N_20311,N_20762);
xnor U22484 (N_22484,N_21780,N_20140);
nor U22485 (N_22485,N_21553,N_21956);
xor U22486 (N_22486,N_21019,N_20184);
or U22487 (N_22487,N_20214,N_21153);
xor U22488 (N_22488,N_20773,N_21482);
and U22489 (N_22489,N_21063,N_21688);
xnor U22490 (N_22490,N_20072,N_20779);
xnor U22491 (N_22491,N_21144,N_20023);
xor U22492 (N_22492,N_20000,N_20223);
or U22493 (N_22493,N_20552,N_20280);
nor U22494 (N_22494,N_20826,N_21215);
xor U22495 (N_22495,N_21946,N_21594);
nor U22496 (N_22496,N_21043,N_20363);
or U22497 (N_22497,N_21428,N_20838);
nor U22498 (N_22498,N_21694,N_20888);
or U22499 (N_22499,N_21995,N_20379);
nand U22500 (N_22500,N_20407,N_21052);
nand U22501 (N_22501,N_21950,N_21293);
nor U22502 (N_22502,N_20040,N_20474);
nand U22503 (N_22503,N_20722,N_21065);
xor U22504 (N_22504,N_20678,N_21491);
nor U22505 (N_22505,N_20213,N_20864);
xor U22506 (N_22506,N_20707,N_20108);
nand U22507 (N_22507,N_20581,N_20629);
xor U22508 (N_22508,N_20967,N_21379);
or U22509 (N_22509,N_20660,N_21554);
and U22510 (N_22510,N_21338,N_21846);
or U22511 (N_22511,N_21661,N_20253);
or U22512 (N_22512,N_21237,N_20317);
xnor U22513 (N_22513,N_20761,N_21259);
or U22514 (N_22514,N_21773,N_21219);
or U22515 (N_22515,N_21193,N_20602);
xnor U22516 (N_22516,N_21140,N_20805);
xor U22517 (N_22517,N_21515,N_20435);
xnor U22518 (N_22518,N_20185,N_20987);
or U22519 (N_22519,N_21146,N_20283);
xnor U22520 (N_22520,N_20002,N_20345);
nand U22521 (N_22521,N_20946,N_21253);
and U22522 (N_22522,N_20092,N_21062);
nor U22523 (N_22523,N_21769,N_21422);
and U22524 (N_22524,N_20929,N_21077);
xor U22525 (N_22525,N_21928,N_21938);
nand U22526 (N_22526,N_21627,N_20701);
xnor U22527 (N_22527,N_21917,N_20093);
and U22528 (N_22528,N_20655,N_20537);
nand U22529 (N_22529,N_20700,N_21086);
and U22530 (N_22530,N_20415,N_21005);
nand U22531 (N_22531,N_20573,N_20301);
xnor U22532 (N_22532,N_21196,N_21071);
xnor U22533 (N_22533,N_21142,N_20203);
or U22534 (N_22534,N_21426,N_21112);
and U22535 (N_22535,N_21471,N_20930);
or U22536 (N_22536,N_20781,N_20691);
and U22537 (N_22537,N_20522,N_20141);
xor U22538 (N_22538,N_21582,N_21399);
xor U22539 (N_22539,N_20361,N_21591);
or U22540 (N_22540,N_20332,N_20369);
and U22541 (N_22541,N_21182,N_21494);
nor U22542 (N_22542,N_21571,N_20308);
xor U22543 (N_22543,N_20479,N_20521);
nand U22544 (N_22544,N_20787,N_21203);
xnor U22545 (N_22545,N_20726,N_21718);
or U22546 (N_22546,N_21798,N_21406);
nor U22547 (N_22547,N_20817,N_20483);
nand U22548 (N_22548,N_20793,N_21075);
and U22549 (N_22549,N_21994,N_20695);
or U22550 (N_22550,N_20768,N_20519);
xnor U22551 (N_22551,N_21914,N_20188);
nor U22552 (N_22552,N_21715,N_21201);
nor U22553 (N_22553,N_20846,N_20938);
xnor U22554 (N_22554,N_20102,N_20588);
nor U22555 (N_22555,N_21139,N_21578);
and U22556 (N_22556,N_21013,N_20948);
xor U22557 (N_22557,N_21881,N_21044);
nand U22558 (N_22558,N_21832,N_20874);
and U22559 (N_22559,N_21748,N_21744);
or U22560 (N_22560,N_20873,N_20439);
nor U22561 (N_22561,N_20858,N_20542);
or U22562 (N_22562,N_21226,N_21243);
or U22563 (N_22563,N_21187,N_20993);
xor U22564 (N_22564,N_21331,N_20859);
nor U22565 (N_22565,N_21601,N_20264);
and U22566 (N_22566,N_20500,N_21222);
nor U22567 (N_22567,N_20503,N_21423);
and U22568 (N_22568,N_20355,N_20318);
nand U22569 (N_22569,N_21296,N_21162);
xnor U22570 (N_22570,N_20758,N_20216);
nand U22571 (N_22571,N_20007,N_21333);
or U22572 (N_22572,N_21658,N_20455);
and U22573 (N_22573,N_20433,N_20980);
nand U22574 (N_22574,N_21903,N_20010);
xnor U22575 (N_22575,N_21936,N_20088);
or U22576 (N_22576,N_20089,N_20215);
xor U22577 (N_22577,N_20044,N_21666);
and U22578 (N_22578,N_20676,N_21159);
and U22579 (N_22579,N_21340,N_21869);
xnor U22580 (N_22580,N_21647,N_21415);
xnor U22581 (N_22581,N_20693,N_21402);
and U22582 (N_22582,N_21301,N_20408);
nand U22583 (N_22583,N_21029,N_20943);
nand U22584 (N_22584,N_20112,N_20981);
nor U22585 (N_22585,N_20517,N_21369);
or U22586 (N_22586,N_21070,N_20716);
xnor U22587 (N_22587,N_21702,N_20034);
and U22588 (N_22588,N_21249,N_20469);
nor U22589 (N_22589,N_21930,N_20499);
nand U22590 (N_22590,N_21766,N_20417);
nor U22591 (N_22591,N_21280,N_21801);
nor U22592 (N_22592,N_21606,N_20689);
or U22593 (N_22593,N_20029,N_21795);
xnor U22594 (N_22594,N_21199,N_20377);
or U22595 (N_22595,N_21972,N_21407);
xnor U22596 (N_22596,N_21434,N_20267);
nor U22597 (N_22597,N_21848,N_21297);
xor U22598 (N_22598,N_20566,N_20282);
or U22599 (N_22599,N_21509,N_20166);
nand U22600 (N_22600,N_20799,N_21456);
xor U22601 (N_22601,N_20157,N_21376);
nand U22602 (N_22602,N_20367,N_21420);
nand U22603 (N_22603,N_21152,N_21592);
xnor U22604 (N_22604,N_21679,N_21939);
xor U22605 (N_22605,N_21667,N_21279);
nor U22606 (N_22606,N_20323,N_20885);
nand U22607 (N_22607,N_21706,N_21608);
xor U22608 (N_22608,N_21525,N_21539);
or U22609 (N_22609,N_20572,N_21864);
xor U22610 (N_22610,N_20992,N_20425);
nand U22611 (N_22611,N_20004,N_21779);
xnor U22612 (N_22612,N_21514,N_21311);
and U22613 (N_22613,N_20634,N_21263);
or U22614 (N_22614,N_21564,N_21110);
xor U22615 (N_22615,N_21932,N_20989);
nand U22616 (N_22616,N_20122,N_21628);
and U22617 (N_22617,N_20996,N_20307);
nand U22618 (N_22618,N_20944,N_21993);
nand U22619 (N_22619,N_21965,N_21244);
nand U22620 (N_22620,N_21211,N_20730);
nor U22621 (N_22621,N_21590,N_21663);
and U22622 (N_22622,N_21002,N_20645);
and U22623 (N_22623,N_21513,N_21378);
xor U22624 (N_22624,N_21815,N_20176);
and U22625 (N_22625,N_20228,N_21317);
nor U22626 (N_22626,N_21217,N_20852);
xnor U22627 (N_22627,N_20568,N_21156);
nand U22628 (N_22628,N_21659,N_21312);
nand U22629 (N_22629,N_21357,N_21343);
nor U22630 (N_22630,N_21677,N_20305);
xnor U22631 (N_22631,N_20728,N_21088);
nor U22632 (N_22632,N_21134,N_20310);
nand U22633 (N_22633,N_20523,N_21095);
nor U22634 (N_22634,N_21326,N_21813);
nand U22635 (N_22635,N_20365,N_21368);
and U22636 (N_22636,N_21665,N_21865);
and U22637 (N_22637,N_20484,N_21765);
and U22638 (N_22638,N_21003,N_21631);
nor U22639 (N_22639,N_21425,N_20711);
nand U22640 (N_22640,N_21195,N_20879);
nand U22641 (N_22641,N_21625,N_21204);
or U22642 (N_22642,N_21091,N_20038);
xor U22643 (N_22643,N_21394,N_21305);
nand U22644 (N_22644,N_20554,N_20790);
nand U22645 (N_22645,N_20478,N_21214);
xor U22646 (N_22646,N_21762,N_20173);
or U22647 (N_22647,N_21820,N_21862);
or U22648 (N_22648,N_21258,N_20821);
and U22649 (N_22649,N_20292,N_21051);
and U22650 (N_22650,N_21235,N_21288);
nand U22651 (N_22651,N_21282,N_21185);
nand U22652 (N_22652,N_21684,N_21884);
or U22653 (N_22653,N_21354,N_21439);
xor U22654 (N_22654,N_21495,N_21926);
nand U22655 (N_22655,N_21499,N_21598);
and U22656 (N_22656,N_20243,N_20738);
xor U22657 (N_22657,N_21449,N_21768);
nand U22658 (N_22658,N_20005,N_20121);
xnor U22659 (N_22659,N_20958,N_21518);
and U22660 (N_22660,N_20792,N_20403);
nor U22661 (N_22661,N_21830,N_21531);
and U22662 (N_22662,N_20589,N_20842);
nand U22663 (N_22663,N_21913,N_21955);
nand U22664 (N_22664,N_21689,N_20065);
nor U22665 (N_22665,N_20120,N_21344);
nand U22666 (N_22666,N_20168,N_21845);
xor U22667 (N_22667,N_21252,N_20898);
nor U22668 (N_22668,N_21821,N_20900);
nor U22669 (N_22669,N_21782,N_20019);
and U22670 (N_22670,N_20857,N_21803);
nor U22671 (N_22671,N_21324,N_21699);
or U22672 (N_22672,N_21256,N_21157);
xor U22673 (N_22673,N_20850,N_21789);
nor U22674 (N_22674,N_20491,N_21447);
or U22675 (N_22675,N_21723,N_21400);
and U22676 (N_22676,N_20511,N_21781);
nand U22677 (N_22677,N_21483,N_21487);
and U22678 (N_22678,N_21602,N_20743);
or U22679 (N_22679,N_20148,N_21870);
nor U22680 (N_22680,N_21777,N_21090);
or U22681 (N_22681,N_20085,N_21004);
or U22682 (N_22682,N_20399,N_21905);
and U22683 (N_22683,N_21167,N_21068);
or U22684 (N_22684,N_21081,N_20945);
xor U22685 (N_22685,N_20442,N_21735);
xor U22686 (N_22686,N_20271,N_20445);
and U22687 (N_22687,N_21284,N_21886);
or U22688 (N_22688,N_21567,N_20153);
nor U22689 (N_22689,N_21319,N_21976);
and U22690 (N_22690,N_20047,N_21534);
and U22691 (N_22691,N_20359,N_21299);
nor U22692 (N_22692,N_21224,N_20536);
or U22693 (N_22693,N_21867,N_20165);
or U22694 (N_22694,N_21336,N_21137);
nor U22695 (N_22695,N_21033,N_21654);
xor U22696 (N_22696,N_20183,N_20239);
nor U22697 (N_22697,N_21074,N_21656);
xor U22698 (N_22698,N_20498,N_20041);
xor U22699 (N_22699,N_21430,N_20833);
nor U22700 (N_22700,N_20510,N_21108);
and U22701 (N_22701,N_20757,N_20715);
nand U22702 (N_22702,N_21000,N_20973);
or U22703 (N_22703,N_21981,N_21115);
nor U22704 (N_22704,N_21968,N_20052);
xor U22705 (N_22705,N_21922,N_21842);
and U22706 (N_22706,N_20950,N_21750);
and U22707 (N_22707,N_20331,N_21294);
and U22708 (N_22708,N_21855,N_20061);
or U22709 (N_22709,N_20229,N_20291);
or U22710 (N_22710,N_20908,N_20413);
and U22711 (N_22711,N_20896,N_20132);
and U22712 (N_22712,N_20013,N_21970);
or U22713 (N_22713,N_20759,N_21589);
nor U22714 (N_22714,N_20823,N_21687);
or U22715 (N_22715,N_20694,N_20835);
nor U22716 (N_22716,N_21462,N_20293);
xnor U22717 (N_22717,N_20130,N_20875);
nor U22718 (N_22718,N_21445,N_21529);
xor U22719 (N_22719,N_21843,N_21920);
or U22720 (N_22720,N_21783,N_21973);
or U22721 (N_22721,N_21892,N_20802);
or U22722 (N_22722,N_21285,N_20668);
and U22723 (N_22723,N_21099,N_21963);
or U22724 (N_22724,N_20481,N_21629);
nand U22725 (N_22725,N_20247,N_20633);
or U22726 (N_22726,N_21009,N_20266);
nand U22727 (N_22727,N_21927,N_21636);
xor U22728 (N_22728,N_20746,N_20745);
or U22729 (N_22729,N_21899,N_20388);
nor U22730 (N_22730,N_20831,N_20960);
or U22731 (N_22731,N_20073,N_20861);
and U22732 (N_22732,N_20026,N_21018);
and U22733 (N_22733,N_20097,N_20397);
and U22734 (N_22734,N_21241,N_20770);
and U22735 (N_22735,N_21008,N_21775);
nor U22736 (N_22736,N_20534,N_21833);
and U22737 (N_22737,N_20351,N_20320);
or U22738 (N_22738,N_20281,N_20995);
xnor U22739 (N_22739,N_21007,N_21953);
or U22740 (N_22740,N_21784,N_20957);
or U22741 (N_22741,N_20724,N_21741);
or U22742 (N_22742,N_21822,N_21912);
xnor U22743 (N_22743,N_21655,N_20212);
nor U22744 (N_22744,N_20974,N_21011);
or U22745 (N_22745,N_20062,N_21130);
xor U22746 (N_22746,N_20346,N_21410);
nand U22747 (N_22747,N_21269,N_20201);
nand U22748 (N_22748,N_20286,N_20335);
and U22749 (N_22749,N_20444,N_20485);
xor U22750 (N_22750,N_21610,N_20493);
or U22751 (N_22751,N_21759,N_21705);
xnor U22752 (N_22752,N_21188,N_21847);
or U22753 (N_22753,N_20255,N_20800);
and U22754 (N_22754,N_20260,N_20279);
or U22755 (N_22755,N_21836,N_20853);
or U22756 (N_22756,N_20543,N_21700);
or U22757 (N_22757,N_20769,N_20863);
xnor U22758 (N_22758,N_21387,N_20105);
nor U22759 (N_22759,N_20330,N_20785);
nor U22760 (N_22760,N_20373,N_20881);
nor U22761 (N_22761,N_20673,N_21904);
xor U22762 (N_22762,N_20677,N_20103);
xnor U22763 (N_22763,N_20254,N_20671);
and U22764 (N_22764,N_20848,N_20654);
or U22765 (N_22765,N_21374,N_20934);
xnor U22766 (N_22766,N_21916,N_21945);
nor U22767 (N_22767,N_20341,N_20133);
nor U22768 (N_22768,N_20066,N_20653);
nand U22769 (N_22769,N_20815,N_21372);
and U22770 (N_22770,N_20349,N_21818);
nand U22771 (N_22771,N_21615,N_21010);
and U22772 (N_22772,N_20322,N_20965);
xor U22773 (N_22773,N_20219,N_20128);
nor U22774 (N_22774,N_21036,N_20494);
nand U22775 (N_22775,N_20270,N_21381);
nor U22776 (N_22776,N_20862,N_21141);
nand U22777 (N_22777,N_20348,N_20328);
or U22778 (N_22778,N_21652,N_21584);
or U22779 (N_22779,N_21524,N_20786);
nor U22780 (N_22780,N_20920,N_21825);
xor U22781 (N_22781,N_20684,N_20149);
xor U22782 (N_22782,N_20932,N_20807);
and U22783 (N_22783,N_21438,N_21347);
xor U22784 (N_22784,N_20375,N_20687);
nor U22785 (N_22785,N_20825,N_21861);
nand U22786 (N_22786,N_20418,N_20454);
and U22787 (N_22787,N_20344,N_21197);
xor U22788 (N_22788,N_21552,N_20376);
nor U22789 (N_22789,N_20194,N_21874);
xnor U22790 (N_22790,N_21952,N_21642);
nor U22791 (N_22791,N_20295,N_21788);
xnor U22792 (N_22792,N_21517,N_20903);
nand U22793 (N_22793,N_21909,N_20189);
nor U22794 (N_22794,N_21686,N_21276);
xor U22795 (N_22795,N_21247,N_20269);
or U22796 (N_22796,N_21990,N_21337);
nand U22797 (N_22797,N_20840,N_20856);
and U22798 (N_22798,N_20698,N_20192);
xnor U22799 (N_22799,N_20497,N_20489);
nor U22800 (N_22800,N_21431,N_21918);
nand U22801 (N_22801,N_20340,N_20275);
nand U22802 (N_22802,N_21691,N_20314);
nand U22803 (N_22803,N_20068,N_21096);
nand U22804 (N_22804,N_21205,N_20947);
nor U22805 (N_22805,N_20170,N_21395);
and U22806 (N_22806,N_21530,N_20294);
xnor U22807 (N_22807,N_21877,N_21806);
nand U22808 (N_22808,N_20705,N_20928);
or U22809 (N_22809,N_21163,N_20506);
nand U22810 (N_22810,N_20570,N_20262);
and U22811 (N_22811,N_20338,N_20252);
nor U22812 (N_22812,N_21595,N_20582);
nand U22813 (N_22813,N_20907,N_21158);
xor U22814 (N_22814,N_21484,N_20652);
xnor U22815 (N_22815,N_21367,N_20636);
xnor U22816 (N_22816,N_21232,N_21949);
and U22817 (N_22817,N_21365,N_20914);
or U22818 (N_22818,N_21712,N_20079);
nor U22819 (N_22819,N_20939,N_20025);
or U22820 (N_22820,N_21648,N_21363);
or U22821 (N_22821,N_20125,N_20525);
nand U22822 (N_22822,N_21512,N_21098);
nor U22823 (N_22823,N_21128,N_20648);
xnor U22824 (N_22824,N_21037,N_21716);
nor U22825 (N_22825,N_20540,N_21322);
nor U22826 (N_22826,N_21985,N_20154);
or U22827 (N_22827,N_21746,N_20644);
or U22828 (N_22828,N_21254,N_21443);
or U22829 (N_22829,N_20845,N_21670);
nor U22830 (N_22830,N_21668,N_20515);
xnor U22831 (N_22831,N_21683,N_20538);
or U22832 (N_22832,N_21361,N_20250);
and U22833 (N_22833,N_20530,N_20393);
xor U22834 (N_22834,N_21059,N_20919);
and U22835 (N_22835,N_20723,N_20238);
nor U22836 (N_22836,N_21161,N_20316);
xnor U22837 (N_22837,N_21545,N_20604);
nand U22838 (N_22838,N_20970,N_20626);
xor U22839 (N_22839,N_21181,N_21458);
and U22840 (N_22840,N_20287,N_21178);
or U22841 (N_22841,N_20622,N_21643);
xor U22842 (N_22842,N_20077,N_21433);
nor U22843 (N_22843,N_20579,N_21852);
xor U22844 (N_22844,N_21941,N_20985);
nor U22845 (N_22845,N_20136,N_21507);
xor U22846 (N_22846,N_21538,N_21771);
xnor U22847 (N_22847,N_21510,N_21907);
nand U22848 (N_22848,N_21238,N_20788);
and U22849 (N_22849,N_20526,N_20954);
and U22850 (N_22850,N_21191,N_20596);
nand U22851 (N_22851,N_21800,N_21585);
or U22852 (N_22852,N_20210,N_20398);
nor U22853 (N_22853,N_21911,N_21747);
nand U22854 (N_22854,N_20548,N_21562);
and U22855 (N_22855,N_20909,N_20087);
or U22856 (N_22856,N_21988,N_20357);
or U22857 (N_22857,N_20027,N_21672);
nor U22858 (N_22858,N_21398,N_21896);
nor U22859 (N_22859,N_20473,N_21793);
nor U22860 (N_22860,N_20709,N_20115);
nand U22861 (N_22861,N_21366,N_20211);
nor U22862 (N_22862,N_21690,N_20150);
or U22863 (N_22863,N_21732,N_21722);
and U22864 (N_22864,N_20551,N_20801);
xor U22865 (N_22865,N_21547,N_21138);
nand U22866 (N_22866,N_21289,N_20868);
and U22867 (N_22867,N_20600,N_21809);
nor U22868 (N_22868,N_20895,N_20585);
and U22869 (N_22869,N_21681,N_21749);
nand U22870 (N_22870,N_20809,N_20756);
xnor U22871 (N_22871,N_20475,N_21079);
nand U22872 (N_22872,N_21786,N_21863);
and U22873 (N_22873,N_20578,N_20977);
nand U22874 (N_22874,N_21511,N_21635);
and U22875 (N_22875,N_20466,N_20234);
and U22876 (N_22876,N_20924,N_21978);
nor U22877 (N_22877,N_20614,N_21049);
and U22878 (N_22878,N_21281,N_20071);
and U22879 (N_22879,N_21332,N_20095);
nor U22880 (N_22880,N_21206,N_20710);
xor U22881 (N_22881,N_20804,N_21490);
or U22882 (N_22882,N_21713,N_20118);
xnor U22883 (N_22883,N_20682,N_20658);
nor U22884 (N_22884,N_21373,N_21058);
nor U22885 (N_22885,N_20949,N_20593);
or U22886 (N_22886,N_20014,N_21857);
or U22887 (N_22887,N_20847,N_20717);
nand U22888 (N_22888,N_20502,N_21557);
xnor U22889 (N_22889,N_21597,N_20669);
nand U22890 (N_22890,N_20535,N_21804);
and U22891 (N_22891,N_20912,N_21823);
or U22892 (N_22892,N_21396,N_20446);
nand U22893 (N_22893,N_20860,N_21323);
nand U22894 (N_22894,N_20775,N_20765);
or U22895 (N_22895,N_21572,N_21565);
nor U22896 (N_22896,N_20647,N_20206);
nand U22897 (N_22897,N_20460,N_21121);
and U22898 (N_22898,N_21502,N_21485);
and U22899 (N_22899,N_21448,N_20146);
xnor U22900 (N_22900,N_20020,N_20753);
nand U22901 (N_22901,N_20527,N_21664);
nor U22902 (N_22902,N_20905,N_21653);
or U22903 (N_22903,N_20968,N_21382);
nor U22904 (N_22904,N_21755,N_21710);
nor U22905 (N_22905,N_20163,N_21570);
nand U22906 (N_22906,N_20450,N_20605);
or U22907 (N_22907,N_21457,N_21799);
and U22908 (N_22908,N_20428,N_21377);
or U22909 (N_22909,N_21951,N_20583);
and U22910 (N_22910,N_21040,N_20380);
nor U22911 (N_22911,N_20222,N_20774);
and U22912 (N_22912,N_21122,N_20035);
nand U22913 (N_22913,N_20866,N_21437);
nand U22914 (N_22914,N_20257,N_21073);
or U22915 (N_22915,N_20923,N_20245);
and U22916 (N_22916,N_20986,N_21295);
and U22917 (N_22917,N_20161,N_21190);
nor U22918 (N_22918,N_20955,N_20683);
nor U22919 (N_22919,N_21834,N_21967);
or U22920 (N_22920,N_21991,N_20042);
nand U22921 (N_22921,N_20158,N_21078);
xor U22922 (N_22922,N_21177,N_20751);
nor U22923 (N_22923,N_20844,N_20518);
nand U22924 (N_22924,N_20175,N_20839);
nor U22925 (N_22925,N_21393,N_20688);
nor U22926 (N_22926,N_21148,N_21291);
nor U22927 (N_22927,N_21754,N_20258);
nor U22928 (N_22928,N_20303,N_20625);
xor U22929 (N_22929,N_21521,N_20226);
xor U22930 (N_22930,N_21887,N_21176);
nor U22931 (N_22931,N_20477,N_21072);
and U22932 (N_22932,N_20449,N_21067);
nand U22933 (N_22933,N_21776,N_20272);
nand U22934 (N_22934,N_20039,N_21408);
nand U22935 (N_22935,N_20350,N_20697);
xnor U22936 (N_22936,N_21302,N_21645);
xor U22937 (N_22937,N_21107,N_21969);
xor U22938 (N_22938,N_21124,N_20911);
nor U22939 (N_22939,N_21891,N_20202);
nor U22940 (N_22940,N_20059,N_21660);
nand U22941 (N_22941,N_21240,N_21327);
nor U22942 (N_22942,N_20598,N_21126);
nand U22943 (N_22943,N_20869,N_21692);
nor U22944 (N_22944,N_20461,N_21364);
xor U22945 (N_22945,N_21465,N_20978);
and U22946 (N_22946,N_20129,N_20256);
xnor U22947 (N_22947,N_21266,N_20162);
and U22948 (N_22948,N_20114,N_20933);
or U22949 (N_22949,N_20739,N_20224);
or U22950 (N_22950,N_21220,N_20675);
or U22951 (N_22951,N_21061,N_20703);
nor U22952 (N_22952,N_20172,N_21189);
nand U22953 (N_22953,N_20824,N_21556);
nand U22954 (N_22954,N_21388,N_20727);
xor U22955 (N_22955,N_20276,N_20513);
nand U22956 (N_22956,N_21729,N_20553);
or U22957 (N_22957,N_20533,N_21872);
nor U22958 (N_22958,N_21150,N_21974);
nand U22959 (N_22959,N_21069,N_20124);
xor U22960 (N_22960,N_20736,N_20080);
nor U22961 (N_22961,N_20456,N_21522);
nand U22962 (N_22962,N_21411,N_20400);
xnor U22963 (N_22963,N_21986,N_21541);
xnor U22964 (N_22964,N_21824,N_21087);
xor U22965 (N_22965,N_20135,N_21342);
nor U22966 (N_22966,N_21308,N_20018);
and U22967 (N_22967,N_20382,N_20457);
nor U22968 (N_22968,N_21925,N_21895);
or U22969 (N_22969,N_20650,N_21186);
or U22970 (N_22970,N_21742,N_20733);
xor U22971 (N_22971,N_21622,N_20789);
or U22972 (N_22972,N_20186,N_21325);
xor U22973 (N_22973,N_20712,N_20334);
xor U22974 (N_22974,N_21262,N_20285);
and U22975 (N_22975,N_21537,N_21349);
or U22976 (N_22976,N_21298,N_21805);
nor U22977 (N_22977,N_21497,N_21283);
and U22978 (N_22978,N_20011,N_21334);
nor U22979 (N_22979,N_20304,N_20830);
nor U22980 (N_22980,N_21581,N_21544);
or U22981 (N_22981,N_21964,N_20412);
and U22982 (N_22982,N_21172,N_20983);
nor U22983 (N_22983,N_20897,N_21734);
and U22984 (N_22984,N_20876,N_20550);
xor U22985 (N_22985,N_20242,N_21519);
and U22986 (N_22986,N_20416,N_21526);
or U22987 (N_22987,N_21048,N_20339);
or U22988 (N_22988,N_21551,N_20343);
and U22989 (N_22989,N_21183,N_21104);
nand U22990 (N_22990,N_20870,N_20431);
nand U22991 (N_22991,N_20764,N_21649);
nand U22992 (N_22992,N_21739,N_21548);
and U22993 (N_22993,N_20640,N_20887);
nand U22994 (N_22994,N_20070,N_20471);
or U22995 (N_22995,N_20352,N_21698);
nor U22996 (N_22996,N_20386,N_20999);
nor U22997 (N_22997,N_21080,N_20387);
nand U22998 (N_22998,N_20798,N_20836);
or U22999 (N_22999,N_21210,N_21838);
or U23000 (N_23000,N_21515,N_20130);
and U23001 (N_23001,N_20341,N_21875);
xor U23002 (N_23002,N_21890,N_21272);
nor U23003 (N_23003,N_21980,N_20696);
nand U23004 (N_23004,N_21923,N_21398);
nor U23005 (N_23005,N_21052,N_20947);
and U23006 (N_23006,N_21787,N_20097);
and U23007 (N_23007,N_20206,N_21622);
or U23008 (N_23008,N_21906,N_20605);
or U23009 (N_23009,N_21359,N_21404);
and U23010 (N_23010,N_20314,N_20939);
and U23011 (N_23011,N_21706,N_21464);
xnor U23012 (N_23012,N_21761,N_20369);
or U23013 (N_23013,N_20016,N_20336);
nand U23014 (N_23014,N_20286,N_20592);
nor U23015 (N_23015,N_20073,N_21165);
xor U23016 (N_23016,N_20165,N_21341);
or U23017 (N_23017,N_21681,N_21501);
and U23018 (N_23018,N_21217,N_20834);
nand U23019 (N_23019,N_21817,N_21913);
and U23020 (N_23020,N_21497,N_20667);
xor U23021 (N_23021,N_21008,N_21127);
xnor U23022 (N_23022,N_20251,N_21837);
nor U23023 (N_23023,N_20695,N_21950);
xnor U23024 (N_23024,N_20318,N_20798);
or U23025 (N_23025,N_21768,N_20846);
nor U23026 (N_23026,N_20992,N_21719);
nor U23027 (N_23027,N_20520,N_21535);
or U23028 (N_23028,N_21152,N_20747);
and U23029 (N_23029,N_21439,N_21846);
nand U23030 (N_23030,N_20410,N_21160);
or U23031 (N_23031,N_21997,N_20262);
or U23032 (N_23032,N_21682,N_21165);
nor U23033 (N_23033,N_20588,N_20405);
xnor U23034 (N_23034,N_20739,N_21593);
or U23035 (N_23035,N_21014,N_20232);
or U23036 (N_23036,N_21142,N_21612);
or U23037 (N_23037,N_20597,N_21131);
nand U23038 (N_23038,N_20886,N_21603);
and U23039 (N_23039,N_21228,N_20878);
and U23040 (N_23040,N_20494,N_20160);
or U23041 (N_23041,N_20512,N_21521);
xnor U23042 (N_23042,N_21236,N_21695);
nand U23043 (N_23043,N_20444,N_20339);
nand U23044 (N_23044,N_20151,N_21507);
xnor U23045 (N_23045,N_21297,N_21805);
or U23046 (N_23046,N_20974,N_21816);
or U23047 (N_23047,N_20418,N_21579);
or U23048 (N_23048,N_20264,N_21708);
nand U23049 (N_23049,N_21816,N_21037);
nor U23050 (N_23050,N_20418,N_21891);
and U23051 (N_23051,N_20260,N_20224);
and U23052 (N_23052,N_21035,N_20919);
or U23053 (N_23053,N_20219,N_20568);
nand U23054 (N_23054,N_20052,N_21002);
xor U23055 (N_23055,N_21058,N_21053);
xor U23056 (N_23056,N_20573,N_21682);
nand U23057 (N_23057,N_21181,N_21733);
nand U23058 (N_23058,N_21356,N_21518);
xor U23059 (N_23059,N_20022,N_20740);
nor U23060 (N_23060,N_20475,N_21364);
or U23061 (N_23061,N_20944,N_21288);
xnor U23062 (N_23062,N_20182,N_20487);
nand U23063 (N_23063,N_20660,N_20237);
and U23064 (N_23064,N_21659,N_20169);
and U23065 (N_23065,N_21267,N_21053);
or U23066 (N_23066,N_21333,N_21634);
xnor U23067 (N_23067,N_20581,N_20215);
nand U23068 (N_23068,N_20508,N_20813);
or U23069 (N_23069,N_20918,N_20687);
xor U23070 (N_23070,N_20213,N_20809);
nand U23071 (N_23071,N_20878,N_21385);
and U23072 (N_23072,N_21720,N_21643);
and U23073 (N_23073,N_20112,N_20435);
and U23074 (N_23074,N_21115,N_20851);
or U23075 (N_23075,N_20217,N_21155);
or U23076 (N_23076,N_20958,N_20451);
and U23077 (N_23077,N_20588,N_21575);
and U23078 (N_23078,N_21296,N_20957);
xnor U23079 (N_23079,N_20393,N_20582);
or U23080 (N_23080,N_21553,N_21238);
nor U23081 (N_23081,N_20075,N_21820);
or U23082 (N_23082,N_20285,N_20939);
and U23083 (N_23083,N_21992,N_20265);
nor U23084 (N_23084,N_21933,N_20401);
xnor U23085 (N_23085,N_21479,N_21270);
nand U23086 (N_23086,N_21440,N_21127);
and U23087 (N_23087,N_21061,N_21316);
or U23088 (N_23088,N_20708,N_20226);
and U23089 (N_23089,N_20260,N_21357);
nand U23090 (N_23090,N_21469,N_21968);
and U23091 (N_23091,N_21006,N_21828);
xor U23092 (N_23092,N_21759,N_21546);
or U23093 (N_23093,N_21303,N_21889);
xnor U23094 (N_23094,N_21956,N_20109);
or U23095 (N_23095,N_21092,N_21269);
nand U23096 (N_23096,N_20293,N_20959);
nand U23097 (N_23097,N_20890,N_20023);
xor U23098 (N_23098,N_21785,N_21846);
or U23099 (N_23099,N_20375,N_20016);
xor U23100 (N_23100,N_21190,N_20685);
or U23101 (N_23101,N_20430,N_20188);
nor U23102 (N_23102,N_20958,N_21409);
nor U23103 (N_23103,N_20448,N_20644);
nor U23104 (N_23104,N_20911,N_21406);
nor U23105 (N_23105,N_20118,N_21007);
nor U23106 (N_23106,N_20873,N_20923);
and U23107 (N_23107,N_21539,N_21591);
and U23108 (N_23108,N_21463,N_21575);
nor U23109 (N_23109,N_20108,N_21113);
nand U23110 (N_23110,N_21944,N_20799);
or U23111 (N_23111,N_21947,N_20527);
or U23112 (N_23112,N_20488,N_20507);
and U23113 (N_23113,N_21459,N_21693);
and U23114 (N_23114,N_21388,N_20835);
xnor U23115 (N_23115,N_21801,N_20257);
and U23116 (N_23116,N_20446,N_21084);
xnor U23117 (N_23117,N_20841,N_21692);
and U23118 (N_23118,N_21434,N_21622);
nor U23119 (N_23119,N_20795,N_20630);
xnor U23120 (N_23120,N_20070,N_20268);
nor U23121 (N_23121,N_20058,N_21520);
nand U23122 (N_23122,N_21639,N_21299);
or U23123 (N_23123,N_21639,N_20858);
xor U23124 (N_23124,N_20028,N_21084);
xnor U23125 (N_23125,N_20566,N_20923);
or U23126 (N_23126,N_21645,N_20802);
or U23127 (N_23127,N_21983,N_21066);
and U23128 (N_23128,N_20774,N_21349);
or U23129 (N_23129,N_20787,N_21907);
nand U23130 (N_23130,N_20199,N_21230);
xor U23131 (N_23131,N_21052,N_21915);
xor U23132 (N_23132,N_20882,N_21309);
xnor U23133 (N_23133,N_21411,N_21603);
or U23134 (N_23134,N_21765,N_21505);
nor U23135 (N_23135,N_20597,N_20932);
and U23136 (N_23136,N_20120,N_21373);
or U23137 (N_23137,N_21581,N_20838);
and U23138 (N_23138,N_21525,N_20486);
and U23139 (N_23139,N_20097,N_21518);
nand U23140 (N_23140,N_21657,N_21819);
nand U23141 (N_23141,N_20626,N_20813);
and U23142 (N_23142,N_20797,N_21133);
nand U23143 (N_23143,N_21712,N_21398);
or U23144 (N_23144,N_21433,N_20779);
nor U23145 (N_23145,N_21077,N_20163);
and U23146 (N_23146,N_20737,N_20822);
nand U23147 (N_23147,N_20169,N_21947);
nand U23148 (N_23148,N_21064,N_21579);
xor U23149 (N_23149,N_21123,N_21917);
or U23150 (N_23150,N_21012,N_21940);
xor U23151 (N_23151,N_20905,N_21207);
xor U23152 (N_23152,N_20141,N_21903);
xor U23153 (N_23153,N_21142,N_20290);
or U23154 (N_23154,N_20217,N_21717);
xnor U23155 (N_23155,N_21914,N_20329);
or U23156 (N_23156,N_21673,N_21636);
xor U23157 (N_23157,N_20567,N_20873);
or U23158 (N_23158,N_20696,N_20749);
nor U23159 (N_23159,N_21583,N_21256);
nand U23160 (N_23160,N_21568,N_20593);
nand U23161 (N_23161,N_20254,N_21011);
xor U23162 (N_23162,N_21539,N_20099);
xor U23163 (N_23163,N_21433,N_20458);
nand U23164 (N_23164,N_21520,N_21831);
nor U23165 (N_23165,N_21705,N_21963);
and U23166 (N_23166,N_20075,N_21811);
nor U23167 (N_23167,N_20423,N_20963);
xnor U23168 (N_23168,N_21865,N_21464);
and U23169 (N_23169,N_21620,N_21177);
nand U23170 (N_23170,N_20480,N_21142);
nand U23171 (N_23171,N_20830,N_21806);
nand U23172 (N_23172,N_20110,N_21432);
nand U23173 (N_23173,N_21629,N_20024);
xnor U23174 (N_23174,N_20606,N_20642);
xor U23175 (N_23175,N_20301,N_20371);
nor U23176 (N_23176,N_20541,N_21330);
nor U23177 (N_23177,N_20775,N_21296);
or U23178 (N_23178,N_20267,N_21445);
nor U23179 (N_23179,N_20453,N_21380);
nand U23180 (N_23180,N_21014,N_20196);
and U23181 (N_23181,N_20315,N_20423);
xnor U23182 (N_23182,N_21824,N_21628);
nor U23183 (N_23183,N_20093,N_20370);
or U23184 (N_23184,N_21316,N_20279);
nor U23185 (N_23185,N_21352,N_21703);
or U23186 (N_23186,N_20958,N_21958);
and U23187 (N_23187,N_21197,N_20991);
and U23188 (N_23188,N_20095,N_20360);
or U23189 (N_23189,N_20235,N_20997);
and U23190 (N_23190,N_21820,N_21671);
xor U23191 (N_23191,N_20774,N_20739);
nor U23192 (N_23192,N_21773,N_21532);
and U23193 (N_23193,N_21067,N_21650);
nand U23194 (N_23194,N_20884,N_20284);
xnor U23195 (N_23195,N_21610,N_21551);
or U23196 (N_23196,N_20825,N_21619);
and U23197 (N_23197,N_20786,N_21076);
nor U23198 (N_23198,N_21039,N_20079);
or U23199 (N_23199,N_21139,N_20374);
xnor U23200 (N_23200,N_21939,N_20639);
nand U23201 (N_23201,N_21232,N_21532);
and U23202 (N_23202,N_21006,N_20282);
nand U23203 (N_23203,N_21861,N_20393);
nand U23204 (N_23204,N_20464,N_21471);
or U23205 (N_23205,N_20474,N_20902);
nand U23206 (N_23206,N_20054,N_20059);
xnor U23207 (N_23207,N_21706,N_20505);
and U23208 (N_23208,N_20506,N_20692);
xnor U23209 (N_23209,N_21831,N_20453);
xor U23210 (N_23210,N_20242,N_21690);
xor U23211 (N_23211,N_21464,N_20303);
nor U23212 (N_23212,N_21086,N_20247);
nor U23213 (N_23213,N_20333,N_20869);
or U23214 (N_23214,N_21028,N_20394);
nor U23215 (N_23215,N_20208,N_20372);
and U23216 (N_23216,N_21574,N_20797);
or U23217 (N_23217,N_20837,N_21573);
nand U23218 (N_23218,N_21161,N_21090);
or U23219 (N_23219,N_20612,N_20953);
nor U23220 (N_23220,N_21615,N_21339);
and U23221 (N_23221,N_20074,N_21389);
xor U23222 (N_23222,N_21981,N_20335);
and U23223 (N_23223,N_20180,N_21912);
xnor U23224 (N_23224,N_20593,N_20626);
nor U23225 (N_23225,N_21808,N_21315);
xnor U23226 (N_23226,N_20820,N_21876);
nor U23227 (N_23227,N_21183,N_21379);
nor U23228 (N_23228,N_21166,N_21869);
or U23229 (N_23229,N_20630,N_21774);
and U23230 (N_23230,N_21538,N_20177);
xor U23231 (N_23231,N_20058,N_20127);
nor U23232 (N_23232,N_21454,N_20203);
nand U23233 (N_23233,N_20780,N_20996);
xor U23234 (N_23234,N_21818,N_21799);
nor U23235 (N_23235,N_20216,N_20255);
nor U23236 (N_23236,N_21855,N_20910);
and U23237 (N_23237,N_21347,N_21714);
xor U23238 (N_23238,N_21109,N_20851);
and U23239 (N_23239,N_20565,N_20146);
and U23240 (N_23240,N_21711,N_20885);
xnor U23241 (N_23241,N_20427,N_20528);
nor U23242 (N_23242,N_20111,N_21922);
nand U23243 (N_23243,N_20244,N_21143);
nand U23244 (N_23244,N_21292,N_21495);
xor U23245 (N_23245,N_20289,N_20183);
or U23246 (N_23246,N_20277,N_20546);
and U23247 (N_23247,N_20576,N_20935);
or U23248 (N_23248,N_21361,N_21962);
nand U23249 (N_23249,N_21967,N_21566);
nand U23250 (N_23250,N_21548,N_20355);
xor U23251 (N_23251,N_20232,N_21343);
nor U23252 (N_23252,N_21146,N_21636);
and U23253 (N_23253,N_21682,N_21875);
and U23254 (N_23254,N_21646,N_20833);
xnor U23255 (N_23255,N_21237,N_20704);
nand U23256 (N_23256,N_21015,N_20078);
nand U23257 (N_23257,N_21970,N_21750);
nor U23258 (N_23258,N_20917,N_21472);
nand U23259 (N_23259,N_21873,N_21397);
or U23260 (N_23260,N_20057,N_21672);
nand U23261 (N_23261,N_21332,N_20044);
nor U23262 (N_23262,N_20524,N_21518);
and U23263 (N_23263,N_21633,N_21147);
nor U23264 (N_23264,N_20134,N_20058);
nand U23265 (N_23265,N_20527,N_21723);
xnor U23266 (N_23266,N_21183,N_20161);
nor U23267 (N_23267,N_20514,N_21076);
or U23268 (N_23268,N_21285,N_21043);
nand U23269 (N_23269,N_20384,N_21357);
nand U23270 (N_23270,N_21289,N_20542);
nand U23271 (N_23271,N_20795,N_20782);
xor U23272 (N_23272,N_21977,N_20010);
nand U23273 (N_23273,N_21501,N_21199);
nand U23274 (N_23274,N_20444,N_20598);
xor U23275 (N_23275,N_20872,N_20911);
nor U23276 (N_23276,N_20764,N_20760);
xnor U23277 (N_23277,N_21189,N_20171);
nand U23278 (N_23278,N_21246,N_21857);
nand U23279 (N_23279,N_20632,N_21115);
xnor U23280 (N_23280,N_20475,N_20077);
nand U23281 (N_23281,N_21307,N_21921);
nor U23282 (N_23282,N_21975,N_20368);
nor U23283 (N_23283,N_20867,N_20388);
or U23284 (N_23284,N_21181,N_20029);
nand U23285 (N_23285,N_20943,N_20034);
xnor U23286 (N_23286,N_20477,N_20385);
nor U23287 (N_23287,N_20060,N_20850);
and U23288 (N_23288,N_21906,N_21533);
or U23289 (N_23289,N_20960,N_20206);
xor U23290 (N_23290,N_21705,N_21348);
and U23291 (N_23291,N_20887,N_21090);
nand U23292 (N_23292,N_20248,N_21535);
nor U23293 (N_23293,N_20559,N_20896);
nand U23294 (N_23294,N_20599,N_21188);
and U23295 (N_23295,N_20880,N_20005);
xnor U23296 (N_23296,N_20674,N_20288);
nand U23297 (N_23297,N_21294,N_21300);
nand U23298 (N_23298,N_21238,N_21532);
nor U23299 (N_23299,N_21937,N_21303);
or U23300 (N_23300,N_21601,N_21714);
xnor U23301 (N_23301,N_20924,N_21603);
and U23302 (N_23302,N_20352,N_21638);
or U23303 (N_23303,N_21639,N_21068);
xor U23304 (N_23304,N_20127,N_20650);
nor U23305 (N_23305,N_21887,N_21789);
and U23306 (N_23306,N_20815,N_21672);
nor U23307 (N_23307,N_21951,N_21591);
and U23308 (N_23308,N_21877,N_21953);
nor U23309 (N_23309,N_20267,N_20786);
nor U23310 (N_23310,N_20203,N_21330);
nor U23311 (N_23311,N_20967,N_20199);
xor U23312 (N_23312,N_21568,N_21461);
or U23313 (N_23313,N_21774,N_21048);
xor U23314 (N_23314,N_21769,N_20985);
or U23315 (N_23315,N_20586,N_21051);
nand U23316 (N_23316,N_20377,N_21911);
xor U23317 (N_23317,N_21065,N_21613);
nor U23318 (N_23318,N_20329,N_21417);
or U23319 (N_23319,N_21581,N_21942);
nand U23320 (N_23320,N_21734,N_20528);
or U23321 (N_23321,N_20485,N_20541);
nand U23322 (N_23322,N_20201,N_20574);
xor U23323 (N_23323,N_20689,N_21839);
or U23324 (N_23324,N_20353,N_20141);
or U23325 (N_23325,N_21037,N_21138);
nor U23326 (N_23326,N_20032,N_20622);
xnor U23327 (N_23327,N_20281,N_20116);
nand U23328 (N_23328,N_21669,N_21883);
and U23329 (N_23329,N_21349,N_20646);
xor U23330 (N_23330,N_20466,N_21347);
xor U23331 (N_23331,N_21062,N_20678);
nand U23332 (N_23332,N_21523,N_20644);
nand U23333 (N_23333,N_20807,N_20850);
or U23334 (N_23334,N_20962,N_20274);
nand U23335 (N_23335,N_21451,N_20230);
nor U23336 (N_23336,N_21267,N_21358);
and U23337 (N_23337,N_21605,N_21703);
xnor U23338 (N_23338,N_20775,N_21450);
nor U23339 (N_23339,N_20974,N_21413);
nor U23340 (N_23340,N_21647,N_21612);
xor U23341 (N_23341,N_21736,N_21352);
and U23342 (N_23342,N_20346,N_20568);
nor U23343 (N_23343,N_21152,N_21154);
and U23344 (N_23344,N_20838,N_21700);
nor U23345 (N_23345,N_20532,N_20251);
nor U23346 (N_23346,N_21296,N_20562);
nand U23347 (N_23347,N_21732,N_21255);
nor U23348 (N_23348,N_20712,N_20677);
nand U23349 (N_23349,N_20754,N_21124);
nor U23350 (N_23350,N_21343,N_20366);
xnor U23351 (N_23351,N_20972,N_20886);
and U23352 (N_23352,N_20576,N_21814);
or U23353 (N_23353,N_20267,N_20256);
nand U23354 (N_23354,N_20808,N_21069);
or U23355 (N_23355,N_20818,N_21070);
and U23356 (N_23356,N_20889,N_20258);
xor U23357 (N_23357,N_20246,N_20458);
nand U23358 (N_23358,N_21640,N_20168);
nor U23359 (N_23359,N_21189,N_20497);
xor U23360 (N_23360,N_21734,N_20495);
nor U23361 (N_23361,N_21937,N_21139);
and U23362 (N_23362,N_20327,N_20013);
or U23363 (N_23363,N_21269,N_20115);
nor U23364 (N_23364,N_21608,N_20221);
and U23365 (N_23365,N_21546,N_20325);
and U23366 (N_23366,N_21085,N_21778);
or U23367 (N_23367,N_20264,N_20048);
nand U23368 (N_23368,N_20166,N_21550);
xor U23369 (N_23369,N_20782,N_20619);
xor U23370 (N_23370,N_20793,N_21353);
and U23371 (N_23371,N_20152,N_20432);
nand U23372 (N_23372,N_21399,N_20407);
xor U23373 (N_23373,N_21808,N_20877);
or U23374 (N_23374,N_21709,N_20739);
and U23375 (N_23375,N_20785,N_21012);
nand U23376 (N_23376,N_21925,N_21410);
and U23377 (N_23377,N_21903,N_20865);
or U23378 (N_23378,N_21338,N_21819);
xor U23379 (N_23379,N_21539,N_20285);
nor U23380 (N_23380,N_21317,N_20377);
and U23381 (N_23381,N_20382,N_20613);
and U23382 (N_23382,N_20660,N_21179);
nor U23383 (N_23383,N_21177,N_20190);
nor U23384 (N_23384,N_21874,N_21953);
or U23385 (N_23385,N_20113,N_21742);
nor U23386 (N_23386,N_21826,N_21151);
or U23387 (N_23387,N_21015,N_20340);
nand U23388 (N_23388,N_20926,N_20798);
nand U23389 (N_23389,N_21469,N_21912);
nor U23390 (N_23390,N_20553,N_21595);
nor U23391 (N_23391,N_21233,N_21476);
and U23392 (N_23392,N_20045,N_21481);
or U23393 (N_23393,N_21086,N_20925);
nand U23394 (N_23394,N_21828,N_21415);
nor U23395 (N_23395,N_20713,N_21200);
nand U23396 (N_23396,N_20404,N_21674);
nand U23397 (N_23397,N_21373,N_21513);
nand U23398 (N_23398,N_21251,N_21727);
nand U23399 (N_23399,N_21121,N_20529);
xnor U23400 (N_23400,N_21651,N_21984);
nand U23401 (N_23401,N_20105,N_21609);
nand U23402 (N_23402,N_20798,N_20908);
nand U23403 (N_23403,N_20542,N_20459);
nand U23404 (N_23404,N_20155,N_20262);
nor U23405 (N_23405,N_21696,N_21204);
nand U23406 (N_23406,N_20095,N_20105);
or U23407 (N_23407,N_21637,N_20427);
nand U23408 (N_23408,N_21850,N_21636);
nand U23409 (N_23409,N_21977,N_21723);
and U23410 (N_23410,N_20589,N_21299);
nor U23411 (N_23411,N_21971,N_21068);
nor U23412 (N_23412,N_20190,N_21790);
nand U23413 (N_23413,N_20125,N_21136);
nor U23414 (N_23414,N_20582,N_21291);
nand U23415 (N_23415,N_21879,N_20562);
or U23416 (N_23416,N_21367,N_20179);
xor U23417 (N_23417,N_21487,N_21077);
xor U23418 (N_23418,N_20588,N_20497);
nand U23419 (N_23419,N_21107,N_21730);
and U23420 (N_23420,N_20485,N_21757);
or U23421 (N_23421,N_21191,N_20931);
xor U23422 (N_23422,N_21810,N_20338);
nor U23423 (N_23423,N_21366,N_20818);
nand U23424 (N_23424,N_20356,N_20128);
and U23425 (N_23425,N_20315,N_20992);
or U23426 (N_23426,N_21647,N_21560);
nor U23427 (N_23427,N_21498,N_20321);
or U23428 (N_23428,N_21782,N_21981);
and U23429 (N_23429,N_20130,N_20293);
nor U23430 (N_23430,N_21757,N_20343);
nor U23431 (N_23431,N_21828,N_21611);
nor U23432 (N_23432,N_21646,N_21283);
and U23433 (N_23433,N_21723,N_21228);
nor U23434 (N_23434,N_20796,N_20076);
xnor U23435 (N_23435,N_21177,N_21173);
nand U23436 (N_23436,N_21114,N_21430);
xor U23437 (N_23437,N_20994,N_21468);
nand U23438 (N_23438,N_21176,N_20573);
or U23439 (N_23439,N_20436,N_20550);
and U23440 (N_23440,N_20026,N_20231);
and U23441 (N_23441,N_20851,N_20241);
nand U23442 (N_23442,N_20103,N_21127);
xor U23443 (N_23443,N_20421,N_20008);
and U23444 (N_23444,N_21038,N_21544);
nor U23445 (N_23445,N_21968,N_20369);
nor U23446 (N_23446,N_21941,N_21805);
nand U23447 (N_23447,N_20616,N_21836);
xor U23448 (N_23448,N_21964,N_20008);
nor U23449 (N_23449,N_20255,N_20521);
and U23450 (N_23450,N_21638,N_20027);
and U23451 (N_23451,N_20196,N_21287);
and U23452 (N_23452,N_20872,N_21352);
xor U23453 (N_23453,N_20650,N_20629);
and U23454 (N_23454,N_21995,N_20046);
and U23455 (N_23455,N_20206,N_20798);
nand U23456 (N_23456,N_21299,N_20162);
nand U23457 (N_23457,N_21353,N_21988);
and U23458 (N_23458,N_21810,N_21174);
nand U23459 (N_23459,N_20391,N_20394);
and U23460 (N_23460,N_21876,N_20492);
and U23461 (N_23461,N_20531,N_20117);
nand U23462 (N_23462,N_21385,N_21668);
xnor U23463 (N_23463,N_20892,N_21920);
xnor U23464 (N_23464,N_20029,N_20098);
xnor U23465 (N_23465,N_20127,N_20093);
and U23466 (N_23466,N_21629,N_20876);
or U23467 (N_23467,N_21392,N_20005);
xor U23468 (N_23468,N_20855,N_21076);
nor U23469 (N_23469,N_20019,N_20058);
nand U23470 (N_23470,N_20323,N_20874);
nor U23471 (N_23471,N_20531,N_20716);
or U23472 (N_23472,N_20900,N_21111);
nand U23473 (N_23473,N_20734,N_21754);
and U23474 (N_23474,N_21847,N_20819);
xnor U23475 (N_23475,N_20756,N_21846);
and U23476 (N_23476,N_21334,N_21298);
or U23477 (N_23477,N_20759,N_20726);
or U23478 (N_23478,N_21157,N_20686);
nand U23479 (N_23479,N_21383,N_21574);
and U23480 (N_23480,N_21535,N_20722);
xor U23481 (N_23481,N_21899,N_20715);
nor U23482 (N_23482,N_21245,N_21362);
nor U23483 (N_23483,N_20423,N_21234);
or U23484 (N_23484,N_20983,N_21220);
xor U23485 (N_23485,N_21537,N_20529);
xnor U23486 (N_23486,N_21463,N_21666);
nand U23487 (N_23487,N_21179,N_20292);
nor U23488 (N_23488,N_21373,N_20100);
and U23489 (N_23489,N_21168,N_21343);
nor U23490 (N_23490,N_21723,N_20394);
nand U23491 (N_23491,N_20766,N_21021);
and U23492 (N_23492,N_21807,N_20822);
or U23493 (N_23493,N_20273,N_20874);
xor U23494 (N_23494,N_21058,N_21366);
nor U23495 (N_23495,N_20921,N_20093);
and U23496 (N_23496,N_20513,N_21630);
or U23497 (N_23497,N_21191,N_20849);
nor U23498 (N_23498,N_21011,N_21838);
xor U23499 (N_23499,N_20147,N_20707);
or U23500 (N_23500,N_21118,N_20561);
nor U23501 (N_23501,N_21741,N_20673);
or U23502 (N_23502,N_20843,N_21433);
nor U23503 (N_23503,N_21714,N_21563);
nor U23504 (N_23504,N_20280,N_21949);
nor U23505 (N_23505,N_20819,N_21027);
or U23506 (N_23506,N_20215,N_21656);
and U23507 (N_23507,N_20299,N_20167);
and U23508 (N_23508,N_21070,N_21454);
nand U23509 (N_23509,N_21623,N_21539);
nand U23510 (N_23510,N_21753,N_21154);
nand U23511 (N_23511,N_21888,N_20099);
xor U23512 (N_23512,N_21496,N_21351);
nor U23513 (N_23513,N_20192,N_20789);
nand U23514 (N_23514,N_21492,N_21190);
xnor U23515 (N_23515,N_20561,N_21433);
and U23516 (N_23516,N_20625,N_20001);
or U23517 (N_23517,N_21978,N_20122);
nor U23518 (N_23518,N_20147,N_20018);
xor U23519 (N_23519,N_20463,N_21780);
or U23520 (N_23520,N_20472,N_21229);
and U23521 (N_23521,N_20701,N_21697);
nor U23522 (N_23522,N_21608,N_21253);
nor U23523 (N_23523,N_20416,N_21152);
nand U23524 (N_23524,N_20653,N_20412);
nand U23525 (N_23525,N_20801,N_21402);
xor U23526 (N_23526,N_21220,N_20086);
nor U23527 (N_23527,N_20338,N_20565);
nor U23528 (N_23528,N_20122,N_20766);
nor U23529 (N_23529,N_20786,N_20401);
nand U23530 (N_23530,N_21564,N_21650);
nand U23531 (N_23531,N_20504,N_21950);
nor U23532 (N_23532,N_21237,N_21674);
or U23533 (N_23533,N_20155,N_20757);
xor U23534 (N_23534,N_20767,N_21543);
nand U23535 (N_23535,N_20356,N_21637);
nand U23536 (N_23536,N_20600,N_21978);
xnor U23537 (N_23537,N_21972,N_21669);
and U23538 (N_23538,N_20414,N_20832);
nand U23539 (N_23539,N_20389,N_21313);
or U23540 (N_23540,N_21286,N_21988);
nand U23541 (N_23541,N_21694,N_21096);
nand U23542 (N_23542,N_21273,N_21929);
and U23543 (N_23543,N_20788,N_21398);
or U23544 (N_23544,N_20686,N_20014);
nand U23545 (N_23545,N_20184,N_20936);
nor U23546 (N_23546,N_20776,N_21363);
and U23547 (N_23547,N_20217,N_20853);
and U23548 (N_23548,N_21470,N_20493);
and U23549 (N_23549,N_21112,N_21057);
nor U23550 (N_23550,N_20252,N_20642);
or U23551 (N_23551,N_20093,N_20069);
xor U23552 (N_23552,N_21731,N_20106);
or U23553 (N_23553,N_20566,N_21168);
and U23554 (N_23554,N_21520,N_20214);
and U23555 (N_23555,N_20844,N_21130);
or U23556 (N_23556,N_21752,N_21017);
or U23557 (N_23557,N_21864,N_21747);
xnor U23558 (N_23558,N_21049,N_20648);
xor U23559 (N_23559,N_21740,N_21143);
and U23560 (N_23560,N_20114,N_20662);
xor U23561 (N_23561,N_20510,N_20935);
nor U23562 (N_23562,N_21805,N_20256);
xor U23563 (N_23563,N_21738,N_20614);
and U23564 (N_23564,N_20939,N_20555);
or U23565 (N_23565,N_21961,N_20476);
or U23566 (N_23566,N_20924,N_21024);
nor U23567 (N_23567,N_21697,N_21373);
or U23568 (N_23568,N_21957,N_21993);
or U23569 (N_23569,N_20533,N_21366);
nand U23570 (N_23570,N_20865,N_21643);
or U23571 (N_23571,N_21128,N_21438);
nor U23572 (N_23572,N_20229,N_21585);
or U23573 (N_23573,N_20683,N_20420);
or U23574 (N_23574,N_20210,N_21522);
nor U23575 (N_23575,N_21593,N_21743);
or U23576 (N_23576,N_20889,N_21695);
or U23577 (N_23577,N_20005,N_21335);
xnor U23578 (N_23578,N_20189,N_20770);
nor U23579 (N_23579,N_21331,N_21412);
and U23580 (N_23580,N_21318,N_21725);
xor U23581 (N_23581,N_20545,N_20846);
xnor U23582 (N_23582,N_21501,N_20198);
nor U23583 (N_23583,N_20768,N_20737);
and U23584 (N_23584,N_20640,N_20881);
and U23585 (N_23585,N_21321,N_20961);
and U23586 (N_23586,N_20899,N_20598);
or U23587 (N_23587,N_21566,N_20973);
xor U23588 (N_23588,N_21033,N_20114);
nand U23589 (N_23589,N_21327,N_20135);
nand U23590 (N_23590,N_21802,N_20649);
or U23591 (N_23591,N_20693,N_20899);
or U23592 (N_23592,N_20595,N_20046);
nor U23593 (N_23593,N_21548,N_21337);
xnor U23594 (N_23594,N_20504,N_21680);
or U23595 (N_23595,N_20912,N_20556);
nor U23596 (N_23596,N_21878,N_20821);
xor U23597 (N_23597,N_20663,N_21657);
xor U23598 (N_23598,N_21716,N_20575);
xor U23599 (N_23599,N_20496,N_20052);
and U23600 (N_23600,N_21568,N_20046);
nor U23601 (N_23601,N_20205,N_21886);
nor U23602 (N_23602,N_21433,N_21892);
xnor U23603 (N_23603,N_21671,N_20734);
nand U23604 (N_23604,N_20800,N_20500);
xor U23605 (N_23605,N_21364,N_21285);
nand U23606 (N_23606,N_21899,N_21916);
or U23607 (N_23607,N_21504,N_21053);
nor U23608 (N_23608,N_21513,N_21969);
xor U23609 (N_23609,N_20626,N_21809);
and U23610 (N_23610,N_20844,N_20041);
and U23611 (N_23611,N_20890,N_20972);
and U23612 (N_23612,N_20337,N_20088);
nor U23613 (N_23613,N_21206,N_20412);
and U23614 (N_23614,N_21384,N_21295);
xor U23615 (N_23615,N_20929,N_21563);
xor U23616 (N_23616,N_20407,N_21686);
nand U23617 (N_23617,N_21279,N_20770);
nor U23618 (N_23618,N_20477,N_20711);
or U23619 (N_23619,N_20448,N_20875);
nor U23620 (N_23620,N_20579,N_20429);
and U23621 (N_23621,N_21056,N_21569);
nand U23622 (N_23622,N_21912,N_21859);
nor U23623 (N_23623,N_20699,N_21757);
nor U23624 (N_23624,N_20383,N_21021);
nand U23625 (N_23625,N_20647,N_20524);
nor U23626 (N_23626,N_21369,N_20114);
nand U23627 (N_23627,N_20956,N_21843);
xor U23628 (N_23628,N_21673,N_21005);
nor U23629 (N_23629,N_20566,N_21813);
and U23630 (N_23630,N_20855,N_21570);
and U23631 (N_23631,N_20639,N_21742);
and U23632 (N_23632,N_21732,N_21499);
xnor U23633 (N_23633,N_20425,N_20073);
nand U23634 (N_23634,N_21740,N_20704);
or U23635 (N_23635,N_21097,N_21991);
nand U23636 (N_23636,N_21194,N_20615);
nor U23637 (N_23637,N_21724,N_20000);
and U23638 (N_23638,N_21216,N_20171);
or U23639 (N_23639,N_20995,N_20703);
nand U23640 (N_23640,N_20916,N_20185);
and U23641 (N_23641,N_20472,N_21033);
nand U23642 (N_23642,N_20250,N_20594);
nand U23643 (N_23643,N_20422,N_20072);
xor U23644 (N_23644,N_21143,N_21253);
nor U23645 (N_23645,N_21812,N_20589);
nor U23646 (N_23646,N_20817,N_21788);
or U23647 (N_23647,N_21842,N_21227);
xor U23648 (N_23648,N_21671,N_21579);
nand U23649 (N_23649,N_21891,N_21512);
xor U23650 (N_23650,N_20115,N_20387);
nand U23651 (N_23651,N_20542,N_21129);
and U23652 (N_23652,N_20108,N_21834);
xor U23653 (N_23653,N_20160,N_21563);
nor U23654 (N_23654,N_21615,N_20430);
nor U23655 (N_23655,N_21319,N_20058);
nor U23656 (N_23656,N_21871,N_21511);
and U23657 (N_23657,N_21288,N_20048);
xor U23658 (N_23658,N_20404,N_20646);
or U23659 (N_23659,N_20303,N_20393);
or U23660 (N_23660,N_21646,N_20042);
or U23661 (N_23661,N_20603,N_20310);
and U23662 (N_23662,N_21062,N_20420);
nand U23663 (N_23663,N_21079,N_21601);
nand U23664 (N_23664,N_20605,N_20377);
nand U23665 (N_23665,N_20021,N_20793);
or U23666 (N_23666,N_21536,N_21442);
nor U23667 (N_23667,N_21792,N_21808);
nor U23668 (N_23668,N_20078,N_21410);
or U23669 (N_23669,N_21890,N_20718);
xor U23670 (N_23670,N_20852,N_20571);
and U23671 (N_23671,N_21239,N_20413);
or U23672 (N_23672,N_21653,N_21904);
nor U23673 (N_23673,N_20704,N_20849);
nand U23674 (N_23674,N_21912,N_21397);
and U23675 (N_23675,N_20757,N_20003);
xnor U23676 (N_23676,N_21471,N_20823);
and U23677 (N_23677,N_21009,N_20752);
or U23678 (N_23678,N_21782,N_20444);
nand U23679 (N_23679,N_21394,N_21854);
and U23680 (N_23680,N_21331,N_20623);
and U23681 (N_23681,N_21623,N_20901);
and U23682 (N_23682,N_20721,N_21193);
nand U23683 (N_23683,N_21442,N_20774);
xnor U23684 (N_23684,N_21757,N_20946);
or U23685 (N_23685,N_21174,N_21036);
xnor U23686 (N_23686,N_20605,N_20237);
xnor U23687 (N_23687,N_20324,N_21324);
xor U23688 (N_23688,N_21526,N_21936);
or U23689 (N_23689,N_20031,N_21645);
nor U23690 (N_23690,N_20111,N_21854);
and U23691 (N_23691,N_20238,N_20550);
nor U23692 (N_23692,N_20530,N_21912);
nand U23693 (N_23693,N_20335,N_20304);
nor U23694 (N_23694,N_21191,N_21034);
nor U23695 (N_23695,N_20327,N_21144);
and U23696 (N_23696,N_21541,N_21427);
and U23697 (N_23697,N_20667,N_21160);
or U23698 (N_23698,N_20844,N_21473);
xnor U23699 (N_23699,N_21853,N_21687);
or U23700 (N_23700,N_21366,N_21614);
nor U23701 (N_23701,N_21564,N_20513);
nand U23702 (N_23702,N_21595,N_20708);
or U23703 (N_23703,N_20259,N_21447);
and U23704 (N_23704,N_20780,N_21791);
or U23705 (N_23705,N_20394,N_20067);
or U23706 (N_23706,N_21057,N_20217);
and U23707 (N_23707,N_20907,N_20750);
or U23708 (N_23708,N_21709,N_20586);
nand U23709 (N_23709,N_20630,N_20613);
and U23710 (N_23710,N_20606,N_20940);
nand U23711 (N_23711,N_20446,N_20498);
xnor U23712 (N_23712,N_21234,N_20977);
nand U23713 (N_23713,N_20339,N_20796);
xnor U23714 (N_23714,N_21212,N_20678);
and U23715 (N_23715,N_21806,N_20894);
and U23716 (N_23716,N_21898,N_21298);
xnor U23717 (N_23717,N_20333,N_21829);
nor U23718 (N_23718,N_21844,N_21986);
nor U23719 (N_23719,N_20388,N_20401);
or U23720 (N_23720,N_20950,N_21367);
and U23721 (N_23721,N_20985,N_20580);
xor U23722 (N_23722,N_21661,N_21564);
xor U23723 (N_23723,N_21342,N_20117);
nand U23724 (N_23724,N_21020,N_20754);
or U23725 (N_23725,N_20310,N_21925);
nor U23726 (N_23726,N_21943,N_21793);
and U23727 (N_23727,N_21424,N_20230);
nand U23728 (N_23728,N_20932,N_21029);
or U23729 (N_23729,N_21907,N_21501);
or U23730 (N_23730,N_20529,N_21999);
xor U23731 (N_23731,N_21812,N_20540);
and U23732 (N_23732,N_21044,N_20141);
nor U23733 (N_23733,N_20603,N_20347);
and U23734 (N_23734,N_20099,N_21133);
nand U23735 (N_23735,N_21266,N_20099);
or U23736 (N_23736,N_20090,N_20301);
or U23737 (N_23737,N_21085,N_20996);
nand U23738 (N_23738,N_20461,N_21564);
and U23739 (N_23739,N_20202,N_20179);
or U23740 (N_23740,N_20346,N_21385);
xnor U23741 (N_23741,N_20784,N_21717);
nand U23742 (N_23742,N_20438,N_20837);
and U23743 (N_23743,N_20218,N_21177);
xnor U23744 (N_23744,N_20617,N_21769);
nor U23745 (N_23745,N_20162,N_21965);
nand U23746 (N_23746,N_21979,N_21718);
and U23747 (N_23747,N_21077,N_21725);
nand U23748 (N_23748,N_20990,N_21429);
nor U23749 (N_23749,N_20903,N_20982);
nand U23750 (N_23750,N_20905,N_21483);
nand U23751 (N_23751,N_21814,N_21204);
xnor U23752 (N_23752,N_21580,N_20833);
or U23753 (N_23753,N_21724,N_21376);
and U23754 (N_23754,N_20398,N_21491);
nand U23755 (N_23755,N_20160,N_20367);
and U23756 (N_23756,N_21261,N_20924);
nor U23757 (N_23757,N_20793,N_20121);
nor U23758 (N_23758,N_21763,N_20723);
or U23759 (N_23759,N_20069,N_21467);
xnor U23760 (N_23760,N_20613,N_21393);
nand U23761 (N_23761,N_20635,N_21349);
nand U23762 (N_23762,N_21400,N_21398);
nor U23763 (N_23763,N_20686,N_21072);
nor U23764 (N_23764,N_20821,N_20011);
or U23765 (N_23765,N_20379,N_21981);
nor U23766 (N_23766,N_21830,N_20999);
nor U23767 (N_23767,N_21556,N_20038);
and U23768 (N_23768,N_21351,N_20623);
and U23769 (N_23769,N_20986,N_21065);
and U23770 (N_23770,N_20513,N_21632);
xor U23771 (N_23771,N_20025,N_20644);
xor U23772 (N_23772,N_20520,N_20278);
xor U23773 (N_23773,N_21331,N_20828);
or U23774 (N_23774,N_20610,N_21474);
nor U23775 (N_23775,N_20437,N_20661);
or U23776 (N_23776,N_21848,N_20421);
and U23777 (N_23777,N_21549,N_21506);
nand U23778 (N_23778,N_21350,N_21433);
or U23779 (N_23779,N_20309,N_20690);
nor U23780 (N_23780,N_20156,N_21732);
and U23781 (N_23781,N_21161,N_21590);
nand U23782 (N_23782,N_21262,N_20693);
xnor U23783 (N_23783,N_20298,N_20223);
and U23784 (N_23784,N_21361,N_21103);
nand U23785 (N_23785,N_21113,N_20173);
and U23786 (N_23786,N_21259,N_20161);
or U23787 (N_23787,N_21085,N_20489);
and U23788 (N_23788,N_21900,N_20396);
nand U23789 (N_23789,N_20985,N_21824);
and U23790 (N_23790,N_20551,N_21626);
xnor U23791 (N_23791,N_21789,N_20715);
or U23792 (N_23792,N_21733,N_20277);
nand U23793 (N_23793,N_21619,N_21053);
and U23794 (N_23794,N_20240,N_21623);
or U23795 (N_23795,N_21284,N_20065);
and U23796 (N_23796,N_20683,N_21823);
and U23797 (N_23797,N_20359,N_20120);
nor U23798 (N_23798,N_21577,N_21712);
and U23799 (N_23799,N_21245,N_20387);
or U23800 (N_23800,N_21753,N_20106);
and U23801 (N_23801,N_20283,N_20099);
and U23802 (N_23802,N_21099,N_21948);
or U23803 (N_23803,N_21265,N_21019);
xnor U23804 (N_23804,N_20289,N_21946);
and U23805 (N_23805,N_20969,N_21854);
and U23806 (N_23806,N_20537,N_21154);
xor U23807 (N_23807,N_20349,N_21187);
and U23808 (N_23808,N_21411,N_21890);
xnor U23809 (N_23809,N_21345,N_20889);
or U23810 (N_23810,N_21834,N_21495);
and U23811 (N_23811,N_21739,N_20973);
or U23812 (N_23812,N_20002,N_20437);
xnor U23813 (N_23813,N_21250,N_21435);
and U23814 (N_23814,N_21496,N_21780);
nand U23815 (N_23815,N_20924,N_20647);
xor U23816 (N_23816,N_21254,N_20310);
and U23817 (N_23817,N_21044,N_21787);
nand U23818 (N_23818,N_21426,N_20459);
or U23819 (N_23819,N_20372,N_20192);
and U23820 (N_23820,N_20578,N_20756);
nor U23821 (N_23821,N_21891,N_20026);
nand U23822 (N_23822,N_20518,N_21703);
nand U23823 (N_23823,N_20050,N_20708);
nand U23824 (N_23824,N_21950,N_20088);
nor U23825 (N_23825,N_20159,N_21911);
xnor U23826 (N_23826,N_20684,N_21376);
xnor U23827 (N_23827,N_21068,N_20624);
nand U23828 (N_23828,N_21522,N_20637);
and U23829 (N_23829,N_20304,N_20298);
nand U23830 (N_23830,N_21850,N_21611);
nand U23831 (N_23831,N_20207,N_20567);
xor U23832 (N_23832,N_21358,N_20473);
nand U23833 (N_23833,N_20644,N_20299);
or U23834 (N_23834,N_20483,N_20708);
nand U23835 (N_23835,N_21637,N_20267);
or U23836 (N_23836,N_20344,N_20932);
and U23837 (N_23837,N_20085,N_20639);
xnor U23838 (N_23838,N_21006,N_21008);
and U23839 (N_23839,N_21439,N_21634);
or U23840 (N_23840,N_21438,N_21921);
nor U23841 (N_23841,N_21908,N_21567);
or U23842 (N_23842,N_20238,N_20968);
nand U23843 (N_23843,N_20260,N_21629);
and U23844 (N_23844,N_21955,N_20806);
xnor U23845 (N_23845,N_20896,N_20536);
nor U23846 (N_23846,N_20096,N_21199);
nor U23847 (N_23847,N_21155,N_20887);
nand U23848 (N_23848,N_20948,N_20017);
xor U23849 (N_23849,N_21456,N_21994);
nand U23850 (N_23850,N_21178,N_20405);
or U23851 (N_23851,N_20460,N_21882);
and U23852 (N_23852,N_21718,N_20221);
nor U23853 (N_23853,N_21833,N_21113);
and U23854 (N_23854,N_20483,N_20703);
nor U23855 (N_23855,N_20771,N_20499);
xnor U23856 (N_23856,N_21723,N_20448);
nor U23857 (N_23857,N_21842,N_20156);
nand U23858 (N_23858,N_21647,N_21566);
and U23859 (N_23859,N_20111,N_21977);
nor U23860 (N_23860,N_20976,N_20008);
and U23861 (N_23861,N_21166,N_20949);
xor U23862 (N_23862,N_21849,N_20783);
nand U23863 (N_23863,N_21919,N_20550);
nor U23864 (N_23864,N_21063,N_21672);
nor U23865 (N_23865,N_21567,N_21902);
and U23866 (N_23866,N_21701,N_21891);
nand U23867 (N_23867,N_21562,N_21851);
or U23868 (N_23868,N_20542,N_20286);
nor U23869 (N_23869,N_21110,N_20954);
xor U23870 (N_23870,N_20645,N_21116);
and U23871 (N_23871,N_21181,N_21573);
nor U23872 (N_23872,N_21624,N_21778);
nor U23873 (N_23873,N_21181,N_20762);
and U23874 (N_23874,N_20288,N_21244);
nand U23875 (N_23875,N_20962,N_21787);
and U23876 (N_23876,N_20356,N_21657);
and U23877 (N_23877,N_21918,N_21138);
nand U23878 (N_23878,N_21832,N_21017);
or U23879 (N_23879,N_21502,N_20670);
nand U23880 (N_23880,N_21844,N_20187);
nand U23881 (N_23881,N_20651,N_20634);
nor U23882 (N_23882,N_20437,N_21880);
or U23883 (N_23883,N_20158,N_21478);
or U23884 (N_23884,N_20298,N_20922);
nand U23885 (N_23885,N_20750,N_20685);
or U23886 (N_23886,N_21229,N_20263);
nand U23887 (N_23887,N_20637,N_21743);
or U23888 (N_23888,N_20762,N_21755);
xnor U23889 (N_23889,N_21258,N_21169);
nor U23890 (N_23890,N_20389,N_21344);
nor U23891 (N_23891,N_21464,N_21334);
or U23892 (N_23892,N_20146,N_20178);
and U23893 (N_23893,N_20475,N_21859);
nor U23894 (N_23894,N_20288,N_21639);
or U23895 (N_23895,N_20933,N_20364);
and U23896 (N_23896,N_21220,N_21228);
xnor U23897 (N_23897,N_20823,N_20016);
and U23898 (N_23898,N_20479,N_20108);
and U23899 (N_23899,N_20861,N_21095);
nor U23900 (N_23900,N_20461,N_20072);
and U23901 (N_23901,N_20368,N_20366);
nor U23902 (N_23902,N_20960,N_21226);
nor U23903 (N_23903,N_20396,N_20962);
nand U23904 (N_23904,N_20528,N_21471);
and U23905 (N_23905,N_21244,N_20637);
xnor U23906 (N_23906,N_20023,N_21410);
xor U23907 (N_23907,N_20657,N_20815);
and U23908 (N_23908,N_20287,N_21281);
xor U23909 (N_23909,N_20579,N_21736);
and U23910 (N_23910,N_20890,N_20668);
nor U23911 (N_23911,N_21897,N_20634);
nor U23912 (N_23912,N_20658,N_20960);
or U23913 (N_23913,N_21925,N_21030);
nor U23914 (N_23914,N_21657,N_20340);
nor U23915 (N_23915,N_20808,N_21792);
or U23916 (N_23916,N_21208,N_21715);
xor U23917 (N_23917,N_20903,N_20893);
nor U23918 (N_23918,N_21449,N_21907);
nor U23919 (N_23919,N_21923,N_21691);
xnor U23920 (N_23920,N_20373,N_20771);
xnor U23921 (N_23921,N_21578,N_21556);
nand U23922 (N_23922,N_21539,N_21627);
nor U23923 (N_23923,N_21984,N_20639);
and U23924 (N_23924,N_20428,N_21537);
and U23925 (N_23925,N_21734,N_20113);
nor U23926 (N_23926,N_20425,N_20699);
and U23927 (N_23927,N_20673,N_21161);
nand U23928 (N_23928,N_21116,N_20730);
xnor U23929 (N_23929,N_20976,N_20813);
nor U23930 (N_23930,N_20142,N_21639);
nand U23931 (N_23931,N_20782,N_21624);
xor U23932 (N_23932,N_21501,N_21723);
xnor U23933 (N_23933,N_21313,N_20523);
and U23934 (N_23934,N_21841,N_21700);
nor U23935 (N_23935,N_21383,N_20490);
or U23936 (N_23936,N_20672,N_20685);
nor U23937 (N_23937,N_21525,N_21242);
xor U23938 (N_23938,N_21039,N_20978);
nand U23939 (N_23939,N_20273,N_20654);
nor U23940 (N_23940,N_21403,N_20256);
or U23941 (N_23941,N_20652,N_21485);
or U23942 (N_23942,N_20580,N_21146);
xor U23943 (N_23943,N_21762,N_21842);
or U23944 (N_23944,N_21873,N_21235);
xnor U23945 (N_23945,N_21148,N_20068);
nor U23946 (N_23946,N_21642,N_20619);
nand U23947 (N_23947,N_21353,N_20487);
and U23948 (N_23948,N_21892,N_21053);
nor U23949 (N_23949,N_21577,N_20623);
or U23950 (N_23950,N_20831,N_20786);
nand U23951 (N_23951,N_20016,N_21023);
or U23952 (N_23952,N_20593,N_20209);
nor U23953 (N_23953,N_20425,N_20179);
xor U23954 (N_23954,N_21043,N_20244);
nand U23955 (N_23955,N_21740,N_20831);
or U23956 (N_23956,N_21262,N_21940);
xnor U23957 (N_23957,N_20927,N_21472);
nand U23958 (N_23958,N_20577,N_21829);
or U23959 (N_23959,N_20794,N_21637);
nand U23960 (N_23960,N_21866,N_20991);
xor U23961 (N_23961,N_21933,N_20846);
xor U23962 (N_23962,N_20451,N_20426);
or U23963 (N_23963,N_21420,N_21602);
or U23964 (N_23964,N_20183,N_20513);
and U23965 (N_23965,N_20985,N_21847);
or U23966 (N_23966,N_20187,N_20478);
xor U23967 (N_23967,N_21645,N_21174);
nor U23968 (N_23968,N_20545,N_21283);
nor U23969 (N_23969,N_21697,N_21832);
and U23970 (N_23970,N_21730,N_20865);
xnor U23971 (N_23971,N_20174,N_20937);
and U23972 (N_23972,N_20376,N_21649);
and U23973 (N_23973,N_21009,N_20497);
xnor U23974 (N_23974,N_20664,N_21591);
and U23975 (N_23975,N_20687,N_20936);
and U23976 (N_23976,N_21225,N_20055);
nand U23977 (N_23977,N_21073,N_21962);
xor U23978 (N_23978,N_20511,N_20372);
xor U23979 (N_23979,N_20218,N_20318);
and U23980 (N_23980,N_20318,N_21694);
or U23981 (N_23981,N_20557,N_20486);
and U23982 (N_23982,N_21968,N_20891);
or U23983 (N_23983,N_21332,N_20093);
and U23984 (N_23984,N_20177,N_20687);
nand U23985 (N_23985,N_21408,N_20694);
nand U23986 (N_23986,N_21169,N_20974);
nor U23987 (N_23987,N_20605,N_21190);
nand U23988 (N_23988,N_21397,N_20908);
or U23989 (N_23989,N_20645,N_20696);
and U23990 (N_23990,N_21048,N_21775);
nor U23991 (N_23991,N_21830,N_20551);
or U23992 (N_23992,N_20871,N_20221);
nor U23993 (N_23993,N_20765,N_21683);
xor U23994 (N_23994,N_21178,N_21294);
nand U23995 (N_23995,N_21861,N_21498);
and U23996 (N_23996,N_20614,N_20587);
nand U23997 (N_23997,N_20037,N_21101);
and U23998 (N_23998,N_20349,N_21958);
nor U23999 (N_23999,N_20489,N_20409);
and U24000 (N_24000,N_23040,N_23518);
nand U24001 (N_24001,N_22972,N_23768);
nor U24002 (N_24002,N_23407,N_22725);
nor U24003 (N_24003,N_22346,N_22527);
and U24004 (N_24004,N_23510,N_23900);
or U24005 (N_24005,N_23125,N_23868);
or U24006 (N_24006,N_23529,N_22571);
nand U24007 (N_24007,N_22007,N_22308);
nand U24008 (N_24008,N_22273,N_23841);
or U24009 (N_24009,N_23416,N_23382);
nor U24010 (N_24010,N_23808,N_23252);
nor U24011 (N_24011,N_22195,N_23314);
nand U24012 (N_24012,N_22604,N_22248);
nor U24013 (N_24013,N_22272,N_22577);
nor U24014 (N_24014,N_23780,N_23654);
nand U24015 (N_24015,N_23751,N_22403);
or U24016 (N_24016,N_22336,N_23219);
nand U24017 (N_24017,N_22239,N_22935);
and U24018 (N_24018,N_23195,N_22772);
or U24019 (N_24019,N_22024,N_23155);
nand U24020 (N_24020,N_23713,N_23482);
or U24021 (N_24021,N_22711,N_22379);
nor U24022 (N_24022,N_23607,N_22019);
nand U24023 (N_24023,N_23235,N_23610);
xor U24024 (N_24024,N_22461,N_23596);
xor U24025 (N_24025,N_22122,N_22191);
or U24026 (N_24026,N_23085,N_22745);
nor U24027 (N_24027,N_23759,N_23464);
and U24028 (N_24028,N_23495,N_22775);
and U24029 (N_24029,N_22919,N_22914);
nand U24030 (N_24030,N_23483,N_22697);
xnor U24031 (N_24031,N_23601,N_22161);
xnor U24032 (N_24032,N_22973,N_22488);
xor U24033 (N_24033,N_22959,N_22908);
xor U24034 (N_24034,N_22767,N_22332);
nor U24035 (N_24035,N_23383,N_23090);
nor U24036 (N_24036,N_22885,N_22438);
or U24037 (N_24037,N_23853,N_23658);
nor U24038 (N_24038,N_23123,N_23865);
and U24039 (N_24039,N_22344,N_23500);
xnor U24040 (N_24040,N_22647,N_23309);
nor U24041 (N_24041,N_22606,N_23203);
or U24042 (N_24042,N_23818,N_23288);
or U24043 (N_24043,N_22646,N_22171);
and U24044 (N_24044,N_23922,N_22644);
and U24045 (N_24045,N_22081,N_22815);
xnor U24046 (N_24046,N_22548,N_23968);
nor U24047 (N_24047,N_23746,N_23068);
nand U24048 (N_24048,N_22754,N_22302);
or U24049 (N_24049,N_22694,N_22559);
or U24050 (N_24050,N_22509,N_22102);
xnor U24051 (N_24051,N_22237,N_23530);
xnor U24052 (N_24052,N_23242,N_22074);
nand U24053 (N_24053,N_22006,N_22194);
nand U24054 (N_24054,N_22947,N_22041);
nor U24055 (N_24055,N_22924,N_22193);
or U24056 (N_24056,N_22693,N_22683);
xor U24057 (N_24057,N_22620,N_22200);
xnor U24058 (N_24058,N_22837,N_22002);
or U24059 (N_24059,N_22372,N_23754);
or U24060 (N_24060,N_22291,N_22627);
and U24061 (N_24061,N_23162,N_23709);
or U24062 (N_24062,N_23347,N_23115);
and U24063 (N_24063,N_23315,N_22840);
or U24064 (N_24064,N_23105,N_23840);
xor U24065 (N_24065,N_22219,N_22893);
nor U24066 (N_24066,N_23683,N_23250);
or U24067 (N_24067,N_22207,N_22317);
and U24068 (N_24068,N_22951,N_22199);
nand U24069 (N_24069,N_22343,N_23706);
and U24070 (N_24070,N_22406,N_22418);
nor U24071 (N_24071,N_23714,N_23629);
or U24072 (N_24072,N_23782,N_22182);
nor U24073 (N_24073,N_22010,N_22226);
nand U24074 (N_24074,N_22466,N_23216);
nand U24075 (N_24075,N_23613,N_22540);
or U24076 (N_24076,N_22516,N_23469);
nor U24077 (N_24077,N_23895,N_22067);
and U24078 (N_24078,N_23661,N_23704);
nand U24079 (N_24079,N_22026,N_23679);
nor U24080 (N_24080,N_22201,N_23667);
nand U24081 (N_24081,N_23797,N_23906);
and U24082 (N_24082,N_22414,N_22356);
xnor U24083 (N_24083,N_22011,N_22501);
and U24084 (N_24084,N_22432,N_22964);
or U24085 (N_24085,N_23997,N_22957);
nand U24086 (N_24086,N_22017,N_22515);
nand U24087 (N_24087,N_23108,N_22234);
xor U24088 (N_24088,N_22728,N_22898);
nor U24089 (N_24089,N_22902,N_23572);
and U24090 (N_24090,N_23860,N_22518);
and U24091 (N_24091,N_22471,N_23342);
nor U24092 (N_24092,N_23415,N_22855);
nand U24093 (N_24093,N_23817,N_23077);
nor U24094 (N_24094,N_23883,N_22611);
nand U24095 (N_24095,N_23862,N_23276);
nand U24096 (N_24096,N_23343,N_23816);
nand U24097 (N_24097,N_23657,N_23786);
and U24098 (N_24098,N_22814,N_22304);
and U24099 (N_24099,N_23515,N_23065);
nand U24100 (N_24100,N_23456,N_22044);
nor U24101 (N_24101,N_23303,N_22116);
or U24102 (N_24102,N_22971,N_23926);
xnor U24103 (N_24103,N_23376,N_23192);
nand U24104 (N_24104,N_23190,N_23512);
and U24105 (N_24105,N_23936,N_22290);
and U24106 (N_24106,N_23438,N_22580);
xor U24107 (N_24107,N_22835,N_23054);
or U24108 (N_24108,N_22779,N_23811);
xnor U24109 (N_24109,N_23005,N_22256);
nand U24110 (N_24110,N_23401,N_22963);
nor U24111 (N_24111,N_22351,N_23381);
and U24112 (N_24112,N_23659,N_22415);
or U24113 (N_24113,N_22663,N_22773);
and U24114 (N_24114,N_23581,N_23813);
nor U24115 (N_24115,N_22053,N_23573);
or U24116 (N_24116,N_22616,N_23268);
nand U24117 (N_24117,N_22051,N_23004);
nor U24118 (N_24118,N_23834,N_22544);
xnor U24119 (N_24119,N_22284,N_22057);
xnor U24120 (N_24120,N_22327,N_23032);
or U24121 (N_24121,N_23145,N_22097);
and U24122 (N_24122,N_22628,N_22532);
xnor U24123 (N_24123,N_22186,N_23437);
xnor U24124 (N_24124,N_23279,N_22521);
and U24125 (N_24125,N_23411,N_22489);
xnor U24126 (N_24126,N_22165,N_23442);
and U24127 (N_24127,N_22369,N_22016);
nand U24128 (N_24128,N_22178,N_23361);
and U24129 (N_24129,N_23474,N_22159);
nor U24130 (N_24130,N_22421,N_22319);
or U24131 (N_24131,N_23103,N_22672);
xnor U24132 (N_24132,N_23267,N_22679);
or U24133 (N_24133,N_22491,N_23019);
nand U24134 (N_24134,N_22744,N_22293);
and U24135 (N_24135,N_23978,N_22554);
xnor U24136 (N_24136,N_23789,N_23349);
nor U24137 (N_24137,N_23890,N_23599);
xnor U24138 (N_24138,N_23735,N_22404);
or U24139 (N_24139,N_22975,N_22792);
nor U24140 (N_24140,N_23119,N_22874);
or U24141 (N_24141,N_23534,N_22196);
or U24142 (N_24142,N_23428,N_22664);
xnor U24143 (N_24143,N_22829,N_23275);
nor U24144 (N_24144,N_22613,N_23163);
nand U24145 (N_24145,N_22798,N_22342);
nor U24146 (N_24146,N_23126,N_23549);
nand U24147 (N_24147,N_23838,N_23293);
nand U24148 (N_24148,N_22790,N_22760);
nand U24149 (N_24149,N_22315,N_23386);
xor U24150 (N_24150,N_22388,N_22054);
nor U24151 (N_24151,N_23101,N_22082);
or U24152 (N_24152,N_23388,N_22668);
nand U24153 (N_24153,N_23033,N_23864);
nor U24154 (N_24154,N_23340,N_22654);
xnor U24155 (N_24155,N_23762,N_22684);
or U24156 (N_24156,N_22891,N_23669);
and U24157 (N_24157,N_23387,N_23747);
and U24158 (N_24158,N_23334,N_23089);
and U24159 (N_24159,N_23966,N_23594);
or U24160 (N_24160,N_23357,N_22522);
nand U24161 (N_24161,N_22166,N_22989);
or U24162 (N_24162,N_23371,N_22791);
and U24163 (N_24163,N_22750,N_22113);
nand U24164 (N_24164,N_22650,N_23589);
nand U24165 (N_24165,N_23588,N_22497);
nand U24166 (N_24166,N_23311,N_22140);
or U24167 (N_24167,N_23419,N_22429);
xnor U24168 (N_24168,N_22478,N_22331);
nor U24169 (N_24169,N_23245,N_22405);
or U24170 (N_24170,N_22085,N_22579);
xnor U24171 (N_24171,N_23053,N_22083);
or U24172 (N_24172,N_23453,N_22637);
nand U24173 (N_24173,N_23225,N_22857);
xnor U24174 (N_24174,N_22175,N_22005);
and U24175 (N_24175,N_23877,N_23194);
and U24176 (N_24176,N_23994,N_22433);
xor U24177 (N_24177,N_22587,N_22378);
and U24178 (N_24178,N_23375,N_22764);
nand U24179 (N_24179,N_22762,N_23698);
nor U24180 (N_24180,N_22955,N_22995);
nand U24181 (N_24181,N_23896,N_22125);
nor U24182 (N_24182,N_22335,N_22546);
and U24183 (N_24183,N_23325,N_22228);
and U24184 (N_24184,N_22245,N_22223);
nor U24185 (N_24185,N_22513,N_22072);
nand U24186 (N_24186,N_22039,N_22842);
or U24187 (N_24187,N_23498,N_22090);
xor U24188 (N_24188,N_22581,N_22354);
xnor U24189 (N_24189,N_22632,N_22820);
xnor U24190 (N_24190,N_23804,N_23645);
nor U24191 (N_24191,N_23973,N_22279);
nand U24192 (N_24192,N_23923,N_22991);
nand U24193 (N_24193,N_23251,N_22472);
nor U24194 (N_24194,N_23409,N_23051);
xnor U24195 (N_24195,N_22148,N_23413);
nor U24196 (N_24196,N_22804,N_23634);
and U24197 (N_24197,N_23370,N_22160);
xnor U24198 (N_24198,N_23977,N_23043);
nand U24199 (N_24199,N_22986,N_22262);
and U24200 (N_24200,N_22813,N_22965);
or U24201 (N_24201,N_23950,N_22751);
nand U24202 (N_24202,N_22251,N_22980);
nor U24203 (N_24203,N_23176,N_23953);
nor U24204 (N_24204,N_22743,N_23335);
xor U24205 (N_24205,N_23322,N_23640);
or U24206 (N_24206,N_23346,N_22662);
nand U24207 (N_24207,N_23856,N_22797);
xnor U24208 (N_24208,N_22271,N_22455);
nand U24209 (N_24209,N_23134,N_23734);
and U24210 (N_24210,N_22312,N_23022);
or U24211 (N_24211,N_23561,N_23109);
or U24212 (N_24212,N_22733,N_23055);
or U24213 (N_24213,N_22392,N_23726);
xor U24214 (N_24214,N_22969,N_23814);
xnor U24215 (N_24215,N_22150,N_22887);
nor U24216 (N_24216,N_23256,N_23258);
nor U24217 (N_24217,N_23663,N_23839);
nand U24218 (N_24218,N_22238,N_23491);
xnor U24219 (N_24219,N_22706,N_22260);
nor U24220 (N_24220,N_23537,N_22297);
nor U24221 (N_24221,N_22961,N_22056);
xor U24222 (N_24222,N_22112,N_22221);
nand U24223 (N_24223,N_23480,N_22204);
or U24224 (N_24224,N_23399,N_23615);
nand U24225 (N_24225,N_22206,N_22707);
nand U24226 (N_24226,N_23405,N_22949);
and U24227 (N_24227,N_22872,N_22323);
xor U24228 (N_24228,N_22292,N_22867);
and U24229 (N_24229,N_23039,N_23948);
nand U24230 (N_24230,N_22249,N_23368);
nand U24231 (N_24231,N_23132,N_23971);
nor U24232 (N_24232,N_23234,N_23644);
xnor U24233 (N_24233,N_22321,N_23133);
xnor U24234 (N_24234,N_22956,N_23815);
and U24235 (N_24235,N_23011,N_23942);
nand U24236 (N_24236,N_22121,N_22446);
and U24237 (N_24237,N_22153,N_23550);
xor U24238 (N_24238,N_22263,N_22583);
or U24239 (N_24239,N_22233,N_22349);
and U24240 (N_24240,N_22731,N_22631);
nor U24241 (N_24241,N_22621,N_22003);
nor U24242 (N_24242,N_23410,N_22868);
or U24243 (N_24243,N_22734,N_23231);
and U24244 (N_24244,N_23801,N_22833);
and U24245 (N_24245,N_22427,N_23633);
nand U24246 (N_24246,N_22720,N_22622);
nor U24247 (N_24247,N_23869,N_23277);
or U24248 (N_24248,N_23114,N_23867);
nor U24249 (N_24249,N_22897,N_22328);
or U24250 (N_24250,N_22769,N_23048);
nand U24251 (N_24251,N_23214,N_23221);
and U24252 (N_24252,N_22596,N_23218);
xor U24253 (N_24253,N_23158,N_22269);
xnor U24254 (N_24254,N_22771,N_22094);
and U24255 (N_24255,N_22475,N_23426);
nand U24256 (N_24256,N_22859,N_22542);
and U24257 (N_24257,N_23450,N_22301);
xor U24258 (N_24258,N_23504,N_23957);
xnor U24259 (N_24259,N_22135,N_23676);
nand U24260 (N_24260,N_22713,N_22740);
and U24261 (N_24261,N_22496,N_23271);
xor U24262 (N_24262,N_22367,N_23847);
and U24263 (N_24263,N_23433,N_23299);
and U24264 (N_24264,N_22757,N_23982);
xnor U24265 (N_24265,N_22643,N_22450);
or U24266 (N_24266,N_23112,N_23648);
nor U24267 (N_24267,N_23725,N_23879);
xor U24268 (N_24268,N_23253,N_22091);
nor U24269 (N_24269,N_22069,N_23720);
nor U24270 (N_24270,N_23765,N_22242);
nand U24271 (N_24271,N_23297,N_23794);
or U24272 (N_24272,N_22374,N_22402);
xor U24273 (N_24273,N_22595,N_23229);
xor U24274 (N_24274,N_22377,N_23030);
nor U24275 (N_24275,N_23859,N_23931);
nor U24276 (N_24276,N_23855,N_23021);
or U24277 (N_24277,N_22574,N_23104);
or U24278 (N_24278,N_23429,N_22983);
nor U24279 (N_24279,N_23711,N_23736);
or U24280 (N_24280,N_22625,N_23833);
nand U24281 (N_24281,N_23603,N_23866);
nand U24282 (N_24282,N_23791,N_23649);
or U24283 (N_24283,N_23960,N_22275);
xor U24284 (N_24284,N_22104,N_23063);
nor U24285 (N_24285,N_23738,N_23673);
xnor U24286 (N_24286,N_22590,N_23631);
nand U24287 (N_24287,N_23542,N_22270);
nand U24288 (N_24288,N_23071,N_23237);
nand U24289 (N_24289,N_22029,N_23008);
and U24290 (N_24290,N_23001,N_22365);
and U24291 (N_24291,N_22950,N_23037);
xnor U24292 (N_24292,N_23580,N_22926);
and U24293 (N_24293,N_22954,N_23878);
nor U24294 (N_24294,N_23183,N_22584);
or U24295 (N_24295,N_22688,N_23702);
or U24296 (N_24296,N_23462,N_23093);
nor U24297 (N_24297,N_22464,N_23637);
nand U24298 (N_24298,N_22468,N_23436);
or U24299 (N_24299,N_22481,N_23511);
nand U24300 (N_24300,N_22451,N_23707);
nor U24301 (N_24301,N_23336,N_23617);
nand U24302 (N_24302,N_23223,N_22075);
and U24303 (N_24303,N_22442,N_22209);
nor U24304 (N_24304,N_23364,N_23752);
nand U24305 (N_24305,N_23424,N_22918);
nor U24306 (N_24306,N_23002,N_22401);
nor U24307 (N_24307,N_23298,N_22189);
xor U24308 (N_24308,N_22203,N_22084);
nor U24309 (N_24309,N_23352,N_23932);
and U24310 (N_24310,N_22676,N_23959);
xnor U24311 (N_24311,N_23576,N_23394);
nand U24312 (N_24312,N_22786,N_23901);
or U24313 (N_24313,N_23822,N_22979);
xnor U24314 (N_24314,N_23286,N_23087);
nand U24315 (N_24315,N_23171,N_23502);
or U24316 (N_24316,N_22132,N_23306);
nor U24317 (N_24317,N_22252,N_22932);
nor U24318 (N_24318,N_22370,N_23151);
nand U24319 (N_24319,N_23798,N_23668);
xor U24320 (N_24320,N_22059,N_22653);
xnor U24321 (N_24321,N_22462,N_22146);
and U24322 (N_24322,N_23898,N_23360);
and U24323 (N_24323,N_22014,N_23174);
nor U24324 (N_24324,N_22858,N_23993);
xor U24325 (N_24325,N_22738,N_22281);
nor U24326 (N_24326,N_23187,N_23984);
nor U24327 (N_24327,N_22708,N_22607);
nor U24328 (N_24328,N_23513,N_23458);
nor U24329 (N_24329,N_22880,N_22741);
nor U24330 (N_24330,N_23076,N_23911);
xnor U24331 (N_24331,N_22819,N_22463);
and U24332 (N_24332,N_23239,N_22753);
xnor U24333 (N_24333,N_23656,N_23208);
or U24334 (N_24334,N_23972,N_23069);
or U24335 (N_24335,N_23965,N_23543);
xor U24336 (N_24336,N_23608,N_22436);
and U24337 (N_24337,N_23992,N_23124);
and U24338 (N_24338,N_22023,N_22528);
nand U24339 (N_24339,N_22334,N_22088);
nand U24340 (N_24340,N_22660,N_22485);
xor U24341 (N_24341,N_22133,N_23312);
or U24342 (N_24342,N_22093,N_23672);
nor U24343 (N_24343,N_22670,N_23374);
nand U24344 (N_24344,N_23991,N_22967);
nor U24345 (N_24345,N_22529,N_22612);
nor U24346 (N_24346,N_22105,N_23585);
or U24347 (N_24347,N_22062,N_22977);
nor U24348 (N_24348,N_23447,N_22123);
and U24349 (N_24349,N_22360,N_23687);
nor U24350 (N_24350,N_23058,N_23116);
nor U24351 (N_24351,N_23820,N_23070);
nor U24352 (N_24352,N_23665,N_22131);
nand U24353 (N_24353,N_22705,N_23283);
and U24354 (N_24354,N_22371,N_23609);
and U24355 (N_24355,N_23691,N_23742);
or U24356 (N_24356,N_22847,N_22289);
xnor U24357 (N_24357,N_23240,N_22530);
or U24358 (N_24358,N_23333,N_22836);
xnor U24359 (N_24359,N_23539,N_23016);
nor U24360 (N_24360,N_22818,N_23630);
or U24361 (N_24361,N_23858,N_23185);
and U24362 (N_24362,N_23472,N_22115);
nor U24363 (N_24363,N_23421,N_23981);
and U24364 (N_24364,N_23044,N_22911);
xor U24365 (N_24365,N_23731,N_23372);
or U24366 (N_24366,N_23882,N_22288);
or U24367 (N_24367,N_22241,N_22445);
xor U24368 (N_24368,N_22338,N_22695);
xor U24369 (N_24369,N_23397,N_22185);
and U24370 (N_24370,N_22994,N_23274);
xnor U24371 (N_24371,N_22848,N_23113);
xnor U24372 (N_24372,N_22064,N_22395);
and U24373 (N_24373,N_22364,N_22357);
and U24374 (N_24374,N_23391,N_22812);
xor U24375 (N_24375,N_23695,N_22032);
nand U24376 (N_24376,N_22061,N_23567);
xor U24377 (N_24377,N_23418,N_23179);
nand U24378 (N_24378,N_22426,N_22156);
nand U24379 (N_24379,N_23307,N_22649);
nor U24380 (N_24380,N_22677,N_22494);
xor U24381 (N_24381,N_23488,N_22507);
xor U24382 (N_24382,N_22990,N_22626);
nor U24383 (N_24383,N_23310,N_23681);
xnor U24384 (N_24384,N_22564,N_23365);
nor U24385 (N_24385,N_22184,N_23781);
and U24386 (N_24386,N_22114,N_23167);
xor U24387 (N_24387,N_22400,N_22851);
nand U24388 (N_24388,N_23774,N_22118);
nor U24389 (N_24389,N_22430,N_23188);
and U24390 (N_24390,N_22366,N_23313);
nor U24391 (N_24391,N_23952,N_23487);
or U24392 (N_24392,N_23344,N_23524);
xnor U24393 (N_24393,N_23639,N_23578);
xor U24394 (N_24394,N_22444,N_23606);
xnor U24395 (N_24395,N_23412,N_22988);
and U24396 (N_24396,N_22952,N_22337);
nand U24397 (N_24397,N_22915,N_22782);
and U24398 (N_24398,N_23503,N_23763);
and U24399 (N_24399,N_23205,N_22800);
xnor U24400 (N_24400,N_23642,N_23122);
nand U24401 (N_24401,N_22520,N_23148);
and U24402 (N_24402,N_22645,N_22998);
nor U24403 (N_24403,N_23574,N_23517);
nor U24404 (N_24404,N_23975,N_22614);
or U24405 (N_24405,N_23930,N_23082);
nor U24406 (N_24406,N_23444,N_22422);
nor U24407 (N_24407,N_23803,N_23558);
xnor U24408 (N_24408,N_23583,N_22929);
xor U24409 (N_24409,N_23292,N_22698);
and U24410 (N_24410,N_23075,N_22941);
nor U24411 (N_24411,N_23540,N_23940);
nor U24412 (N_24412,N_23227,N_23670);
xor U24413 (N_24413,N_23913,N_22098);
and U24414 (N_24414,N_22050,N_23351);
and U24415 (N_24415,N_22139,N_23098);
nand U24416 (N_24416,N_22531,N_22048);
and U24417 (N_24417,N_22552,N_22087);
xor U24418 (N_24418,N_23771,N_22144);
xnor U24419 (N_24419,N_23131,N_23064);
nor U24420 (N_24420,N_23943,N_23243);
nand U24421 (N_24421,N_23775,N_22821);
and U24422 (N_24422,N_23590,N_23497);
and U24423 (N_24423,N_23121,N_23885);
xnor U24424 (N_24424,N_22300,N_23793);
and U24425 (N_24425,N_23743,N_23230);
or U24426 (N_24426,N_23323,N_22883);
and U24427 (N_24427,N_22686,N_22923);
or U24428 (N_24428,N_23262,N_22283);
and U24429 (N_24429,N_23341,N_22250);
nor U24430 (N_24430,N_22788,N_22899);
xor U24431 (N_24431,N_23538,N_22188);
nor U24432 (N_24432,N_23009,N_22657);
nand U24433 (N_24433,N_23431,N_23200);
or U24434 (N_24434,N_23592,N_23985);
nand U24435 (N_24435,N_22827,N_22177);
or U24436 (N_24436,N_22142,N_23699);
and U24437 (N_24437,N_22065,N_23408);
or U24438 (N_24438,N_23577,N_23137);
xor U24439 (N_24439,N_23915,N_22981);
xnor U24440 (N_24440,N_23727,N_22410);
and U24441 (N_24441,N_23827,N_22305);
nand U24442 (N_24442,N_23848,N_23554);
or U24443 (N_24443,N_23619,N_22117);
nor U24444 (N_24444,N_22276,N_22817);
and U24445 (N_24445,N_22440,N_23703);
nor U24446 (N_24446,N_22441,N_22294);
nand U24447 (N_24447,N_22794,N_22452);
nor U24448 (N_24448,N_23324,N_23000);
nor U24449 (N_24449,N_23479,N_23362);
nor U24450 (N_24450,N_22517,N_22839);
nor U24451 (N_24451,N_23976,N_22723);
and U24452 (N_24452,N_23983,N_23091);
and U24453 (N_24453,N_22424,N_22326);
nor U24454 (N_24454,N_22154,N_22149);
or U24455 (N_24455,N_22060,N_23805);
xnor U24456 (N_24456,N_23057,N_22038);
and U24457 (N_24457,N_23398,N_23423);
xor U24458 (N_24458,N_22770,N_23556);
and U24459 (N_24459,N_23184,N_22287);
nand U24460 (N_24460,N_23036,N_22667);
or U24461 (N_24461,N_23800,N_22576);
nand U24462 (N_24462,N_22691,N_23422);
nor U24463 (N_24463,N_23045,N_22480);
nor U24464 (N_24464,N_22838,N_22931);
nand U24465 (N_24465,N_23546,N_22563);
nand U24466 (N_24466,N_22187,N_22145);
nor U24467 (N_24467,N_22070,N_23905);
or U24468 (N_24468,N_22467,N_23593);
xor U24469 (N_24469,N_23248,N_22027);
and U24470 (N_24470,N_23584,N_23933);
nor U24471 (N_24471,N_23169,N_23526);
or U24472 (N_24472,N_23296,N_23118);
or U24473 (N_24473,N_23339,N_22390);
or U24474 (N_24474,N_23400,N_22920);
or U24475 (N_24475,N_22678,N_22465);
xnor U24476 (N_24476,N_22689,N_23326);
xnor U24477 (N_24477,N_22536,N_23460);
and U24478 (N_24478,N_23826,N_22229);
nor U24479 (N_24479,N_23074,N_23935);
or U24480 (N_24480,N_22901,N_22307);
nand U24481 (N_24481,N_23353,N_23689);
xor U24482 (N_24482,N_22639,N_22921);
nor U24483 (N_24483,N_23199,N_22119);
xnor U24484 (N_24484,N_23532,N_23459);
nand U24485 (N_24485,N_23937,N_23259);
nand U24486 (N_24486,N_22970,N_23330);
and U24487 (N_24487,N_23198,N_23023);
nand U24488 (N_24488,N_23652,N_23680);
or U24489 (N_24489,N_22598,N_22916);
xor U24490 (N_24490,N_23481,N_23379);
nor U24491 (N_24491,N_23059,N_23875);
or U24492 (N_24492,N_22533,N_23739);
nor U24493 (N_24493,N_22573,N_22599);
xnor U24494 (N_24494,N_22103,N_22746);
xnor U24495 (N_24495,N_23566,N_22756);
xnor U24496 (N_24496,N_22500,N_22993);
nand U24497 (N_24497,N_23914,N_23284);
and U24498 (N_24498,N_23084,N_23050);
or U24499 (N_24499,N_23963,N_22227);
nand U24500 (N_24500,N_22575,N_23842);
nand U24501 (N_24501,N_22585,N_23903);
nor U24502 (N_24502,N_22162,N_22594);
nor U24503 (N_24503,N_22033,N_23300);
nand U24504 (N_24504,N_23788,N_22387);
nand U24505 (N_24505,N_23136,N_22730);
nor U24506 (N_24506,N_22803,N_22109);
xor U24507 (N_24507,N_23863,N_23210);
nor U24508 (N_24508,N_22748,N_23939);
xor U24509 (N_24509,N_23770,N_22996);
xor U24510 (N_24510,N_23876,N_23152);
nor U24511 (N_24511,N_23917,N_22411);
or U24512 (N_24512,N_23060,N_23066);
and U24513 (N_24513,N_23369,N_23632);
and U24514 (N_24514,N_23378,N_22822);
and U24515 (N_24515,N_23420,N_22447);
nand U24516 (N_24516,N_23180,N_23675);
xnor U24517 (N_24517,N_23260,N_23692);
xor U24518 (N_24518,N_23467,N_22586);
nor U24519 (N_24519,N_22945,N_23732);
nand U24520 (N_24520,N_22569,N_23730);
nand U24521 (N_24521,N_22824,N_22944);
nand U24522 (N_24522,N_23579,N_23189);
and U24523 (N_24523,N_22058,N_23647);
nand U24524 (N_24524,N_22811,N_23570);
and U24525 (N_24525,N_23954,N_22849);
or U24526 (N_24526,N_22439,N_22512);
nand U24527 (N_24527,N_23598,N_23468);
or U24528 (N_24528,N_23565,N_22582);
nand U24529 (N_24529,N_23851,N_23796);
nor U24530 (N_24530,N_22799,N_23861);
or U24531 (N_24531,N_23049,N_23641);
or U24532 (N_24532,N_23332,N_22086);
nand U24533 (N_24533,N_23249,N_22218);
nand U24534 (N_24534,N_22408,N_23988);
nor U24535 (N_24535,N_22147,N_23430);
or U24536 (N_24536,N_23492,N_23521);
nor U24537 (N_24537,N_22020,N_22202);
nor U24538 (N_24538,N_22176,N_22863);
or U24539 (N_24539,N_22550,N_22136);
or U24540 (N_24540,N_22665,N_23197);
or U24541 (N_24541,N_23110,N_22810);
xor U24542 (N_24542,N_22700,N_23305);
nor U24543 (N_24543,N_22047,N_22727);
xor U24544 (N_24544,N_23499,N_22449);
and U24545 (N_24545,N_22348,N_22526);
nor U24546 (N_24546,N_23355,N_23366);
or U24547 (N_24547,N_23384,N_22435);
and U24548 (N_24548,N_23224,N_22128);
and U24549 (N_24549,N_23099,N_22726);
and U24550 (N_24550,N_23772,N_22636);
or U24551 (N_24551,N_23013,N_22505);
nand U24552 (N_24552,N_22942,N_23934);
xnor U24553 (N_24553,N_22232,N_22096);
nor U24554 (N_24554,N_22268,N_22170);
or U24555 (N_24555,N_23626,N_23660);
nor U24556 (N_24556,N_23945,N_23568);
nor U24557 (N_24557,N_22416,N_22001);
nor U24558 (N_24558,N_23666,N_23020);
or U24559 (N_24559,N_23989,N_22458);
xnor U24560 (N_24560,N_22894,N_23918);
or U24561 (N_24561,N_23999,N_23147);
xor U24562 (N_24562,N_22729,N_22854);
nor U24563 (N_24563,N_23027,N_23385);
and U24564 (N_24564,N_23528,N_23244);
xnor U24565 (N_24565,N_22844,N_23716);
nand U24566 (N_24566,N_22490,N_23261);
nor U24567 (N_24567,N_23129,N_23523);
and U24568 (N_24568,N_22443,N_23290);
nor U24569 (N_24569,N_22476,N_23961);
nand U24570 (N_24570,N_23465,N_23186);
xor U24571 (N_24571,N_23471,N_22666);
and U24572 (N_24572,N_23551,N_23165);
and U24573 (N_24573,N_23470,N_23886);
and U24574 (N_24574,N_22295,N_23986);
xnor U24575 (N_24575,N_23729,N_23193);
nor U24576 (N_24576,N_23682,N_22259);
or U24577 (N_24577,N_22420,N_22966);
and U24578 (N_24578,N_23849,N_22905);
or U24579 (N_24579,N_22642,N_23795);
or U24580 (N_24580,N_22167,N_22448);
nor U24581 (N_24581,N_22870,N_22793);
xor U24582 (N_24582,N_22277,N_23273);
nor U24583 (N_24583,N_23081,N_23748);
or U24584 (N_24584,N_22922,N_22523);
nor U24585 (N_24585,N_22777,N_22124);
xor U24586 (N_24586,N_22974,N_23327);
and U24587 (N_24587,N_23741,N_23710);
and U24588 (N_24588,N_22225,N_22469);
nor U24589 (N_24589,N_22843,N_22913);
xor U24590 (N_24590,N_23728,N_23889);
and U24591 (N_24591,N_23201,N_22766);
nor U24592 (N_24592,N_23318,N_22514);
or U24593 (N_24593,N_22566,N_23908);
nor U24594 (N_24594,N_22261,N_23120);
xor U24595 (N_24595,N_22551,N_23078);
xor U24596 (N_24596,N_22934,N_22157);
nor U24597 (N_24597,N_22992,N_23509);
or U24598 (N_24598,N_22608,N_22398);
nand U24599 (N_24599,N_22737,N_22376);
nand U24600 (N_24600,N_22498,N_22025);
or U24601 (N_24601,N_22997,N_23810);
and U24602 (N_24602,N_23496,N_23485);
and U24603 (N_24603,N_22592,N_23773);
and U24604 (N_24604,N_22525,N_23750);
nor U24605 (N_24605,N_23211,N_22049);
nor U24606 (N_24606,N_23182,N_23206);
nor U24607 (N_24607,N_22296,N_22361);
xor U24608 (N_24608,N_23222,N_23393);
or U24609 (N_24609,N_22524,N_23178);
and U24610 (N_24610,N_22886,N_22108);
nor U24611 (N_24611,N_22928,N_22330);
or U24612 (N_24612,N_22381,N_23845);
xnor U24613 (N_24613,N_23263,N_23650);
xor U24614 (N_24614,N_22702,N_23294);
nand U24615 (N_24615,N_22247,N_22669);
xnor U24616 (N_24616,N_23168,N_22254);
and U24617 (N_24617,N_23887,N_23161);
or U24618 (N_24618,N_23338,N_23449);
or U24619 (N_24619,N_23056,N_23144);
and U24620 (N_24620,N_22179,N_22391);
xor U24621 (N_24621,N_22763,N_23541);
nor U24622 (N_24622,N_22417,N_23998);
nor U24623 (N_24623,N_23154,N_22781);
nand U24624 (N_24624,N_22565,N_22701);
or U24625 (N_24625,N_22869,N_23316);
and U24626 (N_24626,N_23345,N_23832);
nand U24627 (N_24627,N_22904,N_22718);
nor U24628 (N_24628,N_23160,N_22823);
or U24629 (N_24629,N_22333,N_22280);
nor U24630 (N_24630,N_23213,N_22311);
xnor U24631 (N_24631,N_23980,N_22946);
xnor U24632 (N_24632,N_23052,N_22013);
or U24633 (N_24633,N_22183,N_23625);
nor U24634 (N_24634,N_23733,N_23622);
nand U24635 (N_24635,N_22224,N_22618);
or U24636 (N_24636,N_23623,N_23696);
or U24637 (N_24637,N_23958,N_22703);
and U24638 (N_24638,N_23287,N_23461);
and U24639 (N_24639,N_22805,N_22742);
or U24640 (N_24640,N_22958,N_23301);
and U24641 (N_24641,N_22888,N_23489);
nand U24642 (N_24642,N_23073,N_22943);
or U24643 (N_24643,N_23220,N_23505);
or U24644 (N_24644,N_23907,N_22724);
nor U24645 (N_24645,N_23836,N_22976);
xnor U24646 (N_24646,N_22784,N_23700);
and U24647 (N_24647,N_23522,N_22345);
and U24648 (N_24648,N_23047,N_23690);
nor U24649 (N_24649,N_23389,N_22036);
xnor U24650 (N_24650,N_22543,N_22004);
xnor U24651 (N_24651,N_23824,N_23484);
xor U24652 (N_24652,N_22470,N_22912);
or U24653 (N_24653,N_23964,N_22508);
and U24654 (N_24654,N_22673,N_23359);
and U24655 (N_24655,N_22562,N_22127);
nor U24656 (N_24656,N_23557,N_22511);
nand U24657 (N_24657,N_23289,N_22197);
nand U24658 (N_24658,N_23046,N_22021);
or U24659 (N_24659,N_22320,N_23938);
and U24660 (N_24660,N_23247,N_22780);
xnor U24661 (N_24661,N_22143,N_23395);
nand U24662 (N_24662,N_23662,N_23026);
and U24663 (N_24663,N_22216,N_23591);
or U24664 (N_24664,N_22557,N_22355);
nor U24665 (N_24665,N_23697,N_23141);
nor U24666 (N_24666,N_23067,N_23514);
and U24667 (N_24667,N_23846,N_22394);
and U24668 (N_24668,N_22925,N_23010);
or U24669 (N_24669,N_23719,N_22937);
or U24670 (N_24670,N_23149,N_23635);
xor U24671 (N_24671,N_23967,N_23403);
nor U24672 (N_24672,N_23321,N_22600);
or U24673 (N_24673,N_22077,N_22431);
or U24674 (N_24674,N_22640,N_22681);
or U24675 (N_24675,N_23646,N_23888);
nor U24676 (N_24676,N_23969,N_22831);
nor U24677 (N_24677,N_22265,N_23767);
nor U24678 (N_24678,N_22875,N_23757);
and U24679 (N_24679,N_22682,N_22318);
nor U24680 (N_24680,N_23925,N_22933);
and U24681 (N_24681,N_22832,N_22138);
xnor U24682 (N_24682,N_23559,N_22399);
or U24683 (N_24683,N_22362,N_23790);
nand U24684 (N_24684,N_23035,N_22787);
nor U24685 (N_24685,N_23701,N_23951);
and U24686 (N_24686,N_22900,N_23486);
nor U24687 (N_24687,N_22968,N_23088);
or U24688 (N_24688,N_23812,N_23024);
or U24689 (N_24689,N_22537,N_23406);
or U24690 (N_24690,N_22078,N_23373);
and U24691 (N_24691,N_23014,N_23029);
or U24692 (N_24692,N_23563,N_22825);
nand U24693 (N_24693,N_22306,N_23871);
or U24694 (N_24694,N_22174,N_23685);
xor U24695 (N_24695,N_22704,N_23620);
or U24696 (N_24696,N_22437,N_23916);
and U24697 (N_24697,N_23562,N_22158);
xnor U24698 (N_24698,N_22412,N_23758);
nand U24699 (N_24699,N_23545,N_23278);
nor U24700 (N_24700,N_23439,N_22641);
nor U24701 (N_24701,N_22110,N_23638);
nor U24702 (N_24702,N_22215,N_23760);
nor U24703 (N_24703,N_22648,N_23434);
and U24704 (N_24704,N_23664,N_23979);
nand U24705 (N_24705,N_22180,N_23544);
nand U24706 (N_24706,N_22483,N_23417);
nor U24707 (N_24707,N_23721,N_22535);
or U24708 (N_24708,N_23226,N_23367);
xnor U24709 (N_24709,N_23457,N_22856);
xnor U24710 (N_24710,N_23874,N_22073);
xor U24711 (N_24711,N_22568,N_22386);
xor U24712 (N_24712,N_23477,N_23507);
nor U24713 (N_24713,N_23377,N_23722);
or U24714 (N_24714,N_23547,N_22938);
xor U24715 (N_24715,N_22940,N_23100);
and U24716 (N_24716,N_23533,N_22423);
nor U24717 (N_24717,N_23478,N_22264);
nor U24718 (N_24718,N_23164,N_23717);
xor U24719 (N_24719,N_22747,N_22765);
xor U24720 (N_24720,N_22063,N_23107);
nand U24721 (N_24721,N_22164,N_22828);
and U24722 (N_24722,N_23694,N_22210);
or U24723 (N_24723,N_22068,N_22601);
xor U24724 (N_24724,N_22603,N_23597);
xor U24725 (N_24725,N_23693,N_22205);
xor U24726 (N_24726,N_22889,N_23092);
nor U24727 (N_24727,N_23829,N_22878);
xnor U24728 (N_24728,N_22137,N_22214);
and U24729 (N_24729,N_23784,N_22659);
xor U24730 (N_24730,N_22322,N_23740);
xor U24731 (N_24731,N_23329,N_22567);
xor U24732 (N_24732,N_22126,N_23337);
and U24733 (N_24733,N_23212,N_22246);
nor U24734 (N_24734,N_23621,N_22860);
and U24735 (N_24735,N_23873,N_22692);
or U24736 (N_24736,N_22895,N_22129);
nor U24737 (N_24737,N_22282,N_23028);
or U24738 (N_24738,N_22962,N_22624);
or U24739 (N_24739,N_22873,N_23902);
or U24740 (N_24740,N_23776,N_22100);
xor U24741 (N_24741,N_23843,N_23232);
or U24742 (N_24742,N_22393,N_23096);
nand U24743 (N_24743,N_22789,N_23844);
xor U24744 (N_24744,N_23018,N_23264);
or U24745 (N_24745,N_22755,N_22473);
and U24746 (N_24746,N_22534,N_22759);
and U24747 (N_24747,N_22230,N_22999);
nor U24748 (N_24748,N_22687,N_22181);
nand U24749 (N_24749,N_22240,N_23872);
nand U24750 (N_24750,N_22015,N_22407);
nand U24751 (N_24751,N_22055,N_23138);
and U24752 (N_24752,N_23575,N_22130);
nor U24753 (N_24753,N_23295,N_22384);
and U24754 (N_24754,N_23783,N_22776);
xor U24755 (N_24755,N_22948,N_23548);
or U24756 (N_24756,N_23285,N_22593);
xnor U24757 (N_24757,N_22816,N_22482);
or U24758 (N_24758,N_22541,N_22709);
nor U24759 (N_24759,N_23586,N_23828);
nor U24760 (N_24760,N_23582,N_22030);
and U24761 (N_24761,N_23358,N_22382);
nand U24762 (N_24762,N_23319,N_23031);
or U24763 (N_24763,N_22208,N_22492);
nor U24764 (N_24764,N_22801,N_23894);
nor U24765 (N_24765,N_23516,N_22696);
and U24766 (N_24766,N_22617,N_22884);
nor U24767 (N_24767,N_22278,N_22578);
nand U24768 (N_24768,N_22783,N_22037);
nor U24769 (N_24769,N_23944,N_23724);
and U24770 (N_24770,N_22419,N_22652);
xor U24771 (N_24771,N_22690,N_22298);
and U24772 (N_24772,N_23929,N_22890);
and U24773 (N_24773,N_22080,N_22008);
or U24774 (N_24774,N_22373,N_23146);
xnor U24775 (N_24775,N_22341,N_22635);
nand U24776 (N_24776,N_23825,N_22752);
or U24777 (N_24777,N_23830,N_22235);
nor U24778 (N_24778,N_23835,N_22198);
or U24779 (N_24779,N_23777,N_22907);
nand U24780 (N_24780,N_23266,N_23688);
xor U24781 (N_24781,N_22043,N_23034);
nor U24782 (N_24782,N_22359,N_23255);
nor U24783 (N_24783,N_23257,N_22807);
nor U24784 (N_24784,N_22749,N_23756);
xnor U24785 (N_24785,N_22099,N_23628);
xnor U24786 (N_24786,N_22152,N_23927);
xor U24787 (N_24787,N_23454,N_23215);
nor U24788 (N_24788,N_22434,N_23463);
nand U24789 (N_24789,N_23012,N_23304);
and U24790 (N_24790,N_23062,N_23535);
xor U24791 (N_24791,N_22651,N_22721);
xnor U24792 (N_24792,N_22809,N_23974);
or U24793 (N_24793,N_22661,N_22739);
or U24794 (N_24794,N_22675,N_23718);
and U24795 (N_24795,N_22556,N_22456);
nor U24796 (N_24796,N_23684,N_22699);
nor U24797 (N_24797,N_23602,N_23350);
or U24798 (N_24798,N_23083,N_22028);
nand U24799 (N_24799,N_23079,N_22046);
nor U24800 (N_24800,N_22826,N_23996);
nand U24801 (N_24801,N_23291,N_22808);
or U24802 (N_24802,N_23928,N_23553);
xnor U24803 (N_24803,N_23924,N_22655);
and U24804 (N_24804,N_23445,N_23837);
and U24805 (N_24805,N_22244,N_22865);
and U24806 (N_24806,N_23616,N_22309);
nand U24807 (N_24807,N_23560,N_22428);
and U24808 (N_24808,N_22685,N_22503);
nor U24809 (N_24809,N_22719,N_23525);
xor U24810 (N_24810,N_22538,N_23715);
xor U24811 (N_24811,N_23097,N_23595);
or U24812 (N_24812,N_22982,N_22845);
nor U24813 (N_24813,N_22506,N_22163);
nor U24814 (N_24814,N_23807,N_22236);
xor U24815 (N_24815,N_22510,N_23269);
or U24816 (N_24816,N_22761,N_22192);
xnor U24817 (N_24817,N_22633,N_22396);
and U24818 (N_24818,N_22168,N_23569);
or U24819 (N_24819,N_23094,N_23166);
nor U24820 (N_24820,N_23792,N_23627);
xnor U24821 (N_24821,N_23241,N_23852);
and U24822 (N_24822,N_22879,N_23272);
or U24823 (N_24823,N_23396,N_23947);
nand U24824 (N_24824,N_23909,N_23156);
or U24825 (N_24825,N_23949,N_23880);
xnor U24826 (N_24826,N_22939,N_22076);
xnor U24827 (N_24827,N_23038,N_23270);
or U24828 (N_24828,N_22561,N_23236);
or U24829 (N_24829,N_23904,N_23128);
xor U24830 (N_24830,N_23555,N_23392);
and U24831 (N_24831,N_22987,N_23604);
and U24832 (N_24832,N_22383,N_23552);
xor U24833 (N_24833,N_22089,N_22358);
or U24834 (N_24834,N_22806,N_23753);
nand U24835 (N_24835,N_22474,N_22397);
xor U24836 (N_24836,N_22680,N_22484);
and U24837 (N_24837,N_23674,N_22299);
or U24838 (N_24838,N_22588,N_22141);
and U24839 (N_24839,N_22834,N_22852);
nand U24840 (N_24840,N_22286,N_22190);
xor U24841 (N_24841,N_22877,N_22519);
and U24842 (N_24842,N_23451,N_22864);
nor U24843 (N_24843,N_22266,N_23893);
nand U24844 (N_24844,N_23041,N_23766);
nand U24845 (N_24845,N_22602,N_23006);
nand U24846 (N_24846,N_22274,N_22012);
and U24847 (N_24847,N_22134,N_23857);
and U24848 (N_24848,N_23102,N_23446);
xnor U24849 (N_24849,N_22339,N_23204);
or U24850 (N_24850,N_22615,N_22917);
nor U24851 (N_24851,N_22910,N_22347);
and U24852 (N_24852,N_22031,N_23228);
or U24853 (N_24853,N_23282,N_22107);
nand U24854 (N_24854,N_22479,N_22502);
and U24855 (N_24855,N_22830,N_22712);
nor U24856 (N_24856,N_23970,N_22425);
or U24857 (N_24857,N_23455,N_23435);
nand U24858 (N_24858,N_22120,N_23003);
nand U24859 (N_24859,N_23170,N_22555);
and U24860 (N_24860,N_22736,N_22066);
nand U24861 (N_24861,N_22984,N_23042);
nand U24862 (N_24862,N_23414,N_23712);
or U24863 (N_24863,N_23990,N_22316);
nor U24864 (N_24864,N_22310,N_23655);
xor U24865 (N_24865,N_22325,N_23624);
or U24866 (N_24866,N_23614,N_23130);
nor U24867 (N_24867,N_22619,N_23519);
and U24868 (N_24868,N_23892,N_22903);
nand U24869 (N_24869,N_22634,N_23308);
nand U24870 (N_24870,N_22092,N_23440);
nand U24871 (N_24871,N_23612,N_23117);
and U24872 (N_24872,N_23785,N_22454);
xor U24873 (N_24873,N_22285,N_23678);
xnor U24874 (N_24874,N_22853,N_22486);
nand U24875 (N_24875,N_23831,N_22710);
nand U24876 (N_24876,N_23520,N_23111);
nor U24877 (N_24877,N_23238,N_23356);
nand U24878 (N_24878,N_23564,N_23432);
xnor U24879 (N_24879,N_23527,N_22212);
nand U24880 (N_24880,N_22169,N_22930);
or U24881 (N_24881,N_22324,N_22253);
xor U24882 (N_24882,N_23265,N_22796);
and U24883 (N_24883,N_22172,N_22040);
nor U24884 (N_24884,N_22363,N_23061);
nand U24885 (N_24885,N_22413,N_23380);
nand U24886 (N_24886,N_23819,N_23140);
nand U24887 (N_24887,N_23209,N_22906);
nor U24888 (N_24888,N_22716,N_22487);
nand U24889 (N_24889,N_22545,N_22785);
nand U24890 (N_24890,N_23919,N_23490);
nand U24891 (N_24891,N_22927,N_23127);
xnor U24892 (N_24892,N_22978,N_23910);
nor U24893 (N_24893,N_23173,N_23427);
nor U24894 (N_24894,N_22213,N_23850);
nor U24895 (N_24895,N_22222,N_23017);
xnor U24896 (N_24896,N_22493,N_23331);
nand U24897 (N_24897,N_23181,N_23823);
nor U24898 (N_24898,N_22881,N_22846);
and U24899 (N_24899,N_22155,N_23080);
xnor U24900 (N_24900,N_22106,N_23363);
and U24901 (N_24901,N_22173,N_23196);
or U24902 (N_24902,N_23799,N_23745);
and U24903 (N_24903,N_22861,N_23671);
nand U24904 (N_24904,N_23254,N_22368);
nor U24905 (N_24905,N_22758,N_22768);
nor U24906 (N_24906,N_23946,N_23233);
nor U24907 (N_24907,N_22560,N_22052);
or U24908 (N_24908,N_22722,N_22960);
and U24909 (N_24909,N_23779,N_22457);
nor U24910 (N_24910,N_23899,N_23508);
and U24911 (N_24911,N_22385,N_23686);
nand U24912 (N_24912,N_22638,N_22231);
and U24913 (N_24913,N_22558,N_23157);
nand U24914 (N_24914,N_22352,N_23881);
nor U24915 (N_24915,N_22034,N_23404);
xnor U24916 (N_24916,N_22018,N_22389);
nand U24917 (N_24917,N_23821,N_23475);
nor U24918 (N_24918,N_22042,N_23302);
nand U24919 (N_24919,N_22079,N_22071);
xnor U24920 (N_24920,N_23159,N_23354);
and U24921 (N_24921,N_23755,N_22892);
nor U24922 (N_24922,N_23501,N_22896);
or U24923 (N_24923,N_23191,N_22610);
xnor U24924 (N_24924,N_23769,N_23636);
or U24925 (N_24925,N_22211,N_23007);
or U24926 (N_24926,N_22499,N_22495);
nand U24927 (N_24927,N_22570,N_22909);
or U24928 (N_24928,N_22409,N_22953);
nor U24929 (N_24929,N_23921,N_22539);
nor U24930 (N_24930,N_23884,N_23348);
xnor U24931 (N_24931,N_22477,N_22314);
nand U24932 (N_24932,N_23425,N_23106);
nor U24933 (N_24933,N_22862,N_22217);
nor U24934 (N_24934,N_22045,N_22459);
or U24935 (N_24935,N_22000,N_22795);
or U24936 (N_24936,N_22774,N_23995);
or U24937 (N_24937,N_22329,N_23443);
nand U24938 (N_24938,N_22630,N_22303);
or U24939 (N_24939,N_23086,N_22866);
nor U24940 (N_24940,N_23506,N_23025);
or U24941 (N_24941,N_22717,N_23150);
or U24942 (N_24942,N_22605,N_23737);
and U24943 (N_24943,N_23787,N_23809);
xnor U24944 (N_24944,N_22876,N_23764);
and U24945 (N_24945,N_23448,N_22597);
nor U24946 (N_24946,N_22715,N_23143);
xor U24947 (N_24947,N_23095,N_23135);
or U24948 (N_24948,N_22101,N_22257);
or U24949 (N_24949,N_23955,N_23723);
nor U24950 (N_24950,N_22629,N_23651);
nor U24951 (N_24951,N_22985,N_22553);
xor U24952 (N_24952,N_23202,N_22375);
and U24953 (N_24953,N_23153,N_23207);
nand U24954 (N_24954,N_23941,N_23280);
xnor U24955 (N_24955,N_22547,N_22732);
nand U24956 (N_24956,N_23920,N_22882);
or U24957 (N_24957,N_22453,N_22802);
and U24958 (N_24958,N_22243,N_23870);
xnor U24959 (N_24959,N_23643,N_23962);
nand U24960 (N_24960,N_23177,N_23677);
nand U24961 (N_24961,N_22623,N_23705);
xor U24962 (N_24962,N_23708,N_22350);
nor U24963 (N_24963,N_23531,N_22095);
xnor U24964 (N_24964,N_23441,N_22572);
nand U24965 (N_24965,N_22871,N_23328);
and U24966 (N_24966,N_23452,N_23571);
nand U24967 (N_24967,N_22609,N_23476);
or U24968 (N_24968,N_22658,N_22549);
xor U24969 (N_24969,N_22313,N_23473);
xor U24970 (N_24970,N_23172,N_23281);
and U24971 (N_24971,N_22589,N_23854);
nor U24972 (N_24972,N_23618,N_23494);
xor U24973 (N_24973,N_23390,N_23912);
nand U24974 (N_24974,N_23217,N_22151);
nand U24975 (N_24975,N_23891,N_23761);
xnor U24976 (N_24976,N_23611,N_22656);
nor U24977 (N_24977,N_22460,N_23587);
nor U24978 (N_24978,N_22220,N_22255);
nor U24979 (N_24979,N_23072,N_22267);
xor U24980 (N_24980,N_23605,N_22714);
xor U24981 (N_24981,N_22936,N_22022);
nor U24982 (N_24982,N_23778,N_22591);
or U24983 (N_24983,N_23987,N_23142);
xor U24984 (N_24984,N_23402,N_22841);
or U24985 (N_24985,N_22778,N_23175);
nor U24986 (N_24986,N_23317,N_22380);
nor U24987 (N_24987,N_23744,N_22671);
or U24988 (N_24988,N_23806,N_22340);
nor U24989 (N_24989,N_22009,N_23015);
nand U24990 (N_24990,N_23139,N_23956);
or U24991 (N_24991,N_22353,N_23802);
nor U24992 (N_24992,N_23536,N_22735);
nor U24993 (N_24993,N_23466,N_23493);
nand U24994 (N_24994,N_22111,N_23600);
and U24995 (N_24995,N_23749,N_23653);
nand U24996 (N_24996,N_23320,N_22850);
or U24997 (N_24997,N_23897,N_22674);
nand U24998 (N_24998,N_22258,N_22035);
xor U24999 (N_24999,N_23246,N_22504);
nor U25000 (N_25000,N_23255,N_22837);
or U25001 (N_25001,N_22285,N_23034);
and U25002 (N_25002,N_22160,N_23619);
and U25003 (N_25003,N_22355,N_23048);
xor U25004 (N_25004,N_22469,N_22602);
or U25005 (N_25005,N_23888,N_22907);
or U25006 (N_25006,N_22360,N_22358);
nor U25007 (N_25007,N_23525,N_22606);
and U25008 (N_25008,N_22288,N_22005);
xnor U25009 (N_25009,N_23519,N_22737);
nor U25010 (N_25010,N_23421,N_23835);
and U25011 (N_25011,N_22696,N_23621);
or U25012 (N_25012,N_23125,N_22685);
nor U25013 (N_25013,N_23513,N_23479);
nor U25014 (N_25014,N_22201,N_22649);
nor U25015 (N_25015,N_23656,N_23468);
nor U25016 (N_25016,N_23225,N_23577);
nor U25017 (N_25017,N_23397,N_22629);
or U25018 (N_25018,N_22646,N_23085);
and U25019 (N_25019,N_23458,N_22800);
or U25020 (N_25020,N_22767,N_23412);
and U25021 (N_25021,N_22134,N_23248);
nand U25022 (N_25022,N_22986,N_22173);
or U25023 (N_25023,N_22887,N_22509);
xor U25024 (N_25024,N_23453,N_22889);
nor U25025 (N_25025,N_22700,N_22501);
and U25026 (N_25026,N_22548,N_23275);
or U25027 (N_25027,N_23944,N_22675);
xor U25028 (N_25028,N_23427,N_22051);
xor U25029 (N_25029,N_23503,N_23719);
xor U25030 (N_25030,N_22158,N_23830);
and U25031 (N_25031,N_23141,N_22097);
nor U25032 (N_25032,N_22654,N_23811);
nor U25033 (N_25033,N_23977,N_22651);
xnor U25034 (N_25034,N_22433,N_22169);
xor U25035 (N_25035,N_22666,N_22053);
nand U25036 (N_25036,N_23417,N_23262);
or U25037 (N_25037,N_23991,N_23089);
nand U25038 (N_25038,N_23078,N_22604);
or U25039 (N_25039,N_23299,N_22736);
and U25040 (N_25040,N_23374,N_23973);
or U25041 (N_25041,N_23907,N_22696);
or U25042 (N_25042,N_22056,N_23907);
or U25043 (N_25043,N_23588,N_22561);
nor U25044 (N_25044,N_23616,N_22179);
or U25045 (N_25045,N_23767,N_22596);
nor U25046 (N_25046,N_22225,N_22753);
nor U25047 (N_25047,N_22907,N_23812);
or U25048 (N_25048,N_23478,N_23829);
nor U25049 (N_25049,N_22790,N_22087);
or U25050 (N_25050,N_23370,N_22783);
or U25051 (N_25051,N_22072,N_22079);
nor U25052 (N_25052,N_23685,N_22268);
xor U25053 (N_25053,N_23076,N_23846);
xor U25054 (N_25054,N_23854,N_23547);
xnor U25055 (N_25055,N_22093,N_23069);
nand U25056 (N_25056,N_23482,N_23488);
or U25057 (N_25057,N_23474,N_22970);
and U25058 (N_25058,N_22893,N_23842);
xnor U25059 (N_25059,N_22148,N_22242);
nor U25060 (N_25060,N_23837,N_22688);
nor U25061 (N_25061,N_22089,N_22284);
nand U25062 (N_25062,N_22888,N_22417);
and U25063 (N_25063,N_22974,N_23370);
xnor U25064 (N_25064,N_22230,N_22775);
xor U25065 (N_25065,N_23865,N_23368);
and U25066 (N_25066,N_22448,N_22427);
nand U25067 (N_25067,N_23960,N_23440);
nor U25068 (N_25068,N_22576,N_23767);
nor U25069 (N_25069,N_22506,N_23526);
and U25070 (N_25070,N_22551,N_22762);
or U25071 (N_25071,N_22354,N_23805);
or U25072 (N_25072,N_22429,N_22959);
xnor U25073 (N_25073,N_22074,N_23602);
nand U25074 (N_25074,N_22193,N_23900);
xor U25075 (N_25075,N_22565,N_22938);
and U25076 (N_25076,N_23189,N_23706);
or U25077 (N_25077,N_22315,N_22444);
xnor U25078 (N_25078,N_23861,N_22819);
nor U25079 (N_25079,N_23381,N_22349);
nor U25080 (N_25080,N_22604,N_23166);
and U25081 (N_25081,N_22929,N_22304);
and U25082 (N_25082,N_22845,N_23136);
xor U25083 (N_25083,N_23020,N_22492);
nand U25084 (N_25084,N_23453,N_22004);
nor U25085 (N_25085,N_23924,N_22392);
nor U25086 (N_25086,N_22334,N_23213);
or U25087 (N_25087,N_23350,N_22615);
nand U25088 (N_25088,N_23723,N_23570);
nor U25089 (N_25089,N_22304,N_22392);
xnor U25090 (N_25090,N_22034,N_22149);
nand U25091 (N_25091,N_23318,N_23346);
or U25092 (N_25092,N_23968,N_22777);
or U25093 (N_25093,N_23351,N_22147);
nor U25094 (N_25094,N_23081,N_22088);
nor U25095 (N_25095,N_22095,N_22619);
or U25096 (N_25096,N_22838,N_22244);
or U25097 (N_25097,N_23006,N_22069);
xor U25098 (N_25098,N_22038,N_23093);
xnor U25099 (N_25099,N_22905,N_23866);
nor U25100 (N_25100,N_23766,N_23983);
nor U25101 (N_25101,N_22918,N_23518);
or U25102 (N_25102,N_22817,N_22477);
and U25103 (N_25103,N_22823,N_22418);
and U25104 (N_25104,N_23568,N_22100);
and U25105 (N_25105,N_22587,N_23545);
or U25106 (N_25106,N_22679,N_22291);
or U25107 (N_25107,N_22369,N_23117);
nor U25108 (N_25108,N_23841,N_23063);
xnor U25109 (N_25109,N_22030,N_23597);
or U25110 (N_25110,N_22922,N_22005);
or U25111 (N_25111,N_23977,N_22890);
nor U25112 (N_25112,N_23211,N_22848);
or U25113 (N_25113,N_22847,N_22492);
xor U25114 (N_25114,N_23047,N_22450);
nor U25115 (N_25115,N_23352,N_22108);
xnor U25116 (N_25116,N_23615,N_22852);
nand U25117 (N_25117,N_23295,N_23191);
xnor U25118 (N_25118,N_23642,N_23543);
xnor U25119 (N_25119,N_23599,N_22861);
xor U25120 (N_25120,N_23991,N_22095);
xor U25121 (N_25121,N_23543,N_23967);
xor U25122 (N_25122,N_22527,N_23643);
xnor U25123 (N_25123,N_22863,N_23985);
nand U25124 (N_25124,N_23559,N_22340);
or U25125 (N_25125,N_23238,N_22410);
nand U25126 (N_25126,N_22396,N_23441);
nand U25127 (N_25127,N_22237,N_23560);
nor U25128 (N_25128,N_22905,N_22525);
and U25129 (N_25129,N_22370,N_22804);
nand U25130 (N_25130,N_23829,N_23095);
xnor U25131 (N_25131,N_22894,N_22314);
nand U25132 (N_25132,N_23519,N_22902);
and U25133 (N_25133,N_22319,N_22982);
nand U25134 (N_25134,N_23130,N_22231);
nor U25135 (N_25135,N_22128,N_22735);
nand U25136 (N_25136,N_23301,N_23286);
nor U25137 (N_25137,N_22842,N_23766);
xor U25138 (N_25138,N_23185,N_22198);
nor U25139 (N_25139,N_23847,N_22605);
xor U25140 (N_25140,N_22643,N_23660);
nand U25141 (N_25141,N_23066,N_22476);
nor U25142 (N_25142,N_22527,N_23367);
xor U25143 (N_25143,N_23314,N_22935);
nor U25144 (N_25144,N_22432,N_23796);
or U25145 (N_25145,N_23466,N_22499);
nor U25146 (N_25146,N_23608,N_22536);
xor U25147 (N_25147,N_22116,N_23150);
xnor U25148 (N_25148,N_23126,N_23129);
xor U25149 (N_25149,N_22684,N_22786);
and U25150 (N_25150,N_22464,N_23644);
xnor U25151 (N_25151,N_23622,N_23144);
nor U25152 (N_25152,N_23143,N_23000);
or U25153 (N_25153,N_23087,N_22845);
xor U25154 (N_25154,N_22677,N_23065);
nand U25155 (N_25155,N_23665,N_22734);
xnor U25156 (N_25156,N_22457,N_22381);
nor U25157 (N_25157,N_23147,N_22161);
nor U25158 (N_25158,N_23978,N_22515);
and U25159 (N_25159,N_23987,N_22541);
or U25160 (N_25160,N_23516,N_23573);
and U25161 (N_25161,N_23298,N_23642);
nor U25162 (N_25162,N_23394,N_22503);
and U25163 (N_25163,N_23888,N_23943);
nor U25164 (N_25164,N_23013,N_22418);
and U25165 (N_25165,N_23638,N_22039);
or U25166 (N_25166,N_23412,N_23385);
xor U25167 (N_25167,N_23312,N_22123);
nand U25168 (N_25168,N_23397,N_23966);
nor U25169 (N_25169,N_22028,N_23412);
or U25170 (N_25170,N_22242,N_22336);
and U25171 (N_25171,N_22789,N_23694);
xor U25172 (N_25172,N_22627,N_23798);
nand U25173 (N_25173,N_22015,N_23940);
xor U25174 (N_25174,N_23194,N_22830);
xor U25175 (N_25175,N_22633,N_23151);
or U25176 (N_25176,N_22968,N_23858);
xor U25177 (N_25177,N_23052,N_23006);
nor U25178 (N_25178,N_23303,N_23732);
nand U25179 (N_25179,N_23391,N_23835);
nand U25180 (N_25180,N_23520,N_23704);
or U25181 (N_25181,N_22492,N_23237);
and U25182 (N_25182,N_22069,N_23817);
nor U25183 (N_25183,N_23338,N_23767);
or U25184 (N_25184,N_23298,N_22489);
and U25185 (N_25185,N_22263,N_23455);
nand U25186 (N_25186,N_23214,N_22071);
nand U25187 (N_25187,N_23559,N_22116);
or U25188 (N_25188,N_23954,N_22369);
nand U25189 (N_25189,N_23742,N_23832);
nand U25190 (N_25190,N_22071,N_22488);
and U25191 (N_25191,N_23736,N_22945);
nor U25192 (N_25192,N_23090,N_22065);
or U25193 (N_25193,N_23531,N_23472);
nor U25194 (N_25194,N_23915,N_23080);
nor U25195 (N_25195,N_23590,N_23588);
and U25196 (N_25196,N_23523,N_22972);
xnor U25197 (N_25197,N_22851,N_23968);
nor U25198 (N_25198,N_22924,N_22005);
nand U25199 (N_25199,N_22017,N_23154);
or U25200 (N_25200,N_22295,N_22488);
nor U25201 (N_25201,N_22548,N_22148);
nor U25202 (N_25202,N_23588,N_22083);
or U25203 (N_25203,N_23262,N_22464);
or U25204 (N_25204,N_22934,N_22714);
nand U25205 (N_25205,N_22314,N_22701);
nor U25206 (N_25206,N_23246,N_22453);
nor U25207 (N_25207,N_22824,N_23835);
or U25208 (N_25208,N_22061,N_23116);
xnor U25209 (N_25209,N_23875,N_22491);
xor U25210 (N_25210,N_23193,N_23024);
nor U25211 (N_25211,N_23758,N_23097);
xor U25212 (N_25212,N_23879,N_22968);
nand U25213 (N_25213,N_23785,N_23471);
xnor U25214 (N_25214,N_22224,N_22175);
or U25215 (N_25215,N_22733,N_22354);
and U25216 (N_25216,N_23331,N_22416);
nand U25217 (N_25217,N_23051,N_22332);
nor U25218 (N_25218,N_23228,N_23118);
nand U25219 (N_25219,N_23908,N_23878);
nor U25220 (N_25220,N_22228,N_22212);
nor U25221 (N_25221,N_22724,N_22570);
nor U25222 (N_25222,N_22301,N_22733);
nor U25223 (N_25223,N_22784,N_22417);
or U25224 (N_25224,N_22341,N_23892);
or U25225 (N_25225,N_22507,N_22703);
xnor U25226 (N_25226,N_23973,N_23223);
or U25227 (N_25227,N_22672,N_22939);
and U25228 (N_25228,N_23370,N_23401);
nand U25229 (N_25229,N_23175,N_22822);
and U25230 (N_25230,N_22608,N_23792);
or U25231 (N_25231,N_23710,N_22231);
or U25232 (N_25232,N_22167,N_23853);
or U25233 (N_25233,N_22744,N_22454);
and U25234 (N_25234,N_22983,N_22063);
nand U25235 (N_25235,N_23989,N_22628);
xor U25236 (N_25236,N_22456,N_23198);
and U25237 (N_25237,N_22741,N_22264);
or U25238 (N_25238,N_23300,N_23501);
or U25239 (N_25239,N_23918,N_22405);
xnor U25240 (N_25240,N_23016,N_23102);
nor U25241 (N_25241,N_22099,N_23546);
nand U25242 (N_25242,N_23579,N_22791);
xnor U25243 (N_25243,N_22743,N_23094);
or U25244 (N_25244,N_23764,N_22346);
or U25245 (N_25245,N_23262,N_23819);
nor U25246 (N_25246,N_23110,N_23686);
nor U25247 (N_25247,N_23671,N_22810);
and U25248 (N_25248,N_22626,N_23542);
or U25249 (N_25249,N_22517,N_22058);
nor U25250 (N_25250,N_23898,N_22174);
and U25251 (N_25251,N_23421,N_23141);
or U25252 (N_25252,N_23561,N_22442);
xor U25253 (N_25253,N_23606,N_23262);
or U25254 (N_25254,N_23314,N_23027);
nand U25255 (N_25255,N_23400,N_23859);
and U25256 (N_25256,N_23984,N_22396);
or U25257 (N_25257,N_22938,N_22092);
and U25258 (N_25258,N_22879,N_22985);
nor U25259 (N_25259,N_23577,N_23022);
and U25260 (N_25260,N_23278,N_23934);
xor U25261 (N_25261,N_23373,N_23921);
nand U25262 (N_25262,N_22707,N_22225);
nor U25263 (N_25263,N_23118,N_22407);
and U25264 (N_25264,N_23597,N_23204);
nor U25265 (N_25265,N_22389,N_23355);
xor U25266 (N_25266,N_22841,N_22020);
and U25267 (N_25267,N_22742,N_23342);
or U25268 (N_25268,N_22489,N_23874);
and U25269 (N_25269,N_22982,N_23450);
nand U25270 (N_25270,N_22540,N_23438);
xnor U25271 (N_25271,N_23304,N_22609);
or U25272 (N_25272,N_22786,N_23287);
nand U25273 (N_25273,N_22431,N_22837);
nor U25274 (N_25274,N_23226,N_22386);
nand U25275 (N_25275,N_22968,N_22684);
nor U25276 (N_25276,N_22347,N_22019);
nand U25277 (N_25277,N_22628,N_23156);
or U25278 (N_25278,N_23608,N_23978);
nand U25279 (N_25279,N_22128,N_23663);
nor U25280 (N_25280,N_23977,N_23862);
nor U25281 (N_25281,N_22902,N_23684);
or U25282 (N_25282,N_23104,N_22095);
xor U25283 (N_25283,N_22433,N_23226);
nor U25284 (N_25284,N_22857,N_23242);
and U25285 (N_25285,N_22534,N_23198);
xor U25286 (N_25286,N_22060,N_22800);
nand U25287 (N_25287,N_23635,N_23837);
nor U25288 (N_25288,N_22746,N_23244);
nand U25289 (N_25289,N_23448,N_23518);
nand U25290 (N_25290,N_22870,N_22136);
or U25291 (N_25291,N_23175,N_23713);
nor U25292 (N_25292,N_22238,N_23249);
nor U25293 (N_25293,N_22281,N_23159);
nor U25294 (N_25294,N_23321,N_22664);
xor U25295 (N_25295,N_22618,N_22920);
nand U25296 (N_25296,N_23031,N_22162);
nand U25297 (N_25297,N_23680,N_22161);
xnor U25298 (N_25298,N_23727,N_23869);
or U25299 (N_25299,N_22703,N_23487);
or U25300 (N_25300,N_22662,N_22011);
nor U25301 (N_25301,N_23956,N_23805);
or U25302 (N_25302,N_22461,N_22896);
or U25303 (N_25303,N_22362,N_23888);
nand U25304 (N_25304,N_22576,N_23921);
nand U25305 (N_25305,N_23869,N_22382);
nand U25306 (N_25306,N_23384,N_22759);
nor U25307 (N_25307,N_22011,N_22100);
and U25308 (N_25308,N_22405,N_22345);
nand U25309 (N_25309,N_23877,N_22978);
or U25310 (N_25310,N_23289,N_22467);
or U25311 (N_25311,N_23206,N_22561);
and U25312 (N_25312,N_22727,N_23459);
or U25313 (N_25313,N_22096,N_22954);
nor U25314 (N_25314,N_22488,N_22775);
nand U25315 (N_25315,N_23371,N_22899);
nand U25316 (N_25316,N_23298,N_23925);
nor U25317 (N_25317,N_22925,N_22612);
xnor U25318 (N_25318,N_23074,N_23830);
xor U25319 (N_25319,N_23779,N_23168);
xor U25320 (N_25320,N_23827,N_23168);
or U25321 (N_25321,N_23522,N_22514);
nor U25322 (N_25322,N_22410,N_22811);
xnor U25323 (N_25323,N_23114,N_22851);
nand U25324 (N_25324,N_22553,N_23246);
and U25325 (N_25325,N_23466,N_23099);
nand U25326 (N_25326,N_22956,N_22001);
nor U25327 (N_25327,N_22141,N_22951);
xnor U25328 (N_25328,N_23539,N_22263);
nand U25329 (N_25329,N_23682,N_22592);
and U25330 (N_25330,N_22056,N_23142);
nor U25331 (N_25331,N_23397,N_23110);
xor U25332 (N_25332,N_22038,N_23676);
nor U25333 (N_25333,N_22115,N_23140);
and U25334 (N_25334,N_23756,N_22342);
nand U25335 (N_25335,N_22282,N_22179);
nor U25336 (N_25336,N_22339,N_22864);
nor U25337 (N_25337,N_22178,N_22827);
and U25338 (N_25338,N_23703,N_23102);
xor U25339 (N_25339,N_22708,N_23634);
and U25340 (N_25340,N_23525,N_22721);
nor U25341 (N_25341,N_22677,N_22004);
nor U25342 (N_25342,N_22701,N_22948);
and U25343 (N_25343,N_23908,N_23219);
nor U25344 (N_25344,N_23728,N_23942);
xnor U25345 (N_25345,N_23158,N_23283);
xor U25346 (N_25346,N_23830,N_23528);
nand U25347 (N_25347,N_23877,N_22969);
nand U25348 (N_25348,N_23647,N_23591);
and U25349 (N_25349,N_22048,N_23151);
xor U25350 (N_25350,N_22062,N_23399);
nand U25351 (N_25351,N_23779,N_22276);
and U25352 (N_25352,N_22627,N_23255);
and U25353 (N_25353,N_22216,N_22122);
and U25354 (N_25354,N_23835,N_22420);
and U25355 (N_25355,N_23698,N_23401);
xnor U25356 (N_25356,N_23292,N_23448);
nand U25357 (N_25357,N_22686,N_22176);
nor U25358 (N_25358,N_23488,N_22293);
nand U25359 (N_25359,N_23238,N_22568);
or U25360 (N_25360,N_23489,N_22253);
nand U25361 (N_25361,N_23862,N_23358);
nor U25362 (N_25362,N_22606,N_22400);
or U25363 (N_25363,N_22354,N_23021);
or U25364 (N_25364,N_22476,N_22067);
xnor U25365 (N_25365,N_23673,N_23396);
nand U25366 (N_25366,N_23829,N_23305);
and U25367 (N_25367,N_23820,N_22338);
nand U25368 (N_25368,N_22543,N_23415);
or U25369 (N_25369,N_23341,N_22416);
xnor U25370 (N_25370,N_23743,N_23988);
xor U25371 (N_25371,N_22140,N_23882);
xnor U25372 (N_25372,N_23767,N_23300);
xor U25373 (N_25373,N_23258,N_23362);
nand U25374 (N_25374,N_23946,N_23213);
or U25375 (N_25375,N_23738,N_23832);
xnor U25376 (N_25376,N_22055,N_23945);
xnor U25377 (N_25377,N_23005,N_22897);
or U25378 (N_25378,N_23359,N_23907);
xnor U25379 (N_25379,N_22098,N_22752);
or U25380 (N_25380,N_23383,N_23810);
xnor U25381 (N_25381,N_22643,N_22302);
nand U25382 (N_25382,N_23059,N_23260);
nand U25383 (N_25383,N_22251,N_23904);
nand U25384 (N_25384,N_22069,N_23406);
xor U25385 (N_25385,N_23369,N_22401);
nor U25386 (N_25386,N_23417,N_23331);
or U25387 (N_25387,N_23637,N_22174);
nor U25388 (N_25388,N_23198,N_22170);
or U25389 (N_25389,N_23585,N_22896);
or U25390 (N_25390,N_23832,N_23781);
nand U25391 (N_25391,N_23505,N_22227);
or U25392 (N_25392,N_22695,N_22818);
xnor U25393 (N_25393,N_23227,N_23727);
nand U25394 (N_25394,N_23974,N_22874);
xnor U25395 (N_25395,N_22702,N_22753);
nor U25396 (N_25396,N_22949,N_22554);
xor U25397 (N_25397,N_23724,N_23308);
nor U25398 (N_25398,N_23612,N_22816);
or U25399 (N_25399,N_23618,N_22078);
nand U25400 (N_25400,N_23291,N_23161);
or U25401 (N_25401,N_22743,N_22731);
or U25402 (N_25402,N_23781,N_22691);
nor U25403 (N_25403,N_23474,N_22854);
and U25404 (N_25404,N_22932,N_23204);
and U25405 (N_25405,N_23828,N_23633);
xor U25406 (N_25406,N_23840,N_23510);
and U25407 (N_25407,N_22782,N_22161);
xor U25408 (N_25408,N_23045,N_23365);
nor U25409 (N_25409,N_23467,N_23294);
xnor U25410 (N_25410,N_22583,N_23107);
nor U25411 (N_25411,N_22962,N_23445);
and U25412 (N_25412,N_23784,N_22558);
or U25413 (N_25413,N_23070,N_22683);
and U25414 (N_25414,N_23890,N_22439);
nand U25415 (N_25415,N_22733,N_23595);
xnor U25416 (N_25416,N_23985,N_23582);
or U25417 (N_25417,N_23370,N_23349);
xnor U25418 (N_25418,N_23840,N_23788);
nor U25419 (N_25419,N_23970,N_23835);
xnor U25420 (N_25420,N_23934,N_22476);
nor U25421 (N_25421,N_23219,N_22810);
nand U25422 (N_25422,N_22268,N_23072);
nand U25423 (N_25423,N_22279,N_22540);
nand U25424 (N_25424,N_23419,N_23368);
and U25425 (N_25425,N_23601,N_23297);
xor U25426 (N_25426,N_23133,N_23936);
nand U25427 (N_25427,N_22461,N_23222);
nor U25428 (N_25428,N_22843,N_23186);
and U25429 (N_25429,N_22067,N_22099);
nand U25430 (N_25430,N_23971,N_22780);
and U25431 (N_25431,N_23298,N_22501);
nor U25432 (N_25432,N_22138,N_22590);
nand U25433 (N_25433,N_23223,N_22702);
and U25434 (N_25434,N_23471,N_23845);
xnor U25435 (N_25435,N_22352,N_23989);
nand U25436 (N_25436,N_22594,N_23012);
xnor U25437 (N_25437,N_23389,N_23296);
nand U25438 (N_25438,N_22113,N_22317);
and U25439 (N_25439,N_23602,N_23686);
and U25440 (N_25440,N_23596,N_23243);
nor U25441 (N_25441,N_22285,N_22631);
and U25442 (N_25442,N_22372,N_22473);
nand U25443 (N_25443,N_22093,N_22903);
nor U25444 (N_25444,N_23649,N_22844);
or U25445 (N_25445,N_23222,N_23175);
xnor U25446 (N_25446,N_22791,N_22781);
or U25447 (N_25447,N_23062,N_23986);
xnor U25448 (N_25448,N_23185,N_23516);
nor U25449 (N_25449,N_22267,N_23709);
nor U25450 (N_25450,N_22246,N_22610);
or U25451 (N_25451,N_23612,N_22307);
xnor U25452 (N_25452,N_22834,N_22577);
nand U25453 (N_25453,N_22647,N_23536);
and U25454 (N_25454,N_23139,N_23765);
and U25455 (N_25455,N_22344,N_22691);
nor U25456 (N_25456,N_23510,N_23277);
and U25457 (N_25457,N_23865,N_23340);
nand U25458 (N_25458,N_23642,N_23550);
nor U25459 (N_25459,N_23485,N_23857);
and U25460 (N_25460,N_22449,N_22696);
or U25461 (N_25461,N_22023,N_23330);
xnor U25462 (N_25462,N_23326,N_22938);
and U25463 (N_25463,N_23566,N_23977);
and U25464 (N_25464,N_22271,N_22280);
nor U25465 (N_25465,N_22152,N_22540);
or U25466 (N_25466,N_22601,N_23166);
and U25467 (N_25467,N_23015,N_23742);
nor U25468 (N_25468,N_23526,N_22101);
or U25469 (N_25469,N_23277,N_22160);
xor U25470 (N_25470,N_22594,N_23311);
nand U25471 (N_25471,N_23805,N_23882);
and U25472 (N_25472,N_22884,N_22959);
nor U25473 (N_25473,N_22414,N_23681);
nor U25474 (N_25474,N_22001,N_22021);
nor U25475 (N_25475,N_22817,N_22175);
nor U25476 (N_25476,N_23314,N_22076);
xor U25477 (N_25477,N_23028,N_22403);
nor U25478 (N_25478,N_23797,N_22614);
xnor U25479 (N_25479,N_23437,N_22907);
and U25480 (N_25480,N_22386,N_23916);
or U25481 (N_25481,N_22494,N_22428);
xor U25482 (N_25482,N_22021,N_23502);
nor U25483 (N_25483,N_22368,N_23303);
or U25484 (N_25484,N_23917,N_23871);
nand U25485 (N_25485,N_23277,N_23640);
nand U25486 (N_25486,N_23021,N_23445);
and U25487 (N_25487,N_22110,N_22252);
nand U25488 (N_25488,N_22059,N_22190);
or U25489 (N_25489,N_23130,N_23437);
and U25490 (N_25490,N_22426,N_22734);
or U25491 (N_25491,N_23598,N_22534);
nand U25492 (N_25492,N_22061,N_22646);
nor U25493 (N_25493,N_22632,N_22406);
xor U25494 (N_25494,N_22325,N_22605);
xor U25495 (N_25495,N_22464,N_23547);
xnor U25496 (N_25496,N_22560,N_23770);
and U25497 (N_25497,N_22082,N_23842);
or U25498 (N_25498,N_23407,N_23558);
xnor U25499 (N_25499,N_23626,N_22650);
and U25500 (N_25500,N_22753,N_23107);
nand U25501 (N_25501,N_23723,N_22740);
xor U25502 (N_25502,N_23973,N_22819);
nand U25503 (N_25503,N_23378,N_22062);
nor U25504 (N_25504,N_22654,N_23174);
xor U25505 (N_25505,N_23169,N_22277);
and U25506 (N_25506,N_23633,N_23273);
and U25507 (N_25507,N_23335,N_22848);
nor U25508 (N_25508,N_23452,N_22277);
nor U25509 (N_25509,N_22218,N_23310);
nor U25510 (N_25510,N_22427,N_23076);
nand U25511 (N_25511,N_22827,N_22346);
or U25512 (N_25512,N_23458,N_22802);
or U25513 (N_25513,N_22342,N_23155);
xnor U25514 (N_25514,N_22729,N_22466);
or U25515 (N_25515,N_22427,N_23036);
nor U25516 (N_25516,N_22042,N_23956);
or U25517 (N_25517,N_22369,N_22354);
xor U25518 (N_25518,N_23771,N_22903);
nor U25519 (N_25519,N_23625,N_23374);
and U25520 (N_25520,N_23798,N_22595);
nor U25521 (N_25521,N_23225,N_23635);
nand U25522 (N_25522,N_23509,N_22061);
or U25523 (N_25523,N_23744,N_22662);
or U25524 (N_25524,N_22392,N_22733);
and U25525 (N_25525,N_23781,N_23739);
xnor U25526 (N_25526,N_22608,N_22227);
nand U25527 (N_25527,N_23321,N_22414);
or U25528 (N_25528,N_23525,N_23655);
or U25529 (N_25529,N_22245,N_23462);
and U25530 (N_25530,N_22344,N_22525);
and U25531 (N_25531,N_23654,N_22914);
nor U25532 (N_25532,N_22740,N_23878);
xnor U25533 (N_25533,N_23549,N_23038);
nor U25534 (N_25534,N_22833,N_22485);
and U25535 (N_25535,N_22841,N_22475);
or U25536 (N_25536,N_23781,N_22693);
nor U25537 (N_25537,N_23381,N_22619);
nand U25538 (N_25538,N_22190,N_23695);
and U25539 (N_25539,N_22037,N_22877);
xor U25540 (N_25540,N_23664,N_23279);
or U25541 (N_25541,N_22966,N_23663);
nor U25542 (N_25542,N_23763,N_23547);
and U25543 (N_25543,N_22412,N_23672);
and U25544 (N_25544,N_23505,N_23787);
nand U25545 (N_25545,N_23301,N_23716);
nand U25546 (N_25546,N_23667,N_22671);
and U25547 (N_25547,N_23380,N_23091);
nand U25548 (N_25548,N_23048,N_22076);
nor U25549 (N_25549,N_23480,N_23112);
and U25550 (N_25550,N_22176,N_22862);
nor U25551 (N_25551,N_22293,N_22414);
and U25552 (N_25552,N_22844,N_23016);
and U25553 (N_25553,N_22357,N_23413);
nor U25554 (N_25554,N_22794,N_23470);
and U25555 (N_25555,N_22533,N_23581);
xor U25556 (N_25556,N_22733,N_22560);
xnor U25557 (N_25557,N_22704,N_23499);
nor U25558 (N_25558,N_22938,N_23773);
and U25559 (N_25559,N_23942,N_22427);
or U25560 (N_25560,N_23624,N_23768);
nor U25561 (N_25561,N_22134,N_22722);
xor U25562 (N_25562,N_22408,N_22787);
nand U25563 (N_25563,N_22973,N_22355);
nor U25564 (N_25564,N_23781,N_22677);
or U25565 (N_25565,N_22237,N_23845);
nor U25566 (N_25566,N_22510,N_22950);
nor U25567 (N_25567,N_23693,N_23132);
nand U25568 (N_25568,N_23466,N_23040);
and U25569 (N_25569,N_23712,N_22445);
xnor U25570 (N_25570,N_22412,N_23357);
nor U25571 (N_25571,N_22040,N_23429);
xor U25572 (N_25572,N_23832,N_22369);
xnor U25573 (N_25573,N_22667,N_23477);
and U25574 (N_25574,N_23697,N_23171);
and U25575 (N_25575,N_22290,N_22116);
or U25576 (N_25576,N_22053,N_22132);
xnor U25577 (N_25577,N_23549,N_23233);
xnor U25578 (N_25578,N_22612,N_23419);
or U25579 (N_25579,N_22496,N_23805);
xnor U25580 (N_25580,N_23446,N_22076);
xor U25581 (N_25581,N_22123,N_22823);
xor U25582 (N_25582,N_23205,N_22890);
nor U25583 (N_25583,N_23791,N_22384);
or U25584 (N_25584,N_23249,N_23273);
and U25585 (N_25585,N_22834,N_23349);
xnor U25586 (N_25586,N_23670,N_22786);
nand U25587 (N_25587,N_23997,N_22614);
nand U25588 (N_25588,N_22511,N_23414);
nand U25589 (N_25589,N_22001,N_23200);
nand U25590 (N_25590,N_22378,N_22957);
xor U25591 (N_25591,N_23588,N_22912);
nor U25592 (N_25592,N_22866,N_22309);
nor U25593 (N_25593,N_22492,N_23886);
nand U25594 (N_25594,N_22279,N_22709);
or U25595 (N_25595,N_23714,N_22447);
nor U25596 (N_25596,N_22579,N_23531);
nor U25597 (N_25597,N_22101,N_23604);
nor U25598 (N_25598,N_23806,N_22030);
nor U25599 (N_25599,N_23215,N_23492);
nor U25600 (N_25600,N_22279,N_23558);
xnor U25601 (N_25601,N_23608,N_23217);
nor U25602 (N_25602,N_22822,N_22705);
xor U25603 (N_25603,N_22821,N_22055);
and U25604 (N_25604,N_23369,N_23966);
xor U25605 (N_25605,N_22183,N_22172);
or U25606 (N_25606,N_23170,N_22263);
xor U25607 (N_25607,N_23907,N_22836);
nor U25608 (N_25608,N_23172,N_23103);
nor U25609 (N_25609,N_22323,N_22253);
nand U25610 (N_25610,N_23988,N_23875);
xor U25611 (N_25611,N_22088,N_23744);
and U25612 (N_25612,N_23642,N_22933);
xor U25613 (N_25613,N_22202,N_22976);
nand U25614 (N_25614,N_23429,N_22991);
xnor U25615 (N_25615,N_22199,N_23215);
and U25616 (N_25616,N_22901,N_22279);
or U25617 (N_25617,N_22133,N_23149);
nand U25618 (N_25618,N_23859,N_22930);
nand U25619 (N_25619,N_22759,N_22764);
or U25620 (N_25620,N_23446,N_22810);
and U25621 (N_25621,N_22713,N_23334);
or U25622 (N_25622,N_23383,N_22829);
nor U25623 (N_25623,N_22140,N_22030);
xor U25624 (N_25624,N_23126,N_23434);
nor U25625 (N_25625,N_23279,N_23980);
or U25626 (N_25626,N_23617,N_23706);
nand U25627 (N_25627,N_23548,N_23490);
or U25628 (N_25628,N_22688,N_22947);
or U25629 (N_25629,N_22849,N_22969);
nand U25630 (N_25630,N_23786,N_23715);
xnor U25631 (N_25631,N_22163,N_23170);
nor U25632 (N_25632,N_23247,N_23533);
or U25633 (N_25633,N_23893,N_23200);
xnor U25634 (N_25634,N_23873,N_22270);
nand U25635 (N_25635,N_22036,N_23593);
or U25636 (N_25636,N_23598,N_23524);
and U25637 (N_25637,N_23049,N_22226);
nand U25638 (N_25638,N_22032,N_22899);
nand U25639 (N_25639,N_23610,N_23704);
nand U25640 (N_25640,N_23520,N_23153);
or U25641 (N_25641,N_22678,N_22200);
nor U25642 (N_25642,N_22564,N_23156);
and U25643 (N_25643,N_23649,N_23997);
xnor U25644 (N_25644,N_22985,N_23794);
or U25645 (N_25645,N_23944,N_23048);
nor U25646 (N_25646,N_22041,N_23543);
or U25647 (N_25647,N_23797,N_22353);
and U25648 (N_25648,N_23632,N_23117);
nand U25649 (N_25649,N_23399,N_22314);
or U25650 (N_25650,N_23507,N_23563);
nor U25651 (N_25651,N_23042,N_23258);
xor U25652 (N_25652,N_22418,N_23100);
and U25653 (N_25653,N_23493,N_23818);
nor U25654 (N_25654,N_22887,N_22034);
nand U25655 (N_25655,N_22710,N_22218);
or U25656 (N_25656,N_23443,N_23290);
xor U25657 (N_25657,N_22287,N_23273);
and U25658 (N_25658,N_22258,N_23045);
nor U25659 (N_25659,N_23444,N_23677);
xnor U25660 (N_25660,N_22456,N_23862);
or U25661 (N_25661,N_22854,N_23813);
nand U25662 (N_25662,N_22926,N_23853);
xnor U25663 (N_25663,N_22159,N_22371);
or U25664 (N_25664,N_22445,N_22496);
or U25665 (N_25665,N_22935,N_23703);
nand U25666 (N_25666,N_23730,N_23147);
or U25667 (N_25667,N_23041,N_23863);
xor U25668 (N_25668,N_23848,N_23908);
nand U25669 (N_25669,N_22333,N_22393);
nand U25670 (N_25670,N_23787,N_23125);
and U25671 (N_25671,N_22511,N_22376);
nor U25672 (N_25672,N_23595,N_22881);
or U25673 (N_25673,N_22478,N_22483);
or U25674 (N_25674,N_22390,N_23275);
xnor U25675 (N_25675,N_23868,N_22741);
nor U25676 (N_25676,N_22516,N_22369);
nor U25677 (N_25677,N_23936,N_22797);
nand U25678 (N_25678,N_23491,N_22853);
and U25679 (N_25679,N_23185,N_22233);
nand U25680 (N_25680,N_22795,N_23077);
nand U25681 (N_25681,N_22959,N_22465);
xnor U25682 (N_25682,N_22995,N_22590);
nor U25683 (N_25683,N_22563,N_22742);
nor U25684 (N_25684,N_22484,N_22661);
nor U25685 (N_25685,N_22929,N_22037);
and U25686 (N_25686,N_23555,N_22485);
xor U25687 (N_25687,N_23323,N_23119);
xor U25688 (N_25688,N_23421,N_23459);
xnor U25689 (N_25689,N_22516,N_23959);
xnor U25690 (N_25690,N_23459,N_22974);
or U25691 (N_25691,N_22649,N_23710);
or U25692 (N_25692,N_22782,N_22081);
and U25693 (N_25693,N_23920,N_22186);
or U25694 (N_25694,N_22130,N_22740);
nand U25695 (N_25695,N_23979,N_23165);
nor U25696 (N_25696,N_23531,N_22454);
nor U25697 (N_25697,N_22053,N_23458);
and U25698 (N_25698,N_22846,N_23889);
nor U25699 (N_25699,N_22444,N_22452);
nor U25700 (N_25700,N_23475,N_22264);
nor U25701 (N_25701,N_22581,N_22678);
xor U25702 (N_25702,N_23803,N_22162);
xor U25703 (N_25703,N_23503,N_22457);
and U25704 (N_25704,N_22030,N_23361);
nor U25705 (N_25705,N_22615,N_22141);
and U25706 (N_25706,N_23126,N_22068);
nor U25707 (N_25707,N_22728,N_22420);
nor U25708 (N_25708,N_23171,N_22164);
nor U25709 (N_25709,N_23624,N_23498);
nand U25710 (N_25710,N_23191,N_22917);
xnor U25711 (N_25711,N_23507,N_23899);
nand U25712 (N_25712,N_23763,N_22386);
nor U25713 (N_25713,N_23569,N_22600);
and U25714 (N_25714,N_23297,N_23146);
nor U25715 (N_25715,N_23643,N_22283);
and U25716 (N_25716,N_22339,N_23037);
and U25717 (N_25717,N_22474,N_22057);
nand U25718 (N_25718,N_23172,N_23159);
or U25719 (N_25719,N_23384,N_23940);
and U25720 (N_25720,N_23438,N_22647);
or U25721 (N_25721,N_22540,N_22291);
xor U25722 (N_25722,N_23289,N_22397);
xnor U25723 (N_25723,N_22223,N_23978);
and U25724 (N_25724,N_22547,N_22587);
and U25725 (N_25725,N_23421,N_22295);
nand U25726 (N_25726,N_23199,N_23891);
and U25727 (N_25727,N_23838,N_22213);
xnor U25728 (N_25728,N_22920,N_22547);
nor U25729 (N_25729,N_22733,N_23610);
and U25730 (N_25730,N_22961,N_23746);
nor U25731 (N_25731,N_22564,N_23519);
or U25732 (N_25732,N_22379,N_22910);
and U25733 (N_25733,N_22278,N_22801);
or U25734 (N_25734,N_22552,N_23029);
xnor U25735 (N_25735,N_23277,N_23771);
and U25736 (N_25736,N_23428,N_23894);
and U25737 (N_25737,N_23112,N_22455);
and U25738 (N_25738,N_23270,N_22458);
xnor U25739 (N_25739,N_22363,N_22229);
nand U25740 (N_25740,N_23316,N_22174);
xor U25741 (N_25741,N_22571,N_22807);
or U25742 (N_25742,N_23145,N_22032);
xnor U25743 (N_25743,N_23526,N_22923);
nor U25744 (N_25744,N_22743,N_22594);
nor U25745 (N_25745,N_22445,N_22069);
nor U25746 (N_25746,N_22468,N_23612);
or U25747 (N_25747,N_22962,N_23687);
or U25748 (N_25748,N_23652,N_23823);
nor U25749 (N_25749,N_22008,N_22175);
or U25750 (N_25750,N_23955,N_23319);
xnor U25751 (N_25751,N_23368,N_22651);
and U25752 (N_25752,N_22983,N_23043);
and U25753 (N_25753,N_22647,N_22580);
nand U25754 (N_25754,N_23666,N_23102);
xnor U25755 (N_25755,N_23872,N_23189);
nor U25756 (N_25756,N_23250,N_23120);
xor U25757 (N_25757,N_22300,N_22880);
or U25758 (N_25758,N_22885,N_23699);
nand U25759 (N_25759,N_23706,N_23012);
nor U25760 (N_25760,N_22738,N_22748);
and U25761 (N_25761,N_23270,N_23088);
nor U25762 (N_25762,N_23069,N_23621);
nand U25763 (N_25763,N_23963,N_22913);
nor U25764 (N_25764,N_22895,N_23020);
or U25765 (N_25765,N_22219,N_23746);
or U25766 (N_25766,N_22802,N_23100);
or U25767 (N_25767,N_22975,N_23160);
nor U25768 (N_25768,N_23048,N_22728);
nand U25769 (N_25769,N_23206,N_23686);
xor U25770 (N_25770,N_22953,N_23194);
or U25771 (N_25771,N_22635,N_23448);
nor U25772 (N_25772,N_23290,N_23045);
nor U25773 (N_25773,N_22429,N_22326);
nand U25774 (N_25774,N_22036,N_22587);
nand U25775 (N_25775,N_23429,N_23761);
nand U25776 (N_25776,N_23952,N_22830);
nor U25777 (N_25777,N_22958,N_22532);
nand U25778 (N_25778,N_23192,N_23892);
nand U25779 (N_25779,N_23960,N_23059);
nor U25780 (N_25780,N_23671,N_23962);
or U25781 (N_25781,N_23792,N_23815);
nor U25782 (N_25782,N_23326,N_22486);
nand U25783 (N_25783,N_23940,N_22887);
or U25784 (N_25784,N_22105,N_23093);
nand U25785 (N_25785,N_23010,N_22821);
or U25786 (N_25786,N_22342,N_22393);
or U25787 (N_25787,N_22741,N_22116);
and U25788 (N_25788,N_22380,N_22930);
nand U25789 (N_25789,N_23928,N_23309);
and U25790 (N_25790,N_22088,N_22462);
nor U25791 (N_25791,N_23628,N_23914);
and U25792 (N_25792,N_23108,N_23208);
and U25793 (N_25793,N_23321,N_22099);
xnor U25794 (N_25794,N_22203,N_23842);
or U25795 (N_25795,N_23970,N_22018);
and U25796 (N_25796,N_22674,N_23099);
and U25797 (N_25797,N_23268,N_22414);
or U25798 (N_25798,N_23128,N_23191);
xnor U25799 (N_25799,N_23902,N_22941);
or U25800 (N_25800,N_22902,N_22102);
xor U25801 (N_25801,N_23799,N_23741);
and U25802 (N_25802,N_22541,N_23290);
xor U25803 (N_25803,N_23089,N_23879);
nand U25804 (N_25804,N_22558,N_23985);
or U25805 (N_25805,N_22162,N_23681);
nor U25806 (N_25806,N_22716,N_22175);
xnor U25807 (N_25807,N_23083,N_22888);
nand U25808 (N_25808,N_22437,N_22440);
nand U25809 (N_25809,N_23886,N_23685);
nand U25810 (N_25810,N_23415,N_22784);
xor U25811 (N_25811,N_23996,N_22817);
xor U25812 (N_25812,N_22844,N_22416);
and U25813 (N_25813,N_23142,N_23904);
and U25814 (N_25814,N_23662,N_23794);
xnor U25815 (N_25815,N_22175,N_23215);
or U25816 (N_25816,N_23546,N_22373);
nand U25817 (N_25817,N_22119,N_23079);
nand U25818 (N_25818,N_23773,N_23096);
xor U25819 (N_25819,N_22529,N_23899);
nand U25820 (N_25820,N_23463,N_22657);
and U25821 (N_25821,N_22475,N_23353);
nor U25822 (N_25822,N_22353,N_22555);
nand U25823 (N_25823,N_22686,N_23120);
xor U25824 (N_25824,N_23927,N_23692);
nand U25825 (N_25825,N_22763,N_22564);
xnor U25826 (N_25826,N_23908,N_23429);
xnor U25827 (N_25827,N_23341,N_23693);
or U25828 (N_25828,N_23556,N_23516);
and U25829 (N_25829,N_23408,N_22836);
or U25830 (N_25830,N_23380,N_22228);
xnor U25831 (N_25831,N_23017,N_22200);
or U25832 (N_25832,N_22994,N_23522);
or U25833 (N_25833,N_23930,N_22885);
xor U25834 (N_25834,N_23613,N_23528);
nor U25835 (N_25835,N_22862,N_22544);
nand U25836 (N_25836,N_23031,N_23109);
and U25837 (N_25837,N_22734,N_23690);
or U25838 (N_25838,N_23582,N_22066);
xnor U25839 (N_25839,N_22551,N_22174);
nor U25840 (N_25840,N_22541,N_23690);
and U25841 (N_25841,N_23607,N_23793);
nand U25842 (N_25842,N_22018,N_22310);
xor U25843 (N_25843,N_23223,N_23990);
and U25844 (N_25844,N_22464,N_22208);
and U25845 (N_25845,N_22220,N_23908);
xor U25846 (N_25846,N_22631,N_22349);
nor U25847 (N_25847,N_23007,N_23277);
nand U25848 (N_25848,N_23943,N_23177);
nor U25849 (N_25849,N_23147,N_22615);
xnor U25850 (N_25850,N_22812,N_23497);
or U25851 (N_25851,N_22529,N_22824);
nand U25852 (N_25852,N_23416,N_23585);
nand U25853 (N_25853,N_23639,N_23524);
and U25854 (N_25854,N_22867,N_23544);
and U25855 (N_25855,N_22014,N_22560);
nor U25856 (N_25856,N_23779,N_22403);
and U25857 (N_25857,N_22720,N_23703);
xnor U25858 (N_25858,N_23175,N_22479);
nor U25859 (N_25859,N_23536,N_23236);
xor U25860 (N_25860,N_23625,N_23400);
xnor U25861 (N_25861,N_23435,N_23244);
nor U25862 (N_25862,N_22599,N_22279);
xnor U25863 (N_25863,N_23868,N_23431);
xor U25864 (N_25864,N_22876,N_22875);
and U25865 (N_25865,N_23923,N_22225);
nand U25866 (N_25866,N_23072,N_23001);
and U25867 (N_25867,N_23122,N_23952);
nor U25868 (N_25868,N_22422,N_22649);
nor U25869 (N_25869,N_22708,N_22097);
nor U25870 (N_25870,N_23924,N_22309);
and U25871 (N_25871,N_23823,N_22596);
and U25872 (N_25872,N_23432,N_23269);
or U25873 (N_25873,N_23292,N_22427);
nand U25874 (N_25874,N_22345,N_22179);
or U25875 (N_25875,N_23304,N_23764);
or U25876 (N_25876,N_23290,N_23062);
or U25877 (N_25877,N_23110,N_22534);
xor U25878 (N_25878,N_22577,N_23146);
xnor U25879 (N_25879,N_23277,N_22291);
and U25880 (N_25880,N_22771,N_23107);
xnor U25881 (N_25881,N_23204,N_22603);
or U25882 (N_25882,N_22914,N_22612);
and U25883 (N_25883,N_23725,N_22654);
xnor U25884 (N_25884,N_23709,N_22460);
or U25885 (N_25885,N_23767,N_23969);
xnor U25886 (N_25886,N_23971,N_22343);
nor U25887 (N_25887,N_23835,N_23633);
and U25888 (N_25888,N_22941,N_22452);
nor U25889 (N_25889,N_23236,N_23370);
nand U25890 (N_25890,N_23180,N_22840);
nor U25891 (N_25891,N_23195,N_23016);
or U25892 (N_25892,N_22922,N_23246);
or U25893 (N_25893,N_23594,N_22524);
nand U25894 (N_25894,N_22155,N_22470);
or U25895 (N_25895,N_22444,N_23305);
nand U25896 (N_25896,N_22380,N_22158);
and U25897 (N_25897,N_23797,N_23438);
or U25898 (N_25898,N_22596,N_23098);
nand U25899 (N_25899,N_22961,N_23196);
xor U25900 (N_25900,N_23515,N_23490);
nor U25901 (N_25901,N_22510,N_23035);
or U25902 (N_25902,N_23761,N_23598);
nor U25903 (N_25903,N_22331,N_22309);
or U25904 (N_25904,N_23957,N_23829);
or U25905 (N_25905,N_23713,N_23850);
xor U25906 (N_25906,N_23402,N_22571);
and U25907 (N_25907,N_22128,N_23414);
nand U25908 (N_25908,N_22204,N_23542);
nor U25909 (N_25909,N_23234,N_23946);
nor U25910 (N_25910,N_22743,N_22387);
or U25911 (N_25911,N_22744,N_22032);
or U25912 (N_25912,N_22392,N_22588);
and U25913 (N_25913,N_23225,N_23662);
nor U25914 (N_25914,N_23756,N_22638);
xnor U25915 (N_25915,N_22040,N_22985);
xnor U25916 (N_25916,N_23543,N_22289);
and U25917 (N_25917,N_22312,N_22980);
nand U25918 (N_25918,N_23538,N_23887);
xnor U25919 (N_25919,N_22834,N_22127);
xnor U25920 (N_25920,N_22523,N_22774);
nor U25921 (N_25921,N_22392,N_23305);
nand U25922 (N_25922,N_22554,N_23340);
and U25923 (N_25923,N_22261,N_22882);
and U25924 (N_25924,N_23310,N_22835);
xnor U25925 (N_25925,N_23954,N_23847);
xnor U25926 (N_25926,N_22938,N_22919);
nor U25927 (N_25927,N_22045,N_23457);
and U25928 (N_25928,N_23616,N_22426);
and U25929 (N_25929,N_22916,N_22261);
nor U25930 (N_25930,N_22557,N_22708);
xor U25931 (N_25931,N_22586,N_23555);
xor U25932 (N_25932,N_22211,N_23877);
xor U25933 (N_25933,N_22092,N_23713);
nand U25934 (N_25934,N_22849,N_22429);
or U25935 (N_25935,N_23382,N_23200);
or U25936 (N_25936,N_22434,N_22862);
and U25937 (N_25937,N_23836,N_23724);
and U25938 (N_25938,N_22333,N_23436);
nand U25939 (N_25939,N_23630,N_22204);
nor U25940 (N_25940,N_23127,N_22541);
xor U25941 (N_25941,N_22222,N_23959);
nand U25942 (N_25942,N_22664,N_22621);
nand U25943 (N_25943,N_22321,N_22582);
or U25944 (N_25944,N_22549,N_23816);
or U25945 (N_25945,N_22108,N_23997);
and U25946 (N_25946,N_22687,N_23517);
nand U25947 (N_25947,N_22660,N_22782);
or U25948 (N_25948,N_23712,N_23599);
nor U25949 (N_25949,N_23629,N_23357);
or U25950 (N_25950,N_23019,N_22941);
xor U25951 (N_25951,N_23780,N_23764);
and U25952 (N_25952,N_22421,N_23550);
and U25953 (N_25953,N_23506,N_23301);
nor U25954 (N_25954,N_23312,N_23631);
or U25955 (N_25955,N_23787,N_22575);
and U25956 (N_25956,N_22050,N_22665);
and U25957 (N_25957,N_22519,N_22932);
xnor U25958 (N_25958,N_23644,N_22295);
nand U25959 (N_25959,N_23583,N_23627);
nand U25960 (N_25960,N_22569,N_23090);
nand U25961 (N_25961,N_22808,N_23423);
nand U25962 (N_25962,N_23035,N_22911);
and U25963 (N_25963,N_23464,N_23403);
or U25964 (N_25964,N_22126,N_23643);
xor U25965 (N_25965,N_22464,N_23719);
nor U25966 (N_25966,N_23272,N_23991);
nand U25967 (N_25967,N_23830,N_22641);
or U25968 (N_25968,N_23259,N_23984);
and U25969 (N_25969,N_23112,N_23651);
and U25970 (N_25970,N_23388,N_22353);
xor U25971 (N_25971,N_23751,N_23048);
nand U25972 (N_25972,N_22642,N_22083);
nor U25973 (N_25973,N_22297,N_22113);
xor U25974 (N_25974,N_23758,N_23947);
nand U25975 (N_25975,N_22877,N_22413);
nor U25976 (N_25976,N_23748,N_22396);
nand U25977 (N_25977,N_22776,N_23936);
nor U25978 (N_25978,N_23043,N_23699);
or U25979 (N_25979,N_22069,N_22580);
nand U25980 (N_25980,N_22557,N_22462);
and U25981 (N_25981,N_23104,N_22666);
and U25982 (N_25982,N_23222,N_23288);
or U25983 (N_25983,N_23986,N_22203);
or U25984 (N_25984,N_22135,N_22213);
xnor U25985 (N_25985,N_23729,N_23607);
and U25986 (N_25986,N_22383,N_23014);
nor U25987 (N_25987,N_22619,N_23335);
and U25988 (N_25988,N_23418,N_23469);
or U25989 (N_25989,N_23780,N_22636);
nor U25990 (N_25990,N_23592,N_23961);
nand U25991 (N_25991,N_23281,N_22264);
or U25992 (N_25992,N_22017,N_22205);
nand U25993 (N_25993,N_23739,N_22470);
nand U25994 (N_25994,N_23043,N_22391);
xor U25995 (N_25995,N_23809,N_22917);
and U25996 (N_25996,N_23998,N_23679);
nand U25997 (N_25997,N_23523,N_22609);
nor U25998 (N_25998,N_23462,N_23178);
nand U25999 (N_25999,N_23904,N_22903);
nand U26000 (N_26000,N_25895,N_24084);
and U26001 (N_26001,N_24381,N_24247);
nand U26002 (N_26002,N_25939,N_24779);
or U26003 (N_26003,N_24044,N_24821);
or U26004 (N_26004,N_24968,N_25248);
nand U26005 (N_26005,N_25308,N_24875);
nor U26006 (N_26006,N_24752,N_24976);
xnor U26007 (N_26007,N_25888,N_25622);
and U26008 (N_26008,N_24059,N_24804);
nand U26009 (N_26009,N_24304,N_24495);
xor U26010 (N_26010,N_25788,N_25272);
nor U26011 (N_26011,N_24532,N_25207);
nor U26012 (N_26012,N_24945,N_25245);
nand U26013 (N_26013,N_24023,N_25063);
and U26014 (N_26014,N_24481,N_24172);
and U26015 (N_26015,N_24053,N_25341);
nor U26016 (N_26016,N_25246,N_25140);
and U26017 (N_26017,N_25877,N_25154);
xor U26018 (N_26018,N_25972,N_24423);
and U26019 (N_26019,N_24042,N_24336);
and U26020 (N_26020,N_24215,N_24556);
nand U26021 (N_26021,N_25813,N_24065);
and U26022 (N_26022,N_24249,N_25894);
and U26023 (N_26023,N_25242,N_24462);
nand U26024 (N_26024,N_24896,N_24045);
xor U26025 (N_26025,N_24699,N_24911);
and U26026 (N_26026,N_25374,N_24468);
or U26027 (N_26027,N_24591,N_25179);
xor U26028 (N_26028,N_25700,N_25468);
and U26029 (N_26029,N_25824,N_24238);
xor U26030 (N_26030,N_24000,N_25965);
xor U26031 (N_26031,N_24349,N_24973);
xor U26032 (N_26032,N_25137,N_25748);
nor U26033 (N_26033,N_24636,N_24576);
nand U26034 (N_26034,N_24110,N_25003);
nand U26035 (N_26035,N_25194,N_25952);
or U26036 (N_26036,N_24477,N_24877);
nand U26037 (N_26037,N_25318,N_25950);
and U26038 (N_26038,N_24957,N_25172);
nand U26039 (N_26039,N_24118,N_24817);
xor U26040 (N_26040,N_24143,N_24288);
or U26041 (N_26041,N_24565,N_25408);
or U26042 (N_26042,N_24054,N_25812);
xor U26043 (N_26043,N_25378,N_24027);
xor U26044 (N_26044,N_25274,N_24775);
and U26045 (N_26045,N_24994,N_24297);
and U26046 (N_26046,N_25560,N_25492);
or U26047 (N_26047,N_24242,N_24272);
nor U26048 (N_26048,N_25232,N_24421);
or U26049 (N_26049,N_24222,N_24912);
and U26050 (N_26050,N_24353,N_24454);
nand U26051 (N_26051,N_24327,N_25552);
nor U26052 (N_26052,N_25696,N_24245);
nor U26053 (N_26053,N_24868,N_25897);
nand U26054 (N_26054,N_25605,N_24796);
or U26055 (N_26055,N_24497,N_25837);
nand U26056 (N_26056,N_25496,N_24401);
nor U26057 (N_26057,N_25528,N_25798);
nor U26058 (N_26058,N_24315,N_25025);
or U26059 (N_26059,N_24364,N_24560);
nor U26060 (N_26060,N_24290,N_25280);
nor U26061 (N_26061,N_24313,N_24774);
nor U26062 (N_26062,N_25311,N_24355);
nor U26063 (N_26063,N_24900,N_24492);
and U26064 (N_26064,N_25505,N_24447);
nand U26065 (N_26065,N_24660,N_25808);
nor U26066 (N_26066,N_24433,N_25029);
xor U26067 (N_26067,N_24521,N_24538);
nor U26068 (N_26068,N_25431,N_24233);
xnor U26069 (N_26069,N_25577,N_24548);
nand U26070 (N_26070,N_24001,N_25754);
and U26071 (N_26071,N_24320,N_24663);
nand U26072 (N_26072,N_24891,N_25987);
and U26073 (N_26073,N_24880,N_24882);
or U26074 (N_26074,N_24700,N_24596);
and U26075 (N_26075,N_24756,N_24113);
xor U26076 (N_26076,N_25529,N_25678);
nor U26077 (N_26077,N_24995,N_24115);
or U26078 (N_26078,N_24562,N_25352);
nand U26079 (N_26079,N_25976,N_24087);
or U26080 (N_26080,N_25629,N_24724);
nand U26081 (N_26081,N_24024,N_24645);
nand U26082 (N_26082,N_24279,N_25327);
nand U26083 (N_26083,N_25466,N_25065);
xor U26084 (N_26084,N_25344,N_24204);
xor U26085 (N_26085,N_25009,N_24936);
xor U26086 (N_26086,N_24533,N_24043);
and U26087 (N_26087,N_25933,N_25078);
xor U26088 (N_26088,N_24793,N_24013);
or U26089 (N_26089,N_24750,N_24616);
and U26090 (N_26090,N_25185,N_24838);
nor U26091 (N_26091,N_24284,N_25237);
and U26092 (N_26092,N_25347,N_25136);
and U26093 (N_26093,N_24913,N_24126);
nor U26094 (N_26094,N_25410,N_24971);
or U26095 (N_26095,N_24039,N_25845);
and U26096 (N_26096,N_25642,N_24346);
and U26097 (N_26097,N_24081,N_24622);
or U26098 (N_26098,N_25566,N_24934);
or U26099 (N_26099,N_25204,N_24812);
and U26100 (N_26100,N_25259,N_24317);
and U26101 (N_26101,N_25491,N_25217);
xor U26102 (N_26102,N_24862,N_24780);
or U26103 (N_26103,N_24630,N_24524);
xor U26104 (N_26104,N_25380,N_24642);
and U26105 (N_26105,N_24685,N_25797);
and U26106 (N_26106,N_25525,N_24374);
xor U26107 (N_26107,N_25776,N_24834);
nand U26108 (N_26108,N_24595,N_25196);
xnor U26109 (N_26109,N_24324,N_25361);
nor U26110 (N_26110,N_25931,N_25511);
xnor U26111 (N_26111,N_24707,N_24475);
nand U26112 (N_26112,N_24487,N_24785);
and U26113 (N_26113,N_24240,N_25129);
nand U26114 (N_26114,N_24369,N_24399);
nand U26115 (N_26115,N_24020,N_24382);
xnor U26116 (N_26116,N_24637,N_25707);
nand U26117 (N_26117,N_24716,N_25602);
nand U26118 (N_26118,N_25085,N_25630);
nor U26119 (N_26119,N_24618,N_25606);
nand U26120 (N_26120,N_24530,N_24305);
nor U26121 (N_26121,N_25626,N_24568);
nand U26122 (N_26122,N_25550,N_25148);
or U26123 (N_26123,N_24255,N_24450);
xnor U26124 (N_26124,N_25252,N_25114);
and U26125 (N_26125,N_25222,N_24489);
nor U26126 (N_26126,N_24280,N_25044);
nor U26127 (N_26127,N_25639,N_24131);
nor U26128 (N_26128,N_25039,N_24795);
nand U26129 (N_26129,N_24907,N_24308);
or U26130 (N_26130,N_25268,N_24014);
nand U26131 (N_26131,N_25495,N_25617);
or U26132 (N_26132,N_25831,N_24747);
nor U26133 (N_26133,N_24544,N_25498);
and U26134 (N_26134,N_24153,N_25735);
or U26135 (N_26135,N_25985,N_25178);
nand U26136 (N_26136,N_25163,N_24649);
nor U26137 (N_26137,N_24947,N_25005);
or U26138 (N_26138,N_25390,N_24119);
nor U26139 (N_26139,N_25142,N_25135);
nand U26140 (N_26140,N_25317,N_24593);
nor U26141 (N_26141,N_24004,N_24250);
nor U26142 (N_26142,N_25239,N_24669);
xor U26143 (N_26143,N_24212,N_25458);
xnor U26144 (N_26144,N_24982,N_25561);
or U26145 (N_26145,N_25184,N_25255);
or U26146 (N_26146,N_24211,N_25611);
xnor U26147 (N_26147,N_24107,N_24347);
or U26148 (N_26148,N_25806,N_25388);
nand U26149 (N_26149,N_24389,N_24564);
nand U26150 (N_26150,N_24363,N_25227);
and U26151 (N_26151,N_24810,N_25929);
xor U26152 (N_26152,N_24464,N_24186);
nor U26153 (N_26153,N_25143,N_25333);
or U26154 (N_26154,N_24155,N_24070);
or U26155 (N_26155,N_25126,N_24469);
and U26156 (N_26156,N_24999,N_24935);
nand U26157 (N_26157,N_25462,N_24668);
and U26158 (N_26158,N_25102,N_24169);
xnor U26159 (N_26159,N_24848,N_24268);
nand U26160 (N_26160,N_25805,N_24960);
nor U26161 (N_26161,N_24439,N_25067);
nand U26162 (N_26162,N_24323,N_25998);
nand U26163 (N_26163,N_25463,N_24986);
or U26164 (N_26164,N_25166,N_25192);
xor U26165 (N_26165,N_25328,N_25307);
nand U26166 (N_26166,N_24626,N_24015);
nor U26167 (N_26167,N_25835,N_25319);
nor U26168 (N_26168,N_25923,N_24712);
nor U26169 (N_26169,N_24166,N_25963);
nor U26170 (N_26170,N_24078,N_24152);
xnor U26171 (N_26171,N_24306,N_25335);
nor U26172 (N_26172,N_25337,N_24176);
and U26173 (N_26173,N_25524,N_24441);
or U26174 (N_26174,N_25077,N_24377);
xor U26175 (N_26175,N_25910,N_24102);
nand U26176 (N_26176,N_25241,N_24016);
xnor U26177 (N_26177,N_24444,N_24763);
or U26178 (N_26178,N_25989,N_24585);
or U26179 (N_26179,N_25489,N_25718);
xor U26180 (N_26180,N_25594,N_24011);
or U26181 (N_26181,N_24844,N_24525);
and U26182 (N_26182,N_24594,N_25784);
xor U26183 (N_26183,N_25739,N_24683);
or U26184 (N_26184,N_24270,N_25969);
xor U26185 (N_26185,N_24569,N_24792);
xor U26186 (N_26186,N_24566,N_25325);
and U26187 (N_26187,N_25761,N_25116);
xor U26188 (N_26188,N_25714,N_24640);
or U26189 (N_26189,N_25072,N_24436);
or U26190 (N_26190,N_25330,N_25257);
nor U26191 (N_26191,N_24002,N_24652);
xnor U26192 (N_26192,N_24767,N_24979);
and U26193 (N_26193,N_25370,N_25690);
nor U26194 (N_26194,N_24460,N_24856);
xor U26195 (N_26195,N_24728,N_24607);
nand U26196 (N_26196,N_24772,N_25467);
nand U26197 (N_26197,N_24701,N_25814);
nor U26198 (N_26198,N_24170,N_25850);
or U26199 (N_26199,N_25375,N_25609);
nand U26200 (N_26200,N_25663,N_25538);
and U26201 (N_26201,N_24650,N_25225);
and U26202 (N_26202,N_24505,N_24356);
or U26203 (N_26203,N_24326,N_24582);
nand U26204 (N_26204,N_24943,N_24855);
and U26205 (N_26205,N_25915,N_24427);
xor U26206 (N_26206,N_24851,N_24758);
nor U26207 (N_26207,N_25269,N_24037);
xor U26208 (N_26208,N_24828,N_24406);
nand U26209 (N_26209,N_25656,N_24952);
xnor U26210 (N_26210,N_25113,N_24151);
xnor U26211 (N_26211,N_24679,N_24402);
nand U26212 (N_26212,N_25559,N_25381);
or U26213 (N_26213,N_25454,N_25809);
and U26214 (N_26214,N_25376,N_24908);
nand U26215 (N_26215,N_25180,N_24335);
xnor U26216 (N_26216,N_25612,N_24511);
nand U26217 (N_26217,N_25900,N_25125);
nor U26218 (N_26218,N_24930,N_25093);
nor U26219 (N_26219,N_25292,N_25149);
nand U26220 (N_26220,N_24062,N_24634);
or U26221 (N_26221,N_25296,N_24412);
nor U26222 (N_26222,N_25816,N_25913);
or U26223 (N_26223,N_25428,N_24905);
or U26224 (N_26224,N_24112,N_24442);
nand U26225 (N_26225,N_24416,N_25437);
nor U26226 (N_26226,N_25916,N_24476);
xor U26227 (N_26227,N_24019,N_24512);
or U26228 (N_26228,N_25421,N_25710);
nor U26229 (N_26229,N_25956,N_24127);
and U26230 (N_26230,N_25397,N_25064);
nor U26231 (N_26231,N_25434,N_25018);
or U26232 (N_26232,N_24414,N_25017);
nor U26233 (N_26233,N_25951,N_25726);
nand U26234 (N_26234,N_24061,N_25023);
xnor U26235 (N_26235,N_25088,N_24498);
nor U26236 (N_26236,N_25389,N_25062);
nor U26237 (N_26237,N_25342,N_25363);
or U26238 (N_26238,N_25106,N_24185);
xnor U26239 (N_26239,N_24052,N_24098);
and U26240 (N_26240,N_24354,N_25298);
xor U26241 (N_26241,N_25999,N_25262);
nor U26242 (N_26242,N_25980,N_25219);
nand U26243 (N_26243,N_24285,N_25476);
or U26244 (N_26244,N_25264,N_25068);
and U26245 (N_26245,N_24437,N_25941);
xnor U26246 (N_26246,N_24064,N_24182);
xor U26247 (N_26247,N_24651,N_24967);
nand U26248 (N_26248,N_25815,N_25619);
nand U26249 (N_26249,N_25351,N_25155);
xor U26250 (N_26250,N_24195,N_24309);
and U26251 (N_26251,N_24673,N_24730);
and U26252 (N_26252,N_25087,N_24220);
nor U26253 (N_26253,N_24299,N_25182);
xnor U26254 (N_26254,N_24551,N_24040);
and U26255 (N_26255,N_24643,N_25984);
xnor U26256 (N_26256,N_24571,N_24573);
and U26257 (N_26257,N_25305,N_25213);
nand U26258 (N_26258,N_25562,N_25852);
and U26259 (N_26259,N_25066,N_25299);
or U26260 (N_26260,N_24764,N_24429);
nand U26261 (N_26261,N_25478,N_24262);
and U26262 (N_26262,N_24431,N_24760);
and U26263 (N_26263,N_24937,N_25756);
xor U26264 (N_26264,N_24214,N_25653);
xnor U26265 (N_26265,N_25302,N_24748);
nand U26266 (N_26266,N_25127,N_25197);
nor U26267 (N_26267,N_25287,N_25953);
and U26268 (N_26268,N_25654,N_25418);
and U26269 (N_26269,N_25392,N_24659);
nor U26270 (N_26270,N_24101,N_25345);
nor U26271 (N_26271,N_24430,N_24587);
nand U26272 (N_26272,N_24733,N_24738);
nand U26273 (N_26273,N_25395,N_25975);
and U26274 (N_26274,N_25481,N_24762);
nand U26275 (N_26275,N_25506,N_25230);
nor U26276 (N_26276,N_24675,N_24311);
xnor U26277 (N_26277,N_24410,N_24149);
xnor U26278 (N_26278,N_25535,N_24395);
and U26279 (N_26279,N_24588,N_25387);
or U26280 (N_26280,N_24623,N_24619);
nor U26281 (N_26281,N_24067,N_24422);
or U26282 (N_26282,N_24765,N_25156);
nor U26283 (N_26283,N_24403,N_24373);
xor U26284 (N_26284,N_25541,N_24895);
and U26285 (N_26285,N_25668,N_25384);
and U26286 (N_26286,N_25310,N_25445);
and U26287 (N_26287,N_24134,N_24835);
or U26288 (N_26288,N_24229,N_24372);
nor U26289 (N_26289,N_24289,N_25666);
or U26290 (N_26290,N_25260,N_25021);
and U26291 (N_26291,N_24889,N_25537);
xor U26292 (N_26292,N_24193,N_24578);
and U26293 (N_26293,N_25157,N_24682);
or U26294 (N_26294,N_24209,N_24876);
nor U26295 (N_26295,N_25205,N_25024);
nand U26296 (N_26296,N_25743,N_25847);
or U26297 (N_26297,N_25719,N_24869);
and U26298 (N_26298,N_24150,N_25680);
or U26299 (N_26299,N_25540,N_25867);
nor U26300 (N_26300,N_24671,N_25440);
or U26301 (N_26301,N_25176,N_25215);
xor U26302 (N_26302,N_25443,N_24329);
and U26303 (N_26303,N_24041,N_25636);
nor U26304 (N_26304,N_24513,N_25669);
or U26305 (N_26305,N_24114,N_24605);
xnor U26306 (N_26306,N_25439,N_24391);
and U26307 (N_26307,N_25919,N_25794);
or U26308 (N_26308,N_24488,N_24225);
nor U26309 (N_26309,N_24096,N_24567);
nor U26310 (N_26310,N_25322,N_25187);
nor U26311 (N_26311,N_25638,N_24598);
nand U26312 (N_26312,N_25240,N_25997);
xnor U26313 (N_26313,N_24358,N_24163);
nand U26314 (N_26314,N_24165,N_25134);
nor U26315 (N_26315,N_24853,N_25061);
or U26316 (N_26316,N_25303,N_24589);
nor U26317 (N_26317,N_25927,N_25493);
and U26318 (N_26318,N_25047,N_24337);
xor U26319 (N_26319,N_24390,N_24946);
and U26320 (N_26320,N_25879,N_24864);
nand U26321 (N_26321,N_24725,N_25214);
and U26322 (N_26322,N_25405,N_24648);
and U26323 (N_26323,N_24520,N_24333);
and U26324 (N_26324,N_25357,N_24731);
or U26325 (N_26325,N_24552,N_25403);
xor U26326 (N_26326,N_24610,N_24580);
nand U26327 (N_26327,N_24319,N_24539);
nor U26328 (N_26328,N_25071,N_25684);
and U26329 (N_26329,N_25667,N_24926);
nand U26330 (N_26330,N_24396,N_24987);
and U26331 (N_26331,N_25741,N_24426);
and U26332 (N_26332,N_25682,N_25730);
xnor U26333 (N_26333,N_24639,N_25243);
nor U26334 (N_26334,N_24802,N_24997);
nand U26335 (N_26335,N_24076,N_25278);
nand U26336 (N_26336,N_24768,N_24375);
nor U26337 (N_26337,N_25253,N_25271);
and U26338 (N_26338,N_25247,N_25946);
and U26339 (N_26339,N_24196,N_25530);
nor U26340 (N_26340,N_24890,N_24108);
nand U26341 (N_26341,N_25470,N_25206);
nor U26342 (N_26342,N_24490,N_24226);
and U26343 (N_26343,N_24665,N_24507);
or U26344 (N_26344,N_25261,N_24867);
or U26345 (N_26345,N_24583,N_25059);
xor U26346 (N_26346,N_25050,N_24345);
xnor U26347 (N_26347,N_24074,N_25738);
or U26348 (N_26348,N_25613,N_25258);
nor U26349 (N_26349,N_25881,N_25935);
xor U26350 (N_26350,N_24380,N_24807);
and U26351 (N_26351,N_25717,N_24627);
nor U26352 (N_26352,N_25692,N_25886);
or U26353 (N_26353,N_25709,N_24722);
nor U26354 (N_26354,N_25169,N_25429);
or U26355 (N_26355,N_25882,N_25906);
nand U26356 (N_26356,N_24811,N_24068);
xor U26357 (N_26357,N_24504,N_24717);
and U26358 (N_26358,N_24252,N_24388);
nor U26359 (N_26359,N_25460,N_25905);
xnor U26360 (N_26360,N_25315,N_24048);
xor U26361 (N_26361,N_25829,N_25548);
or U26362 (N_26362,N_25645,N_25507);
or U26363 (N_26363,N_25627,N_25546);
and U26364 (N_26364,N_25358,N_24090);
xnor U26365 (N_26365,N_24342,N_25751);
xor U26366 (N_26366,N_25851,N_24428);
nand U26367 (N_26367,N_25160,N_25819);
nor U26368 (N_26368,N_25990,N_24711);
or U26369 (N_26369,N_25728,N_24473);
xnor U26370 (N_26370,N_24137,N_25830);
or U26371 (N_26371,N_25008,N_25041);
nand U26372 (N_26372,N_24813,N_24620);
or U26373 (N_26373,N_25796,N_25393);
xnor U26374 (N_26374,N_24357,N_24534);
xor U26375 (N_26375,N_24678,N_25516);
or U26376 (N_26376,N_25949,N_24897);
and U26377 (N_26377,N_24254,N_24094);
nand U26378 (N_26378,N_25121,N_25607);
nand U26379 (N_26379,N_24799,N_24558);
or U26380 (N_26380,N_25109,N_25379);
xor U26381 (N_26381,N_25871,N_25509);
or U26382 (N_26382,N_24018,N_24561);
and U26383 (N_26383,N_24050,N_25080);
xor U26384 (N_26384,N_25360,N_25051);
or U26385 (N_26385,N_25817,N_25450);
nor U26386 (N_26386,N_25785,N_24379);
and U26387 (N_26387,N_25288,N_25229);
nand U26388 (N_26388,N_25779,N_25677);
nor U26389 (N_26389,N_24443,N_25356);
nor U26390 (N_26390,N_25111,N_25448);
or U26391 (N_26391,N_24085,N_25563);
xnor U26392 (N_26392,N_25407,N_24049);
nand U26393 (N_26393,N_24542,N_24261);
nand U26394 (N_26394,N_24737,N_25840);
and U26395 (N_26395,N_24129,N_24122);
or U26396 (N_26396,N_25049,N_25485);
or U26397 (N_26397,N_24958,N_24281);
xor U26398 (N_26398,N_24694,N_25766);
or U26399 (N_26399,N_24362,N_24842);
nand U26400 (N_26400,N_24025,N_25279);
and U26401 (N_26401,N_24072,N_25856);
nand U26402 (N_26402,N_24051,N_24258);
xnor U26403 (N_26403,N_25526,N_25235);
xnor U26404 (N_26404,N_25747,N_25593);
nand U26405 (N_26405,N_24208,N_24797);
nand U26406 (N_26406,N_24601,N_25555);
nor U26407 (N_26407,N_24194,N_25267);
and U26408 (N_26408,N_25820,N_25420);
nand U26409 (N_26409,N_25903,N_24871);
and U26410 (N_26410,N_24922,N_25876);
nor U26411 (N_26411,N_24420,N_24283);
and U26412 (N_26412,N_24740,N_24291);
or U26413 (N_26413,N_24502,N_25020);
nor U26414 (N_26414,N_24241,N_25772);
xnor U26415 (N_26415,N_25917,N_24575);
and U26416 (N_26416,N_24961,N_24332);
nor U26417 (N_26417,N_25283,N_25446);
xor U26418 (N_26418,N_25899,N_24003);
or U26419 (N_26419,N_25010,N_24608);
xor U26420 (N_26420,N_25054,N_24878);
xnor U26421 (N_26421,N_25866,N_24839);
nand U26422 (N_26422,N_24597,N_24641);
and U26423 (N_26423,N_24782,N_25254);
nor U26424 (N_26424,N_25734,N_25661);
or U26425 (N_26425,N_25281,N_25263);
or U26426 (N_26426,N_24501,N_25821);
nor U26427 (N_26427,N_25101,N_24452);
nor U26428 (N_26428,N_24784,N_24621);
nor U26429 (N_26429,N_24778,N_24234);
xor U26430 (N_26430,N_25918,N_25843);
and U26431 (N_26431,N_24263,N_25786);
nor U26432 (N_26432,N_24145,N_24535);
nor U26433 (N_26433,N_25273,N_24017);
or U26434 (N_26434,N_25986,N_25032);
xnor U26435 (N_26435,N_24162,N_24998);
xor U26436 (N_26436,N_25174,N_24378);
nand U26437 (N_26437,N_24135,N_25732);
nand U26438 (N_26438,N_25763,N_24223);
and U26439 (N_26439,N_25623,N_25233);
or U26440 (N_26440,N_24713,N_25861);
nor U26441 (N_26441,N_24798,N_24554);
xor U26442 (N_26442,N_24188,N_25727);
nor U26443 (N_26443,N_25256,N_24055);
and U26444 (N_26444,N_25171,N_24510);
nor U26445 (N_26445,N_25650,N_24631);
xor U26446 (N_26446,N_25013,N_25790);
nor U26447 (N_26447,N_24965,N_25465);
and U26448 (N_26448,N_24457,N_25146);
nand U26449 (N_26449,N_24328,N_25573);
nor U26450 (N_26450,N_25745,N_24586);
or U26451 (N_26451,N_25947,N_24235);
nand U26452 (N_26452,N_24187,N_25614);
and U26453 (N_26453,N_25801,N_24365);
nand U26454 (N_26454,N_24167,N_24874);
or U26455 (N_26455,N_25477,N_25596);
and U26456 (N_26456,N_24509,N_24298);
xnor U26457 (N_26457,N_24924,N_25368);
nand U26458 (N_26458,N_25725,N_24825);
xnor U26459 (N_26459,N_24761,N_25838);
xnor U26460 (N_26460,N_24914,N_24644);
nor U26461 (N_26461,N_25777,N_24351);
and U26462 (N_26462,N_24277,N_24517);
nand U26463 (N_26463,N_25570,N_25221);
nand U26464 (N_26464,N_25652,N_25729);
xnor U26465 (N_26465,N_25499,N_25996);
xor U26466 (N_26466,N_24939,N_24425);
xnor U26467 (N_26467,N_25015,N_24786);
and U26468 (N_26468,N_24231,N_24352);
nand U26469 (N_26469,N_24046,N_25189);
or U26470 (N_26470,N_24549,N_25715);
or U26471 (N_26471,N_24557,N_24692);
and U26472 (N_26472,N_24334,N_25430);
xnor U26473 (N_26473,N_25175,N_25521);
nand U26474 (N_26474,N_24948,N_25469);
nand U26475 (N_26475,N_25519,N_24350);
and U26476 (N_26476,N_25438,N_25633);
and U26477 (N_26477,N_25123,N_24066);
nand U26478 (N_26478,N_25670,N_25904);
and U26479 (N_26479,N_24977,N_24244);
xor U26480 (N_26480,N_24739,N_24177);
nor U26481 (N_26481,N_24815,N_25048);
nor U26482 (N_26482,N_25783,N_25592);
nor U26483 (N_26483,N_25236,N_24901);
or U26484 (N_26484,N_25402,N_25052);
and U26485 (N_26485,N_24499,N_25089);
or U26486 (N_26486,N_25100,N_24527);
nand U26487 (N_26487,N_25757,N_24360);
nand U26488 (N_26488,N_24563,N_24927);
or U26489 (N_26489,N_24392,N_25539);
nor U26490 (N_26490,N_25648,N_24680);
or U26491 (N_26491,N_24984,N_25664);
xnor U26492 (N_26492,N_24030,N_25971);
nor U26493 (N_26493,N_25115,N_24274);
and U26494 (N_26494,N_24988,N_24951);
and U26495 (N_26495,N_25896,N_25191);
nor U26496 (N_26496,N_25334,N_24695);
nor U26497 (N_26497,N_25959,N_24148);
nand U26498 (N_26498,N_25604,N_25084);
or U26499 (N_26499,N_24325,N_24886);
or U26500 (N_26500,N_25314,N_24693);
or U26501 (N_26501,N_24033,N_25177);
nand U26502 (N_26502,N_25060,N_25512);
or U26503 (N_26503,N_24654,N_25713);
nand U26504 (N_26504,N_25366,N_24691);
and U26505 (N_26505,N_25731,N_24829);
nand U26506 (N_26506,N_25875,N_24031);
nand U26507 (N_26507,N_25449,N_25750);
nor U26508 (N_26508,N_24006,N_24057);
nand U26509 (N_26509,N_24133,N_24376);
nand U26510 (N_26510,N_25687,N_24664);
nor U26511 (N_26511,N_24029,N_25083);
xor U26512 (N_26512,N_25250,N_24095);
nand U26513 (N_26513,N_24746,N_25551);
nand U26514 (N_26514,N_24791,N_24230);
nor U26515 (N_26515,N_25228,N_25800);
nor U26516 (N_26516,N_24918,N_25073);
nor U26517 (N_26517,N_25892,N_25587);
xor U26518 (N_26518,N_24453,N_24415);
nand U26519 (N_26519,N_24371,N_24941);
or U26520 (N_26520,N_25581,N_24833);
xor U26521 (N_26521,N_24674,N_25802);
nand U26522 (N_26522,N_24805,N_25275);
xor U26523 (N_26523,N_24446,N_24522);
nor U26524 (N_26524,N_24111,N_24899);
nand U26525 (N_26525,N_25471,N_24269);
nand U26526 (N_26526,N_25936,N_25752);
or U26527 (N_26527,N_25276,N_25208);
and U26528 (N_26528,N_25647,N_25658);
nand U26529 (N_26529,N_24175,N_25686);
nor U26530 (N_26530,N_24814,N_24236);
or U26531 (N_26531,N_25868,N_25167);
nor U26532 (N_26532,N_25497,N_25295);
and U26533 (N_26533,N_24228,N_25170);
nor U26534 (N_26534,N_25858,N_24827);
and U26535 (N_26535,N_24486,N_25842);
nand U26536 (N_26536,N_24547,N_24950);
xor U26537 (N_26537,N_25567,N_25472);
xnor U26538 (N_26538,N_25038,N_25873);
xnor U26539 (N_26539,N_24032,N_25122);
nand U26540 (N_26540,N_24092,N_25007);
nor U26541 (N_26541,N_24603,N_25855);
and U26542 (N_26542,N_25016,N_24574);
nor U26543 (N_26543,N_25394,N_24843);
nand U26544 (N_26544,N_24720,N_24993);
or U26545 (N_26545,N_25442,N_25928);
xor U26546 (N_26546,N_25957,N_25755);
or U26547 (N_26547,N_24590,N_25810);
and U26548 (N_26548,N_24800,N_25545);
nor U26549 (N_26549,N_24847,N_25771);
nor U26550 (N_26550,N_24859,N_24923);
nand U26551 (N_26551,N_24438,N_25026);
nand U26552 (N_26552,N_25720,N_24227);
xnor U26553 (N_26553,N_24197,N_25967);
xnor U26554 (N_26554,N_24777,N_25354);
or U26555 (N_26555,N_24808,N_25398);
and U26556 (N_26556,N_25893,N_24852);
xor U26557 (N_26557,N_24955,N_24005);
nor U26558 (N_26558,N_25435,N_25451);
or U26559 (N_26559,N_24161,N_25510);
nand U26560 (N_26560,N_24519,N_25640);
nand U26561 (N_26561,N_24077,N_25326);
nor U26562 (N_26562,N_25436,N_25128);
or U26563 (N_26563,N_24954,N_25503);
or U26564 (N_26564,N_25076,N_24572);
xnor U26565 (N_26565,N_25413,N_24735);
nor U26566 (N_26566,N_25937,N_24972);
or U26567 (N_26567,N_24218,N_25694);
xnor U26568 (N_26568,N_24705,N_24205);
nand U26569 (N_26569,N_25099,N_24173);
and U26570 (N_26570,N_25331,N_25883);
or U26571 (N_26571,N_24259,N_24790);
xor U26572 (N_26572,N_24966,N_25557);
or U26573 (N_26573,N_25070,N_24826);
xnor U26574 (N_26574,N_25572,N_25396);
nand U26575 (N_26575,N_24123,N_25635);
or U26576 (N_26576,N_24992,N_25834);
nor U26577 (N_26577,N_24466,N_25721);
and U26578 (N_26578,N_24060,N_24904);
xnor U26579 (N_26579,N_25371,N_25644);
xnor U26580 (N_26580,N_24500,N_25908);
or U26581 (N_26581,N_24888,N_24666);
or U26582 (N_26582,N_24806,N_24559);
and U26583 (N_26583,N_24910,N_24393);
and U26584 (N_26584,N_24872,N_24472);
xor U26585 (N_26585,N_24278,N_25453);
or U26586 (N_26586,N_24408,N_24266);
xnor U26587 (N_26587,N_24863,N_24749);
nor U26588 (N_26588,N_24138,N_25671);
or U26589 (N_26589,N_24689,N_24818);
xor U26590 (N_26590,N_25926,N_24903);
and U26591 (N_26591,N_24082,N_24892);
nor U26592 (N_26592,N_25461,N_24609);
and U26593 (N_26593,N_24160,N_24154);
and U26594 (N_26594,N_25474,N_24103);
or U26595 (N_26595,N_25220,N_25827);
or U26596 (N_26596,N_25523,N_25266);
and U26597 (N_26597,N_25419,N_24271);
nor U26598 (N_26598,N_24384,N_25854);
and U26599 (N_26599,N_25699,N_25676);
xor U26600 (N_26600,N_24788,N_24206);
nand U26601 (N_26601,N_24969,N_25958);
xor U26602 (N_26602,N_24387,N_25200);
xor U26603 (N_26603,N_25056,N_25569);
nor U26604 (N_26604,N_25890,N_24570);
or U26605 (N_26605,N_25037,N_24088);
nand U26606 (N_26606,N_25618,N_24543);
nor U26607 (N_26607,N_25444,N_25103);
xor U26608 (N_26608,N_25968,N_24385);
nor U26609 (N_26609,N_24203,N_25074);
and U26610 (N_26610,N_25857,N_25464);
and U26611 (N_26611,N_24677,N_24893);
or U26612 (N_26612,N_25028,N_25432);
nor U26613 (N_26613,N_25770,N_25329);
nor U26614 (N_26614,N_24766,N_24413);
xor U26615 (N_26615,N_24755,N_25490);
xnor U26616 (N_26616,N_25234,N_25832);
and U26617 (N_26617,N_25597,N_25508);
and U26618 (N_26618,N_25536,N_25672);
nor U26619 (N_26619,N_25902,N_24100);
nor U26620 (N_26620,N_24656,N_24794);
xor U26621 (N_26621,N_24198,N_25313);
xnor U26622 (N_26622,N_25921,N_25058);
or U26623 (N_26623,N_25359,N_24734);
and U26624 (N_26624,N_24021,N_24909);
and U26625 (N_26625,N_25962,N_24368);
nand U26626 (N_26626,N_24465,N_24661);
xnor U26627 (N_26627,N_25712,N_25954);
or U26628 (N_26628,N_24459,N_24493);
nor U26629 (N_26629,N_25300,N_24885);
and U26630 (N_26630,N_25836,N_25145);
nor U26631 (N_26631,N_24273,N_25774);
xnor U26632 (N_26632,N_25579,N_25620);
nand U26633 (N_26633,N_24411,N_25673);
nor U26634 (N_26634,N_24293,N_24404);
nand U26635 (N_26635,N_24754,N_25270);
or U26636 (N_26636,N_25657,N_25198);
nor U26637 (N_26637,N_25702,N_25591);
xnor U26638 (N_26638,N_25138,N_24959);
and U26639 (N_26639,N_25423,N_25584);
xor U26640 (N_26640,N_24832,N_24091);
xor U26641 (N_26641,N_24638,N_25369);
and U26642 (N_26642,N_25404,N_24120);
nor U26643 (N_26643,N_24089,N_24850);
nand U26644 (N_26644,N_25165,N_24584);
or U26645 (N_26645,N_24310,N_25841);
and U26646 (N_26646,N_25377,N_25104);
nor U26647 (N_26647,N_25425,N_24253);
and U26648 (N_26648,N_24348,N_24265);
and U26649 (N_26649,N_25681,N_25683);
nand U26650 (N_26650,N_25789,N_24116);
or U26651 (N_26651,N_25600,N_25616);
nand U26652 (N_26652,N_24751,N_24434);
and U26653 (N_26653,N_25487,N_25632);
nand U26654 (N_26654,N_24732,N_25889);
xnor U26655 (N_26655,N_25382,N_25865);
and U26656 (N_26656,N_24260,N_25674);
and U26657 (N_26657,N_25309,N_24267);
and U26658 (N_26658,N_25768,N_25571);
xnor U26659 (N_26659,N_24397,N_24956);
xnor U26660 (N_26660,N_24613,N_24056);
nor U26661 (N_26661,N_24929,N_25679);
xnor U26662 (N_26662,N_24461,N_24451);
xnor U26663 (N_26663,N_25595,N_24991);
nand U26664 (N_26664,N_25575,N_25787);
nor U26665 (N_26665,N_25869,N_24742);
nor U26666 (N_26666,N_25350,N_25117);
nand U26667 (N_26667,N_25848,N_25568);
or U26668 (N_26668,N_25320,N_24884);
xnor U26669 (N_26669,N_25543,N_24687);
nand U26670 (N_26670,N_24721,N_24190);
nor U26671 (N_26671,N_24727,N_25373);
xor U26672 (N_26672,N_25685,N_24295);
xnor U26673 (N_26673,N_24816,N_25482);
xor U26674 (N_26674,N_24316,N_24147);
and U26675 (N_26675,N_24028,N_25870);
and U26676 (N_26676,N_24770,N_24830);
or U26677 (N_26677,N_25286,N_25580);
and U26678 (N_26678,N_24047,N_24781);
and U26679 (N_26679,N_25249,N_24849);
nor U26680 (N_26680,N_25799,N_24330);
and U26681 (N_26681,N_24743,N_25339);
nand U26682 (N_26682,N_25586,N_24156);
and U26683 (N_26683,N_24606,N_25480);
nand U26684 (N_26684,N_25181,N_24836);
or U26685 (N_26685,N_24612,N_24553);
xor U26686 (N_26686,N_25291,N_25703);
or U26687 (N_26687,N_24482,N_24824);
or U26688 (N_26688,N_25792,N_25033);
nand U26689 (N_26689,N_24710,N_24318);
and U26690 (N_26690,N_24210,N_24474);
xnor U26691 (N_26691,N_25190,N_25108);
nor U26692 (N_26692,N_25705,N_24773);
xnor U26693 (N_26693,N_25304,N_24080);
or U26694 (N_26694,N_25457,N_24518);
nand U26695 (N_26695,N_25651,N_24823);
and U26696 (N_26696,N_24142,N_24820);
and U26697 (N_26697,N_24990,N_25367);
xor U26698 (N_26698,N_25706,N_24819);
nand U26699 (N_26699,N_25991,N_25459);
and U26700 (N_26700,N_24383,N_25500);
nand U26701 (N_26701,N_25891,N_25982);
and U26702 (N_26702,N_24370,N_25878);
xor U26703 (N_26703,N_25934,N_25150);
and U26704 (N_26704,N_24635,N_24484);
xnor U26705 (N_26705,N_25637,N_24109);
or U26706 (N_26706,N_24729,N_25043);
and U26707 (N_26707,N_25399,N_25701);
xnor U26708 (N_26708,N_25634,N_25513);
or U26709 (N_26709,N_25961,N_24783);
nand U26710 (N_26710,N_25574,N_25040);
nand U26711 (N_26711,N_24657,N_25086);
nand U26712 (N_26712,N_25960,N_24480);
nor U26713 (N_26713,N_25193,N_24314);
nor U26714 (N_26714,N_24703,N_24906);
nor U26715 (N_26715,N_25907,N_25203);
xnor U26716 (N_26716,N_24628,N_25769);
nand U26717 (N_26717,N_25911,N_25940);
xnor U26718 (N_26718,N_24219,N_25601);
nor U26719 (N_26719,N_24776,N_24702);
xnor U26720 (N_26720,N_25212,N_25722);
nor U26721 (N_26721,N_25930,N_24706);
nor U26722 (N_26722,N_25695,N_24925);
and U26723 (N_26723,N_24629,N_24200);
nor U26724 (N_26724,N_25483,N_24653);
nand U26725 (N_26725,N_24938,N_24232);
xnor U26726 (N_26726,N_24684,N_25807);
nor U26727 (N_26727,N_24916,N_25427);
nand U26728 (N_26728,N_25826,N_24494);
xor U26729 (N_26729,N_25764,N_25042);
nor U26730 (N_26730,N_25767,N_25152);
nor U26731 (N_26731,N_24440,N_25833);
or U26732 (N_26732,N_25226,N_24071);
nor U26733 (N_26733,N_25301,N_25818);
and U26734 (N_26734,N_25306,N_24286);
or U26735 (N_26735,N_24418,N_24978);
xor U26736 (N_26736,N_24624,N_25689);
xnor U26737 (N_26737,N_24405,N_24184);
xor U26738 (N_26738,N_24861,N_25452);
and U26739 (N_26739,N_25124,N_24010);
and U26740 (N_26740,N_24130,N_25992);
or U26741 (N_26741,N_25055,N_24841);
nor U26742 (N_26742,N_25416,N_25621);
xnor U26743 (N_26743,N_24007,N_24550);
xnor U26744 (N_26744,N_25284,N_24448);
nand U26745 (N_26745,N_24321,N_25321);
xnor U26746 (N_26746,N_25932,N_25297);
or U26747 (N_26747,N_24745,N_25348);
and U26748 (N_26748,N_25034,N_25515);
and U26749 (N_26749,N_25518,N_25553);
nor U26750 (N_26750,N_24920,N_25983);
xnor U26751 (N_26751,N_24932,N_25479);
nand U26752 (N_26752,N_24338,N_24592);
nand U26753 (N_26753,N_25885,N_25825);
xnor U26754 (N_26754,N_24708,N_25014);
nor U26755 (N_26755,N_25365,N_24515);
nor U26756 (N_26756,N_24026,N_25736);
and U26757 (N_26757,N_25153,N_24456);
or U26758 (N_26758,N_25708,N_24614);
xnor U26759 (N_26759,N_24667,N_25583);
or U26760 (N_26760,N_25655,N_24523);
or U26761 (N_26761,N_24467,N_24698);
or U26762 (N_26762,N_25139,N_25979);
or U26763 (N_26763,N_24419,N_25455);
or U26764 (N_26764,N_25092,N_24136);
or U26765 (N_26765,N_25183,N_24726);
xnor U26766 (N_26766,N_25544,N_24546);
or U26767 (N_26767,N_25486,N_25094);
nor U26768 (N_26768,N_24191,N_24599);
xor U26769 (N_26769,N_24845,N_25978);
and U26770 (N_26770,N_24038,N_25588);
nor U26771 (N_26771,N_24340,N_25780);
xnor U26772 (N_26772,N_24361,N_24540);
xor U26773 (N_26773,N_24579,N_24471);
nand U26774 (N_26774,N_25909,N_25758);
xnor U26775 (N_26775,N_24617,N_25641);
nand U26776 (N_26776,N_25920,N_24217);
and U26777 (N_26777,N_25791,N_25624);
and U26778 (N_26778,N_24140,N_25282);
nand U26779 (N_26779,N_24256,N_25312);
xnor U26780 (N_26780,N_25542,N_24615);
nand U26781 (N_26781,N_24012,N_24359);
and U26782 (N_26782,N_24697,N_25001);
and U26783 (N_26783,N_25643,N_25608);
nand U26784 (N_26784,N_25988,N_24894);
xor U26785 (N_26785,N_24201,N_25533);
xor U26786 (N_26786,N_25740,N_25091);
and U26787 (N_26787,N_25662,N_25164);
nand U26788 (N_26788,N_24394,N_25859);
xnor U26789 (N_26789,N_25133,N_24164);
and U26790 (N_26790,N_25285,N_25585);
nand U26791 (N_26791,N_25000,N_24541);
and U26792 (N_26792,N_25846,N_24715);
or U26793 (N_26793,N_24980,N_24887);
xor U26794 (N_26794,N_25346,N_24409);
nor U26795 (N_26795,N_25186,N_25188);
nor U26796 (N_26796,N_25795,N_25144);
nor U26797 (N_26797,N_24251,N_25793);
xor U26798 (N_26798,N_25293,N_24516);
nand U26799 (N_26799,N_25576,N_24207);
xnor U26800 (N_26800,N_25475,N_25244);
or U26801 (N_26801,N_25970,N_25781);
and U26802 (N_26802,N_25141,N_24063);
and U26803 (N_26803,N_24344,N_25290);
xnor U26804 (N_26804,N_24168,N_25202);
nand U26805 (N_26805,N_25456,N_25131);
or U26806 (N_26806,N_24902,N_24008);
nor U26807 (N_26807,N_24822,N_24216);
xor U26808 (N_26808,N_25874,N_24366);
and U26809 (N_26809,N_25534,N_24662);
and U26810 (N_26810,N_25011,N_25504);
xnor U26811 (N_26811,N_24144,N_25386);
or U26812 (N_26812,N_25132,N_24128);
xnor U26813 (N_26813,N_25414,N_25353);
xor U26814 (N_26814,N_25022,N_24831);
xor U26815 (N_26815,N_24696,N_24099);
nor U26816 (N_26816,N_25880,N_24917);
and U26817 (N_26817,N_25006,N_25097);
or U26818 (N_26818,N_24171,N_25659);
or U26819 (N_26819,N_25554,N_25765);
xor U26820 (N_26820,N_24121,N_25955);
nor U26821 (N_26821,N_25522,N_24022);
nand U26822 (N_26822,N_24944,N_25716);
nand U26823 (N_26823,N_25925,N_25343);
xnor U26824 (N_26824,N_25338,N_24919);
nor U26825 (N_26825,N_25811,N_25942);
xnor U26826 (N_26826,N_24239,N_25424);
xor U26827 (N_26827,N_25981,N_25294);
or U26828 (N_26828,N_25628,N_25473);
and U26829 (N_26829,N_24483,N_24491);
or U26830 (N_26830,N_25411,N_25406);
xor U26831 (N_26831,N_25578,N_24276);
or U26832 (N_26832,N_25046,N_25173);
nand U26833 (N_26833,N_25589,N_25075);
nor U26834 (N_26834,N_25417,N_25822);
or U26835 (N_26835,N_24146,N_24275);
and U26836 (N_26836,N_24581,N_24331);
nor U26837 (N_26837,N_24105,N_25549);
xor U26838 (N_26838,N_24753,N_24339);
or U26839 (N_26839,N_25966,N_25053);
and U26840 (N_26840,N_25517,N_24600);
xor U26841 (N_26841,N_25973,N_24714);
xnor U26842 (N_26842,N_25316,N_24221);
and U26843 (N_26843,N_25603,N_25195);
and U26844 (N_26844,N_25383,N_25804);
nand U26845 (N_26845,N_24723,N_24180);
nand U26846 (N_26846,N_24928,N_24343);
or U26847 (N_26847,N_25323,N_25598);
or U26848 (N_26848,N_24555,N_25839);
or U26849 (N_26849,N_25090,N_25782);
nand U26850 (N_26850,N_24478,N_25218);
and U26851 (N_26851,N_24237,N_25336);
nand U26852 (N_26852,N_24681,N_24736);
xnor U26853 (N_26853,N_24224,N_25547);
nand U26854 (N_26854,N_25625,N_25803);
and U26855 (N_26855,N_24974,N_25147);
or U26856 (N_26856,N_24771,N_25898);
or U26857 (N_26857,N_25733,N_25158);
nor U26858 (N_26858,N_25400,N_24529);
nor U26859 (N_26859,N_25974,N_24528);
nand U26860 (N_26860,N_25362,N_25045);
xor U26861 (N_26861,N_25531,N_24075);
nand U26862 (N_26862,N_25161,N_25105);
xor U26863 (N_26863,N_24672,N_24302);
nand U26864 (N_26864,N_25631,N_24989);
nor U26865 (N_26865,N_24470,N_25409);
nor U26866 (N_26866,N_25223,N_24857);
nand U26867 (N_26867,N_24449,N_25887);
and U26868 (N_26868,N_25211,N_24301);
xnor U26869 (N_26869,N_24809,N_25760);
nand U26870 (N_26870,N_24503,N_24300);
nor U26871 (N_26871,N_24719,N_24690);
nor U26872 (N_26872,N_25385,N_25872);
nand U26873 (N_26873,N_24981,N_25391);
nand U26874 (N_26874,N_25964,N_25565);
nand U26875 (N_26875,N_24307,N_25823);
nor U26876 (N_26876,N_25697,N_25558);
or U26877 (N_26877,N_25251,N_25520);
xnor U26878 (N_26878,N_25762,N_24647);
xor U26879 (N_26879,N_25977,N_24514);
xor U26880 (N_26880,N_24837,N_24132);
or U26881 (N_26881,N_25488,N_25494);
and U26882 (N_26882,N_24536,N_24009);
nand U26883 (N_26883,N_24179,N_24983);
xor U26884 (N_26884,N_25095,N_25199);
xnor U26885 (N_26885,N_25002,N_24398);
nand U26886 (N_26886,N_25019,N_24178);
and U26887 (N_26887,N_24117,N_24537);
or U26888 (N_26888,N_24192,N_25724);
xnor U26889 (N_26889,N_25433,N_25216);
or U26890 (N_26890,N_25422,N_24545);
nor U26891 (N_26891,N_24846,N_24531);
nand U26892 (N_26892,N_25231,N_24093);
xnor U26893 (N_26893,N_25556,N_25691);
xnor U26894 (N_26894,N_24704,N_25035);
nand U26895 (N_26895,N_24282,N_25112);
nand U26896 (N_26896,N_24676,N_25030);
nand U26897 (N_26897,N_24432,N_24485);
and U26898 (N_26898,N_25412,N_25994);
nor U26899 (N_26899,N_25527,N_24199);
nand U26900 (N_26900,N_24322,N_24069);
nor U26901 (N_26901,N_25610,N_24933);
nor U26902 (N_26902,N_25415,N_25737);
xnor U26903 (N_26903,N_25447,N_25340);
xor U26904 (N_26904,N_25289,N_25704);
nand U26905 (N_26905,N_25004,N_24296);
nor U26906 (N_26906,N_25944,N_24158);
nor U26907 (N_26907,N_24602,N_24940);
or U26908 (N_26908,N_25759,N_24246);
nand U26909 (N_26909,N_25938,N_25441);
and U26910 (N_26910,N_24801,N_25082);
or U26911 (N_26911,N_25901,N_24159);
or U26912 (N_26912,N_24125,N_24526);
nand U26913 (N_26913,N_25277,N_24870);
xor U26914 (N_26914,N_25711,N_24860);
and U26915 (N_26915,N_25355,N_25209);
or U26916 (N_26916,N_24367,N_25031);
xnor U26917 (N_26917,N_25828,N_25484);
xnor U26918 (N_26918,N_24058,N_24455);
nor U26919 (N_26919,N_24757,N_24921);
and U26920 (N_26920,N_24287,N_25349);
nor U26921 (N_26921,N_25564,N_24931);
or U26922 (N_26922,N_25096,N_25159);
xnor U26923 (N_26923,N_24883,N_24034);
and U26924 (N_26924,N_24970,N_25590);
or U26925 (N_26925,N_24744,N_25778);
or U26926 (N_26926,N_25844,N_24181);
nand U26927 (N_26927,N_24400,N_24508);
nand U26928 (N_26928,N_24840,N_25693);
nand U26929 (N_26929,N_25036,N_24202);
or U26930 (N_26930,N_24312,N_25864);
xnor U26931 (N_26931,N_25401,N_24035);
and U26932 (N_26932,N_25646,N_24506);
and U26933 (N_26933,N_24709,N_25201);
nor U26934 (N_26934,N_25853,N_25069);
nand U26935 (N_26935,N_24124,N_24086);
nor U26936 (N_26936,N_25688,N_24688);
xor U26937 (N_26937,N_24741,N_25426);
nor U26938 (N_26938,N_25675,N_25665);
and U26939 (N_26939,N_25615,N_24386);
and U26940 (N_26940,N_24881,N_24803);
and U26941 (N_26941,N_25168,N_24633);
and U26942 (N_26942,N_25995,N_25753);
nand U26943 (N_26943,N_25372,N_25107);
xor U26944 (N_26944,N_25332,N_25860);
xor U26945 (N_26945,N_25027,N_24769);
xnor U26946 (N_26946,N_24975,N_25723);
xnor U26947 (N_26947,N_24718,N_24879);
nand U26948 (N_26948,N_25849,N_25862);
xor U26949 (N_26949,N_24139,N_25945);
nor U26950 (N_26950,N_24083,N_24658);
xor U26951 (N_26951,N_24858,N_25742);
xnor U26952 (N_26952,N_25599,N_24479);
or U26953 (N_26953,N_24964,N_25081);
and U26954 (N_26954,N_25649,N_24417);
nand U26955 (N_26955,N_24183,N_24963);
and U26956 (N_26956,N_24213,N_24942);
and U26957 (N_26957,N_24079,N_24949);
nand U26958 (N_26958,N_25943,N_25912);
nor U26959 (N_26959,N_25948,N_24243);
xor U26960 (N_26960,N_24496,N_24435);
nand U26961 (N_26961,N_25118,N_25884);
nor U26962 (N_26962,N_25079,N_24670);
nor U26963 (N_26963,N_24036,N_24604);
nand U26964 (N_26964,N_25582,N_24189);
nor U26965 (N_26965,N_24157,N_25012);
nand U26966 (N_26966,N_25532,N_24097);
xnor U26967 (N_26967,N_24962,N_25119);
xor U26968 (N_26968,N_25130,N_24898);
nor U26969 (N_26969,N_25224,N_24264);
xor U26970 (N_26970,N_25993,N_24303);
and U26971 (N_26971,N_25057,N_25746);
and U26972 (N_26972,N_25238,N_24611);
and U26973 (N_26973,N_24915,N_25744);
nor U26974 (N_26974,N_25660,N_24257);
and U26975 (N_26975,N_24759,N_25098);
nand U26976 (N_26976,N_24341,N_24445);
nor U26977 (N_26977,N_25502,N_24953);
nand U26978 (N_26978,N_24646,N_24996);
xor U26979 (N_26979,N_24106,N_24985);
and U26980 (N_26980,N_24407,N_25110);
xnor U26981 (N_26981,N_25265,N_24104);
or U26982 (N_26982,N_25501,N_24866);
nand U26983 (N_26983,N_24292,N_24787);
nor U26984 (N_26984,N_25210,N_25749);
and U26985 (N_26985,N_25364,N_25698);
and U26986 (N_26986,N_24789,N_24873);
nor U26987 (N_26987,N_25924,N_24248);
nor U26988 (N_26988,N_24458,N_24073);
nand U26989 (N_26989,N_25514,N_24141);
xnor U26990 (N_26990,N_24854,N_24577);
xor U26991 (N_26991,N_24625,N_25162);
nor U26992 (N_26992,N_25922,N_24686);
nand U26993 (N_26993,N_24865,N_24424);
nand U26994 (N_26994,N_25324,N_24632);
xnor U26995 (N_26995,N_24294,N_25914);
or U26996 (N_26996,N_25775,N_25863);
xnor U26997 (N_26997,N_24655,N_25773);
xnor U26998 (N_26998,N_25120,N_24463);
nor U26999 (N_26999,N_25151,N_24174);
and U27000 (N_27000,N_25641,N_25427);
xor U27001 (N_27001,N_25172,N_24181);
or U27002 (N_27002,N_25476,N_25292);
or U27003 (N_27003,N_24905,N_25489);
nor U27004 (N_27004,N_24697,N_24126);
xor U27005 (N_27005,N_25061,N_25657);
nor U27006 (N_27006,N_25554,N_24949);
xnor U27007 (N_27007,N_25402,N_25819);
and U27008 (N_27008,N_25982,N_25406);
or U27009 (N_27009,N_24338,N_24603);
xor U27010 (N_27010,N_25331,N_25717);
nand U27011 (N_27011,N_24196,N_25720);
nand U27012 (N_27012,N_24770,N_24322);
nor U27013 (N_27013,N_25628,N_24949);
or U27014 (N_27014,N_24554,N_25408);
xor U27015 (N_27015,N_24880,N_25494);
and U27016 (N_27016,N_24065,N_24870);
nor U27017 (N_27017,N_25214,N_25361);
or U27018 (N_27018,N_24060,N_24639);
xnor U27019 (N_27019,N_24118,N_24336);
and U27020 (N_27020,N_24856,N_24211);
nand U27021 (N_27021,N_24317,N_24532);
nand U27022 (N_27022,N_25483,N_25653);
and U27023 (N_27023,N_24594,N_24008);
and U27024 (N_27024,N_25289,N_25724);
and U27025 (N_27025,N_24326,N_25200);
or U27026 (N_27026,N_25010,N_24209);
nand U27027 (N_27027,N_24547,N_25337);
nand U27028 (N_27028,N_24485,N_24113);
nor U27029 (N_27029,N_24190,N_25639);
and U27030 (N_27030,N_25478,N_25878);
nor U27031 (N_27031,N_24984,N_24499);
nor U27032 (N_27032,N_24543,N_25553);
xnor U27033 (N_27033,N_24726,N_24352);
and U27034 (N_27034,N_25846,N_25408);
xnor U27035 (N_27035,N_25031,N_24703);
xnor U27036 (N_27036,N_25553,N_24561);
and U27037 (N_27037,N_24102,N_25234);
nand U27038 (N_27038,N_24366,N_25622);
and U27039 (N_27039,N_24534,N_25502);
or U27040 (N_27040,N_24254,N_24713);
or U27041 (N_27041,N_24730,N_25848);
xor U27042 (N_27042,N_25248,N_24330);
xor U27043 (N_27043,N_25216,N_25991);
or U27044 (N_27044,N_24900,N_25305);
xor U27045 (N_27045,N_25006,N_24054);
nand U27046 (N_27046,N_25117,N_25054);
nor U27047 (N_27047,N_24296,N_24366);
nand U27048 (N_27048,N_25191,N_25146);
nor U27049 (N_27049,N_25977,N_25851);
and U27050 (N_27050,N_25655,N_24350);
xor U27051 (N_27051,N_25981,N_24059);
or U27052 (N_27052,N_25051,N_25455);
nor U27053 (N_27053,N_25248,N_25808);
nor U27054 (N_27054,N_25627,N_24084);
xor U27055 (N_27055,N_25473,N_24624);
nand U27056 (N_27056,N_24914,N_24438);
nand U27057 (N_27057,N_25100,N_25325);
xnor U27058 (N_27058,N_25856,N_25639);
and U27059 (N_27059,N_24300,N_25941);
and U27060 (N_27060,N_24566,N_25754);
nor U27061 (N_27061,N_24891,N_24464);
and U27062 (N_27062,N_25654,N_24766);
xor U27063 (N_27063,N_25684,N_25391);
nand U27064 (N_27064,N_24548,N_24820);
xor U27065 (N_27065,N_25931,N_25482);
xnor U27066 (N_27066,N_25155,N_25718);
nor U27067 (N_27067,N_25868,N_25958);
xnor U27068 (N_27068,N_25954,N_24565);
or U27069 (N_27069,N_25455,N_25805);
and U27070 (N_27070,N_25472,N_24312);
nor U27071 (N_27071,N_24897,N_24600);
xor U27072 (N_27072,N_24629,N_25004);
nand U27073 (N_27073,N_24394,N_25106);
xor U27074 (N_27074,N_25234,N_25970);
nand U27075 (N_27075,N_25490,N_24305);
nor U27076 (N_27076,N_25633,N_25677);
or U27077 (N_27077,N_25337,N_24916);
xnor U27078 (N_27078,N_25992,N_24721);
nor U27079 (N_27079,N_24036,N_25585);
or U27080 (N_27080,N_25951,N_24419);
and U27081 (N_27081,N_24149,N_25848);
xor U27082 (N_27082,N_24097,N_24816);
xor U27083 (N_27083,N_25490,N_25289);
and U27084 (N_27084,N_25149,N_25700);
nor U27085 (N_27085,N_25821,N_25677);
and U27086 (N_27086,N_24854,N_24889);
nand U27087 (N_27087,N_25967,N_25653);
and U27088 (N_27088,N_24579,N_25527);
nand U27089 (N_27089,N_25687,N_25970);
or U27090 (N_27090,N_25572,N_24305);
xnor U27091 (N_27091,N_24953,N_25086);
xnor U27092 (N_27092,N_24192,N_24509);
or U27093 (N_27093,N_24213,N_25598);
and U27094 (N_27094,N_24579,N_25324);
nand U27095 (N_27095,N_24822,N_24534);
nor U27096 (N_27096,N_24339,N_25873);
or U27097 (N_27097,N_25128,N_25024);
nand U27098 (N_27098,N_25036,N_24738);
nor U27099 (N_27099,N_24527,N_24494);
or U27100 (N_27100,N_25568,N_25730);
and U27101 (N_27101,N_24453,N_24061);
nor U27102 (N_27102,N_24852,N_25124);
nor U27103 (N_27103,N_25770,N_25646);
or U27104 (N_27104,N_25892,N_25807);
or U27105 (N_27105,N_25642,N_24383);
nor U27106 (N_27106,N_24994,N_24959);
nand U27107 (N_27107,N_24001,N_25113);
and U27108 (N_27108,N_24276,N_24138);
xor U27109 (N_27109,N_24775,N_25468);
nor U27110 (N_27110,N_24058,N_25599);
nand U27111 (N_27111,N_24142,N_24738);
or U27112 (N_27112,N_25129,N_25856);
or U27113 (N_27113,N_25287,N_25504);
and U27114 (N_27114,N_25279,N_24633);
nand U27115 (N_27115,N_24982,N_25327);
xnor U27116 (N_27116,N_25426,N_25526);
or U27117 (N_27117,N_24466,N_25722);
nand U27118 (N_27118,N_24812,N_25370);
or U27119 (N_27119,N_24600,N_25870);
nor U27120 (N_27120,N_25733,N_24974);
nor U27121 (N_27121,N_25982,N_25181);
nor U27122 (N_27122,N_24518,N_25257);
nor U27123 (N_27123,N_24714,N_24295);
xnor U27124 (N_27124,N_24983,N_25958);
xor U27125 (N_27125,N_25425,N_25201);
nor U27126 (N_27126,N_25062,N_25358);
xnor U27127 (N_27127,N_24547,N_25816);
nand U27128 (N_27128,N_25575,N_24875);
nor U27129 (N_27129,N_24309,N_24293);
or U27130 (N_27130,N_24038,N_24826);
nor U27131 (N_27131,N_25070,N_24582);
nor U27132 (N_27132,N_25789,N_25215);
nand U27133 (N_27133,N_25087,N_25410);
and U27134 (N_27134,N_24054,N_25476);
nand U27135 (N_27135,N_25989,N_25593);
and U27136 (N_27136,N_25349,N_24513);
nor U27137 (N_27137,N_24182,N_25218);
nand U27138 (N_27138,N_24048,N_24031);
nor U27139 (N_27139,N_25821,N_24042);
xnor U27140 (N_27140,N_24591,N_25192);
nand U27141 (N_27141,N_24995,N_24769);
or U27142 (N_27142,N_24594,N_25891);
xnor U27143 (N_27143,N_24770,N_24297);
and U27144 (N_27144,N_24034,N_25661);
nor U27145 (N_27145,N_25762,N_25725);
and U27146 (N_27146,N_24221,N_24043);
nand U27147 (N_27147,N_24639,N_25432);
nor U27148 (N_27148,N_25653,N_24031);
nor U27149 (N_27149,N_25902,N_24381);
xor U27150 (N_27150,N_24298,N_25587);
xor U27151 (N_27151,N_24383,N_24607);
nand U27152 (N_27152,N_24237,N_24325);
xnor U27153 (N_27153,N_25267,N_24714);
nor U27154 (N_27154,N_25658,N_24771);
nor U27155 (N_27155,N_25012,N_24263);
or U27156 (N_27156,N_24873,N_25808);
and U27157 (N_27157,N_24463,N_25594);
nor U27158 (N_27158,N_24891,N_24589);
and U27159 (N_27159,N_25913,N_25586);
nor U27160 (N_27160,N_24608,N_24928);
or U27161 (N_27161,N_25961,N_24026);
nor U27162 (N_27162,N_25870,N_24996);
or U27163 (N_27163,N_25529,N_25590);
nor U27164 (N_27164,N_25049,N_25228);
or U27165 (N_27165,N_25610,N_25339);
or U27166 (N_27166,N_24397,N_24986);
nand U27167 (N_27167,N_24036,N_25849);
nor U27168 (N_27168,N_24791,N_25461);
and U27169 (N_27169,N_25186,N_24937);
or U27170 (N_27170,N_24246,N_24707);
or U27171 (N_27171,N_24960,N_25264);
or U27172 (N_27172,N_25621,N_24538);
xor U27173 (N_27173,N_25551,N_25546);
nor U27174 (N_27174,N_24997,N_25411);
nor U27175 (N_27175,N_24209,N_25053);
and U27176 (N_27176,N_25396,N_24017);
nor U27177 (N_27177,N_24299,N_24504);
xor U27178 (N_27178,N_24841,N_25805);
nor U27179 (N_27179,N_25426,N_24104);
and U27180 (N_27180,N_25182,N_25502);
nand U27181 (N_27181,N_25827,N_25792);
and U27182 (N_27182,N_24166,N_25767);
nor U27183 (N_27183,N_25052,N_24593);
and U27184 (N_27184,N_24157,N_24467);
or U27185 (N_27185,N_24410,N_24236);
or U27186 (N_27186,N_25376,N_24974);
nand U27187 (N_27187,N_25873,N_24117);
or U27188 (N_27188,N_24179,N_25943);
and U27189 (N_27189,N_25567,N_24178);
nor U27190 (N_27190,N_25855,N_24595);
nand U27191 (N_27191,N_24138,N_24619);
and U27192 (N_27192,N_25004,N_25054);
nand U27193 (N_27193,N_25913,N_25155);
xor U27194 (N_27194,N_24947,N_25641);
xor U27195 (N_27195,N_24642,N_24522);
or U27196 (N_27196,N_24633,N_25961);
and U27197 (N_27197,N_25142,N_25995);
or U27198 (N_27198,N_24271,N_24621);
xnor U27199 (N_27199,N_24342,N_25873);
and U27200 (N_27200,N_24734,N_24135);
or U27201 (N_27201,N_25406,N_24485);
nor U27202 (N_27202,N_25162,N_24680);
nor U27203 (N_27203,N_25348,N_25251);
nand U27204 (N_27204,N_25807,N_24933);
xnor U27205 (N_27205,N_24502,N_25006);
nor U27206 (N_27206,N_25247,N_24909);
xor U27207 (N_27207,N_24994,N_24081);
xor U27208 (N_27208,N_24954,N_25197);
and U27209 (N_27209,N_25016,N_24639);
xnor U27210 (N_27210,N_25010,N_25654);
xnor U27211 (N_27211,N_24907,N_24811);
xnor U27212 (N_27212,N_24123,N_25414);
or U27213 (N_27213,N_25147,N_25032);
or U27214 (N_27214,N_24898,N_25820);
nand U27215 (N_27215,N_24177,N_25865);
or U27216 (N_27216,N_25383,N_25975);
xor U27217 (N_27217,N_24462,N_24093);
nor U27218 (N_27218,N_25866,N_25035);
or U27219 (N_27219,N_25456,N_25461);
and U27220 (N_27220,N_25780,N_24288);
nand U27221 (N_27221,N_25762,N_24904);
xnor U27222 (N_27222,N_24959,N_25261);
nor U27223 (N_27223,N_25212,N_24744);
xnor U27224 (N_27224,N_24322,N_25242);
xor U27225 (N_27225,N_25545,N_24007);
xnor U27226 (N_27226,N_25840,N_25766);
nor U27227 (N_27227,N_25017,N_24071);
xnor U27228 (N_27228,N_24277,N_25461);
nor U27229 (N_27229,N_24500,N_24034);
xnor U27230 (N_27230,N_24486,N_24028);
nor U27231 (N_27231,N_24118,N_24789);
or U27232 (N_27232,N_24413,N_25482);
nor U27233 (N_27233,N_25159,N_25059);
and U27234 (N_27234,N_24925,N_25442);
nand U27235 (N_27235,N_25479,N_25282);
or U27236 (N_27236,N_24406,N_24673);
nand U27237 (N_27237,N_24914,N_25570);
xnor U27238 (N_27238,N_25897,N_24068);
xnor U27239 (N_27239,N_24394,N_24529);
or U27240 (N_27240,N_24662,N_24073);
nor U27241 (N_27241,N_24040,N_24520);
or U27242 (N_27242,N_25664,N_24916);
nor U27243 (N_27243,N_24538,N_24492);
nand U27244 (N_27244,N_25465,N_24540);
xor U27245 (N_27245,N_25541,N_24851);
or U27246 (N_27246,N_24106,N_25342);
nor U27247 (N_27247,N_24461,N_25518);
nand U27248 (N_27248,N_25258,N_25888);
or U27249 (N_27249,N_25681,N_25021);
xnor U27250 (N_27250,N_24150,N_24804);
xnor U27251 (N_27251,N_25546,N_25780);
xor U27252 (N_27252,N_24431,N_24065);
nand U27253 (N_27253,N_25844,N_24017);
xor U27254 (N_27254,N_24802,N_24823);
or U27255 (N_27255,N_24032,N_24173);
and U27256 (N_27256,N_24251,N_25576);
nand U27257 (N_27257,N_24076,N_24434);
nand U27258 (N_27258,N_24950,N_24001);
nand U27259 (N_27259,N_25384,N_24070);
nand U27260 (N_27260,N_24175,N_25421);
or U27261 (N_27261,N_24839,N_24615);
and U27262 (N_27262,N_25381,N_24055);
xnor U27263 (N_27263,N_24517,N_25106);
and U27264 (N_27264,N_25591,N_25294);
or U27265 (N_27265,N_24399,N_25776);
xor U27266 (N_27266,N_25734,N_24473);
xnor U27267 (N_27267,N_24957,N_25064);
and U27268 (N_27268,N_24198,N_24181);
nand U27269 (N_27269,N_25995,N_24724);
xor U27270 (N_27270,N_25482,N_25503);
xor U27271 (N_27271,N_24694,N_24916);
nand U27272 (N_27272,N_24143,N_24113);
nor U27273 (N_27273,N_25565,N_24669);
and U27274 (N_27274,N_24195,N_24319);
xnor U27275 (N_27275,N_24960,N_24913);
and U27276 (N_27276,N_24022,N_25520);
or U27277 (N_27277,N_25243,N_24790);
and U27278 (N_27278,N_24669,N_25696);
xor U27279 (N_27279,N_25018,N_25294);
or U27280 (N_27280,N_24655,N_24962);
xnor U27281 (N_27281,N_25819,N_25162);
nand U27282 (N_27282,N_24057,N_24565);
or U27283 (N_27283,N_25903,N_24940);
and U27284 (N_27284,N_24150,N_25124);
nor U27285 (N_27285,N_24993,N_24814);
and U27286 (N_27286,N_25177,N_25536);
nand U27287 (N_27287,N_24858,N_25445);
or U27288 (N_27288,N_24373,N_24110);
xnor U27289 (N_27289,N_24857,N_25470);
nor U27290 (N_27290,N_25302,N_24650);
xor U27291 (N_27291,N_25342,N_24833);
or U27292 (N_27292,N_25640,N_24842);
or U27293 (N_27293,N_25505,N_24830);
nor U27294 (N_27294,N_24262,N_25558);
xnor U27295 (N_27295,N_24724,N_25479);
and U27296 (N_27296,N_25113,N_24505);
xnor U27297 (N_27297,N_25044,N_25339);
or U27298 (N_27298,N_25809,N_25974);
nand U27299 (N_27299,N_24291,N_24363);
or U27300 (N_27300,N_25117,N_25049);
xor U27301 (N_27301,N_24035,N_25926);
nor U27302 (N_27302,N_24876,N_24133);
nor U27303 (N_27303,N_25117,N_25968);
and U27304 (N_27304,N_24652,N_24396);
nand U27305 (N_27305,N_25875,N_25060);
nor U27306 (N_27306,N_25187,N_24701);
or U27307 (N_27307,N_25186,N_25641);
or U27308 (N_27308,N_24602,N_25116);
or U27309 (N_27309,N_25518,N_25459);
or U27310 (N_27310,N_25028,N_25739);
or U27311 (N_27311,N_25512,N_24051);
or U27312 (N_27312,N_24957,N_25564);
or U27313 (N_27313,N_24375,N_25407);
nor U27314 (N_27314,N_24472,N_24865);
xnor U27315 (N_27315,N_24660,N_25875);
xor U27316 (N_27316,N_24538,N_24519);
or U27317 (N_27317,N_25981,N_24504);
or U27318 (N_27318,N_24754,N_25157);
nand U27319 (N_27319,N_24986,N_24794);
nand U27320 (N_27320,N_25992,N_24640);
nand U27321 (N_27321,N_24069,N_25566);
and U27322 (N_27322,N_24498,N_25477);
and U27323 (N_27323,N_25931,N_25995);
and U27324 (N_27324,N_24926,N_25203);
and U27325 (N_27325,N_25547,N_25135);
nor U27326 (N_27326,N_24841,N_24286);
nor U27327 (N_27327,N_24687,N_25174);
nand U27328 (N_27328,N_25071,N_25593);
and U27329 (N_27329,N_25183,N_25885);
and U27330 (N_27330,N_25389,N_24623);
nor U27331 (N_27331,N_25991,N_25402);
nand U27332 (N_27332,N_24989,N_24387);
xnor U27333 (N_27333,N_24572,N_24395);
and U27334 (N_27334,N_24765,N_24929);
xor U27335 (N_27335,N_24293,N_24941);
nor U27336 (N_27336,N_24039,N_25543);
nor U27337 (N_27337,N_24853,N_24680);
or U27338 (N_27338,N_24895,N_25640);
and U27339 (N_27339,N_25745,N_25030);
xor U27340 (N_27340,N_25129,N_25051);
and U27341 (N_27341,N_24519,N_24764);
and U27342 (N_27342,N_25718,N_25372);
nor U27343 (N_27343,N_25235,N_24031);
nand U27344 (N_27344,N_25241,N_24137);
nand U27345 (N_27345,N_25613,N_24714);
nor U27346 (N_27346,N_25051,N_25021);
and U27347 (N_27347,N_24139,N_24178);
nand U27348 (N_27348,N_25051,N_25512);
nor U27349 (N_27349,N_25963,N_25519);
nand U27350 (N_27350,N_25095,N_24671);
or U27351 (N_27351,N_24896,N_24978);
xor U27352 (N_27352,N_24676,N_24213);
nor U27353 (N_27353,N_24686,N_24875);
nor U27354 (N_27354,N_25086,N_24676);
and U27355 (N_27355,N_25973,N_24229);
and U27356 (N_27356,N_24819,N_24062);
and U27357 (N_27357,N_24253,N_24603);
or U27358 (N_27358,N_24315,N_24629);
nand U27359 (N_27359,N_25751,N_24486);
and U27360 (N_27360,N_24509,N_24617);
or U27361 (N_27361,N_24689,N_25647);
nor U27362 (N_27362,N_25420,N_24744);
nor U27363 (N_27363,N_24166,N_24542);
and U27364 (N_27364,N_25628,N_24828);
nand U27365 (N_27365,N_24068,N_24229);
or U27366 (N_27366,N_24905,N_25811);
xnor U27367 (N_27367,N_25914,N_25580);
xor U27368 (N_27368,N_25016,N_24117);
and U27369 (N_27369,N_25410,N_24695);
nand U27370 (N_27370,N_24584,N_25522);
nand U27371 (N_27371,N_24791,N_25454);
and U27372 (N_27372,N_24419,N_24841);
nor U27373 (N_27373,N_25503,N_25310);
and U27374 (N_27374,N_24513,N_25429);
nand U27375 (N_27375,N_24209,N_24236);
or U27376 (N_27376,N_25197,N_24395);
nand U27377 (N_27377,N_25487,N_24900);
xor U27378 (N_27378,N_24982,N_25256);
nor U27379 (N_27379,N_25186,N_24341);
or U27380 (N_27380,N_25197,N_25040);
nand U27381 (N_27381,N_24656,N_24522);
and U27382 (N_27382,N_24553,N_25366);
nor U27383 (N_27383,N_24700,N_25051);
xnor U27384 (N_27384,N_25776,N_25761);
nand U27385 (N_27385,N_25101,N_24600);
nor U27386 (N_27386,N_24176,N_24082);
nand U27387 (N_27387,N_24311,N_24104);
nand U27388 (N_27388,N_25510,N_25519);
and U27389 (N_27389,N_25333,N_25740);
xnor U27390 (N_27390,N_25673,N_24201);
xor U27391 (N_27391,N_24833,N_25850);
nand U27392 (N_27392,N_25674,N_24104);
and U27393 (N_27393,N_25315,N_24469);
nor U27394 (N_27394,N_24091,N_25877);
nand U27395 (N_27395,N_25397,N_24262);
or U27396 (N_27396,N_25077,N_24301);
or U27397 (N_27397,N_24299,N_25123);
xnor U27398 (N_27398,N_24475,N_24209);
nand U27399 (N_27399,N_25008,N_24328);
nor U27400 (N_27400,N_24721,N_25747);
or U27401 (N_27401,N_24875,N_24244);
nand U27402 (N_27402,N_25445,N_24641);
and U27403 (N_27403,N_24380,N_25575);
or U27404 (N_27404,N_25271,N_24902);
nor U27405 (N_27405,N_24977,N_25464);
or U27406 (N_27406,N_24425,N_25451);
xor U27407 (N_27407,N_24078,N_24781);
or U27408 (N_27408,N_24978,N_24374);
nor U27409 (N_27409,N_25699,N_25961);
and U27410 (N_27410,N_25320,N_25962);
and U27411 (N_27411,N_25308,N_25821);
nand U27412 (N_27412,N_24223,N_24542);
nor U27413 (N_27413,N_24138,N_24315);
nor U27414 (N_27414,N_24726,N_25088);
or U27415 (N_27415,N_24001,N_24331);
or U27416 (N_27416,N_25069,N_25929);
nand U27417 (N_27417,N_25244,N_25605);
nand U27418 (N_27418,N_24699,N_24437);
or U27419 (N_27419,N_24042,N_24117);
nand U27420 (N_27420,N_24423,N_25306);
nand U27421 (N_27421,N_25076,N_25393);
and U27422 (N_27422,N_25039,N_24319);
and U27423 (N_27423,N_25240,N_24212);
or U27424 (N_27424,N_25186,N_24706);
or U27425 (N_27425,N_24465,N_25394);
xnor U27426 (N_27426,N_25940,N_24013);
xnor U27427 (N_27427,N_24449,N_24973);
and U27428 (N_27428,N_25050,N_25005);
nor U27429 (N_27429,N_24957,N_25807);
or U27430 (N_27430,N_24558,N_24794);
nand U27431 (N_27431,N_24389,N_24290);
or U27432 (N_27432,N_24692,N_24041);
or U27433 (N_27433,N_25506,N_24855);
nand U27434 (N_27434,N_24368,N_24774);
xor U27435 (N_27435,N_24686,N_25014);
or U27436 (N_27436,N_24679,N_25271);
or U27437 (N_27437,N_25307,N_24871);
xor U27438 (N_27438,N_25790,N_25185);
nor U27439 (N_27439,N_24681,N_25212);
nand U27440 (N_27440,N_24829,N_25193);
xor U27441 (N_27441,N_24787,N_25563);
and U27442 (N_27442,N_25695,N_24811);
nor U27443 (N_27443,N_24983,N_25667);
xnor U27444 (N_27444,N_25950,N_24349);
nor U27445 (N_27445,N_24493,N_24081);
and U27446 (N_27446,N_25752,N_24423);
nand U27447 (N_27447,N_25036,N_25509);
nand U27448 (N_27448,N_25953,N_24198);
and U27449 (N_27449,N_25940,N_24846);
nor U27450 (N_27450,N_25680,N_24056);
nor U27451 (N_27451,N_24331,N_24587);
xnor U27452 (N_27452,N_25376,N_25995);
nand U27453 (N_27453,N_24534,N_24573);
nand U27454 (N_27454,N_24260,N_24206);
xor U27455 (N_27455,N_24292,N_24247);
or U27456 (N_27456,N_24789,N_24360);
nor U27457 (N_27457,N_24934,N_24910);
xor U27458 (N_27458,N_25399,N_25518);
xnor U27459 (N_27459,N_24734,N_25321);
nor U27460 (N_27460,N_25118,N_24857);
or U27461 (N_27461,N_24432,N_24885);
and U27462 (N_27462,N_25369,N_25855);
nand U27463 (N_27463,N_24679,N_25367);
or U27464 (N_27464,N_24929,N_25280);
xnor U27465 (N_27465,N_25083,N_25904);
and U27466 (N_27466,N_25975,N_25781);
xnor U27467 (N_27467,N_24193,N_25018);
and U27468 (N_27468,N_24875,N_24540);
nor U27469 (N_27469,N_24804,N_24638);
and U27470 (N_27470,N_24598,N_25459);
nand U27471 (N_27471,N_24095,N_24244);
xor U27472 (N_27472,N_24184,N_25339);
nor U27473 (N_27473,N_24711,N_24784);
nor U27474 (N_27474,N_25621,N_25383);
nor U27475 (N_27475,N_25852,N_25840);
xnor U27476 (N_27476,N_24820,N_25725);
and U27477 (N_27477,N_24485,N_25089);
nand U27478 (N_27478,N_24299,N_24175);
and U27479 (N_27479,N_25499,N_25678);
and U27480 (N_27480,N_25546,N_24986);
or U27481 (N_27481,N_25735,N_25512);
or U27482 (N_27482,N_25919,N_25303);
xor U27483 (N_27483,N_24038,N_24126);
or U27484 (N_27484,N_24152,N_24920);
or U27485 (N_27485,N_25527,N_25072);
nor U27486 (N_27486,N_25128,N_25098);
xor U27487 (N_27487,N_25050,N_24154);
nand U27488 (N_27488,N_24256,N_25636);
nand U27489 (N_27489,N_24692,N_24903);
nand U27490 (N_27490,N_24389,N_25616);
xor U27491 (N_27491,N_25144,N_25975);
xor U27492 (N_27492,N_25770,N_25866);
or U27493 (N_27493,N_24789,N_25318);
or U27494 (N_27494,N_25290,N_24787);
and U27495 (N_27495,N_25270,N_25929);
nor U27496 (N_27496,N_24969,N_24569);
nor U27497 (N_27497,N_24753,N_25709);
nand U27498 (N_27498,N_24107,N_24993);
nand U27499 (N_27499,N_25516,N_25483);
nor U27500 (N_27500,N_24591,N_25964);
nor U27501 (N_27501,N_25787,N_25701);
and U27502 (N_27502,N_24973,N_24594);
or U27503 (N_27503,N_24982,N_25942);
and U27504 (N_27504,N_24847,N_24170);
nor U27505 (N_27505,N_24771,N_25807);
nand U27506 (N_27506,N_24513,N_24269);
or U27507 (N_27507,N_25593,N_24583);
or U27508 (N_27508,N_24143,N_24259);
or U27509 (N_27509,N_25866,N_25087);
nand U27510 (N_27510,N_25211,N_24934);
nor U27511 (N_27511,N_24242,N_25503);
or U27512 (N_27512,N_25785,N_25214);
or U27513 (N_27513,N_25962,N_25176);
and U27514 (N_27514,N_24261,N_24942);
xnor U27515 (N_27515,N_25231,N_24494);
nand U27516 (N_27516,N_24220,N_24651);
or U27517 (N_27517,N_24246,N_25926);
nand U27518 (N_27518,N_25756,N_24967);
nor U27519 (N_27519,N_25449,N_25419);
nand U27520 (N_27520,N_25049,N_24592);
or U27521 (N_27521,N_25992,N_25402);
or U27522 (N_27522,N_25008,N_25546);
or U27523 (N_27523,N_25441,N_24263);
nand U27524 (N_27524,N_24633,N_24910);
nand U27525 (N_27525,N_25034,N_24722);
nand U27526 (N_27526,N_24811,N_25301);
xnor U27527 (N_27527,N_25760,N_25547);
or U27528 (N_27528,N_24617,N_25648);
nor U27529 (N_27529,N_24923,N_24076);
nor U27530 (N_27530,N_25946,N_25677);
nand U27531 (N_27531,N_25431,N_24325);
or U27532 (N_27532,N_24480,N_24508);
nor U27533 (N_27533,N_24266,N_24374);
xor U27534 (N_27534,N_24997,N_24127);
nand U27535 (N_27535,N_24959,N_25435);
nor U27536 (N_27536,N_25345,N_25879);
and U27537 (N_27537,N_25014,N_24254);
nand U27538 (N_27538,N_24485,N_24423);
xor U27539 (N_27539,N_24266,N_24976);
nand U27540 (N_27540,N_25514,N_25652);
or U27541 (N_27541,N_24015,N_25863);
and U27542 (N_27542,N_24364,N_24515);
nand U27543 (N_27543,N_24226,N_24044);
xor U27544 (N_27544,N_25669,N_24285);
nor U27545 (N_27545,N_25292,N_24027);
xor U27546 (N_27546,N_24326,N_24669);
or U27547 (N_27547,N_25185,N_25044);
and U27548 (N_27548,N_24484,N_25526);
nor U27549 (N_27549,N_25779,N_25318);
xor U27550 (N_27550,N_24298,N_24312);
nand U27551 (N_27551,N_24852,N_25053);
xor U27552 (N_27552,N_24407,N_24854);
nand U27553 (N_27553,N_24358,N_24806);
and U27554 (N_27554,N_25889,N_25401);
xor U27555 (N_27555,N_25548,N_25418);
nand U27556 (N_27556,N_25296,N_24909);
nor U27557 (N_27557,N_25474,N_25770);
xnor U27558 (N_27558,N_25268,N_24719);
xnor U27559 (N_27559,N_25014,N_25902);
nor U27560 (N_27560,N_24394,N_25656);
nand U27561 (N_27561,N_25133,N_25426);
nand U27562 (N_27562,N_24948,N_24980);
xor U27563 (N_27563,N_24059,N_25267);
nand U27564 (N_27564,N_25818,N_24647);
nor U27565 (N_27565,N_25936,N_25680);
nor U27566 (N_27566,N_25944,N_24421);
and U27567 (N_27567,N_25682,N_25856);
and U27568 (N_27568,N_25862,N_25968);
nand U27569 (N_27569,N_25753,N_25478);
and U27570 (N_27570,N_25746,N_24709);
nor U27571 (N_27571,N_24081,N_25178);
and U27572 (N_27572,N_25127,N_25135);
xnor U27573 (N_27573,N_25736,N_24761);
nor U27574 (N_27574,N_25106,N_25290);
or U27575 (N_27575,N_24463,N_24983);
nand U27576 (N_27576,N_25794,N_24787);
and U27577 (N_27577,N_24499,N_24881);
xnor U27578 (N_27578,N_24221,N_25813);
xor U27579 (N_27579,N_24615,N_24899);
and U27580 (N_27580,N_25532,N_24459);
and U27581 (N_27581,N_25771,N_24538);
or U27582 (N_27582,N_24551,N_25710);
xnor U27583 (N_27583,N_24142,N_25934);
xnor U27584 (N_27584,N_24763,N_25057);
xnor U27585 (N_27585,N_24303,N_25395);
xor U27586 (N_27586,N_24419,N_25923);
and U27587 (N_27587,N_24291,N_25331);
nand U27588 (N_27588,N_24532,N_24400);
nand U27589 (N_27589,N_25416,N_25329);
nor U27590 (N_27590,N_24162,N_25409);
xnor U27591 (N_27591,N_25773,N_25169);
or U27592 (N_27592,N_25988,N_24593);
and U27593 (N_27593,N_25863,N_25048);
nand U27594 (N_27594,N_24455,N_25949);
nor U27595 (N_27595,N_25508,N_25836);
nand U27596 (N_27596,N_25584,N_25608);
and U27597 (N_27597,N_24209,N_24523);
or U27598 (N_27598,N_25165,N_24736);
xnor U27599 (N_27599,N_24802,N_25701);
nand U27600 (N_27600,N_25199,N_24267);
nand U27601 (N_27601,N_25441,N_24420);
nor U27602 (N_27602,N_25113,N_25347);
nand U27603 (N_27603,N_25962,N_25267);
or U27604 (N_27604,N_25169,N_25798);
nand U27605 (N_27605,N_24983,N_24549);
and U27606 (N_27606,N_24422,N_24830);
or U27607 (N_27607,N_25432,N_25874);
and U27608 (N_27608,N_25655,N_25402);
nor U27609 (N_27609,N_24069,N_24920);
and U27610 (N_27610,N_25190,N_25179);
xnor U27611 (N_27611,N_24648,N_25940);
nor U27612 (N_27612,N_25988,N_25135);
and U27613 (N_27613,N_24527,N_24897);
nor U27614 (N_27614,N_25202,N_25054);
and U27615 (N_27615,N_24690,N_25544);
nand U27616 (N_27616,N_24892,N_25968);
nor U27617 (N_27617,N_25619,N_25358);
nor U27618 (N_27618,N_24152,N_24868);
and U27619 (N_27619,N_25213,N_24997);
nand U27620 (N_27620,N_25379,N_25941);
or U27621 (N_27621,N_25918,N_24315);
xnor U27622 (N_27622,N_25889,N_25659);
xnor U27623 (N_27623,N_25479,N_24960);
nand U27624 (N_27624,N_24148,N_24371);
xnor U27625 (N_27625,N_24696,N_25322);
xnor U27626 (N_27626,N_25081,N_25260);
nand U27627 (N_27627,N_25444,N_24226);
and U27628 (N_27628,N_24818,N_25970);
xnor U27629 (N_27629,N_25829,N_24028);
nor U27630 (N_27630,N_24410,N_24466);
xor U27631 (N_27631,N_25259,N_24822);
xnor U27632 (N_27632,N_24819,N_25879);
xnor U27633 (N_27633,N_25896,N_25354);
xnor U27634 (N_27634,N_25985,N_24436);
and U27635 (N_27635,N_25019,N_24487);
or U27636 (N_27636,N_25400,N_25195);
nor U27637 (N_27637,N_24245,N_25743);
nand U27638 (N_27638,N_25819,N_25233);
nor U27639 (N_27639,N_24511,N_24676);
nor U27640 (N_27640,N_24340,N_24693);
and U27641 (N_27641,N_25764,N_25185);
nand U27642 (N_27642,N_25657,N_24134);
nand U27643 (N_27643,N_24860,N_25569);
and U27644 (N_27644,N_25461,N_25222);
nand U27645 (N_27645,N_25960,N_25991);
nand U27646 (N_27646,N_25045,N_24764);
xnor U27647 (N_27647,N_24760,N_24021);
or U27648 (N_27648,N_25717,N_24405);
or U27649 (N_27649,N_25052,N_25983);
nand U27650 (N_27650,N_24755,N_24426);
nand U27651 (N_27651,N_24996,N_25355);
nor U27652 (N_27652,N_24726,N_25246);
nand U27653 (N_27653,N_24758,N_25559);
xnor U27654 (N_27654,N_24859,N_24342);
nand U27655 (N_27655,N_24763,N_24396);
and U27656 (N_27656,N_24343,N_24648);
xnor U27657 (N_27657,N_25085,N_24889);
xnor U27658 (N_27658,N_25948,N_24285);
and U27659 (N_27659,N_25477,N_24704);
xor U27660 (N_27660,N_24148,N_24146);
and U27661 (N_27661,N_24088,N_25228);
nor U27662 (N_27662,N_25224,N_24448);
nor U27663 (N_27663,N_24380,N_24327);
nor U27664 (N_27664,N_24663,N_25807);
nor U27665 (N_27665,N_25309,N_24487);
nor U27666 (N_27666,N_24281,N_24235);
or U27667 (N_27667,N_25720,N_24782);
or U27668 (N_27668,N_25033,N_24133);
or U27669 (N_27669,N_25186,N_24512);
nor U27670 (N_27670,N_24461,N_24147);
nand U27671 (N_27671,N_24436,N_24176);
nand U27672 (N_27672,N_24775,N_25204);
nand U27673 (N_27673,N_25974,N_25166);
nor U27674 (N_27674,N_24360,N_25487);
nor U27675 (N_27675,N_25583,N_24835);
nor U27676 (N_27676,N_25982,N_24708);
nand U27677 (N_27677,N_25030,N_24696);
xnor U27678 (N_27678,N_24831,N_24700);
nand U27679 (N_27679,N_25670,N_24671);
xor U27680 (N_27680,N_24483,N_25231);
xnor U27681 (N_27681,N_24335,N_24777);
or U27682 (N_27682,N_24120,N_25707);
nor U27683 (N_27683,N_24040,N_24405);
nor U27684 (N_27684,N_25996,N_25741);
and U27685 (N_27685,N_24130,N_25234);
or U27686 (N_27686,N_24067,N_25876);
nand U27687 (N_27687,N_24382,N_24057);
and U27688 (N_27688,N_25812,N_25210);
and U27689 (N_27689,N_24121,N_24620);
xnor U27690 (N_27690,N_25401,N_24173);
or U27691 (N_27691,N_24665,N_24018);
nand U27692 (N_27692,N_25898,N_24418);
and U27693 (N_27693,N_25338,N_25292);
xor U27694 (N_27694,N_25382,N_24000);
or U27695 (N_27695,N_25227,N_24428);
nand U27696 (N_27696,N_25403,N_24610);
or U27697 (N_27697,N_24149,N_25500);
nand U27698 (N_27698,N_25843,N_25107);
nor U27699 (N_27699,N_24236,N_25729);
or U27700 (N_27700,N_25339,N_24812);
and U27701 (N_27701,N_24268,N_24723);
and U27702 (N_27702,N_25476,N_25345);
nand U27703 (N_27703,N_24750,N_25492);
xor U27704 (N_27704,N_24512,N_24105);
xor U27705 (N_27705,N_24166,N_25172);
nor U27706 (N_27706,N_24687,N_24278);
xor U27707 (N_27707,N_24942,N_24702);
or U27708 (N_27708,N_25059,N_25097);
nand U27709 (N_27709,N_25602,N_24867);
or U27710 (N_27710,N_24107,N_24482);
nor U27711 (N_27711,N_25216,N_25777);
xor U27712 (N_27712,N_25336,N_25350);
nor U27713 (N_27713,N_24634,N_24425);
xor U27714 (N_27714,N_25373,N_24703);
or U27715 (N_27715,N_25717,N_24057);
xnor U27716 (N_27716,N_24149,N_24208);
nor U27717 (N_27717,N_25541,N_25786);
and U27718 (N_27718,N_25737,N_24825);
nand U27719 (N_27719,N_25601,N_24202);
xor U27720 (N_27720,N_25809,N_25191);
or U27721 (N_27721,N_24255,N_24311);
nor U27722 (N_27722,N_25785,N_25614);
xnor U27723 (N_27723,N_24994,N_24803);
nor U27724 (N_27724,N_25254,N_24560);
nor U27725 (N_27725,N_25431,N_24674);
and U27726 (N_27726,N_25794,N_24780);
and U27727 (N_27727,N_24949,N_25519);
or U27728 (N_27728,N_25731,N_24511);
nand U27729 (N_27729,N_25996,N_25021);
nand U27730 (N_27730,N_25448,N_25896);
nor U27731 (N_27731,N_24131,N_24545);
nand U27732 (N_27732,N_24290,N_25098);
and U27733 (N_27733,N_25744,N_25844);
nand U27734 (N_27734,N_25132,N_25424);
and U27735 (N_27735,N_24877,N_24628);
nor U27736 (N_27736,N_25673,N_25724);
and U27737 (N_27737,N_24916,N_24508);
nor U27738 (N_27738,N_25859,N_24916);
nand U27739 (N_27739,N_25394,N_24033);
and U27740 (N_27740,N_24814,N_25096);
and U27741 (N_27741,N_24334,N_25594);
nor U27742 (N_27742,N_25302,N_24064);
and U27743 (N_27743,N_25595,N_25813);
nor U27744 (N_27744,N_24518,N_24931);
nand U27745 (N_27745,N_25178,N_25222);
and U27746 (N_27746,N_25287,N_25211);
nor U27747 (N_27747,N_24754,N_24019);
nor U27748 (N_27748,N_24170,N_24618);
nand U27749 (N_27749,N_25404,N_24282);
or U27750 (N_27750,N_25444,N_25282);
xor U27751 (N_27751,N_25301,N_24938);
and U27752 (N_27752,N_25552,N_24576);
nand U27753 (N_27753,N_24313,N_25444);
and U27754 (N_27754,N_24780,N_25318);
or U27755 (N_27755,N_25431,N_24704);
and U27756 (N_27756,N_24842,N_24458);
nand U27757 (N_27757,N_24622,N_25720);
nand U27758 (N_27758,N_25556,N_24015);
or U27759 (N_27759,N_25725,N_25708);
or U27760 (N_27760,N_25186,N_24271);
and U27761 (N_27761,N_25624,N_24244);
or U27762 (N_27762,N_25689,N_25612);
nor U27763 (N_27763,N_25446,N_25898);
nor U27764 (N_27764,N_24731,N_24910);
xor U27765 (N_27765,N_24778,N_24533);
and U27766 (N_27766,N_24416,N_25064);
xnor U27767 (N_27767,N_24241,N_24510);
and U27768 (N_27768,N_25354,N_24491);
nor U27769 (N_27769,N_25368,N_25951);
or U27770 (N_27770,N_25645,N_25154);
or U27771 (N_27771,N_25331,N_25080);
or U27772 (N_27772,N_24822,N_25101);
and U27773 (N_27773,N_25311,N_24365);
or U27774 (N_27774,N_24152,N_25505);
nand U27775 (N_27775,N_25900,N_25737);
xor U27776 (N_27776,N_24049,N_24896);
nor U27777 (N_27777,N_25845,N_24940);
nor U27778 (N_27778,N_24241,N_25289);
and U27779 (N_27779,N_24881,N_24005);
nor U27780 (N_27780,N_24821,N_24695);
nor U27781 (N_27781,N_25347,N_24343);
nor U27782 (N_27782,N_25099,N_25346);
xor U27783 (N_27783,N_25807,N_24928);
xor U27784 (N_27784,N_25248,N_25165);
or U27785 (N_27785,N_24542,N_25953);
nand U27786 (N_27786,N_25523,N_25326);
or U27787 (N_27787,N_24835,N_24269);
and U27788 (N_27788,N_25390,N_24808);
and U27789 (N_27789,N_24270,N_24791);
nor U27790 (N_27790,N_25396,N_25033);
nand U27791 (N_27791,N_25044,N_25810);
or U27792 (N_27792,N_25204,N_24068);
xor U27793 (N_27793,N_24185,N_24757);
or U27794 (N_27794,N_25326,N_24243);
nand U27795 (N_27795,N_25619,N_25242);
and U27796 (N_27796,N_25619,N_24675);
xnor U27797 (N_27797,N_24632,N_24747);
xnor U27798 (N_27798,N_24311,N_25545);
and U27799 (N_27799,N_24458,N_24393);
nand U27800 (N_27800,N_24245,N_25737);
xnor U27801 (N_27801,N_24254,N_25974);
or U27802 (N_27802,N_24512,N_25626);
nand U27803 (N_27803,N_25131,N_24521);
and U27804 (N_27804,N_24958,N_25357);
nand U27805 (N_27805,N_24310,N_24121);
xnor U27806 (N_27806,N_24554,N_25017);
xnor U27807 (N_27807,N_24712,N_25862);
and U27808 (N_27808,N_25707,N_25411);
xnor U27809 (N_27809,N_24685,N_25527);
nand U27810 (N_27810,N_25864,N_25849);
xor U27811 (N_27811,N_24703,N_25780);
xor U27812 (N_27812,N_25961,N_25231);
nand U27813 (N_27813,N_24478,N_24574);
and U27814 (N_27814,N_24002,N_24000);
or U27815 (N_27815,N_25091,N_25112);
nand U27816 (N_27816,N_24518,N_24422);
and U27817 (N_27817,N_24442,N_25528);
nand U27818 (N_27818,N_24889,N_24672);
nand U27819 (N_27819,N_24531,N_24841);
xnor U27820 (N_27820,N_24103,N_24946);
or U27821 (N_27821,N_25697,N_24892);
or U27822 (N_27822,N_25209,N_24674);
nand U27823 (N_27823,N_24184,N_25374);
xnor U27824 (N_27824,N_24436,N_24150);
nor U27825 (N_27825,N_24814,N_24414);
nor U27826 (N_27826,N_25944,N_24772);
nand U27827 (N_27827,N_24113,N_25084);
nand U27828 (N_27828,N_24457,N_25068);
or U27829 (N_27829,N_24701,N_25488);
xnor U27830 (N_27830,N_24563,N_24214);
or U27831 (N_27831,N_25369,N_24424);
or U27832 (N_27832,N_25000,N_25066);
nand U27833 (N_27833,N_24532,N_25292);
nand U27834 (N_27834,N_25119,N_24071);
nand U27835 (N_27835,N_24837,N_24731);
and U27836 (N_27836,N_25467,N_24263);
nor U27837 (N_27837,N_25938,N_25633);
xnor U27838 (N_27838,N_25671,N_24085);
or U27839 (N_27839,N_24770,N_25467);
xor U27840 (N_27840,N_24744,N_24054);
nor U27841 (N_27841,N_25182,N_24388);
or U27842 (N_27842,N_25631,N_24971);
xnor U27843 (N_27843,N_24301,N_25954);
nand U27844 (N_27844,N_25047,N_24239);
xor U27845 (N_27845,N_24692,N_25016);
or U27846 (N_27846,N_24489,N_24001);
xnor U27847 (N_27847,N_25474,N_25561);
and U27848 (N_27848,N_24897,N_24576);
and U27849 (N_27849,N_24155,N_25142);
nand U27850 (N_27850,N_25989,N_24604);
nor U27851 (N_27851,N_24636,N_25258);
nand U27852 (N_27852,N_24297,N_24632);
nor U27853 (N_27853,N_24181,N_24672);
and U27854 (N_27854,N_25959,N_24505);
xnor U27855 (N_27855,N_25410,N_25248);
xor U27856 (N_27856,N_24941,N_25809);
nand U27857 (N_27857,N_24261,N_24359);
or U27858 (N_27858,N_25392,N_24086);
xor U27859 (N_27859,N_24377,N_25908);
or U27860 (N_27860,N_24092,N_25731);
and U27861 (N_27861,N_24352,N_24205);
nor U27862 (N_27862,N_25592,N_25015);
xor U27863 (N_27863,N_24677,N_25189);
nand U27864 (N_27864,N_25352,N_25576);
nor U27865 (N_27865,N_25473,N_25119);
xor U27866 (N_27866,N_25463,N_25250);
or U27867 (N_27867,N_24353,N_25634);
nand U27868 (N_27868,N_25028,N_24231);
and U27869 (N_27869,N_24086,N_24449);
nor U27870 (N_27870,N_24449,N_24823);
xor U27871 (N_27871,N_25309,N_25164);
nor U27872 (N_27872,N_25242,N_24804);
xor U27873 (N_27873,N_24934,N_24418);
or U27874 (N_27874,N_24733,N_25731);
and U27875 (N_27875,N_25736,N_25533);
xor U27876 (N_27876,N_24880,N_25523);
nor U27877 (N_27877,N_25303,N_25458);
nor U27878 (N_27878,N_24157,N_24062);
and U27879 (N_27879,N_24126,N_24193);
or U27880 (N_27880,N_25833,N_24650);
nand U27881 (N_27881,N_24259,N_24978);
nand U27882 (N_27882,N_25004,N_24748);
nand U27883 (N_27883,N_25945,N_24058);
or U27884 (N_27884,N_24836,N_24589);
or U27885 (N_27885,N_24720,N_25950);
nor U27886 (N_27886,N_25457,N_25254);
nor U27887 (N_27887,N_24216,N_25435);
nand U27888 (N_27888,N_25796,N_24678);
nor U27889 (N_27889,N_25148,N_24045);
xor U27890 (N_27890,N_25507,N_25151);
nand U27891 (N_27891,N_24058,N_24153);
nor U27892 (N_27892,N_25044,N_24722);
xor U27893 (N_27893,N_24152,N_25849);
xor U27894 (N_27894,N_25136,N_24453);
or U27895 (N_27895,N_24720,N_25560);
xnor U27896 (N_27896,N_24966,N_25887);
xor U27897 (N_27897,N_24158,N_24915);
or U27898 (N_27898,N_25950,N_25056);
and U27899 (N_27899,N_25138,N_25264);
or U27900 (N_27900,N_25528,N_25998);
and U27901 (N_27901,N_25057,N_25277);
and U27902 (N_27902,N_25538,N_24113);
or U27903 (N_27903,N_25919,N_25569);
xor U27904 (N_27904,N_25495,N_25218);
nand U27905 (N_27905,N_25683,N_25951);
nand U27906 (N_27906,N_25112,N_25904);
nand U27907 (N_27907,N_25415,N_25707);
nor U27908 (N_27908,N_24898,N_24972);
and U27909 (N_27909,N_25615,N_25298);
nand U27910 (N_27910,N_25328,N_25204);
nand U27911 (N_27911,N_24945,N_25093);
nor U27912 (N_27912,N_25903,N_25973);
xnor U27913 (N_27913,N_24537,N_25168);
nor U27914 (N_27914,N_24114,N_25369);
nor U27915 (N_27915,N_24989,N_25859);
and U27916 (N_27916,N_25920,N_25996);
xor U27917 (N_27917,N_24786,N_25524);
and U27918 (N_27918,N_25575,N_24678);
nand U27919 (N_27919,N_25029,N_24673);
and U27920 (N_27920,N_25989,N_25623);
and U27921 (N_27921,N_24587,N_24633);
nor U27922 (N_27922,N_25149,N_24086);
xor U27923 (N_27923,N_24433,N_25276);
and U27924 (N_27924,N_25035,N_25557);
and U27925 (N_27925,N_25098,N_25379);
and U27926 (N_27926,N_25029,N_24426);
or U27927 (N_27927,N_24162,N_24582);
nand U27928 (N_27928,N_25404,N_25646);
xor U27929 (N_27929,N_25655,N_25296);
nor U27930 (N_27930,N_25955,N_25864);
nor U27931 (N_27931,N_25877,N_25816);
nand U27932 (N_27932,N_25997,N_25130);
xor U27933 (N_27933,N_24213,N_25997);
and U27934 (N_27934,N_25720,N_25847);
nor U27935 (N_27935,N_25291,N_25089);
or U27936 (N_27936,N_25329,N_25836);
nand U27937 (N_27937,N_24816,N_25334);
xnor U27938 (N_27938,N_24836,N_24700);
nor U27939 (N_27939,N_24081,N_24632);
or U27940 (N_27940,N_24200,N_25417);
or U27941 (N_27941,N_24114,N_25248);
and U27942 (N_27942,N_24494,N_25557);
and U27943 (N_27943,N_25507,N_24336);
and U27944 (N_27944,N_25791,N_25421);
xor U27945 (N_27945,N_25105,N_24797);
and U27946 (N_27946,N_24380,N_24128);
nand U27947 (N_27947,N_24035,N_24424);
xor U27948 (N_27948,N_24512,N_25846);
xnor U27949 (N_27949,N_25135,N_25518);
xor U27950 (N_27950,N_24014,N_24332);
or U27951 (N_27951,N_24467,N_24485);
and U27952 (N_27952,N_25320,N_25155);
xnor U27953 (N_27953,N_25082,N_25939);
xnor U27954 (N_27954,N_24160,N_25458);
xnor U27955 (N_27955,N_25213,N_24153);
or U27956 (N_27956,N_25602,N_25413);
nor U27957 (N_27957,N_25023,N_25829);
and U27958 (N_27958,N_25254,N_25236);
nand U27959 (N_27959,N_25846,N_24030);
xnor U27960 (N_27960,N_25683,N_25412);
xnor U27961 (N_27961,N_24175,N_24885);
nand U27962 (N_27962,N_25514,N_25322);
xor U27963 (N_27963,N_25358,N_24204);
nor U27964 (N_27964,N_24575,N_25427);
and U27965 (N_27965,N_25635,N_25674);
xor U27966 (N_27966,N_25099,N_24672);
nor U27967 (N_27967,N_25073,N_24614);
xor U27968 (N_27968,N_24187,N_24221);
xnor U27969 (N_27969,N_25587,N_24817);
nand U27970 (N_27970,N_24582,N_24361);
nor U27971 (N_27971,N_25674,N_24881);
xor U27972 (N_27972,N_25835,N_25779);
nor U27973 (N_27973,N_25797,N_24259);
xnor U27974 (N_27974,N_24494,N_25856);
nand U27975 (N_27975,N_24216,N_24853);
and U27976 (N_27976,N_24247,N_25206);
xnor U27977 (N_27977,N_24647,N_25866);
and U27978 (N_27978,N_25739,N_25947);
nand U27979 (N_27979,N_25627,N_24743);
xnor U27980 (N_27980,N_25333,N_25063);
xor U27981 (N_27981,N_24119,N_25874);
nand U27982 (N_27982,N_24610,N_25253);
and U27983 (N_27983,N_24219,N_25056);
nand U27984 (N_27984,N_24449,N_25523);
or U27985 (N_27985,N_24210,N_24999);
xor U27986 (N_27986,N_24518,N_25917);
and U27987 (N_27987,N_25269,N_24786);
xor U27988 (N_27988,N_24062,N_24094);
xnor U27989 (N_27989,N_24903,N_24508);
nand U27990 (N_27990,N_25551,N_25853);
and U27991 (N_27991,N_25373,N_25098);
nor U27992 (N_27992,N_25868,N_24910);
nand U27993 (N_27993,N_24743,N_25479);
nand U27994 (N_27994,N_24798,N_24344);
nor U27995 (N_27995,N_25142,N_25127);
xnor U27996 (N_27996,N_25278,N_24784);
nand U27997 (N_27997,N_24745,N_25854);
nor U27998 (N_27998,N_25846,N_25447);
or U27999 (N_27999,N_24304,N_25437);
or U28000 (N_28000,N_26960,N_26671);
xnor U28001 (N_28001,N_26182,N_27222);
nand U28002 (N_28002,N_26279,N_26870);
or U28003 (N_28003,N_26504,N_27395);
and U28004 (N_28004,N_27279,N_27541);
or U28005 (N_28005,N_27420,N_26029);
nor U28006 (N_28006,N_27740,N_27250);
xor U28007 (N_28007,N_26146,N_27717);
or U28008 (N_28008,N_26933,N_27559);
nor U28009 (N_28009,N_27406,N_27366);
nand U28010 (N_28010,N_27630,N_26784);
xnor U28011 (N_28011,N_26667,N_26977);
xnor U28012 (N_28012,N_26908,N_27381);
nand U28013 (N_28013,N_26253,N_27453);
xnor U28014 (N_28014,N_26650,N_27493);
nor U28015 (N_28015,N_26570,N_26392);
nor U28016 (N_28016,N_26345,N_27735);
xnor U28017 (N_28017,N_27842,N_26724);
nor U28018 (N_28018,N_27326,N_26987);
nand U28019 (N_28019,N_27462,N_26705);
nand U28020 (N_28020,N_27027,N_26357);
or U28021 (N_28021,N_27747,N_27286);
xnor U28022 (N_28022,N_26626,N_27751);
xor U28023 (N_28023,N_27107,N_27074);
xnor U28024 (N_28024,N_27860,N_26301);
xor U28025 (N_28025,N_27321,N_27430);
xor U28026 (N_28026,N_26553,N_27861);
xor U28027 (N_28027,N_27772,N_27543);
or U28028 (N_28028,N_26482,N_26444);
nor U28029 (N_28029,N_27606,N_27376);
xnor U28030 (N_28030,N_27216,N_27020);
nor U28031 (N_28031,N_27973,N_27203);
or U28032 (N_28032,N_27716,N_26600);
xnor U28033 (N_28033,N_26715,N_26419);
nor U28034 (N_28034,N_27707,N_27007);
nor U28035 (N_28035,N_26965,N_27658);
nand U28036 (N_28036,N_27583,N_27648);
nand U28037 (N_28037,N_27136,N_27334);
or U28038 (N_28038,N_26718,N_26922);
xnor U28039 (N_28039,N_26354,N_27210);
nor U28040 (N_28040,N_27387,N_27417);
or U28041 (N_28041,N_26223,N_27053);
xor U28042 (N_28042,N_27487,N_27498);
nor U28043 (N_28043,N_26390,N_27758);
xnor U28044 (N_28044,N_27674,N_26575);
nor U28045 (N_28045,N_27356,N_26101);
and U28046 (N_28046,N_26951,N_26537);
nor U28047 (N_28047,N_26347,N_27358);
nor U28048 (N_28048,N_26231,N_27185);
nor U28049 (N_28049,N_26215,N_26610);
or U28050 (N_28050,N_26837,N_27383);
xnor U28051 (N_28051,N_27433,N_27613);
nor U28052 (N_28052,N_27525,N_27838);
or U28053 (N_28053,N_26308,N_26814);
nand U28054 (N_28054,N_27934,N_26596);
nand U28055 (N_28055,N_27299,N_26425);
xnor U28056 (N_28056,N_26720,N_27204);
or U28057 (N_28057,N_26636,N_27470);
nand U28058 (N_28058,N_27284,N_26020);
nand U28059 (N_28059,N_26561,N_27260);
nand U28060 (N_28060,N_27659,N_26394);
or U28061 (N_28061,N_27983,N_27783);
nor U28062 (N_28062,N_27790,N_26976);
and U28063 (N_28063,N_26689,N_26435);
or U28064 (N_28064,N_26080,N_26518);
nor U28065 (N_28065,N_27837,N_26205);
and U28066 (N_28066,N_27705,N_27480);
nand U28067 (N_28067,N_27925,N_26142);
nand U28068 (N_28068,N_27815,N_26663);
nand U28069 (N_28069,N_27598,N_27290);
nand U28070 (N_28070,N_27845,N_26361);
and U28071 (N_28071,N_26487,N_27823);
xor U28072 (N_28072,N_26500,N_27155);
or U28073 (N_28073,N_27930,N_26754);
or U28074 (N_28074,N_26240,N_26796);
and U28075 (N_28075,N_26386,N_27411);
xor U28076 (N_28076,N_26370,N_26547);
nand U28077 (N_28077,N_26203,N_26753);
or U28078 (N_28078,N_26676,N_27414);
nor U28079 (N_28079,N_27229,N_27832);
and U28080 (N_28080,N_27856,N_27643);
xor U28081 (N_28081,N_26198,N_26767);
nor U28082 (N_28082,N_27288,N_27004);
xnor U28083 (N_28083,N_27562,N_26298);
nand U28084 (N_28084,N_26766,N_26191);
or U28085 (N_28085,N_26768,N_26373);
xnor U28086 (N_28086,N_26700,N_27574);
xor U28087 (N_28087,N_27786,N_26632);
nand U28088 (N_28088,N_26092,N_27446);
or U28089 (N_28089,N_27901,N_26963);
nor U28090 (N_28090,N_27087,N_26611);
nand U28091 (N_28091,N_26804,N_27197);
nand U28092 (N_28092,N_27324,N_26272);
and U28093 (N_28093,N_27784,N_26004);
xnor U28094 (N_28094,N_26103,N_27548);
nand U28095 (N_28095,N_27370,N_27371);
nand U28096 (N_28096,N_26929,N_27465);
or U28097 (N_28097,N_26845,N_26384);
nand U28098 (N_28098,N_27443,N_26986);
nor U28099 (N_28099,N_26839,N_27103);
xor U28100 (N_28100,N_27367,N_27677);
and U28101 (N_28101,N_27173,N_27967);
and U28102 (N_28102,N_26809,N_26056);
nand U28103 (N_28103,N_26590,N_27280);
and U28104 (N_28104,N_27137,N_27424);
xor U28105 (N_28105,N_26218,N_27228);
or U28106 (N_28106,N_27911,N_26902);
nand U28107 (N_28107,N_26260,N_27187);
nor U28108 (N_28108,N_27265,N_27186);
or U28109 (N_28109,N_26037,N_26116);
nor U28110 (N_28110,N_27746,N_26434);
or U28111 (N_28111,N_26359,N_27866);
xor U28112 (N_28112,N_26981,N_27209);
nor U28113 (N_28113,N_27850,N_26888);
nand U28114 (N_28114,N_26675,N_27252);
nor U28115 (N_28115,N_26057,N_26463);
and U28116 (N_28116,N_26199,N_26014);
nor U28117 (N_28117,N_26395,N_26009);
xnor U28118 (N_28118,N_26582,N_26498);
xnor U28119 (N_28119,N_27890,N_27205);
xor U28120 (N_28120,N_26196,N_26466);
xnor U28121 (N_28121,N_26710,N_26073);
or U28122 (N_28122,N_27078,N_26880);
or U28123 (N_28123,N_26366,N_27932);
or U28124 (N_28124,N_26916,N_26643);
and U28125 (N_28125,N_27661,N_27870);
nand U28126 (N_28126,N_26488,N_27323);
or U28127 (N_28127,N_26524,N_27322);
or U28128 (N_28128,N_26085,N_26641);
nor U28129 (N_28129,N_27935,N_26138);
or U28130 (N_28130,N_26033,N_27234);
nor U28131 (N_28131,N_27499,N_26712);
xor U28132 (N_28132,N_27627,N_27211);
xnor U28133 (N_28133,N_27615,N_27245);
xor U28134 (N_28134,N_27879,N_26648);
nand U28135 (N_28135,N_26040,N_27949);
and U28136 (N_28136,N_27928,N_26564);
xor U28137 (N_28137,N_26858,N_26380);
and U28138 (N_28138,N_26584,N_27361);
and U28139 (N_28139,N_26213,N_26343);
nor U28140 (N_28140,N_27695,N_26999);
nand U28141 (N_28141,N_26782,N_27782);
nor U28142 (N_28142,N_27638,N_26789);
nand U28143 (N_28143,N_27828,N_26525);
nand U28144 (N_28144,N_27343,N_27033);
or U28145 (N_28145,N_26065,N_27120);
nor U28146 (N_28146,N_26995,N_26304);
nor U28147 (N_28147,N_26252,N_27877);
and U28148 (N_28148,N_26911,N_27202);
and U28149 (N_28149,N_26521,N_27475);
nand U28150 (N_28150,N_26688,N_26467);
and U28151 (N_28151,N_26595,N_27984);
nand U28152 (N_28152,N_26744,N_27628);
nor U28153 (N_28153,N_26277,N_27864);
and U28154 (N_28154,N_27161,N_27089);
and U28155 (N_28155,N_26907,N_27626);
and U28156 (N_28156,N_27633,N_26083);
nand U28157 (N_28157,N_26428,N_27251);
nor U28158 (N_28158,N_26098,N_26447);
xnor U28159 (N_28159,N_26980,N_26456);
nor U28160 (N_28160,N_26638,N_27226);
or U28161 (N_28161,N_27671,N_27513);
or U28162 (N_28162,N_26137,N_26317);
xnor U28163 (N_28163,N_26257,N_26674);
xnor U28164 (N_28164,N_26235,N_26315);
xnor U28165 (N_28165,N_27408,N_27987);
nand U28166 (N_28166,N_27486,N_27409);
nor U28167 (N_28167,N_27594,N_26574);
nor U28168 (N_28168,N_26226,N_27821);
or U28169 (N_28169,N_27804,N_26221);
xnor U28170 (N_28170,N_27785,N_27913);
and U28171 (N_28171,N_26740,N_27142);
nor U28172 (N_28172,N_27360,N_27494);
xnor U28173 (N_28173,N_27457,N_27561);
xor U28174 (N_28174,N_26531,N_27311);
nand U28175 (N_28175,N_26241,N_27773);
and U28176 (N_28176,N_27884,N_26850);
nand U28177 (N_28177,N_26925,N_27237);
nand U28178 (N_28178,N_27188,N_26418);
xnor U28179 (N_28179,N_26751,N_27725);
and U28180 (N_28180,N_26312,N_27506);
nand U28181 (N_28181,N_27015,N_26421);
and U28182 (N_28182,N_26602,N_27741);
nor U28183 (N_28183,N_27581,N_26285);
nand U28184 (N_28184,N_27254,N_27176);
nand U28185 (N_28185,N_26451,N_26422);
nand U28186 (N_28186,N_27110,N_26687);
or U28187 (N_28187,N_26058,N_27421);
xor U28188 (N_28188,N_26708,N_26681);
or U28189 (N_28189,N_27143,N_26779);
and U28190 (N_28190,N_26352,N_27950);
nor U28191 (N_28191,N_27082,N_27545);
or U28192 (N_28192,N_27327,N_27748);
xor U28193 (N_28193,N_26350,N_26338);
or U28194 (N_28194,N_26802,N_27029);
or U28195 (N_28195,N_27955,N_27490);
xor U28196 (N_28196,N_26015,N_26480);
nand U28197 (N_28197,N_26898,N_27900);
nand U28198 (N_28198,N_26332,N_27578);
xnor U28199 (N_28199,N_26016,N_26893);
and U28200 (N_28200,N_26078,N_26549);
or U28201 (N_28201,N_26398,N_27129);
nand U28202 (N_28202,N_27798,N_26661);
nand U28203 (N_28203,N_26598,N_27501);
and U28204 (N_28204,N_27463,N_27080);
nor U28205 (N_28205,N_26454,N_27511);
nand U28206 (N_28206,N_27744,N_27102);
and U28207 (N_28207,N_26256,N_26120);
or U28208 (N_28208,N_26523,N_26145);
and U28209 (N_28209,N_27841,N_27694);
xor U28210 (N_28210,N_27704,N_26091);
xnor U28211 (N_28211,N_26382,N_26325);
and U28212 (N_28212,N_26051,N_26852);
xor U28213 (N_28213,N_26946,N_26917);
or U28214 (N_28214,N_27824,N_27172);
xnor U28215 (N_28215,N_27047,N_27055);
nor U28216 (N_28216,N_26247,N_26473);
xnor U28217 (N_28217,N_27422,N_26416);
and U28218 (N_28218,N_27320,N_26627);
nor U28219 (N_28219,N_27384,N_27392);
nand U28220 (N_28220,N_27862,N_26490);
nor U28221 (N_28221,N_26771,N_27757);
or U28222 (N_28222,N_26479,N_26635);
nand U28223 (N_28223,N_26812,N_27650);
nor U28224 (N_28224,N_27914,N_26420);
or U28225 (N_28225,N_26732,N_27907);
or U28226 (N_28226,N_26964,N_26528);
and U28227 (N_28227,N_26748,N_27703);
nand U28228 (N_28228,N_27612,N_27571);
xor U28229 (N_28229,N_26872,N_27374);
and U28230 (N_28230,N_27997,N_26403);
or U28231 (N_28231,N_27912,N_26426);
nand U28232 (N_28232,N_26143,N_26476);
xor U28233 (N_28233,N_26472,N_27607);
nand U28234 (N_28234,N_27037,N_27419);
nor U28235 (N_28235,N_27792,N_26507);
xnor U28236 (N_28236,N_27231,N_26573);
xor U28237 (N_28237,N_26654,N_26792);
nand U28238 (N_28238,N_27039,N_26055);
nor U28239 (N_28239,N_27156,N_27401);
or U28240 (N_28240,N_26956,N_26932);
xor U28241 (N_28241,N_27728,N_26179);
and U28242 (N_28242,N_27602,N_27160);
xnor U28243 (N_28243,N_26329,N_26129);
and U28244 (N_28244,N_27413,N_27774);
xnor U28245 (N_28245,N_27993,N_26777);
nand U28246 (N_28246,N_27968,N_26721);
nand U28247 (N_28247,N_27466,N_26555);
nor U28248 (N_28248,N_26013,N_26897);
xnor U28249 (N_28249,N_27031,N_27567);
and U28250 (N_28250,N_27464,N_27379);
xor U28251 (N_28251,N_27255,N_27981);
nand U28252 (N_28252,N_27675,N_26026);
nand U28253 (N_28253,N_26873,N_27179);
nor U28254 (N_28254,N_26307,N_27362);
or U28255 (N_28255,N_27939,N_27244);
and U28256 (N_28256,N_27817,N_27781);
or U28257 (N_28257,N_27022,N_26316);
or U28258 (N_28258,N_26012,N_26536);
nor U28259 (N_28259,N_27769,N_27897);
xor U28260 (N_28260,N_26994,N_27236);
and U28261 (N_28261,N_27305,N_26903);
and U28262 (N_28262,N_26548,N_27090);
xor U28263 (N_28263,N_27770,N_26867);
or U28264 (N_28264,N_26268,N_27839);
or U28265 (N_28265,N_27503,N_27721);
nand U28266 (N_28266,N_27831,N_27294);
xnor U28267 (N_28267,N_27846,N_27982);
nand U28268 (N_28268,N_27714,N_27732);
or U28269 (N_28269,N_26238,N_26499);
xnor U28270 (N_28270,N_27584,N_26188);
nor U28271 (N_28271,N_27009,N_26757);
xor U28272 (N_28272,N_27686,N_27833);
and U28273 (N_28273,N_27492,N_27335);
or U28274 (N_28274,N_26758,N_27274);
or U28275 (N_28275,N_26112,N_26209);
xnor U28276 (N_28276,N_26156,N_26857);
nor U28277 (N_28277,N_27921,N_27620);
and U28278 (N_28278,N_27980,N_26614);
nand U28279 (N_28279,N_26431,N_27262);
nor U28280 (N_28280,N_27801,N_27233);
xor U28281 (N_28281,N_26152,N_26323);
or U28282 (N_28282,N_27182,N_27200);
nand U28283 (N_28283,N_26230,N_26429);
nor U28284 (N_28284,N_26794,N_26175);
or U28285 (N_28285,N_27946,N_27611);
nand U28286 (N_28286,N_27127,N_27796);
xor U28287 (N_28287,N_26220,N_26023);
and U28288 (N_28288,N_27162,N_27777);
and U28289 (N_28289,N_27070,N_27601);
nor U28290 (N_28290,N_26599,N_26511);
xor U28291 (N_28291,N_26168,N_26618);
xnor U28292 (N_28292,N_26334,N_26204);
nor U28293 (N_28293,N_27380,N_27342);
and U28294 (N_28294,N_27296,N_26578);
xnor U28295 (N_28295,N_26242,N_27372);
xor U28296 (N_28296,N_27230,N_26335);
or U28297 (N_28297,N_27952,N_27969);
and U28298 (N_28298,N_27235,N_27552);
and U28299 (N_28299,N_27397,N_27868);
and U28300 (N_28300,N_26750,N_27793);
or U28301 (N_28301,N_27818,N_26605);
xor U28302 (N_28302,N_27257,N_26569);
nor U28303 (N_28303,N_27719,N_27359);
nand U28304 (N_28304,N_26642,N_26066);
or U28305 (N_28305,N_26633,N_26512);
or U28306 (N_28306,N_26214,N_26666);
nor U28307 (N_28307,N_27592,N_26342);
and U28308 (N_28308,N_27608,N_27038);
nand U28309 (N_28309,N_26344,N_27123);
xor U28310 (N_28310,N_26087,N_27302);
and U28311 (N_28311,N_26228,N_26973);
nand U28312 (N_28312,N_26053,N_26442);
or U28313 (N_28313,N_26491,N_26719);
and U28314 (N_28314,N_27779,N_27437);
nand U28315 (N_28315,N_26704,N_26022);
and U28316 (N_28316,N_27948,N_27460);
nand U28317 (N_28317,N_26990,N_27775);
nor U28318 (N_28318,N_27750,N_27600);
or U28319 (N_28319,N_26699,N_26800);
nand U28320 (N_28320,N_27963,N_27125);
nor U28321 (N_28321,N_27780,N_26515);
or U28322 (N_28322,N_27789,N_27167);
and U28323 (N_28323,N_26864,N_27622);
and U28324 (N_28324,N_26278,N_27242);
nand U28325 (N_28325,N_27263,N_26952);
xor U28326 (N_28326,N_26982,N_27099);
nor U28327 (N_28327,N_27436,N_26362);
xnor U28328 (N_28328,N_27636,N_27440);
and U28329 (N_28329,N_26117,N_26159);
nor U28330 (N_28330,N_27546,N_26935);
and U28331 (N_28331,N_27269,N_26140);
xor U28332 (N_28332,N_27352,N_27206);
and U28333 (N_28333,N_26604,N_26464);
or U28334 (N_28334,N_26538,N_26725);
and U28335 (N_28335,N_27149,N_26974);
or U28336 (N_28336,N_26251,N_26743);
and U28337 (N_28337,N_26969,N_27550);
xor U28338 (N_28338,N_26397,N_26224);
nor U28339 (N_28339,N_27880,N_27905);
nor U28340 (N_28340,N_27666,N_26032);
or U28341 (N_28341,N_27524,N_26904);
nor U28342 (N_28342,N_26207,N_26572);
and U28343 (N_28343,N_27876,N_27962);
nor U28344 (N_28344,N_27005,N_26079);
and U28345 (N_28345,N_26601,N_26664);
or U28346 (N_28346,N_26381,N_27544);
nor U28347 (N_28347,N_26926,N_27063);
nand U28348 (N_28348,N_26659,N_26727);
and U28349 (N_28349,N_27412,N_26271);
or U28350 (N_28350,N_27599,N_27995);
nand U28351 (N_28351,N_26878,N_27131);
nor U28352 (N_28352,N_27227,N_26449);
xor U28353 (N_28353,N_27644,N_27985);
or U28354 (N_28354,N_27391,N_27405);
and U28355 (N_28355,N_26532,N_26527);
and U28356 (N_28356,N_27504,N_27016);
and U28357 (N_28357,N_27259,N_26539);
or U28358 (N_28358,N_27189,N_26943);
and U28359 (N_28359,N_27509,N_27141);
and U28360 (N_28360,N_26589,N_26625);
nor U28361 (N_28361,N_27892,N_27882);
or U28362 (N_28362,N_26645,N_27520);
nor U28363 (N_28363,N_26901,N_27069);
nor U28364 (N_28364,N_26594,N_26270);
xnor U28365 (N_28365,N_27517,N_26562);
nor U28366 (N_28366,N_26047,N_27761);
nor U28367 (N_28367,N_26383,N_26516);
nor U28368 (N_28368,N_26246,N_27469);
nand U28369 (N_28369,N_26002,N_27183);
and U28370 (N_28370,N_27332,N_27402);
or U28371 (N_28371,N_26509,N_27711);
nor U28372 (N_28372,N_26297,N_26764);
nand U28373 (N_28373,N_26808,N_26723);
or U28374 (N_28374,N_26036,N_27766);
nor U28375 (N_28375,N_27726,N_27811);
and U28376 (N_28376,N_26593,N_27134);
nand U28377 (N_28377,N_26707,N_26164);
nand U28378 (N_28378,N_27118,N_26163);
nor U28379 (N_28379,N_27526,N_26035);
or U28380 (N_28380,N_27333,N_27762);
nand U28381 (N_28381,N_26501,N_26025);
nand U28382 (N_28382,N_26623,N_27529);
or U28383 (N_28383,N_26673,N_26187);
or U28384 (N_28384,N_26680,N_27927);
and U28385 (N_28385,N_26286,N_26160);
and U28386 (N_28386,N_26759,N_26206);
or U28387 (N_28387,N_26127,N_26640);
xnor U28388 (N_28388,N_26303,N_27688);
and U28389 (N_28389,N_26722,N_26389);
and U28390 (N_28390,N_27858,N_26662);
or U28391 (N_28391,N_27166,N_26807);
nor U28392 (N_28392,N_26942,N_26798);
nor U28393 (N_28393,N_26010,N_27906);
and U28394 (N_28394,N_27192,N_27283);
and U28395 (N_28395,N_27642,N_26519);
and U28396 (N_28396,N_27135,N_26559);
nor U28397 (N_28397,N_26401,N_27249);
nand U28398 (N_28398,N_26517,N_27776);
and U28399 (N_28399,N_26086,N_26842);
or U28400 (N_28400,N_27903,N_26311);
nand U28401 (N_28401,N_26302,N_26408);
xor U28402 (N_28402,N_27656,N_27247);
or U28403 (N_28403,N_27522,N_26749);
nor U28404 (N_28404,N_26510,N_27219);
nor U28405 (N_28405,N_27094,N_26195);
nor U28406 (N_28406,N_27330,N_26906);
xnor U28407 (N_28407,N_27241,N_26027);
or U28408 (N_28408,N_27316,N_26379);
or U28409 (N_28409,N_26736,N_27554);
or U28410 (N_28410,N_27692,N_27690);
xnor U28411 (N_28411,N_26905,N_26606);
nand U28412 (N_28412,N_26915,N_27428);
nand U28413 (N_28413,N_26745,N_27347);
and U28414 (N_28414,N_26031,N_26630);
xnor U28415 (N_28415,N_27351,N_27393);
nand U28416 (N_28416,N_27113,N_26044);
xnor U28417 (N_28417,N_26210,N_27024);
and U28418 (N_28418,N_26243,N_27220);
nand U28419 (N_28419,N_26496,N_27451);
or U28420 (N_28420,N_26998,N_26436);
nor U28421 (N_28421,N_26495,N_26529);
or U28422 (N_28422,N_27036,N_26245);
and U28423 (N_28423,N_26938,N_26848);
xnor U28424 (N_28424,N_27085,N_26502);
or U28425 (N_28425,N_26294,N_26828);
or U28426 (N_28426,N_27415,N_27797);
nand U28427 (N_28427,N_27052,N_26781);
nor U28428 (N_28428,N_27570,N_26678);
nand U28429 (N_28429,N_27590,N_27291);
nand U28430 (N_28430,N_26114,N_27878);
nor U28431 (N_28431,N_27275,N_26043);
nor U28432 (N_28432,N_27043,N_27497);
xor U28433 (N_28433,N_27496,N_27479);
nor U28434 (N_28434,N_27528,N_26717);
and U28435 (N_28435,N_27065,N_26690);
nand U28436 (N_28436,N_26697,N_27178);
nor U28437 (N_28437,N_26150,N_27706);
nor U28438 (N_28438,N_27959,N_26000);
nand U28439 (N_28439,N_26949,N_26062);
nand U28440 (N_28440,N_27276,N_27998);
xor U28441 (N_28441,N_27001,N_26534);
and U28442 (N_28442,N_26692,N_27763);
nor U28443 (N_28443,N_27083,N_26471);
and U28444 (N_28444,N_26233,N_26563);
or U28445 (N_28445,N_26095,N_26513);
nor U28446 (N_28446,N_27278,N_26739);
nor U28447 (N_28447,N_26264,N_27605);
and U28448 (N_28448,N_27681,N_26585);
nand U28449 (N_28449,N_27034,N_26176);
nand U28450 (N_28450,N_26263,N_27488);
nand U28451 (N_28451,N_27426,N_27683);
nor U28452 (N_28452,N_27300,N_26876);
nor U28453 (N_28453,N_26470,N_26111);
xor U28454 (N_28454,N_26968,N_26669);
nor U28455 (N_28455,N_26437,N_26983);
nor U28456 (N_28456,N_27325,N_26856);
and U28457 (N_28457,N_26076,N_27273);
or U28458 (N_28458,N_26412,N_27565);
nand U28459 (N_28459,N_27697,N_27104);
and U28460 (N_28460,N_27558,N_27964);
or U28461 (N_28461,N_27191,N_26369);
nand U28462 (N_28462,N_26822,N_27699);
or U28463 (N_28463,N_27947,N_27101);
and U28464 (N_28464,N_27086,N_26445);
or U28465 (N_28465,N_27084,N_27768);
xnor U28466 (N_28466,N_27631,N_27502);
nor U28467 (N_28467,N_27657,N_27986);
nand U28468 (N_28468,N_27282,N_26752);
xnor U28469 (N_28469,N_26291,N_26686);
or U28470 (N_28470,N_26762,N_27268);
or U28471 (N_28471,N_26468,N_26365);
and U28472 (N_28472,N_26577,N_27215);
xor U28473 (N_28473,N_26832,N_27795);
nand U28474 (N_28474,N_27992,N_26346);
nor U28475 (N_28475,N_27093,N_26877);
and U28476 (N_28476,N_26282,N_26695);
xnor U28477 (N_28477,N_26306,N_26970);
and U28478 (N_28478,N_27212,N_26193);
or U28479 (N_28479,N_26107,N_27536);
nor U28480 (N_28480,N_27046,N_27224);
or U28481 (N_28481,N_26934,N_26580);
nor U28482 (N_28482,N_26992,N_26797);
xnor U28483 (N_28483,N_27875,N_26360);
xor U28484 (N_28484,N_26249,N_27549);
nor U28485 (N_28485,N_27434,N_27957);
nor U28486 (N_28486,N_27072,N_26147);
nand U28487 (N_28487,N_27645,N_27679);
nor U28488 (N_28488,N_27385,N_27566);
and U28489 (N_28489,N_27910,N_27708);
and U28490 (N_28490,N_27050,N_26321);
xor U28491 (N_28491,N_26406,N_26774);
or U28492 (N_28492,N_26289,N_27954);
and U28493 (N_28493,N_27685,N_26928);
xnor U28494 (N_28494,N_27163,N_27739);
nand U28495 (N_28495,N_26371,N_27867);
and U28496 (N_28496,N_26871,N_26860);
xor U28497 (N_28497,N_27532,N_26399);
nand U28498 (N_28498,N_26778,N_26219);
nor U28499 (N_28499,N_26813,N_26829);
nor U28500 (N_28500,N_27344,N_27432);
and U28501 (N_28501,N_27115,N_26139);
nor U28502 (N_28502,N_27853,N_26082);
nor U28503 (N_28503,N_26333,N_26967);
or U28504 (N_28504,N_26455,N_27266);
xor U28505 (N_28505,N_27822,N_26192);
and U28506 (N_28506,N_27632,N_26180);
or U28507 (N_28507,N_27647,N_27791);
or U28508 (N_28508,N_27132,N_27338);
xnor U28509 (N_28509,N_27835,N_27159);
and U28510 (N_28510,N_27151,N_27452);
and U28511 (N_28511,N_27665,N_27629);
xor U28512 (N_28512,N_26481,N_26293);
nand U28513 (N_28513,N_26806,N_27336);
or U28514 (N_28514,N_27759,N_27195);
or U28515 (N_28515,N_26733,N_26166);
xor U28516 (N_28516,N_27482,N_26647);
and U28517 (N_28517,N_27427,N_27042);
nor U28518 (N_28518,N_26126,N_27410);
and U28519 (N_28519,N_26071,N_26728);
xor U28520 (N_28520,N_27836,N_27938);
nand U28521 (N_28521,N_26693,N_26831);
and U28522 (N_28522,N_26244,N_26151);
nor U28523 (N_28523,N_27971,N_27157);
xnor U28524 (N_28524,N_26950,N_27701);
or U28525 (N_28525,N_26296,N_27616);
nor U28526 (N_28526,N_27328,N_26446);
or U28527 (N_28527,N_26318,N_26088);
and U28528 (N_28528,N_26072,N_27095);
nand U28529 (N_28529,N_27730,N_27902);
nand U28530 (N_28530,N_27495,N_27002);
nor U28531 (N_28531,N_27794,N_27331);
nor U28532 (N_28532,N_27749,N_26194);
xor U28533 (N_28533,N_26568,N_26713);
nor U28534 (N_28534,N_26656,N_27597);
and U28535 (N_28535,N_27896,N_26830);
or U28536 (N_28536,N_26859,N_26737);
and U28537 (N_28537,N_26125,N_27060);
nand U28538 (N_28538,N_27540,N_27576);
and U28539 (N_28539,N_27456,N_27547);
nor U28540 (N_28540,N_27641,N_26007);
or U28541 (N_28541,N_26824,N_26966);
xnor U28542 (N_28542,N_26869,N_27041);
nor U28543 (N_28543,N_26612,N_26567);
or U28544 (N_28544,N_26646,N_26694);
or U28545 (N_28545,N_27551,N_26543);
xnor U28546 (N_28546,N_26462,N_27976);
nand U28547 (N_28547,N_26227,N_26677);
and U28548 (N_28548,N_26785,N_26154);
or U28549 (N_28549,N_27175,N_26503);
xor U28550 (N_28550,N_27154,N_27908);
nand U28551 (N_28551,N_27945,N_26801);
nor U28552 (N_28552,N_27731,N_26775);
nand U28553 (N_28553,N_26927,N_26339);
xor U28554 (N_28554,N_27915,N_26841);
nor U28555 (N_28555,N_27140,N_27662);
nand U28556 (N_28556,N_27088,N_26735);
nor U28557 (N_28557,N_27979,N_26835);
and U28558 (N_28558,N_26174,N_26059);
or U28559 (N_28559,N_26439,N_26823);
nor U28560 (N_28560,N_27377,N_26328);
xor U28561 (N_28561,N_26374,N_26288);
xnor U28562 (N_28562,N_27718,N_26330);
xor U28563 (N_28563,N_26658,N_26324);
and U28564 (N_28564,N_26660,N_27396);
xnor U28565 (N_28565,N_27449,N_26319);
xor U28566 (N_28566,N_27313,N_27258);
nor U28567 (N_28567,N_27312,N_27058);
nor U28568 (N_28568,N_27217,N_26128);
xnor U28569 (N_28569,N_27614,N_27329);
nand U28570 (N_28570,N_27148,N_26616);
or U28571 (N_28571,N_26919,N_27589);
nand U28572 (N_28572,N_27285,N_26077);
nand U28573 (N_28573,N_27109,N_27277);
nor U28574 (N_28574,N_26975,N_27181);
nand U28575 (N_28575,N_26701,N_27560);
and U28576 (N_28576,N_27586,N_27221);
or U28577 (N_28577,N_27006,N_26836);
nor U28578 (N_28578,N_27678,N_26273);
and U28579 (N_28579,N_27165,N_26119);
xnor U28580 (N_28580,N_27068,N_27256);
and U28581 (N_28581,N_26396,N_27729);
xor U28582 (N_28582,N_26874,N_26696);
nor U28583 (N_28583,N_26755,N_27057);
nand U28584 (N_28584,N_26084,N_27895);
nand U28585 (N_28585,N_26947,N_27026);
nor U28586 (N_28586,N_26351,N_26565);
or U28587 (N_28587,N_27106,N_26787);
xor U28588 (N_28588,N_27557,N_27021);
or U28589 (N_28589,N_26665,N_26327);
nand U28590 (N_28590,N_26581,N_26448);
nand U28591 (N_28591,N_27514,N_26889);
and U28592 (N_28592,N_27840,N_26409);
xor U28593 (N_28593,N_27128,N_26008);
or U28594 (N_28594,N_26820,N_27147);
nor U28595 (N_28595,N_27940,N_27609);
and U28596 (N_28596,N_26108,N_26716);
nor U28597 (N_28597,N_27438,N_27894);
and U28598 (N_28598,N_26423,N_26202);
nand U28599 (N_28599,N_27812,N_26854);
and U28600 (N_28600,N_26483,N_26292);
xor U28601 (N_28601,N_27778,N_27720);
and U28602 (N_28602,N_26216,N_27363);
xnor U28603 (N_28603,N_27516,N_26440);
and U28604 (N_28604,N_26619,N_26651);
nor U28605 (N_28605,N_26123,N_26001);
or U28606 (N_28606,N_27919,N_27297);
and U28607 (N_28607,N_27872,N_26937);
nand U28608 (N_28608,N_26225,N_26941);
or U28609 (N_28609,N_27152,N_26054);
xor U28610 (N_28610,N_26287,N_27542);
xnor U28611 (N_28611,N_27130,N_26478);
xnor U28612 (N_28612,N_27429,N_26505);
xnor U28613 (N_28613,N_26372,N_26799);
nand U28614 (N_28614,N_27960,N_27929);
nand U28615 (N_28615,N_27164,N_27399);
nor U28616 (N_28616,N_26038,N_27956);
nor U28617 (N_28617,N_26212,N_26019);
xor U28618 (N_28618,N_26795,N_26817);
nor U28619 (N_28619,N_27318,N_27000);
and U28620 (N_28620,N_26954,N_26962);
or U28621 (N_28621,N_26104,N_27298);
xnor U28622 (N_28622,N_26254,N_26587);
nand U28623 (N_28623,N_26060,N_27308);
xnor U28624 (N_28624,N_27349,N_27353);
or U28625 (N_28625,N_27756,N_27174);
or U28626 (N_28626,N_26554,N_26081);
nor U28627 (N_28627,N_27849,N_27826);
nor U28628 (N_28628,N_27441,N_26684);
nand U28629 (N_28629,N_26391,N_27639);
xnor U28630 (N_28630,N_27289,N_27303);
or U28631 (N_28631,N_27569,N_27484);
or U28632 (N_28632,N_26178,N_26237);
and U28633 (N_28633,N_26295,N_26522);
xor U28634 (N_28634,N_27937,N_26588);
nand U28635 (N_28635,N_27958,N_26438);
xor U28636 (N_28636,N_27049,N_27400);
or U28637 (N_28637,N_26541,N_27885);
xnor U28638 (N_28638,N_27032,N_26441);
nor U28639 (N_28639,N_26356,N_27579);
and U28640 (N_28640,N_26430,N_26706);
nand U28641 (N_28641,N_27170,N_27687);
and U28642 (N_28642,N_27595,N_26236);
xor U28643 (N_28643,N_27184,N_27168);
or U28644 (N_28644,N_26484,N_26017);
xor U28645 (N_28645,N_26711,N_27802);
xnor U28646 (N_28646,N_26414,N_26050);
nand U28647 (N_28647,N_27990,N_26791);
nor U28648 (N_28648,N_26494,N_27712);
or U28649 (N_28649,N_26912,N_27619);
or U28650 (N_28650,N_27727,N_27388);
nor U28651 (N_28651,N_26691,N_27012);
or U28652 (N_28652,N_26644,N_26506);
or U28653 (N_28653,N_27883,N_26655);
and U28654 (N_28654,N_27028,N_26861);
and U28655 (N_28655,N_27523,N_27287);
nor U28656 (N_28656,N_27996,N_27500);
or U28657 (N_28657,N_26566,N_27680);
xor U28658 (N_28658,N_27253,N_27755);
nand U28659 (N_28659,N_27481,N_27246);
and U28660 (N_28660,N_26475,N_26991);
xnor U28661 (N_28661,N_26052,N_26900);
xor U28662 (N_28662,N_26530,N_27489);
or U28663 (N_28663,N_26988,N_27888);
or U28664 (N_28664,N_27760,N_27931);
and U28665 (N_28665,N_27067,N_27458);
and U28666 (N_28666,N_27306,N_27723);
nor U28667 (N_28667,N_27076,N_26551);
xnor U28668 (N_28668,N_26229,N_27933);
and U28669 (N_28669,N_26161,N_27267);
and U28670 (N_28670,N_27243,N_27851);
and U28671 (N_28671,N_27669,N_27098);
xnor U28672 (N_28672,N_26776,N_26089);
nor U28673 (N_28673,N_27899,N_27364);
xor U28674 (N_28674,N_26557,N_27061);
nor U28675 (N_28675,N_26913,N_26450);
nand U28676 (N_28676,N_26064,N_27920);
nand U28677 (N_28677,N_26067,N_27389);
nand U28678 (N_28678,N_26742,N_27893);
xnor U28679 (N_28679,N_27752,N_26115);
or U28680 (N_28680,N_26134,N_27240);
or U28681 (N_28681,N_26895,N_27369);
nand U28682 (N_28682,N_26560,N_27814);
nor U28683 (N_28683,N_27909,N_27339);
nand U28684 (N_28684,N_27693,N_26849);
or U28685 (N_28685,N_26309,N_26939);
and U28686 (N_28686,N_26825,N_27468);
nand U28687 (N_28687,N_27942,N_27459);
and U28688 (N_28688,N_27261,N_27307);
and U28689 (N_28689,N_27010,N_27505);
and U28690 (N_28690,N_27350,N_26124);
nand U28691 (N_28691,N_26746,N_27218);
nand U28692 (N_28692,N_27898,N_27119);
xor U28693 (N_28693,N_26281,N_26730);
and U28694 (N_28694,N_26894,N_27111);
or U28695 (N_28695,N_27403,N_27568);
or U28696 (N_28696,N_26550,N_27651);
and U28697 (N_28697,N_27738,N_26868);
and U28698 (N_28698,N_27951,N_26657);
and U28699 (N_28699,N_26094,N_27941);
nor U28700 (N_28700,N_26881,N_26979);
nor U28701 (N_28701,N_26427,N_27035);
and U28702 (N_28702,N_27225,N_27295);
nor U28703 (N_28703,N_26514,N_26048);
nor U28704 (N_28704,N_27972,N_26652);
xor U28705 (N_28705,N_26355,N_27442);
nor U28706 (N_28706,N_26780,N_27977);
nor U28707 (N_28707,N_27625,N_27515);
or U28708 (N_28708,N_27304,N_27476);
or U28709 (N_28709,N_27617,N_27077);
or U28710 (N_28710,N_26393,N_26410);
or U28711 (N_28711,N_26816,N_26714);
and U28712 (N_28712,N_26989,N_26953);
nor U28713 (N_28713,N_26248,N_26886);
nor U28714 (N_28714,N_27454,N_27048);
or U28715 (N_28715,N_27827,N_27518);
nand U28716 (N_28716,N_27710,N_26322);
nand U28717 (N_28717,N_26533,N_26432);
or U28718 (N_28718,N_26793,N_27357);
and U28719 (N_28719,N_26405,N_26284);
or U28720 (N_28720,N_26526,N_27869);
nand U28721 (N_28721,N_26452,N_27820);
nand U28722 (N_28722,N_27407,N_26552);
xnor U28723 (N_28723,N_26863,N_27117);
or U28724 (N_28724,N_27753,N_26818);
and U28725 (N_28725,N_26914,N_26063);
and U28726 (N_28726,N_27742,N_27450);
xor U28727 (N_28727,N_26540,N_27354);
nand U28728 (N_28728,N_27765,N_26634);
and U28729 (N_28729,N_27975,N_27974);
nor U28730 (N_28730,N_27844,N_27045);
and U28731 (N_28731,N_26341,N_26261);
or U28732 (N_28732,N_26844,N_26402);
xnor U28733 (N_28733,N_27924,N_26763);
nand U28734 (N_28734,N_27572,N_26299);
or U28735 (N_28735,N_27382,N_26805);
xnor U28736 (N_28736,N_27834,N_27825);
and U28737 (N_28737,N_26683,N_26955);
nor U28738 (N_28738,N_26883,N_26090);
nor U28739 (N_28739,N_27754,N_26788);
and U28740 (N_28740,N_27474,N_26021);
xor U28741 (N_28741,N_26586,N_26469);
and U28742 (N_28742,N_26136,N_27859);
nand U28743 (N_28743,N_27857,N_27097);
and U28744 (N_28744,N_26821,N_26096);
nand U28745 (N_28745,N_26313,N_27023);
and U28746 (N_28746,N_27887,N_26269);
nor U28747 (N_28747,N_26121,N_27510);
xor U28748 (N_28748,N_26703,N_27431);
and U28749 (N_28749,N_27623,N_26603);
nor U28750 (N_28750,N_26443,N_26702);
nor U28751 (N_28751,N_27577,N_27668);
or U28752 (N_28752,N_26041,N_27610);
nand U28753 (N_28753,N_26834,N_27310);
xnor U28754 (N_28754,N_26424,N_27999);
and U28755 (N_28755,N_27564,N_26668);
nor U28756 (N_28756,N_26909,N_27477);
and U28757 (N_28757,N_27114,N_26865);
or U28758 (N_28758,N_26275,N_27139);
xor U28759 (N_28759,N_27961,N_27314);
nand U28760 (N_28760,N_26118,N_26637);
or U28761 (N_28761,N_26153,N_27345);
xor U28762 (N_28762,N_27507,N_26413);
xnor U28763 (N_28763,N_26364,N_26544);
nor U28764 (N_28764,N_26185,N_27116);
xor U28765 (N_28765,N_26337,N_26069);
nor U28766 (N_28766,N_27788,N_27588);
or U28767 (N_28767,N_27150,N_26545);
nor U28768 (N_28768,N_27691,N_26579);
nor U28769 (N_28769,N_27003,N_27365);
or U28770 (N_28770,N_26149,N_27530);
and U28771 (N_28771,N_26485,N_27375);
nor U28772 (N_28772,N_26314,N_27854);
or U28773 (N_28773,N_26239,N_26385);
xor U28774 (N_28774,N_26122,N_26046);
nor U28775 (N_28775,N_27966,N_26415);
nor U28776 (N_28776,N_27865,N_27670);
and U28777 (N_28777,N_26459,N_27563);
nor U28778 (N_28778,N_26885,N_26772);
and U28779 (N_28779,N_27292,N_26377);
and U28780 (N_28780,N_26018,N_27640);
nand U28781 (N_28781,N_27593,N_26508);
or U28782 (N_28782,N_27891,N_27051);
and U28783 (N_28783,N_27208,N_26158);
xnor U28784 (N_28784,N_26197,N_27096);
or U28785 (N_28785,N_26891,N_27199);
nor U28786 (N_28786,N_27852,N_27535);
or U28787 (N_28787,N_26765,N_27471);
and U28788 (N_28788,N_26698,N_26945);
or U28789 (N_28789,N_26617,N_26959);
or U28790 (N_28790,N_27444,N_26331);
xnor U28791 (N_28791,N_26591,N_26376);
nand U28792 (N_28792,N_27926,N_26996);
xnor U28793 (N_28793,N_27373,N_27238);
and U28794 (N_28794,N_27653,N_26786);
nand U28795 (N_28795,N_27816,N_27075);
nand U28796 (N_28796,N_27805,N_27944);
or U28797 (N_28797,N_27124,N_27508);
or U28798 (N_28798,N_27056,N_26924);
nor U28799 (N_28799,N_26571,N_26971);
nor U28800 (N_28800,N_26931,N_27013);
nand U28801 (N_28801,N_26961,N_26984);
or U28802 (N_28802,N_27017,N_27485);
nor U28803 (N_28803,N_26157,N_27819);
or U28804 (N_28804,N_26773,N_26672);
nand U28805 (N_28805,N_26070,N_27635);
or U28806 (N_28806,N_27994,N_27539);
or U28807 (N_28807,N_26305,N_26709);
xnor U28808 (N_28808,N_26486,N_27071);
nor U28809 (N_28809,N_26367,N_26866);
nand U28810 (N_28810,N_27555,N_26133);
xor U28811 (N_28811,N_27715,N_26769);
nor U28812 (N_28812,N_27767,N_27100);
or U28813 (N_28813,N_26592,N_26896);
and U28814 (N_28814,N_27418,N_26899);
nor U28815 (N_28815,N_26097,N_26375);
nor U28816 (N_28816,N_26855,N_27709);
and U28817 (N_28817,N_27177,N_27953);
and U28818 (N_28818,N_27232,N_26760);
nand U28819 (N_28819,N_27146,N_26113);
or U28820 (N_28820,N_26110,N_27153);
nand U28821 (N_28821,N_27281,N_26474);
or U28822 (N_28822,N_27054,N_26320);
and U28823 (N_28823,N_27404,N_26940);
or U28824 (N_28824,N_27603,N_27713);
and U28825 (N_28825,N_26170,N_26729);
and U28826 (N_28826,N_27138,N_27223);
nor U28827 (N_28827,N_26433,N_26387);
xnor U28828 (N_28828,N_27527,N_27848);
nor U28829 (N_28829,N_27596,N_27917);
or U28830 (N_28830,N_27724,N_27272);
xor U28831 (N_28831,N_27066,N_27734);
and U28832 (N_28832,N_26879,N_26102);
and U28833 (N_28833,N_27064,N_27348);
xor U28834 (N_28834,N_27337,N_27133);
nor U28835 (N_28835,N_27180,N_26492);
nand U28836 (N_28836,N_27473,N_26266);
or U28837 (N_28837,N_26685,N_26653);
or U28838 (N_28838,N_26006,N_26882);
nor U28839 (N_28839,N_26189,N_27040);
or U28840 (N_28840,N_26542,N_27582);
xor U28841 (N_28841,N_26211,N_26790);
and U28842 (N_28842,N_27467,N_26597);
and U28843 (N_28843,N_26535,N_26489);
nand U28844 (N_28844,N_27655,N_26105);
or U28845 (N_28845,N_26607,N_26731);
xor U28846 (N_28846,N_26682,N_26833);
or U28847 (N_28847,N_27621,N_27702);
nor U28848 (N_28848,N_27700,N_26144);
and U28849 (N_28849,N_27682,N_26756);
nor U28850 (N_28850,N_27573,N_27008);
nor U28851 (N_28851,N_26628,N_26726);
or U28852 (N_28852,N_27575,N_26132);
nor U28853 (N_28853,N_26747,N_27585);
or U28854 (N_28854,N_27904,N_26738);
or U28855 (N_28855,N_27416,N_26417);
or U28856 (N_28856,N_26853,N_26135);
and U28857 (N_28857,N_27293,N_27386);
and U28858 (N_28858,N_27194,N_27652);
or U28859 (N_28859,N_26100,N_27810);
or U28860 (N_28860,N_27315,N_26148);
nand U28861 (N_28861,N_27991,N_27301);
nand U28862 (N_28862,N_26155,N_26944);
or U28863 (N_28863,N_27239,N_27689);
xnor U28864 (N_28864,N_27787,N_26400);
nand U28865 (N_28865,N_27309,N_26336);
nand U28866 (N_28866,N_26679,N_26613);
and U28867 (N_28867,N_26887,N_26049);
nand U28868 (N_28868,N_26958,N_26173);
and U28869 (N_28869,N_26363,N_26921);
xnor U28870 (N_28870,N_27696,N_26280);
nand U28871 (N_28871,N_27745,N_26920);
and U28872 (N_28872,N_26283,N_26093);
or U28873 (N_28873,N_27807,N_27144);
xnor U28874 (N_28874,N_26171,N_26250);
or U28875 (N_28875,N_26255,N_27886);
or U28876 (N_28876,N_27922,N_26840);
nor U28877 (N_28877,N_26649,N_26190);
nor U28878 (N_28878,N_26034,N_27743);
xnor U28879 (N_28879,N_27059,N_27843);
and U28880 (N_28880,N_27445,N_27145);
nand U28881 (N_28881,N_26109,N_27684);
or U28882 (N_28882,N_27472,N_26826);
or U28883 (N_28883,N_26045,N_26130);
nand U28884 (N_28884,N_27207,N_27813);
and U28885 (N_28885,N_27271,N_26340);
or U28886 (N_28886,N_26183,N_27108);
or U28887 (N_28887,N_27660,N_26348);
xnor U28888 (N_28888,N_26222,N_27881);
nand U28889 (N_28889,N_27044,N_27855);
or U28890 (N_28890,N_27847,N_26310);
nand U28891 (N_28891,N_26910,N_27637);
or U28892 (N_28892,N_27672,N_27014);
or U28893 (N_28893,N_26368,N_27447);
nand U28894 (N_28894,N_27341,N_27519);
xnor U28895 (N_28895,N_27190,N_27533);
nor U28896 (N_28896,N_26629,N_26061);
xor U28897 (N_28897,N_26234,N_26985);
nor U28898 (N_28898,N_27368,N_27248);
nor U28899 (N_28899,N_26558,N_27664);
xnor U28900 (N_28900,N_26267,N_26005);
nand U28901 (N_28901,N_26639,N_26042);
nor U28902 (N_28902,N_27439,N_27158);
nand U28903 (N_28903,N_27062,N_26265);
nand U28904 (N_28904,N_26276,N_26162);
or U28905 (N_28905,N_27455,N_26326);
nor U28906 (N_28906,N_27025,N_27081);
nor U28907 (N_28907,N_26075,N_27978);
nand U28908 (N_28908,N_26290,N_26583);
nor U28909 (N_28909,N_27512,N_26936);
or U28910 (N_28910,N_27916,N_27483);
or U28911 (N_28911,N_26520,N_26024);
nor U28912 (N_28912,N_26167,N_26181);
nor U28913 (N_28913,N_27649,N_26493);
nor U28914 (N_28914,N_26258,N_27537);
nor U28915 (N_28915,N_26358,N_26200);
xor U28916 (N_28916,N_27829,N_27340);
and U28917 (N_28917,N_27435,N_26622);
nor U28918 (N_28918,N_27989,N_26411);
and U28919 (N_28919,N_27534,N_27733);
and U28920 (N_28920,N_26404,N_26259);
or U28921 (N_28921,N_27830,N_27018);
and U28922 (N_28922,N_26274,N_27531);
or U28923 (N_28923,N_26875,N_26620);
xor U28924 (N_28924,N_27799,N_27196);
and U28925 (N_28925,N_26621,N_27604);
or U28926 (N_28926,N_26177,N_26827);
and U28927 (N_28927,N_26030,N_26997);
xor U28928 (N_28928,N_26923,N_27676);
xnor U28929 (N_28929,N_26734,N_27722);
or U28930 (N_28930,N_27809,N_26847);
nor U28931 (N_28931,N_26003,N_27553);
or U28932 (N_28932,N_26631,N_27808);
and U28933 (N_28933,N_27394,N_26556);
xnor U28934 (N_28934,N_26232,N_26609);
xnor U28935 (N_28935,N_26993,N_27126);
nand U28936 (N_28936,N_27091,N_27965);
nor U28937 (N_28937,N_27591,N_27736);
or U28938 (N_28938,N_27461,N_27355);
nand U28939 (N_28939,N_26141,N_26811);
and U28940 (N_28940,N_26862,N_27806);
or U28941 (N_28941,N_26884,N_27425);
nand U28942 (N_28942,N_26453,N_26843);
and U28943 (N_28943,N_26106,N_27889);
nor U28944 (N_28944,N_27580,N_27019);
and U28945 (N_28945,N_26039,N_27646);
xor U28946 (N_28946,N_27654,N_27079);
nand U28947 (N_28947,N_27346,N_26608);
nand U28948 (N_28948,N_27803,N_27398);
and U28949 (N_28949,N_26068,N_26074);
xnor U28950 (N_28950,N_26624,N_27011);
and U28951 (N_28951,N_27169,N_26957);
or U28952 (N_28952,N_26497,N_27521);
nor U28953 (N_28953,N_27270,N_27030);
and U28954 (N_28954,N_26184,N_27936);
and U28955 (N_28955,N_26407,N_27873);
and U28956 (N_28956,N_26978,N_26208);
nand U28957 (N_28957,N_26011,N_27923);
and U28958 (N_28958,N_26169,N_26217);
xnor U28959 (N_28959,N_27918,N_27213);
xor U28960 (N_28960,N_27198,N_26918);
or U28961 (N_28961,N_26349,N_26819);
nor U28962 (N_28962,N_27943,N_27378);
xor U28963 (N_28963,N_27319,N_27112);
nor U28964 (N_28964,N_26761,N_27193);
nand U28965 (N_28965,N_27478,N_26576);
or U28966 (N_28966,N_27092,N_26615);
nor U28967 (N_28967,N_27423,N_26972);
or U28968 (N_28968,N_27667,N_27863);
nor U28969 (N_28969,N_27264,N_26783);
nand U28970 (N_28970,N_26172,N_27214);
or U28971 (N_28971,N_27871,N_26741);
nor U28972 (N_28972,N_26892,N_27737);
or U28973 (N_28973,N_27673,N_27171);
and U28974 (N_28974,N_27764,N_26803);
or U28975 (N_28975,N_26838,N_26028);
and U28976 (N_28976,N_27800,N_26201);
nor U28977 (N_28977,N_26770,N_26186);
and U28978 (N_28978,N_26131,N_27874);
nand U28979 (N_28979,N_26461,N_26948);
or U28980 (N_28980,N_27317,N_26458);
nor U28981 (N_28981,N_26262,N_27390);
and U28982 (N_28982,N_27698,N_26300);
or U28983 (N_28983,N_27073,N_26810);
nand U28984 (N_28984,N_26670,N_26465);
xnor U28985 (N_28985,N_26099,N_26457);
nor U28986 (N_28986,N_27618,N_26378);
or U28987 (N_28987,N_26546,N_26353);
nand U28988 (N_28988,N_27105,N_27556);
and U28989 (N_28989,N_27634,N_26460);
or U28990 (N_28990,N_26890,N_27587);
or U28991 (N_28991,N_26477,N_27663);
xnor U28992 (N_28992,N_26930,N_26815);
xnor U28993 (N_28993,N_26851,N_26165);
or U28994 (N_28994,N_27970,N_27538);
or U28995 (N_28995,N_27122,N_26388);
or U28996 (N_28996,N_27491,N_27771);
nor U28997 (N_28997,N_27988,N_26846);
xnor U28998 (N_28998,N_27624,N_27448);
nand U28999 (N_28999,N_27201,N_27121);
nor U29000 (N_29000,N_27399,N_27864);
nand U29001 (N_29001,N_27223,N_26886);
xor U29002 (N_29002,N_26160,N_26435);
xnor U29003 (N_29003,N_27901,N_26515);
or U29004 (N_29004,N_27270,N_27132);
nor U29005 (N_29005,N_27224,N_27797);
nor U29006 (N_29006,N_26229,N_27965);
or U29007 (N_29007,N_26500,N_26676);
or U29008 (N_29008,N_27051,N_27510);
xnor U29009 (N_29009,N_27927,N_26437);
xor U29010 (N_29010,N_27270,N_26136);
xnor U29011 (N_29011,N_27434,N_26409);
or U29012 (N_29012,N_27759,N_27712);
or U29013 (N_29013,N_26155,N_27934);
nor U29014 (N_29014,N_27002,N_27288);
nor U29015 (N_29015,N_26847,N_26352);
and U29016 (N_29016,N_26241,N_27165);
and U29017 (N_29017,N_27539,N_27342);
xor U29018 (N_29018,N_26781,N_26243);
xnor U29019 (N_29019,N_26793,N_27382);
and U29020 (N_29020,N_26276,N_27898);
nor U29021 (N_29021,N_27740,N_26945);
nor U29022 (N_29022,N_26586,N_27166);
and U29023 (N_29023,N_26185,N_26302);
nor U29024 (N_29024,N_26248,N_27440);
nand U29025 (N_29025,N_26298,N_27727);
nand U29026 (N_29026,N_27143,N_27799);
xnor U29027 (N_29027,N_26652,N_26324);
nor U29028 (N_29028,N_26837,N_27090);
nand U29029 (N_29029,N_26613,N_26419);
xor U29030 (N_29030,N_26265,N_26436);
or U29031 (N_29031,N_27443,N_27228);
xnor U29032 (N_29032,N_27379,N_26269);
and U29033 (N_29033,N_27240,N_26681);
nand U29034 (N_29034,N_26948,N_26510);
and U29035 (N_29035,N_26875,N_27525);
nand U29036 (N_29036,N_26152,N_27340);
and U29037 (N_29037,N_26078,N_26826);
and U29038 (N_29038,N_26447,N_27698);
nand U29039 (N_29039,N_26714,N_26056);
nor U29040 (N_29040,N_26151,N_27555);
xor U29041 (N_29041,N_27001,N_27153);
nand U29042 (N_29042,N_26310,N_26852);
nor U29043 (N_29043,N_26542,N_26674);
xor U29044 (N_29044,N_26613,N_26432);
nand U29045 (N_29045,N_26329,N_26526);
and U29046 (N_29046,N_27001,N_26383);
nor U29047 (N_29047,N_26073,N_26762);
or U29048 (N_29048,N_26667,N_27526);
and U29049 (N_29049,N_27697,N_26727);
nand U29050 (N_29050,N_26343,N_26011);
nand U29051 (N_29051,N_27835,N_26971);
nand U29052 (N_29052,N_26509,N_26409);
nand U29053 (N_29053,N_26397,N_26811);
nor U29054 (N_29054,N_27367,N_27566);
nand U29055 (N_29055,N_26228,N_26066);
xnor U29056 (N_29056,N_26508,N_26619);
nand U29057 (N_29057,N_26456,N_26703);
or U29058 (N_29058,N_27839,N_26377);
nand U29059 (N_29059,N_27097,N_27484);
nor U29060 (N_29060,N_27515,N_27066);
and U29061 (N_29061,N_26782,N_27406);
nor U29062 (N_29062,N_27425,N_26597);
xor U29063 (N_29063,N_27417,N_26722);
nor U29064 (N_29064,N_26567,N_27075);
xnor U29065 (N_29065,N_26612,N_26599);
nand U29066 (N_29066,N_26649,N_27117);
nand U29067 (N_29067,N_26600,N_26413);
nand U29068 (N_29068,N_26828,N_26092);
nor U29069 (N_29069,N_26879,N_27687);
nor U29070 (N_29070,N_26424,N_26696);
xor U29071 (N_29071,N_26185,N_27676);
and U29072 (N_29072,N_26208,N_26113);
and U29073 (N_29073,N_27217,N_26852);
xor U29074 (N_29074,N_27466,N_27698);
nor U29075 (N_29075,N_27968,N_27550);
and U29076 (N_29076,N_27935,N_27302);
or U29077 (N_29077,N_26097,N_27972);
xnor U29078 (N_29078,N_27867,N_26039);
nand U29079 (N_29079,N_26677,N_27485);
and U29080 (N_29080,N_27426,N_27653);
and U29081 (N_29081,N_27804,N_26710);
nor U29082 (N_29082,N_27405,N_27914);
nor U29083 (N_29083,N_26026,N_26892);
xnor U29084 (N_29084,N_27198,N_26919);
and U29085 (N_29085,N_27699,N_26012);
nor U29086 (N_29086,N_26351,N_27456);
or U29087 (N_29087,N_27330,N_27162);
and U29088 (N_29088,N_26029,N_26251);
or U29089 (N_29089,N_27196,N_26725);
and U29090 (N_29090,N_26824,N_27395);
and U29091 (N_29091,N_26283,N_26295);
nor U29092 (N_29092,N_26205,N_27970);
nor U29093 (N_29093,N_26272,N_27325);
nor U29094 (N_29094,N_26273,N_26037);
nand U29095 (N_29095,N_27201,N_26304);
and U29096 (N_29096,N_26057,N_27582);
nor U29097 (N_29097,N_26959,N_26210);
and U29098 (N_29098,N_27028,N_26144);
nor U29099 (N_29099,N_27564,N_26705);
nor U29100 (N_29100,N_26218,N_26097);
nand U29101 (N_29101,N_26635,N_26988);
nor U29102 (N_29102,N_27597,N_26816);
nand U29103 (N_29103,N_26210,N_27815);
nand U29104 (N_29104,N_27575,N_27023);
nor U29105 (N_29105,N_27437,N_27520);
or U29106 (N_29106,N_27884,N_27841);
nor U29107 (N_29107,N_26149,N_27529);
nor U29108 (N_29108,N_27762,N_27811);
nor U29109 (N_29109,N_26831,N_26512);
nor U29110 (N_29110,N_27433,N_27280);
nand U29111 (N_29111,N_27403,N_26045);
nand U29112 (N_29112,N_27669,N_26168);
nand U29113 (N_29113,N_27914,N_26472);
xor U29114 (N_29114,N_27568,N_26592);
nor U29115 (N_29115,N_27680,N_26544);
or U29116 (N_29116,N_27917,N_26673);
nand U29117 (N_29117,N_27329,N_27090);
and U29118 (N_29118,N_26487,N_27396);
xor U29119 (N_29119,N_26062,N_27929);
xor U29120 (N_29120,N_27503,N_27120);
and U29121 (N_29121,N_27566,N_26354);
nand U29122 (N_29122,N_26577,N_26267);
nand U29123 (N_29123,N_26006,N_27906);
nor U29124 (N_29124,N_27170,N_27126);
nor U29125 (N_29125,N_27356,N_26552);
nor U29126 (N_29126,N_27339,N_27070);
and U29127 (N_29127,N_26812,N_26338);
xor U29128 (N_29128,N_26235,N_27044);
or U29129 (N_29129,N_26673,N_26398);
or U29130 (N_29130,N_26427,N_26337);
nand U29131 (N_29131,N_27086,N_27381);
xor U29132 (N_29132,N_27396,N_26065);
nor U29133 (N_29133,N_27143,N_27756);
xnor U29134 (N_29134,N_27140,N_26395);
and U29135 (N_29135,N_27496,N_27422);
nand U29136 (N_29136,N_26541,N_27200);
xor U29137 (N_29137,N_27894,N_26008);
nand U29138 (N_29138,N_27808,N_26892);
nand U29139 (N_29139,N_27265,N_26306);
xor U29140 (N_29140,N_27430,N_27178);
nor U29141 (N_29141,N_27036,N_26393);
nor U29142 (N_29142,N_27584,N_26624);
xor U29143 (N_29143,N_27324,N_26047);
nand U29144 (N_29144,N_27790,N_26144);
and U29145 (N_29145,N_26908,N_26256);
nor U29146 (N_29146,N_27572,N_26476);
nor U29147 (N_29147,N_26484,N_27142);
nor U29148 (N_29148,N_26210,N_27406);
nand U29149 (N_29149,N_27122,N_27820);
nor U29150 (N_29150,N_26520,N_26762);
nand U29151 (N_29151,N_26642,N_26549);
nor U29152 (N_29152,N_26933,N_26675);
nand U29153 (N_29153,N_27922,N_26870);
or U29154 (N_29154,N_27668,N_26472);
nor U29155 (N_29155,N_26521,N_27875);
or U29156 (N_29156,N_26048,N_27494);
xor U29157 (N_29157,N_26404,N_26713);
nand U29158 (N_29158,N_27405,N_26760);
or U29159 (N_29159,N_27707,N_27504);
nor U29160 (N_29160,N_26185,N_26040);
xor U29161 (N_29161,N_27956,N_26236);
nand U29162 (N_29162,N_26812,N_26862);
nand U29163 (N_29163,N_26576,N_27103);
nor U29164 (N_29164,N_26223,N_26010);
or U29165 (N_29165,N_27313,N_26922);
xnor U29166 (N_29166,N_27682,N_26385);
or U29167 (N_29167,N_27118,N_27103);
nor U29168 (N_29168,N_26305,N_26801);
nor U29169 (N_29169,N_26139,N_27544);
or U29170 (N_29170,N_27169,N_27326);
and U29171 (N_29171,N_26357,N_26355);
xnor U29172 (N_29172,N_27130,N_27272);
or U29173 (N_29173,N_27014,N_27092);
nor U29174 (N_29174,N_26800,N_26172);
xor U29175 (N_29175,N_27282,N_26111);
xnor U29176 (N_29176,N_27744,N_27216);
and U29177 (N_29177,N_26053,N_27121);
and U29178 (N_29178,N_26363,N_27907);
and U29179 (N_29179,N_26310,N_27880);
and U29180 (N_29180,N_27733,N_26194);
nor U29181 (N_29181,N_27147,N_27124);
nand U29182 (N_29182,N_26216,N_26084);
and U29183 (N_29183,N_27365,N_27463);
and U29184 (N_29184,N_26646,N_27242);
xnor U29185 (N_29185,N_27267,N_27336);
or U29186 (N_29186,N_26266,N_27104);
xnor U29187 (N_29187,N_27384,N_27163);
nand U29188 (N_29188,N_26342,N_26811);
or U29189 (N_29189,N_27177,N_26102);
nor U29190 (N_29190,N_26536,N_27124);
nand U29191 (N_29191,N_27339,N_27254);
nand U29192 (N_29192,N_27779,N_26305);
and U29193 (N_29193,N_26469,N_26559);
xor U29194 (N_29194,N_27713,N_26649);
nor U29195 (N_29195,N_26939,N_27571);
or U29196 (N_29196,N_26170,N_27366);
xnor U29197 (N_29197,N_26495,N_26863);
xor U29198 (N_29198,N_26045,N_27162);
or U29199 (N_29199,N_27161,N_26846);
nor U29200 (N_29200,N_27944,N_26584);
or U29201 (N_29201,N_26543,N_27658);
and U29202 (N_29202,N_27987,N_26306);
xnor U29203 (N_29203,N_26223,N_26244);
xor U29204 (N_29204,N_26673,N_26876);
nand U29205 (N_29205,N_26554,N_26232);
and U29206 (N_29206,N_27347,N_27339);
nand U29207 (N_29207,N_27781,N_27465);
nand U29208 (N_29208,N_26191,N_26638);
and U29209 (N_29209,N_27259,N_26578);
nor U29210 (N_29210,N_26011,N_27056);
nand U29211 (N_29211,N_27152,N_26954);
xor U29212 (N_29212,N_27959,N_26144);
xor U29213 (N_29213,N_26500,N_26873);
or U29214 (N_29214,N_26142,N_27562);
nand U29215 (N_29215,N_26314,N_26718);
xor U29216 (N_29216,N_26880,N_27933);
xor U29217 (N_29217,N_27859,N_27585);
nand U29218 (N_29218,N_27142,N_26958);
xor U29219 (N_29219,N_27195,N_27575);
nand U29220 (N_29220,N_27142,N_27494);
nand U29221 (N_29221,N_27845,N_26861);
nor U29222 (N_29222,N_26633,N_27148);
nand U29223 (N_29223,N_27176,N_27449);
or U29224 (N_29224,N_27327,N_26093);
or U29225 (N_29225,N_27360,N_27747);
or U29226 (N_29226,N_27678,N_27756);
and U29227 (N_29227,N_26466,N_26431);
or U29228 (N_29228,N_27597,N_27013);
and U29229 (N_29229,N_26729,N_26239);
nand U29230 (N_29230,N_26977,N_27224);
nand U29231 (N_29231,N_26970,N_27335);
and U29232 (N_29232,N_27505,N_27704);
xnor U29233 (N_29233,N_27780,N_26684);
and U29234 (N_29234,N_26086,N_27123);
nor U29235 (N_29235,N_26517,N_27436);
or U29236 (N_29236,N_26541,N_26327);
xnor U29237 (N_29237,N_26270,N_26942);
and U29238 (N_29238,N_27404,N_26963);
nor U29239 (N_29239,N_27091,N_26177);
nand U29240 (N_29240,N_26923,N_26329);
nand U29241 (N_29241,N_26300,N_27010);
and U29242 (N_29242,N_27267,N_27847);
nand U29243 (N_29243,N_26649,N_26179);
or U29244 (N_29244,N_27180,N_26447);
and U29245 (N_29245,N_27911,N_27665);
nand U29246 (N_29246,N_27184,N_26614);
xor U29247 (N_29247,N_27390,N_27978);
xor U29248 (N_29248,N_27087,N_27768);
nand U29249 (N_29249,N_26220,N_27403);
xor U29250 (N_29250,N_27431,N_27567);
and U29251 (N_29251,N_27820,N_26269);
xor U29252 (N_29252,N_26463,N_26823);
xor U29253 (N_29253,N_27943,N_27258);
nand U29254 (N_29254,N_26702,N_27894);
or U29255 (N_29255,N_26922,N_26093);
nor U29256 (N_29256,N_26701,N_26742);
xor U29257 (N_29257,N_26387,N_26050);
nor U29258 (N_29258,N_27422,N_26391);
xnor U29259 (N_29259,N_27731,N_26889);
and U29260 (N_29260,N_27014,N_26310);
and U29261 (N_29261,N_27697,N_26060);
nor U29262 (N_29262,N_27871,N_27424);
or U29263 (N_29263,N_27415,N_26223);
xor U29264 (N_29264,N_27666,N_27235);
xnor U29265 (N_29265,N_27451,N_26643);
and U29266 (N_29266,N_26687,N_27428);
nor U29267 (N_29267,N_26087,N_26367);
nor U29268 (N_29268,N_26944,N_27280);
nand U29269 (N_29269,N_26579,N_27756);
or U29270 (N_29270,N_27207,N_26334);
or U29271 (N_29271,N_27011,N_27333);
nand U29272 (N_29272,N_26718,N_27479);
nand U29273 (N_29273,N_26131,N_27760);
xor U29274 (N_29274,N_27134,N_27660);
and U29275 (N_29275,N_27247,N_26421);
and U29276 (N_29276,N_26042,N_27933);
nand U29277 (N_29277,N_26218,N_26540);
nand U29278 (N_29278,N_27145,N_27825);
and U29279 (N_29279,N_27060,N_27935);
nand U29280 (N_29280,N_27990,N_26488);
nand U29281 (N_29281,N_27382,N_27877);
or U29282 (N_29282,N_26798,N_26241);
and U29283 (N_29283,N_27526,N_27660);
nor U29284 (N_29284,N_26553,N_26281);
or U29285 (N_29285,N_26220,N_27834);
or U29286 (N_29286,N_26489,N_27920);
or U29287 (N_29287,N_26242,N_26601);
and U29288 (N_29288,N_27687,N_27986);
nand U29289 (N_29289,N_27635,N_27920);
or U29290 (N_29290,N_27307,N_26173);
and U29291 (N_29291,N_26408,N_27454);
nor U29292 (N_29292,N_26625,N_26893);
xor U29293 (N_29293,N_27814,N_26024);
and U29294 (N_29294,N_26089,N_27093);
and U29295 (N_29295,N_26414,N_27015);
nand U29296 (N_29296,N_27533,N_26804);
and U29297 (N_29297,N_26246,N_27754);
and U29298 (N_29298,N_26226,N_26735);
nand U29299 (N_29299,N_27847,N_27578);
nand U29300 (N_29300,N_26368,N_27660);
nor U29301 (N_29301,N_27661,N_27876);
xnor U29302 (N_29302,N_27084,N_27087);
nor U29303 (N_29303,N_26378,N_27465);
nor U29304 (N_29304,N_27195,N_26505);
nor U29305 (N_29305,N_27401,N_26268);
and U29306 (N_29306,N_27257,N_27357);
nor U29307 (N_29307,N_26218,N_26528);
or U29308 (N_29308,N_26022,N_27004);
or U29309 (N_29309,N_26499,N_26576);
nor U29310 (N_29310,N_27060,N_27910);
nand U29311 (N_29311,N_26157,N_26033);
nor U29312 (N_29312,N_26057,N_26588);
nor U29313 (N_29313,N_26083,N_26411);
and U29314 (N_29314,N_26644,N_27414);
nand U29315 (N_29315,N_27727,N_26606);
nor U29316 (N_29316,N_26957,N_26554);
or U29317 (N_29317,N_27549,N_26465);
xnor U29318 (N_29318,N_27407,N_26610);
or U29319 (N_29319,N_26531,N_26813);
or U29320 (N_29320,N_27460,N_27475);
nand U29321 (N_29321,N_27856,N_26660);
nand U29322 (N_29322,N_27559,N_27290);
xnor U29323 (N_29323,N_26392,N_27395);
and U29324 (N_29324,N_27134,N_26800);
nor U29325 (N_29325,N_26663,N_26189);
nor U29326 (N_29326,N_27253,N_26775);
xnor U29327 (N_29327,N_26021,N_27745);
nand U29328 (N_29328,N_27363,N_26264);
and U29329 (N_29329,N_26244,N_27478);
and U29330 (N_29330,N_27790,N_26455);
nand U29331 (N_29331,N_27203,N_27955);
or U29332 (N_29332,N_27275,N_26581);
and U29333 (N_29333,N_26482,N_27333);
xnor U29334 (N_29334,N_27179,N_27426);
nor U29335 (N_29335,N_27897,N_27945);
nor U29336 (N_29336,N_26241,N_26054);
nand U29337 (N_29337,N_26159,N_26418);
or U29338 (N_29338,N_27786,N_26541);
nor U29339 (N_29339,N_27012,N_26679);
and U29340 (N_29340,N_26215,N_27029);
or U29341 (N_29341,N_27176,N_26660);
xor U29342 (N_29342,N_26205,N_27754);
or U29343 (N_29343,N_27095,N_26543);
or U29344 (N_29344,N_27700,N_26256);
and U29345 (N_29345,N_27970,N_27124);
nand U29346 (N_29346,N_27865,N_26391);
or U29347 (N_29347,N_27923,N_27983);
nand U29348 (N_29348,N_26884,N_27240);
xor U29349 (N_29349,N_26326,N_27173);
or U29350 (N_29350,N_27350,N_27124);
nand U29351 (N_29351,N_26231,N_26594);
nor U29352 (N_29352,N_27027,N_26155);
or U29353 (N_29353,N_26589,N_27285);
and U29354 (N_29354,N_27149,N_27650);
xnor U29355 (N_29355,N_27500,N_26738);
nor U29356 (N_29356,N_27083,N_26248);
or U29357 (N_29357,N_27163,N_26053);
nand U29358 (N_29358,N_26346,N_27218);
xnor U29359 (N_29359,N_26230,N_26091);
nor U29360 (N_29360,N_27645,N_26638);
xor U29361 (N_29361,N_26006,N_26196);
xor U29362 (N_29362,N_27013,N_27872);
or U29363 (N_29363,N_27596,N_27631);
or U29364 (N_29364,N_27436,N_26882);
xor U29365 (N_29365,N_26884,N_27093);
and U29366 (N_29366,N_26610,N_26137);
nor U29367 (N_29367,N_26630,N_26014);
or U29368 (N_29368,N_26707,N_27184);
xnor U29369 (N_29369,N_27066,N_26043);
nor U29370 (N_29370,N_27719,N_27806);
xnor U29371 (N_29371,N_27698,N_27451);
or U29372 (N_29372,N_26079,N_26359);
and U29373 (N_29373,N_26741,N_27420);
or U29374 (N_29374,N_26375,N_26972);
and U29375 (N_29375,N_27663,N_26686);
and U29376 (N_29376,N_26350,N_26890);
nor U29377 (N_29377,N_26334,N_26656);
xnor U29378 (N_29378,N_26420,N_26590);
nor U29379 (N_29379,N_27643,N_26869);
or U29380 (N_29380,N_26783,N_27157);
nor U29381 (N_29381,N_27121,N_26204);
and U29382 (N_29382,N_27682,N_26956);
nor U29383 (N_29383,N_26266,N_27489);
xnor U29384 (N_29384,N_27320,N_27911);
and U29385 (N_29385,N_26754,N_27801);
nor U29386 (N_29386,N_27486,N_26802);
nor U29387 (N_29387,N_27709,N_27838);
and U29388 (N_29388,N_26385,N_26903);
nand U29389 (N_29389,N_26702,N_27269);
nand U29390 (N_29390,N_27000,N_26886);
nand U29391 (N_29391,N_26670,N_26259);
or U29392 (N_29392,N_27127,N_26664);
xor U29393 (N_29393,N_27729,N_27992);
nor U29394 (N_29394,N_26835,N_26889);
and U29395 (N_29395,N_27544,N_27656);
or U29396 (N_29396,N_27559,N_27135);
xnor U29397 (N_29397,N_27705,N_26659);
and U29398 (N_29398,N_27749,N_26948);
xor U29399 (N_29399,N_27093,N_26658);
or U29400 (N_29400,N_26924,N_26216);
and U29401 (N_29401,N_27240,N_26741);
and U29402 (N_29402,N_26894,N_26425);
xor U29403 (N_29403,N_27244,N_26428);
nand U29404 (N_29404,N_27825,N_26709);
xor U29405 (N_29405,N_27012,N_26423);
xnor U29406 (N_29406,N_27436,N_26806);
xnor U29407 (N_29407,N_27168,N_27145);
nand U29408 (N_29408,N_27185,N_27340);
xor U29409 (N_29409,N_26881,N_26159);
xor U29410 (N_29410,N_26004,N_27292);
nor U29411 (N_29411,N_27348,N_27507);
nor U29412 (N_29412,N_27559,N_26862);
nor U29413 (N_29413,N_27006,N_26569);
nand U29414 (N_29414,N_27188,N_26948);
nand U29415 (N_29415,N_27718,N_26633);
xnor U29416 (N_29416,N_26895,N_26384);
xor U29417 (N_29417,N_26232,N_26738);
nor U29418 (N_29418,N_26812,N_27109);
and U29419 (N_29419,N_27788,N_27767);
or U29420 (N_29420,N_26553,N_26015);
nor U29421 (N_29421,N_26023,N_26458);
nand U29422 (N_29422,N_26180,N_26905);
nand U29423 (N_29423,N_27432,N_26496);
nand U29424 (N_29424,N_26578,N_26646);
nor U29425 (N_29425,N_27296,N_27974);
nand U29426 (N_29426,N_26240,N_26515);
nor U29427 (N_29427,N_26731,N_26324);
nor U29428 (N_29428,N_26327,N_27871);
nand U29429 (N_29429,N_27204,N_26486);
xor U29430 (N_29430,N_27878,N_27755);
and U29431 (N_29431,N_27437,N_26389);
and U29432 (N_29432,N_26538,N_26383);
nor U29433 (N_29433,N_26841,N_27837);
xnor U29434 (N_29434,N_27219,N_26932);
xor U29435 (N_29435,N_26685,N_27246);
xor U29436 (N_29436,N_26304,N_26766);
or U29437 (N_29437,N_26388,N_26905);
and U29438 (N_29438,N_27313,N_26981);
nor U29439 (N_29439,N_27855,N_26742);
xnor U29440 (N_29440,N_27721,N_27049);
xor U29441 (N_29441,N_27306,N_26965);
or U29442 (N_29442,N_26902,N_27566);
nand U29443 (N_29443,N_26263,N_26333);
and U29444 (N_29444,N_26874,N_27643);
and U29445 (N_29445,N_26048,N_27127);
or U29446 (N_29446,N_26121,N_26370);
xnor U29447 (N_29447,N_26796,N_26897);
or U29448 (N_29448,N_27177,N_26412);
and U29449 (N_29449,N_27262,N_27977);
or U29450 (N_29450,N_26921,N_27068);
nor U29451 (N_29451,N_27922,N_27016);
xnor U29452 (N_29452,N_26934,N_27546);
nor U29453 (N_29453,N_27178,N_26245);
and U29454 (N_29454,N_27489,N_26820);
and U29455 (N_29455,N_27183,N_26999);
and U29456 (N_29456,N_27166,N_26910);
xnor U29457 (N_29457,N_26436,N_27478);
nor U29458 (N_29458,N_26164,N_27339);
nand U29459 (N_29459,N_27159,N_27083);
xnor U29460 (N_29460,N_26502,N_26467);
nand U29461 (N_29461,N_26790,N_27379);
nor U29462 (N_29462,N_27025,N_26107);
or U29463 (N_29463,N_26310,N_26557);
nor U29464 (N_29464,N_27191,N_27359);
nand U29465 (N_29465,N_26971,N_27643);
nor U29466 (N_29466,N_27566,N_26881);
nand U29467 (N_29467,N_27948,N_26385);
xnor U29468 (N_29468,N_26853,N_27581);
nor U29469 (N_29469,N_27127,N_26277);
nand U29470 (N_29470,N_26462,N_27579);
nand U29471 (N_29471,N_26370,N_26969);
or U29472 (N_29472,N_27464,N_26798);
xor U29473 (N_29473,N_27271,N_27053);
and U29474 (N_29474,N_26464,N_26502);
and U29475 (N_29475,N_26874,N_27345);
nor U29476 (N_29476,N_27718,N_26127);
or U29477 (N_29477,N_27484,N_26509);
or U29478 (N_29478,N_26532,N_27097);
or U29479 (N_29479,N_26714,N_27866);
and U29480 (N_29480,N_26125,N_27973);
nand U29481 (N_29481,N_26450,N_27356);
and U29482 (N_29482,N_26121,N_27253);
nor U29483 (N_29483,N_26587,N_27753);
nand U29484 (N_29484,N_26956,N_26548);
and U29485 (N_29485,N_27305,N_27849);
and U29486 (N_29486,N_27922,N_26638);
xnor U29487 (N_29487,N_27263,N_26375);
nand U29488 (N_29488,N_26523,N_27572);
nand U29489 (N_29489,N_27086,N_26675);
nor U29490 (N_29490,N_27765,N_26258);
nor U29491 (N_29491,N_26682,N_27975);
nor U29492 (N_29492,N_27722,N_27347);
xor U29493 (N_29493,N_27648,N_26720);
and U29494 (N_29494,N_26092,N_26969);
nand U29495 (N_29495,N_26539,N_27271);
nand U29496 (N_29496,N_26903,N_26102);
nand U29497 (N_29497,N_26508,N_27702);
and U29498 (N_29498,N_26543,N_27627);
nor U29499 (N_29499,N_27068,N_26842);
xor U29500 (N_29500,N_27525,N_27902);
nor U29501 (N_29501,N_27674,N_26781);
nor U29502 (N_29502,N_26395,N_26193);
or U29503 (N_29503,N_27459,N_26475);
nand U29504 (N_29504,N_26659,N_27429);
and U29505 (N_29505,N_27323,N_27568);
nor U29506 (N_29506,N_27035,N_27277);
nor U29507 (N_29507,N_26045,N_26469);
nand U29508 (N_29508,N_26099,N_27962);
or U29509 (N_29509,N_27819,N_26458);
xnor U29510 (N_29510,N_26798,N_26011);
and U29511 (N_29511,N_26639,N_27721);
nor U29512 (N_29512,N_27090,N_26042);
and U29513 (N_29513,N_26233,N_27807);
nor U29514 (N_29514,N_26505,N_26671);
xnor U29515 (N_29515,N_27533,N_27813);
or U29516 (N_29516,N_26211,N_27798);
nand U29517 (N_29517,N_26226,N_27490);
or U29518 (N_29518,N_26207,N_26919);
xor U29519 (N_29519,N_27990,N_26449);
and U29520 (N_29520,N_26833,N_27111);
and U29521 (N_29521,N_27023,N_27113);
or U29522 (N_29522,N_26543,N_26442);
nand U29523 (N_29523,N_26027,N_26923);
and U29524 (N_29524,N_27200,N_26872);
xor U29525 (N_29525,N_26186,N_26305);
xor U29526 (N_29526,N_26517,N_27990);
and U29527 (N_29527,N_27040,N_26520);
xnor U29528 (N_29528,N_26387,N_26920);
or U29529 (N_29529,N_27637,N_26977);
nand U29530 (N_29530,N_26452,N_26248);
nand U29531 (N_29531,N_27910,N_26010);
or U29532 (N_29532,N_27625,N_27829);
or U29533 (N_29533,N_27732,N_27266);
or U29534 (N_29534,N_27076,N_26277);
or U29535 (N_29535,N_27076,N_27325);
xor U29536 (N_29536,N_26025,N_27332);
xor U29537 (N_29537,N_27175,N_26054);
nor U29538 (N_29538,N_26070,N_27479);
and U29539 (N_29539,N_26984,N_26999);
nand U29540 (N_29540,N_27773,N_27374);
xnor U29541 (N_29541,N_26999,N_27847);
and U29542 (N_29542,N_27706,N_27470);
xnor U29543 (N_29543,N_26587,N_26514);
xor U29544 (N_29544,N_26202,N_26431);
or U29545 (N_29545,N_26738,N_26900);
nand U29546 (N_29546,N_26903,N_26875);
nand U29547 (N_29547,N_27776,N_27930);
nand U29548 (N_29548,N_26327,N_27135);
xor U29549 (N_29549,N_26916,N_26487);
nand U29550 (N_29550,N_27698,N_27650);
nor U29551 (N_29551,N_27214,N_26383);
and U29552 (N_29552,N_27908,N_27654);
xnor U29553 (N_29553,N_26322,N_26021);
or U29554 (N_29554,N_26705,N_27733);
nand U29555 (N_29555,N_26324,N_27208);
xnor U29556 (N_29556,N_27665,N_27324);
xor U29557 (N_29557,N_26729,N_27121);
and U29558 (N_29558,N_26837,N_27405);
and U29559 (N_29559,N_27938,N_26808);
nand U29560 (N_29560,N_27366,N_27007);
nor U29561 (N_29561,N_27575,N_26023);
xor U29562 (N_29562,N_26862,N_27283);
or U29563 (N_29563,N_26390,N_27560);
xnor U29564 (N_29564,N_26278,N_26563);
nor U29565 (N_29565,N_27409,N_27673);
nand U29566 (N_29566,N_26829,N_27391);
or U29567 (N_29567,N_27214,N_27710);
xor U29568 (N_29568,N_27456,N_26659);
nand U29569 (N_29569,N_26218,N_27312);
nor U29570 (N_29570,N_27252,N_26205);
and U29571 (N_29571,N_26624,N_26967);
nand U29572 (N_29572,N_26720,N_27537);
or U29573 (N_29573,N_26282,N_26031);
and U29574 (N_29574,N_26961,N_27931);
xor U29575 (N_29575,N_27005,N_27174);
xnor U29576 (N_29576,N_26113,N_26668);
nand U29577 (N_29577,N_26189,N_27187);
and U29578 (N_29578,N_27841,N_27628);
xnor U29579 (N_29579,N_26068,N_27282);
or U29580 (N_29580,N_26525,N_27869);
and U29581 (N_29581,N_26430,N_27368);
nor U29582 (N_29582,N_26807,N_26488);
or U29583 (N_29583,N_27948,N_27882);
xor U29584 (N_29584,N_27208,N_26916);
and U29585 (N_29585,N_27711,N_26014);
xor U29586 (N_29586,N_26980,N_27962);
and U29587 (N_29587,N_27478,N_27298);
or U29588 (N_29588,N_26787,N_26218);
nand U29589 (N_29589,N_27973,N_26120);
xor U29590 (N_29590,N_27112,N_27404);
and U29591 (N_29591,N_26761,N_27710);
and U29592 (N_29592,N_27642,N_26556);
nor U29593 (N_29593,N_27563,N_26076);
nor U29594 (N_29594,N_27066,N_27183);
and U29595 (N_29595,N_26899,N_27320);
nor U29596 (N_29596,N_26125,N_26902);
or U29597 (N_29597,N_27958,N_26815);
nand U29598 (N_29598,N_27126,N_27314);
xor U29599 (N_29599,N_27111,N_27026);
or U29600 (N_29600,N_27957,N_27230);
or U29601 (N_29601,N_26204,N_27850);
nor U29602 (N_29602,N_26621,N_26142);
and U29603 (N_29603,N_26329,N_27521);
xnor U29604 (N_29604,N_26900,N_27821);
nand U29605 (N_29605,N_26108,N_27357);
xnor U29606 (N_29606,N_26914,N_26669);
nor U29607 (N_29607,N_27713,N_26696);
or U29608 (N_29608,N_27131,N_27988);
nand U29609 (N_29609,N_27570,N_26223);
nor U29610 (N_29610,N_26267,N_27292);
xor U29611 (N_29611,N_26109,N_26457);
or U29612 (N_29612,N_27673,N_26356);
nor U29613 (N_29613,N_27008,N_27482);
and U29614 (N_29614,N_26256,N_26931);
xor U29615 (N_29615,N_27643,N_26343);
xnor U29616 (N_29616,N_27822,N_27295);
or U29617 (N_29617,N_27988,N_27294);
nand U29618 (N_29618,N_26136,N_26350);
nand U29619 (N_29619,N_26442,N_27337);
xnor U29620 (N_29620,N_27102,N_26425);
xor U29621 (N_29621,N_26448,N_26121);
xor U29622 (N_29622,N_27842,N_27766);
or U29623 (N_29623,N_26245,N_26286);
nor U29624 (N_29624,N_27339,N_27012);
or U29625 (N_29625,N_27313,N_26018);
nor U29626 (N_29626,N_26520,N_27783);
xor U29627 (N_29627,N_27131,N_26639);
or U29628 (N_29628,N_26562,N_27505);
nor U29629 (N_29629,N_27508,N_26783);
nand U29630 (N_29630,N_27935,N_26637);
nand U29631 (N_29631,N_27274,N_26420);
nor U29632 (N_29632,N_26994,N_27530);
or U29633 (N_29633,N_27058,N_27381);
and U29634 (N_29634,N_27059,N_27261);
nor U29635 (N_29635,N_26992,N_27162);
and U29636 (N_29636,N_26182,N_26842);
and U29637 (N_29637,N_27541,N_26290);
nor U29638 (N_29638,N_26306,N_27896);
xnor U29639 (N_29639,N_27119,N_26673);
nand U29640 (N_29640,N_26839,N_27871);
and U29641 (N_29641,N_26865,N_26691);
and U29642 (N_29642,N_26637,N_27887);
xnor U29643 (N_29643,N_27884,N_27946);
and U29644 (N_29644,N_27712,N_27319);
or U29645 (N_29645,N_27418,N_27218);
nor U29646 (N_29646,N_27883,N_27172);
nand U29647 (N_29647,N_27206,N_27613);
and U29648 (N_29648,N_27000,N_27643);
or U29649 (N_29649,N_26068,N_26783);
and U29650 (N_29650,N_26534,N_27204);
xnor U29651 (N_29651,N_26984,N_26153);
nand U29652 (N_29652,N_27115,N_27991);
xor U29653 (N_29653,N_27213,N_27816);
xor U29654 (N_29654,N_27857,N_27513);
and U29655 (N_29655,N_26749,N_26302);
or U29656 (N_29656,N_26801,N_26976);
xnor U29657 (N_29657,N_26772,N_27457);
xor U29658 (N_29658,N_26872,N_26054);
or U29659 (N_29659,N_26561,N_26801);
xor U29660 (N_29660,N_27711,N_27487);
nand U29661 (N_29661,N_26515,N_26961);
and U29662 (N_29662,N_27343,N_27752);
nor U29663 (N_29663,N_26578,N_26117);
or U29664 (N_29664,N_26045,N_27275);
nand U29665 (N_29665,N_26346,N_27275);
and U29666 (N_29666,N_27213,N_26442);
and U29667 (N_29667,N_27114,N_26347);
and U29668 (N_29668,N_27840,N_26034);
nand U29669 (N_29669,N_27110,N_27396);
xor U29670 (N_29670,N_26777,N_26841);
or U29671 (N_29671,N_26023,N_26814);
nand U29672 (N_29672,N_26045,N_26601);
and U29673 (N_29673,N_26329,N_26558);
nand U29674 (N_29674,N_26188,N_27724);
or U29675 (N_29675,N_26494,N_26198);
or U29676 (N_29676,N_26512,N_26795);
nand U29677 (N_29677,N_26237,N_26386);
xnor U29678 (N_29678,N_27308,N_26647);
nor U29679 (N_29679,N_26347,N_27658);
nand U29680 (N_29680,N_26870,N_26729);
or U29681 (N_29681,N_27923,N_27818);
xor U29682 (N_29682,N_27109,N_27735);
and U29683 (N_29683,N_27673,N_27964);
and U29684 (N_29684,N_26207,N_27721);
nand U29685 (N_29685,N_26036,N_26307);
and U29686 (N_29686,N_27767,N_26935);
and U29687 (N_29687,N_26556,N_27007);
xor U29688 (N_29688,N_26244,N_27446);
nor U29689 (N_29689,N_27026,N_27768);
xor U29690 (N_29690,N_27560,N_26781);
or U29691 (N_29691,N_26784,N_27336);
or U29692 (N_29692,N_27939,N_27024);
or U29693 (N_29693,N_26453,N_27293);
xor U29694 (N_29694,N_27892,N_26957);
nand U29695 (N_29695,N_26538,N_27500);
xnor U29696 (N_29696,N_26575,N_26297);
and U29697 (N_29697,N_27161,N_26471);
xor U29698 (N_29698,N_27244,N_27253);
or U29699 (N_29699,N_26952,N_26967);
or U29700 (N_29700,N_27554,N_27516);
nand U29701 (N_29701,N_27850,N_27969);
or U29702 (N_29702,N_27455,N_26129);
or U29703 (N_29703,N_27126,N_26532);
xnor U29704 (N_29704,N_26310,N_26745);
and U29705 (N_29705,N_27589,N_27951);
nor U29706 (N_29706,N_26009,N_27756);
and U29707 (N_29707,N_26459,N_26543);
nor U29708 (N_29708,N_26944,N_27644);
and U29709 (N_29709,N_26828,N_26023);
xnor U29710 (N_29710,N_27611,N_27643);
or U29711 (N_29711,N_27559,N_26550);
nor U29712 (N_29712,N_27137,N_26993);
xnor U29713 (N_29713,N_26622,N_26118);
xnor U29714 (N_29714,N_26227,N_26893);
and U29715 (N_29715,N_27019,N_26653);
nor U29716 (N_29716,N_26497,N_26013);
and U29717 (N_29717,N_27177,N_27940);
nand U29718 (N_29718,N_26830,N_26790);
or U29719 (N_29719,N_27910,N_27791);
nand U29720 (N_29720,N_26024,N_26653);
nand U29721 (N_29721,N_26553,N_26362);
nand U29722 (N_29722,N_27590,N_27468);
nor U29723 (N_29723,N_26765,N_26111);
and U29724 (N_29724,N_26296,N_26859);
nor U29725 (N_29725,N_27562,N_27404);
xnor U29726 (N_29726,N_27529,N_26320);
nor U29727 (N_29727,N_26097,N_27459);
xor U29728 (N_29728,N_27162,N_26950);
nand U29729 (N_29729,N_27612,N_26429);
nor U29730 (N_29730,N_26547,N_27460);
and U29731 (N_29731,N_26968,N_27643);
or U29732 (N_29732,N_26227,N_27958);
and U29733 (N_29733,N_26890,N_27275);
and U29734 (N_29734,N_26469,N_26075);
nand U29735 (N_29735,N_26337,N_26820);
xor U29736 (N_29736,N_26047,N_27984);
nand U29737 (N_29737,N_26539,N_26633);
or U29738 (N_29738,N_27098,N_26818);
xnor U29739 (N_29739,N_27282,N_27780);
nand U29740 (N_29740,N_27453,N_27442);
xor U29741 (N_29741,N_27802,N_26186);
or U29742 (N_29742,N_27677,N_26165);
nand U29743 (N_29743,N_26154,N_26553);
and U29744 (N_29744,N_27815,N_26268);
or U29745 (N_29745,N_26404,N_27696);
xnor U29746 (N_29746,N_27771,N_27026);
nor U29747 (N_29747,N_26697,N_27773);
nor U29748 (N_29748,N_27849,N_26866);
and U29749 (N_29749,N_26238,N_26336);
nand U29750 (N_29750,N_27807,N_26977);
and U29751 (N_29751,N_26659,N_26345);
xor U29752 (N_29752,N_27734,N_26983);
or U29753 (N_29753,N_26533,N_26944);
nand U29754 (N_29754,N_26283,N_26575);
or U29755 (N_29755,N_27417,N_26168);
xnor U29756 (N_29756,N_26721,N_26637);
xor U29757 (N_29757,N_26662,N_27713);
or U29758 (N_29758,N_26417,N_26457);
nor U29759 (N_29759,N_27986,N_27304);
nand U29760 (N_29760,N_26309,N_26776);
and U29761 (N_29761,N_26345,N_27396);
or U29762 (N_29762,N_26590,N_26453);
xnor U29763 (N_29763,N_26562,N_27493);
or U29764 (N_29764,N_26345,N_27263);
or U29765 (N_29765,N_27883,N_26502);
xnor U29766 (N_29766,N_27805,N_26681);
or U29767 (N_29767,N_26189,N_27024);
and U29768 (N_29768,N_26324,N_26599);
nand U29769 (N_29769,N_27427,N_27912);
or U29770 (N_29770,N_27616,N_27721);
or U29771 (N_29771,N_27355,N_27460);
and U29772 (N_29772,N_26324,N_27110);
nand U29773 (N_29773,N_27173,N_27788);
or U29774 (N_29774,N_26785,N_26261);
or U29775 (N_29775,N_26292,N_27044);
and U29776 (N_29776,N_27815,N_27857);
or U29777 (N_29777,N_27736,N_26942);
and U29778 (N_29778,N_26854,N_27276);
nand U29779 (N_29779,N_27129,N_26603);
nor U29780 (N_29780,N_27757,N_27468);
or U29781 (N_29781,N_26186,N_26136);
nor U29782 (N_29782,N_26601,N_27768);
nand U29783 (N_29783,N_27892,N_26647);
or U29784 (N_29784,N_27401,N_27830);
nand U29785 (N_29785,N_26267,N_26704);
and U29786 (N_29786,N_26140,N_26118);
xnor U29787 (N_29787,N_26475,N_27495);
nand U29788 (N_29788,N_27356,N_27415);
and U29789 (N_29789,N_27876,N_27425);
nor U29790 (N_29790,N_27183,N_26636);
xnor U29791 (N_29791,N_26287,N_26619);
xor U29792 (N_29792,N_27420,N_27367);
nand U29793 (N_29793,N_27667,N_26549);
xnor U29794 (N_29794,N_27637,N_27350);
or U29795 (N_29795,N_27628,N_26999);
xnor U29796 (N_29796,N_26399,N_26739);
and U29797 (N_29797,N_27679,N_26701);
xor U29798 (N_29798,N_26427,N_27024);
and U29799 (N_29799,N_26081,N_26416);
xor U29800 (N_29800,N_26447,N_26448);
xnor U29801 (N_29801,N_27363,N_27931);
and U29802 (N_29802,N_26980,N_26904);
nand U29803 (N_29803,N_26403,N_26574);
nand U29804 (N_29804,N_27237,N_26265);
and U29805 (N_29805,N_26723,N_27665);
nor U29806 (N_29806,N_26425,N_27217);
and U29807 (N_29807,N_26703,N_27941);
nor U29808 (N_29808,N_26921,N_27351);
nand U29809 (N_29809,N_26763,N_26025);
or U29810 (N_29810,N_26808,N_26857);
nor U29811 (N_29811,N_27974,N_27437);
xnor U29812 (N_29812,N_26814,N_26503);
nand U29813 (N_29813,N_26127,N_26548);
nand U29814 (N_29814,N_27093,N_26954);
xor U29815 (N_29815,N_27422,N_27620);
and U29816 (N_29816,N_26648,N_27073);
xnor U29817 (N_29817,N_27595,N_26542);
xor U29818 (N_29818,N_27411,N_26738);
nand U29819 (N_29819,N_26992,N_26215);
and U29820 (N_29820,N_27571,N_26608);
xnor U29821 (N_29821,N_27276,N_26134);
xor U29822 (N_29822,N_26855,N_26103);
or U29823 (N_29823,N_26275,N_26875);
and U29824 (N_29824,N_26032,N_26571);
xnor U29825 (N_29825,N_26290,N_27899);
nand U29826 (N_29826,N_27666,N_26605);
and U29827 (N_29827,N_27728,N_27357);
and U29828 (N_29828,N_26797,N_26226);
or U29829 (N_29829,N_27725,N_27651);
nor U29830 (N_29830,N_27938,N_27200);
nor U29831 (N_29831,N_27223,N_27192);
xor U29832 (N_29832,N_27631,N_26987);
nand U29833 (N_29833,N_26512,N_27110);
nor U29834 (N_29834,N_26513,N_27662);
nor U29835 (N_29835,N_26860,N_26381);
nand U29836 (N_29836,N_26750,N_26960);
xnor U29837 (N_29837,N_26954,N_26632);
xor U29838 (N_29838,N_27979,N_27840);
xnor U29839 (N_29839,N_26820,N_26545);
and U29840 (N_29840,N_26032,N_27379);
xnor U29841 (N_29841,N_26030,N_27454);
xor U29842 (N_29842,N_26733,N_27622);
nor U29843 (N_29843,N_27008,N_27702);
or U29844 (N_29844,N_26489,N_27061);
nor U29845 (N_29845,N_26120,N_26562);
or U29846 (N_29846,N_26161,N_26079);
xor U29847 (N_29847,N_27647,N_27460);
nor U29848 (N_29848,N_26139,N_27242);
or U29849 (N_29849,N_27076,N_27641);
xor U29850 (N_29850,N_26908,N_27546);
xnor U29851 (N_29851,N_27500,N_26849);
nand U29852 (N_29852,N_26174,N_26690);
xor U29853 (N_29853,N_27157,N_26210);
xor U29854 (N_29854,N_27494,N_27720);
nand U29855 (N_29855,N_26429,N_27486);
nand U29856 (N_29856,N_26901,N_27349);
xor U29857 (N_29857,N_26226,N_26560);
nand U29858 (N_29858,N_26351,N_26580);
and U29859 (N_29859,N_27855,N_27308);
and U29860 (N_29860,N_27658,N_26323);
or U29861 (N_29861,N_26989,N_26542);
or U29862 (N_29862,N_27182,N_26496);
or U29863 (N_29863,N_27808,N_27880);
xnor U29864 (N_29864,N_26131,N_27403);
and U29865 (N_29865,N_26826,N_27343);
nand U29866 (N_29866,N_27308,N_26346);
or U29867 (N_29867,N_27705,N_27675);
nor U29868 (N_29868,N_26340,N_26209);
or U29869 (N_29869,N_26659,N_26606);
nor U29870 (N_29870,N_27461,N_26210);
nand U29871 (N_29871,N_27017,N_27460);
or U29872 (N_29872,N_27067,N_27621);
and U29873 (N_29873,N_27347,N_27534);
nand U29874 (N_29874,N_27343,N_26515);
nand U29875 (N_29875,N_26864,N_26336);
xor U29876 (N_29876,N_27306,N_27473);
nand U29877 (N_29877,N_26162,N_27814);
xnor U29878 (N_29878,N_26651,N_26654);
and U29879 (N_29879,N_26375,N_26490);
xor U29880 (N_29880,N_26916,N_26892);
xnor U29881 (N_29881,N_26583,N_27657);
nor U29882 (N_29882,N_27366,N_26610);
xnor U29883 (N_29883,N_26454,N_27234);
and U29884 (N_29884,N_26744,N_27698);
nor U29885 (N_29885,N_27850,N_26043);
nand U29886 (N_29886,N_27720,N_26703);
xor U29887 (N_29887,N_26180,N_26395);
nor U29888 (N_29888,N_27320,N_26482);
xor U29889 (N_29889,N_26872,N_26649);
and U29890 (N_29890,N_26800,N_27934);
xnor U29891 (N_29891,N_27849,N_26132);
nand U29892 (N_29892,N_27131,N_27150);
nand U29893 (N_29893,N_27206,N_26541);
and U29894 (N_29894,N_27016,N_26884);
nor U29895 (N_29895,N_26736,N_27366);
nand U29896 (N_29896,N_27001,N_27561);
and U29897 (N_29897,N_27148,N_27333);
xor U29898 (N_29898,N_27600,N_27513);
or U29899 (N_29899,N_27592,N_27658);
or U29900 (N_29900,N_27829,N_27028);
nor U29901 (N_29901,N_26971,N_27984);
nand U29902 (N_29902,N_27118,N_26481);
xnor U29903 (N_29903,N_27921,N_26467);
nor U29904 (N_29904,N_26397,N_26947);
and U29905 (N_29905,N_26337,N_26126);
and U29906 (N_29906,N_26682,N_26935);
nand U29907 (N_29907,N_27179,N_26636);
and U29908 (N_29908,N_27193,N_27244);
nor U29909 (N_29909,N_27538,N_26932);
nor U29910 (N_29910,N_27235,N_27614);
and U29911 (N_29911,N_27472,N_26040);
xor U29912 (N_29912,N_26097,N_26517);
nand U29913 (N_29913,N_26599,N_27743);
nand U29914 (N_29914,N_27150,N_26604);
xnor U29915 (N_29915,N_26884,N_27187);
nor U29916 (N_29916,N_26585,N_27005);
or U29917 (N_29917,N_27754,N_26079);
or U29918 (N_29918,N_26778,N_26606);
and U29919 (N_29919,N_26119,N_27459);
nor U29920 (N_29920,N_26663,N_26470);
nand U29921 (N_29921,N_27076,N_27607);
and U29922 (N_29922,N_27859,N_27553);
and U29923 (N_29923,N_27895,N_27361);
or U29924 (N_29924,N_26969,N_27572);
or U29925 (N_29925,N_26311,N_27679);
and U29926 (N_29926,N_26284,N_26775);
nor U29927 (N_29927,N_27336,N_27352);
nor U29928 (N_29928,N_26451,N_26014);
or U29929 (N_29929,N_27047,N_27874);
or U29930 (N_29930,N_27972,N_26724);
nor U29931 (N_29931,N_27720,N_26539);
nor U29932 (N_29932,N_26125,N_26832);
nor U29933 (N_29933,N_27496,N_27180);
xor U29934 (N_29934,N_27728,N_26599);
or U29935 (N_29935,N_26488,N_26774);
nor U29936 (N_29936,N_27780,N_27963);
nor U29937 (N_29937,N_27703,N_27139);
and U29938 (N_29938,N_27157,N_27347);
or U29939 (N_29939,N_27853,N_26383);
nand U29940 (N_29940,N_27619,N_27223);
or U29941 (N_29941,N_26681,N_27058);
nor U29942 (N_29942,N_26377,N_27190);
nand U29943 (N_29943,N_26779,N_26766);
and U29944 (N_29944,N_26625,N_27995);
nand U29945 (N_29945,N_26480,N_27042);
or U29946 (N_29946,N_26575,N_26994);
xor U29947 (N_29947,N_27729,N_27385);
or U29948 (N_29948,N_26640,N_27054);
xnor U29949 (N_29949,N_26743,N_26459);
nand U29950 (N_29950,N_26346,N_27646);
and U29951 (N_29951,N_26722,N_26577);
xor U29952 (N_29952,N_27839,N_27034);
or U29953 (N_29953,N_26166,N_26785);
or U29954 (N_29954,N_27653,N_26207);
xor U29955 (N_29955,N_27579,N_26460);
nand U29956 (N_29956,N_27696,N_26044);
and U29957 (N_29957,N_26196,N_26506);
and U29958 (N_29958,N_26157,N_27575);
xor U29959 (N_29959,N_27743,N_26781);
xor U29960 (N_29960,N_26503,N_27976);
or U29961 (N_29961,N_26804,N_27700);
nor U29962 (N_29962,N_27979,N_26459);
nand U29963 (N_29963,N_27540,N_27610);
xnor U29964 (N_29964,N_27330,N_26735);
xor U29965 (N_29965,N_26425,N_26971);
nand U29966 (N_29966,N_26304,N_26929);
or U29967 (N_29967,N_26960,N_26880);
or U29968 (N_29968,N_26391,N_27075);
nor U29969 (N_29969,N_27909,N_27464);
and U29970 (N_29970,N_26455,N_26052);
xnor U29971 (N_29971,N_26144,N_27431);
and U29972 (N_29972,N_27945,N_27204);
nor U29973 (N_29973,N_26312,N_27796);
and U29974 (N_29974,N_26812,N_26934);
nor U29975 (N_29975,N_27921,N_27730);
nand U29976 (N_29976,N_27171,N_27677);
nand U29977 (N_29977,N_27728,N_27843);
or U29978 (N_29978,N_27123,N_27310);
or U29979 (N_29979,N_27015,N_26534);
nor U29980 (N_29980,N_26361,N_26685);
or U29981 (N_29981,N_26233,N_26309);
or U29982 (N_29982,N_26634,N_27503);
and U29983 (N_29983,N_27809,N_26001);
xor U29984 (N_29984,N_27963,N_27323);
or U29985 (N_29985,N_26393,N_27501);
xor U29986 (N_29986,N_26604,N_26537);
nand U29987 (N_29987,N_26281,N_26865);
nand U29988 (N_29988,N_27819,N_27107);
nand U29989 (N_29989,N_26927,N_27617);
or U29990 (N_29990,N_26785,N_27846);
nand U29991 (N_29991,N_27371,N_26082);
nand U29992 (N_29992,N_26173,N_27952);
nand U29993 (N_29993,N_27751,N_27396);
nand U29994 (N_29994,N_26534,N_27372);
xnor U29995 (N_29995,N_27806,N_26472);
and U29996 (N_29996,N_26911,N_27130);
or U29997 (N_29997,N_27109,N_26440);
or U29998 (N_29998,N_26815,N_26507);
and U29999 (N_29999,N_27393,N_27861);
and U30000 (N_30000,N_29829,N_29609);
xor U30001 (N_30001,N_28606,N_28626);
or U30002 (N_30002,N_29864,N_28137);
nor U30003 (N_30003,N_28037,N_28923);
xor U30004 (N_30004,N_29557,N_28162);
nand U30005 (N_30005,N_29811,N_29241);
and U30006 (N_30006,N_29381,N_29880);
nor U30007 (N_30007,N_28552,N_28382);
nand U30008 (N_30008,N_29098,N_29224);
nand U30009 (N_30009,N_28328,N_28012);
and U30010 (N_30010,N_29531,N_28129);
and U30011 (N_30011,N_29397,N_28106);
xnor U30012 (N_30012,N_28995,N_28958);
nand U30013 (N_30013,N_29756,N_29147);
or U30014 (N_30014,N_29968,N_29665);
xnor U30015 (N_30015,N_28721,N_29136);
nand U30016 (N_30016,N_29010,N_29475);
xor U30017 (N_30017,N_28863,N_29998);
xor U30018 (N_30018,N_29121,N_28185);
or U30019 (N_30019,N_28718,N_29799);
nand U30020 (N_30020,N_29697,N_28864);
or U30021 (N_30021,N_28160,N_28984);
and U30022 (N_30022,N_29419,N_29584);
or U30023 (N_30023,N_28269,N_28642);
xnor U30024 (N_30024,N_29912,N_28372);
nand U30025 (N_30025,N_28108,N_29384);
and U30026 (N_30026,N_29644,N_28885);
xor U30027 (N_30027,N_29634,N_29480);
or U30028 (N_30028,N_28837,N_29863);
nand U30029 (N_30029,N_28409,N_28332);
nand U30030 (N_30030,N_28579,N_28344);
or U30031 (N_30031,N_29095,N_29738);
xnor U30032 (N_30032,N_28595,N_29960);
xnor U30033 (N_30033,N_28479,N_28002);
and U30034 (N_30034,N_29619,N_28508);
and U30035 (N_30035,N_28191,N_28125);
xnor U30036 (N_30036,N_29306,N_29698);
nor U30037 (N_30037,N_29303,N_28456);
and U30038 (N_30038,N_29356,N_28325);
or U30039 (N_30039,N_29153,N_29656);
or U30040 (N_30040,N_28932,N_29714);
xor U30041 (N_30041,N_28458,N_29749);
nor U30042 (N_30042,N_28820,N_28169);
and U30043 (N_30043,N_28460,N_29739);
nand U30044 (N_30044,N_28340,N_28588);
or U30045 (N_30045,N_28273,N_29175);
nor U30046 (N_30046,N_29130,N_28555);
and U30047 (N_30047,N_28636,N_28951);
xnor U30048 (N_30048,N_28693,N_28940);
nand U30049 (N_30049,N_29393,N_28713);
nand U30050 (N_30050,N_28445,N_28838);
or U30051 (N_30051,N_28538,N_29786);
nand U30052 (N_30052,N_29598,N_29457);
and U30053 (N_30053,N_28462,N_29509);
or U30054 (N_30054,N_28289,N_28966);
or U30055 (N_30055,N_29802,N_28893);
xor U30056 (N_30056,N_29637,N_29294);
nor U30057 (N_30057,N_29783,N_29488);
or U30058 (N_30058,N_29309,N_29441);
xnor U30059 (N_30059,N_28985,N_28607);
and U30060 (N_30060,N_28979,N_28374);
nor U30061 (N_30061,N_28840,N_28824);
or U30062 (N_30062,N_28154,N_29345);
or U30063 (N_30063,N_28926,N_29617);
nor U30064 (N_30064,N_29624,N_29431);
or U30065 (N_30065,N_29769,N_29360);
nand U30066 (N_30066,N_28829,N_28878);
xor U30067 (N_30067,N_28298,N_28691);
and U30068 (N_30068,N_29128,N_28706);
and U30069 (N_30069,N_29784,N_29501);
nand U30070 (N_30070,N_28165,N_29762);
xnor U30071 (N_30071,N_28876,N_28723);
xnor U30072 (N_30072,N_29366,N_29329);
nor U30073 (N_30073,N_29975,N_29026);
and U30074 (N_30074,N_29442,N_28288);
xor U30075 (N_30075,N_28021,N_29704);
or U30076 (N_30076,N_28050,N_28174);
and U30077 (N_30077,N_28381,N_28939);
xor U30078 (N_30078,N_28076,N_28310);
and U30079 (N_30079,N_28234,N_29641);
xor U30080 (N_30080,N_28114,N_28099);
nor U30081 (N_30081,N_28272,N_28069);
nor U30082 (N_30082,N_29801,N_28687);
or U30083 (N_30083,N_28354,N_28390);
and U30084 (N_30084,N_29422,N_29909);
nand U30085 (N_30085,N_28350,N_29196);
nor U30086 (N_30086,N_29893,N_29974);
nand U30087 (N_30087,N_28625,N_29058);
nor U30088 (N_30088,N_28281,N_28361);
xnor U30089 (N_30089,N_28004,N_28360);
nor U30090 (N_30090,N_28639,N_28250);
xor U30091 (N_30091,N_28241,N_29823);
or U30092 (N_30092,N_28286,N_29396);
and U30093 (N_30093,N_29293,N_28919);
xor U30094 (N_30094,N_29179,N_29340);
nor U30095 (N_30095,N_28722,N_29161);
xor U30096 (N_30096,N_29251,N_28148);
nand U30097 (N_30097,N_29227,N_29141);
or U30098 (N_30098,N_28735,N_29857);
nor U30099 (N_30099,N_28854,N_29590);
xor U30100 (N_30100,N_28578,N_28535);
and U30101 (N_30101,N_28484,N_29220);
xnor U30102 (N_30102,N_28425,N_28686);
and U30103 (N_30103,N_28637,N_28983);
nand U30104 (N_30104,N_29674,N_28957);
nand U30105 (N_30105,N_28355,N_29253);
or U30106 (N_30106,N_29677,N_29006);
xor U30107 (N_30107,N_28821,N_29032);
nand U30108 (N_30108,N_29803,N_28223);
and U30109 (N_30109,N_29187,N_29159);
nand U30110 (N_30110,N_29407,N_29699);
and U30111 (N_30111,N_29625,N_29773);
nor U30112 (N_30112,N_29341,N_28244);
or U30113 (N_30113,N_29719,N_29631);
nand U30114 (N_30114,N_29229,N_28378);
or U30115 (N_30115,N_28600,N_28225);
or U30116 (N_30116,N_29533,N_28815);
xor U30117 (N_30117,N_29449,N_29069);
nand U30118 (N_30118,N_28717,N_29410);
and U30119 (N_30119,N_29920,N_28008);
nand U30120 (N_30120,N_29458,N_28480);
nand U30121 (N_30121,N_29482,N_29554);
and U30122 (N_30122,N_29589,N_28377);
xnor U30123 (N_30123,N_29859,N_28442);
xnor U30124 (N_30124,N_29603,N_29020);
or U30125 (N_30125,N_29398,N_29191);
and U30126 (N_30126,N_29537,N_29242);
nand U30127 (N_30127,N_28605,N_28113);
nor U30128 (N_30128,N_29160,N_28653);
and U30129 (N_30129,N_28331,N_28088);
nand U30130 (N_30130,N_29831,N_28300);
nand U30131 (N_30131,N_29945,N_29670);
nand U30132 (N_30132,N_29099,N_29135);
or U30133 (N_30133,N_28565,N_28036);
xor U30134 (N_30134,N_28173,N_28924);
or U30135 (N_30135,N_29074,N_28655);
nor U30136 (N_30136,N_28909,N_28765);
or U30137 (N_30137,N_29228,N_29133);
xnor U30138 (N_30138,N_28055,N_28439);
xnor U30139 (N_30139,N_29922,N_29065);
nor U30140 (N_30140,N_29225,N_28093);
nand U30141 (N_30141,N_29205,N_28776);
nor U30142 (N_30142,N_28391,N_28194);
nand U30143 (N_30143,N_28187,N_29914);
or U30144 (N_30144,N_29351,N_28712);
nand U30145 (N_30145,N_28715,N_29226);
nand U30146 (N_30146,N_29182,N_29260);
nand U30147 (N_30147,N_28451,N_29266);
xnor U30148 (N_30148,N_29737,N_29887);
nor U30149 (N_30149,N_28965,N_29497);
nand U30150 (N_30150,N_29888,N_28074);
or U30151 (N_30151,N_28942,N_28949);
or U30152 (N_30152,N_28168,N_28058);
nand U30153 (N_30153,N_28911,N_28211);
nor U30154 (N_30154,N_28816,N_29275);
and U30155 (N_30155,N_29576,N_29889);
nand U30156 (N_30156,N_29519,N_29639);
nor U30157 (N_30157,N_28976,N_29597);
nand U30158 (N_30158,N_29499,N_29405);
xnor U30159 (N_30159,N_29729,N_29392);
xnor U30160 (N_30160,N_28163,N_28351);
nor U30161 (N_30161,N_29595,N_29828);
nor U30162 (N_30162,N_29165,N_28769);
nand U30163 (N_30163,N_29038,N_29152);
nor U30164 (N_30164,N_28515,N_29621);
or U30165 (N_30165,N_29461,N_28930);
or U30166 (N_30166,N_29800,N_29292);
and U30167 (N_30167,N_29459,N_28753);
xor U30168 (N_30168,N_28539,N_28574);
nor U30169 (N_30169,N_29472,N_28231);
nand U30170 (N_30170,N_29940,N_28054);
xor U30171 (N_30171,N_29751,N_29297);
or U30172 (N_30172,N_29666,N_29939);
and U30173 (N_30173,N_28516,N_28274);
xnor U30174 (N_30174,N_29653,N_29562);
nand U30175 (N_30175,N_28373,N_28233);
nand U30176 (N_30176,N_28592,N_29463);
and U30177 (N_30177,N_28570,N_29898);
nor U30178 (N_30178,N_29701,N_28857);
nand U30179 (N_30179,N_29223,N_28399);
xnor U30180 (N_30180,N_28665,N_28183);
nand U30181 (N_30181,N_28363,N_28386);
or U30182 (N_30182,N_29417,N_28748);
or U30183 (N_30183,N_28556,N_28783);
or U30184 (N_30184,N_29148,N_28963);
nor U30185 (N_30185,N_28064,N_28464);
nor U30186 (N_30186,N_29623,N_29996);
nand U30187 (N_30187,N_29155,N_28259);
and U30188 (N_30188,N_28469,N_29250);
nor U30189 (N_30189,N_28400,N_29834);
xnor U30190 (N_30190,N_29540,N_29782);
or U30191 (N_30191,N_29365,N_29296);
nor U30192 (N_30192,N_29234,N_29416);
xor U30193 (N_30193,N_29096,N_28964);
xnor U30194 (N_30194,N_28337,N_28405);
nor U30195 (N_30195,N_29307,N_28827);
nor U30196 (N_30196,N_28845,N_28703);
nor U30197 (N_30197,N_28950,N_29087);
nand U30198 (N_30198,N_29401,N_29913);
nand U30199 (N_30199,N_28034,N_29308);
nor U30200 (N_30200,N_29336,N_28887);
nand U30201 (N_30201,N_28334,N_28192);
xnor U30202 (N_30202,N_28773,N_28726);
nand U30203 (N_30203,N_29288,N_29832);
xnor U30204 (N_30204,N_29156,N_29890);
xnor U30205 (N_30205,N_29273,N_28629);
nor U30206 (N_30206,N_29197,N_28052);
or U30207 (N_30207,N_29511,N_28415);
nor U30208 (N_30208,N_29916,N_29867);
xor U30209 (N_30209,N_29077,N_29319);
nor U30210 (N_30210,N_29040,N_28678);
and U30211 (N_30211,N_29048,N_28254);
or U30212 (N_30212,N_28151,N_29219);
and U30213 (N_30213,N_28253,N_28448);
or U30214 (N_30214,N_28784,N_29648);
nor U30215 (N_30215,N_29795,N_28772);
and U30216 (N_30216,N_29917,N_28463);
xor U30217 (N_30217,N_28610,N_29851);
nand U30218 (N_30218,N_28802,N_29462);
nand U30219 (N_30219,N_28696,N_28246);
nand U30220 (N_30220,N_29139,N_28920);
nor U30221 (N_30221,N_29185,N_29728);
nand U30222 (N_30222,N_28514,N_29490);
and U30223 (N_30223,N_28850,N_28537);
nor U30224 (N_30224,N_29777,N_28486);
nand U30225 (N_30225,N_28488,N_28195);
and U30226 (N_30226,N_29532,N_28754);
nand U30227 (N_30227,N_28471,N_28338);
and U30228 (N_30228,N_28710,N_29715);
nor U30229 (N_30229,N_28856,N_28228);
nand U30230 (N_30230,N_29189,N_29173);
or U30231 (N_30231,N_28811,N_29243);
and U30232 (N_30232,N_28212,N_28482);
xor U30233 (N_30233,N_28157,N_29259);
nand U30234 (N_30234,N_28658,N_28199);
nor U30235 (N_30235,N_29053,N_29723);
xor U30236 (N_30236,N_28063,N_28413);
nor U30237 (N_30237,N_29316,N_29444);
nor U30238 (N_30238,N_29702,N_29211);
xor U30239 (N_30239,N_28743,N_29051);
and U30240 (N_30240,N_29369,N_28520);
nand U30241 (N_30241,N_28899,N_28265);
or U30242 (N_30242,N_28644,N_28872);
and U30243 (N_30243,N_29808,N_29836);
or U30244 (N_30244,N_28329,N_29201);
and U30245 (N_30245,N_28559,N_28522);
nor U30246 (N_30246,N_29796,N_29233);
nor U30247 (N_30247,N_29947,N_28420);
nand U30248 (N_30248,N_28181,N_28683);
nor U30249 (N_30249,N_29549,N_28819);
or U30250 (N_30250,N_28379,N_28098);
nor U30251 (N_30251,N_28122,N_28356);
xor U30252 (N_30252,N_28201,N_28142);
nor U30253 (N_30253,N_29334,N_28299);
xnor U30254 (N_30254,N_28789,N_28818);
or U30255 (N_30255,N_29385,N_29951);
and U30256 (N_30256,N_28204,N_29108);
or U30257 (N_30257,N_29843,N_28348);
nand U30258 (N_30258,N_29237,N_28842);
nor U30259 (N_30259,N_28944,N_28708);
nor U30260 (N_30260,N_28364,N_28190);
or U30261 (N_30261,N_29391,N_29055);
and U30262 (N_30262,N_29302,N_28466);
nor U30263 (N_30263,N_28280,N_29199);
or U30264 (N_30264,N_28068,N_29232);
and U30265 (N_30265,N_29818,N_28673);
nand U30266 (N_30266,N_28057,N_29717);
nand U30267 (N_30267,N_29082,N_28627);
or U30268 (N_30268,N_28022,N_29630);
or U30269 (N_30269,N_28918,N_29587);
xnor U30270 (N_30270,N_29981,N_28970);
nor U30271 (N_30271,N_28764,N_28719);
nor U30272 (N_30272,N_28621,N_29426);
nand U30273 (N_30273,N_28436,N_29412);
and U30274 (N_30274,N_28327,N_29269);
nor U30275 (N_30275,N_28132,N_29992);
nor U30276 (N_30276,N_28105,N_29985);
nand U30277 (N_30277,N_29477,N_29815);
nand U30278 (N_30278,N_28035,N_29989);
xnor U30279 (N_30279,N_28198,N_28188);
or U30280 (N_30280,N_29097,N_29467);
nand U30281 (N_30281,N_28871,N_28407);
nor U30282 (N_30282,N_28575,N_28264);
xor U30283 (N_30283,N_29868,N_28224);
nand U30284 (N_30284,N_28144,N_28416);
nand U30285 (N_30285,N_29675,N_28504);
and U30286 (N_30286,N_28603,N_28127);
nand U30287 (N_30287,N_28077,N_29740);
or U30288 (N_30288,N_29725,N_29635);
or U30289 (N_30289,N_28345,N_29807);
and U30290 (N_30290,N_28015,N_29395);
nand U30291 (N_30291,N_29325,N_29057);
xnor U30292 (N_30292,N_29854,N_29983);
xnor U30293 (N_30293,N_28741,N_28524);
xor U30294 (N_30294,N_28503,N_29708);
or U30295 (N_30295,N_28179,N_28905);
and U30296 (N_30296,N_28852,N_29484);
nor U30297 (N_30297,N_28526,N_29137);
and U30298 (N_30298,N_28116,N_29797);
nor U30299 (N_30299,N_28807,N_28397);
nor U30300 (N_30300,N_28252,N_28271);
or U30301 (N_30301,N_28525,N_29936);
nand U30302 (N_30302,N_28548,N_28060);
and U30303 (N_30303,N_28417,N_29346);
nor U30304 (N_30304,N_29037,N_29169);
nand U30305 (N_30305,N_28581,N_28357);
or U30306 (N_30306,N_29882,N_28270);
nand U30307 (N_30307,N_28256,N_29453);
nor U30308 (N_30308,N_28751,N_28564);
xor U30309 (N_30309,N_29314,N_28682);
and U30310 (N_30310,N_29892,N_29886);
nor U30311 (N_30311,N_28330,N_28608);
xnor U30312 (N_30312,N_29869,N_29036);
and U30313 (N_30313,N_28041,N_29663);
or U30314 (N_30314,N_29425,N_28907);
or U30315 (N_30315,N_29208,N_29215);
xor U30316 (N_30316,N_28306,N_29937);
nand U30317 (N_30317,N_29620,N_28883);
nor U30318 (N_30318,N_28779,N_28652);
or U30319 (N_30319,N_28229,N_29387);
nand U30320 (N_30320,N_29944,N_29256);
nand U30321 (N_30321,N_29279,N_29154);
xor U30322 (N_30322,N_28346,N_29669);
xnor U30323 (N_30323,N_29004,N_28571);
or U30324 (N_30324,N_28701,N_28793);
xor U30325 (N_30325,N_28146,N_28990);
and U30326 (N_30326,N_28029,N_28688);
or U30327 (N_30327,N_28534,N_29041);
or U30328 (N_30328,N_28095,N_28103);
or U30329 (N_30329,N_29235,N_29700);
xor U30330 (N_30330,N_28238,N_29768);
and U30331 (N_30331,N_29967,N_29984);
xor U30332 (N_30332,N_29206,N_28955);
xnor U30333 (N_30333,N_28669,N_29849);
nor U30334 (N_30334,N_28728,N_29817);
or U30335 (N_30335,N_28855,N_29632);
nor U30336 (N_30336,N_28066,N_28744);
xor U30337 (N_30337,N_28203,N_29638);
nand U30338 (N_30338,N_28962,N_29753);
and U30339 (N_30339,N_28999,N_28171);
or U30340 (N_30340,N_29861,N_28900);
xor U30341 (N_30341,N_28767,N_29907);
and U30342 (N_30342,N_28075,N_29933);
nor U30343 (N_30343,N_29517,N_28178);
xor U30344 (N_30344,N_28542,N_29915);
and U30345 (N_30345,N_28205,N_28236);
nor U30346 (N_30346,N_29645,N_28953);
or U30347 (N_30347,N_29493,N_29918);
xnor U30348 (N_30348,N_29627,N_28489);
xor U30349 (N_30349,N_28470,N_29195);
nand U30350 (N_30350,N_29021,N_28841);
nor U30351 (N_30351,N_28695,N_29473);
nand U30352 (N_30352,N_28287,N_29448);
nor U30353 (N_30353,N_29932,N_28319);
or U30354 (N_30354,N_29962,N_29485);
xor U30355 (N_30355,N_28352,N_28938);
nor U30356 (N_30356,N_29776,N_29420);
nand U30357 (N_30357,N_28597,N_28267);
nor U30358 (N_30358,N_29840,N_29774);
nor U30359 (N_30359,N_29327,N_29418);
or U30360 (N_30360,N_28993,N_29378);
nor U30361 (N_30361,N_29508,N_28646);
nand U30362 (N_30362,N_28822,N_29093);
and U30363 (N_30363,N_29551,N_28017);
xnor U30364 (N_30364,N_28278,N_28622);
nand U30365 (N_30365,N_29899,N_29368);
nor U30366 (N_30366,N_29231,N_28320);
nand U30367 (N_30367,N_29804,N_28517);
nor U30368 (N_30368,N_29607,N_29498);
nor U30369 (N_30369,N_28768,N_29982);
and U30370 (N_30370,N_28509,N_29359);
and U30371 (N_30371,N_28609,N_29186);
nor U30372 (N_30372,N_29837,N_28813);
xor U30373 (N_30373,N_29112,N_28974);
nor U30374 (N_30374,N_28086,N_28175);
and U30375 (N_30375,N_28679,N_28312);
nor U30376 (N_30376,N_29657,N_29612);
nand U30377 (N_30377,N_29094,N_29436);
nor U30378 (N_30378,N_29122,N_28189);
nand U30379 (N_30379,N_29556,N_29820);
and U30380 (N_30380,N_29927,N_29027);
xnor U30381 (N_30381,N_28014,N_29692);
or U30382 (N_30382,N_28851,N_29568);
or U30383 (N_30383,N_29317,N_28638);
or U30384 (N_30384,N_28112,N_29144);
nor U30385 (N_30385,N_29794,N_29954);
nand U30386 (N_30386,N_29980,N_29878);
xor U30387 (N_30387,N_28670,N_28121);
nor U30388 (N_30388,N_29658,N_28573);
nand U30389 (N_30389,N_29895,N_29901);
or U30390 (N_30390,N_28365,N_28794);
nor U30391 (N_30391,N_29299,N_29813);
nand U30392 (N_30392,N_29247,N_29158);
and U30393 (N_30393,N_28933,N_29850);
nand U30394 (N_30394,N_29421,N_29403);
nor U30395 (N_30395,N_28643,N_29236);
nor U30396 (N_30396,N_29295,N_28619);
nand U30397 (N_30397,N_29758,N_29547);
or U30398 (N_30398,N_29879,N_28011);
nor U30399 (N_30399,N_28598,N_29548);
nand U30400 (N_30400,N_28847,N_29044);
and U30401 (N_30401,N_28888,N_29078);
nand U30402 (N_30402,N_29382,N_29732);
and U30403 (N_30403,N_29827,N_29125);
nor U30404 (N_30404,N_29935,N_29957);
or U30405 (N_30405,N_29846,N_28560);
nand U30406 (N_30406,N_28586,N_28410);
xor U30407 (N_30407,N_28694,N_28587);
nor U30408 (N_30408,N_28633,N_28197);
nor U30409 (N_30409,N_28967,N_28874);
xor U30410 (N_30410,N_28785,N_29290);
nor U30411 (N_30411,N_29443,N_28868);
or U30412 (N_30412,N_29263,N_29118);
or U30413 (N_30413,N_28159,N_28833);
or U30414 (N_30414,N_28620,N_28936);
xor U30415 (N_30415,N_29566,N_28533);
nand U30416 (N_30416,N_29860,N_29386);
xor U30417 (N_30417,N_29583,N_29924);
xnor U30418 (N_30418,N_28946,N_28875);
nand U30419 (N_30419,N_29103,N_29522);
and U30420 (N_30420,N_29676,N_29202);
or U30421 (N_30421,N_28853,N_29791);
and U30422 (N_30422,N_29973,N_28156);
nor U30423 (N_30423,N_28446,N_29281);
nand U30424 (N_30424,N_28831,N_28495);
and U30425 (N_30425,N_29560,N_29976);
and U30426 (N_30426,N_28155,N_29427);
nor U30427 (N_30427,N_29249,N_28294);
nor U30428 (N_30428,N_29865,N_28707);
xor U30429 (N_30429,N_28640,N_29798);
and U30430 (N_30430,N_28368,N_28040);
nand U30431 (N_30431,N_29614,N_29724);
nor U30432 (N_30432,N_28681,N_29505);
nor U30433 (N_30433,N_29399,N_28805);
and U30434 (N_30434,N_29239,N_28677);
and U30435 (N_30435,N_29706,N_29287);
and U30436 (N_30436,N_29034,N_28759);
or U30437 (N_30437,N_29582,N_28832);
and U30438 (N_30438,N_29476,N_28865);
and U30439 (N_30439,N_28322,N_29563);
and U30440 (N_30440,N_28038,N_29184);
and U30441 (N_30441,N_29544,N_28049);
xor U30442 (N_30442,N_28929,N_28649);
xor U30443 (N_30443,N_29323,N_28553);
nand U30444 (N_30444,N_28998,N_28947);
or U30445 (N_30445,N_29993,N_29622);
and U30446 (N_30446,N_28227,N_29528);
and U30447 (N_30447,N_28859,N_28825);
and U30448 (N_30448,N_29602,N_28921);
xnor U30449 (N_30449,N_28800,N_28161);
nand U30450 (N_30450,N_28455,N_29321);
or U30451 (N_30451,N_28523,N_29902);
nand U30452 (N_30452,N_29163,N_28120);
nor U30453 (N_30453,N_29730,N_28787);
and U30454 (N_30454,N_28910,N_28795);
nand U30455 (N_30455,N_28797,N_28616);
nor U30456 (N_30456,N_28690,N_28725);
xor U30457 (N_30457,N_29240,N_29885);
xnor U30458 (N_30458,N_28437,N_29580);
xor U30459 (N_30459,N_28305,N_28081);
xor U30460 (N_30460,N_29372,N_28654);
and U30461 (N_30461,N_28981,N_29310);
xor U30462 (N_30462,N_28362,N_29322);
nand U30463 (N_30463,N_28762,N_28303);
and U30464 (N_30464,N_28558,N_29601);
or U30465 (N_30465,N_28782,N_28136);
or U30466 (N_30466,N_29066,N_28492);
nor U30467 (N_30467,N_29212,N_28118);
and U30468 (N_30468,N_29031,N_29304);
and U30469 (N_30469,N_29111,N_28884);
or U30470 (N_30470,N_28430,N_28182);
nand U30471 (N_30471,N_28485,N_28353);
nor U30472 (N_30472,N_28546,N_28247);
nand U30473 (N_30473,N_28001,N_29763);
xnor U30474 (N_30474,N_29991,N_29588);
or U30475 (N_30475,N_28528,N_28554);
nor U30476 (N_30476,N_29192,N_28072);
nor U30477 (N_30477,N_29514,N_28367);
or U30478 (N_30478,N_28333,N_28343);
or U30479 (N_30479,N_28803,N_29842);
or U30480 (N_30480,N_28576,N_29636);
and U30481 (N_30481,N_28734,N_29157);
or U30482 (N_30482,N_28006,N_29883);
or U30483 (N_30483,N_29324,N_29605);
xnor U30484 (N_30484,N_29571,N_28497);
or U30485 (N_30485,N_28843,N_29358);
xnor U30486 (N_30486,N_29995,N_29780);
nand U30487 (N_30487,N_29106,N_28214);
nand U30488 (N_30488,N_29862,N_29997);
or U30489 (N_30489,N_29305,N_28674);
and U30490 (N_30490,N_29084,N_28230);
or U30491 (N_30491,N_29838,N_29592);
or U30492 (N_30492,N_28781,N_28218);
nor U30493 (N_30493,N_28452,N_28704);
nor U30494 (N_30494,N_29203,N_29207);
nand U30495 (N_30495,N_28295,N_28048);
nor U30496 (N_30496,N_28697,N_29526);
xor U30497 (N_30497,N_28501,N_29090);
and U30498 (N_30498,N_28323,N_28000);
nand U30499 (N_30499,N_29971,N_29143);
nor U30500 (N_30500,N_29142,N_29017);
nand U30501 (N_30501,N_29440,N_29565);
and U30502 (N_30502,N_29874,N_28235);
nor U30503 (N_30503,N_28078,N_28483);
nor U30504 (N_30504,N_29703,N_28758);
nor U30505 (N_30505,N_28167,N_29705);
or U30506 (N_30506,N_28097,N_28315);
or U30507 (N_30507,N_28044,N_29897);
nor U30508 (N_30508,N_29925,N_29694);
or U30509 (N_30509,N_29711,N_29331);
or U30510 (N_30510,N_28019,N_28358);
or U30511 (N_30511,N_28130,N_29109);
or U30512 (N_30512,N_28913,N_29257);
or U30513 (N_30513,N_28262,N_28716);
nand U30514 (N_30514,N_28711,N_29848);
xnor U30515 (N_30515,N_28336,N_29423);
nand U30516 (N_30516,N_29138,N_28196);
xnor U30517 (N_30517,N_29437,N_29262);
xnor U30518 (N_30518,N_28749,N_29651);
xor U30519 (N_30519,N_29948,N_28059);
or U30520 (N_30520,N_28904,N_29001);
or U30521 (N_30521,N_28651,N_29367);
or U30522 (N_30522,N_29569,N_29685);
and U30523 (N_30523,N_29682,N_29131);
or U30524 (N_30524,N_28527,N_29743);
or U30525 (N_30525,N_29687,N_29478);
nand U30526 (N_30526,N_29012,N_29668);
nor U30527 (N_30527,N_28213,N_29516);
and U30528 (N_30528,N_28429,N_29966);
nand U30529 (N_30529,N_29835,N_28172);
or U30530 (N_30530,N_28792,N_29767);
and U30531 (N_30531,N_28302,N_29626);
or U30532 (N_30532,N_28561,N_29083);
xnor U30533 (N_30533,N_29910,N_29999);
xnor U30534 (N_30534,N_29429,N_28170);
and U30535 (N_30535,N_29722,N_28285);
and U30536 (N_30536,N_28209,N_29267);
xor U30537 (N_30537,N_29552,N_29650);
and U30538 (N_30538,N_28870,N_28659);
or U30539 (N_30539,N_28317,N_29013);
xor U30540 (N_30540,N_28613,N_29350);
nand U30541 (N_30541,N_28176,N_28449);
or U30542 (N_30542,N_28860,N_29896);
xor U30543 (N_30543,N_29190,N_29390);
or U30544 (N_30544,N_29430,N_29370);
and U30545 (N_30545,N_28304,N_29757);
xor U30546 (N_30546,N_29716,N_28771);
or U30547 (N_30547,N_28432,N_28612);
or U30548 (N_30548,N_28505,N_29222);
xnor U30549 (N_30549,N_28177,N_29613);
nor U30550 (N_30550,N_29943,N_29755);
nor U30551 (N_30551,N_29474,N_28258);
nor U30552 (N_30552,N_29546,N_28729);
nor U30553 (N_30553,N_29271,N_28914);
nand U30554 (N_30554,N_29481,N_28567);
nor U30555 (N_30555,N_29465,N_29075);
xnor U30556 (N_30556,N_29919,N_28882);
xnor U30557 (N_30557,N_28839,N_28275);
nand U30558 (N_30558,N_28020,N_29760);
xnor U30559 (N_30559,N_28318,N_29789);
xor U30560 (N_30560,N_28786,N_28994);
nand U30561 (N_30561,N_29752,N_29091);
nand U30562 (N_30562,N_28846,N_28518);
nand U30563 (N_30563,N_29718,N_29400);
nand U30564 (N_30564,N_28934,N_29002);
or U30565 (N_30565,N_28880,N_29050);
xnor U30566 (N_30566,N_28817,N_29357);
xnor U30567 (N_30567,N_29105,N_28917);
and U30568 (N_30568,N_29447,N_29388);
nand U30569 (N_30569,N_29956,N_28061);
nor U30570 (N_30570,N_29332,N_29347);
xor U30571 (N_30571,N_28084,N_28110);
and U30572 (N_30572,N_29438,N_29567);
nand U30573 (N_30573,N_28065,N_28242);
nand U30574 (N_30574,N_29364,N_29979);
xor U30575 (N_30575,N_29963,N_28208);
nand U30576 (N_30576,N_29853,N_29339);
nand U30577 (N_30577,N_28540,N_29335);
or U30578 (N_30578,N_28996,N_29214);
nor U30579 (N_30579,N_29486,N_29023);
nor U30580 (N_30580,N_28263,N_28309);
and U30581 (N_30581,N_29502,N_28862);
or U30582 (N_30582,N_29894,N_28891);
nand U30583 (N_30583,N_29553,N_29949);
and U30584 (N_30584,N_28507,N_28487);
or U30585 (N_30585,N_29671,N_29830);
nand U30586 (N_30586,N_28389,N_28062);
and U30587 (N_30587,N_29469,N_28873);
and U30588 (N_30588,N_28277,N_29129);
and U30589 (N_30589,N_28740,N_29535);
nand U30590 (N_30590,N_28780,N_29527);
and U30591 (N_30591,N_28790,N_29140);
nor U30592 (N_30592,N_29745,N_29466);
nand U30593 (N_30593,N_29070,N_28268);
nand U30594 (N_30594,N_29080,N_28869);
nand U30595 (N_30595,N_29348,N_29930);
nand U30596 (N_30596,N_28153,N_29411);
and U30597 (N_30597,N_29404,N_28543);
nand U30598 (N_30598,N_29283,N_29043);
and U30599 (N_30599,N_29286,N_29424);
and U30600 (N_30600,N_28519,N_29060);
or U30601 (N_30601,N_28510,N_28801);
xnor U30602 (N_30602,N_29819,N_29629);
or U30603 (N_30603,N_29904,N_29270);
nand U30604 (N_30604,N_28849,N_29633);
xnor U30605 (N_30605,N_29076,N_29394);
xor U30606 (N_30606,N_29679,N_29510);
or U30607 (N_30607,N_28039,N_28927);
nor U30608 (N_30608,N_28491,N_29117);
nor U30609 (N_30609,N_28394,N_28890);
xor U30610 (N_30610,N_29726,N_28474);
nor U30611 (N_30611,N_29151,N_28745);
nor U30612 (N_30612,N_28667,N_28809);
nand U30613 (N_30613,N_29759,N_28023);
xnor U30614 (N_30614,N_28698,N_29355);
and U30615 (N_30615,N_28844,N_29019);
or U30616 (N_30616,N_29712,N_28089);
nor U30617 (N_30617,N_28757,N_28594);
nand U30618 (N_30618,N_28147,N_29389);
xor U30619 (N_30619,N_29529,N_29961);
nor U30620 (N_30620,N_29684,N_28403);
or U30621 (N_30621,N_28671,N_28080);
and U30622 (N_30622,N_29343,N_28447);
nand U30623 (N_30623,N_28433,N_29825);
xor U30624 (N_30624,N_29809,N_28016);
or U30625 (N_30625,N_28541,N_29216);
or U30626 (N_30626,N_28450,N_28796);
xnor U30627 (N_30627,N_28428,N_29284);
or U30628 (N_30628,N_28814,N_28755);
and U30629 (N_30629,N_29072,N_28714);
nand U30630 (N_30630,N_28443,N_29011);
nor U30631 (N_30631,N_28370,N_28836);
xnor U30632 (N_30632,N_29471,N_28980);
nand U30633 (N_30633,N_29744,N_29866);
nor U30634 (N_30634,N_29772,N_28421);
nand U30635 (N_30635,N_29406,N_29217);
and U30636 (N_30636,N_28968,N_28043);
nand U30637 (N_30637,N_28408,N_29661);
or U30638 (N_30638,N_29127,N_28435);
and U30639 (N_30639,N_29362,N_28107);
nand U30640 (N_30640,N_29258,N_29870);
or U30641 (N_30641,N_28138,N_28326);
xnor U30642 (N_30642,N_28385,N_28550);
or U30643 (N_30643,N_29643,N_28210);
and U30644 (N_30644,N_28676,N_28478);
and U30645 (N_30645,N_28134,N_28584);
or U30646 (N_30646,N_29988,N_28858);
or U30647 (N_30647,N_28473,N_28426);
or U30648 (N_30648,N_28375,N_28135);
xnor U30649 (N_30649,N_29068,N_28580);
nor U30650 (N_30650,N_28908,N_29787);
nand U30651 (N_30651,N_28255,N_28207);
or U30652 (N_30652,N_28812,N_28730);
nor U30653 (N_30653,N_29180,N_29007);
nor U30654 (N_30654,N_29734,N_29649);
nor U30655 (N_30655,N_29454,N_28788);
and U30656 (N_30656,N_29433,N_28623);
xnor U30657 (N_30657,N_29747,N_28959);
and U30658 (N_30658,N_29518,N_28454);
nor U30659 (N_30659,N_29047,N_28047);
or U30660 (N_30660,N_28952,N_28477);
xnor U30661 (N_30661,N_28997,N_29841);
and U30662 (N_30662,N_29145,N_28948);
nand U30663 (N_30663,N_29503,N_28733);
xnor U30664 (N_30664,N_28232,N_28028);
nor U30665 (N_30665,N_28453,N_28736);
and U30666 (N_30666,N_29512,N_28532);
nand U30667 (N_30667,N_28341,N_29733);
nor U30668 (N_30668,N_28007,N_28219);
or U30669 (N_30669,N_29964,N_28261);
nand U30670 (N_30670,N_29972,N_28401);
nand U30671 (N_30671,N_29683,N_29168);
nand U30672 (N_30672,N_28513,N_29054);
xor U30673 (N_30673,N_29167,N_28239);
or U30674 (N_30674,N_28599,N_29600);
nand U30675 (N_30675,N_28422,N_28051);
xnor U30676 (N_30676,N_29881,N_29494);
and U30677 (N_30677,N_29707,N_29495);
nor U30678 (N_30678,N_29543,N_28104);
or U30679 (N_30679,N_29451,N_28313);
nand U30680 (N_30680,N_29025,N_28775);
nor U30681 (N_30681,N_29452,N_28631);
or U30682 (N_30682,N_28925,N_28660);
or U30683 (N_30683,N_28545,N_29855);
and U30684 (N_30684,N_28954,N_28257);
and U30685 (N_30685,N_29200,N_29790);
nand U30686 (N_30686,N_28424,N_29210);
or U30687 (N_30687,N_28664,N_28321);
nand U30688 (N_30688,N_29278,N_29455);
and U30689 (N_30689,N_28376,N_29063);
nor U30690 (N_30690,N_28987,N_29073);
nor U30691 (N_30691,N_28481,N_29470);
or U30692 (N_30692,N_29931,N_29170);
xnor U30693 (N_30693,N_28411,N_29298);
xor U30694 (N_30694,N_28648,N_28202);
nand U30695 (N_30695,N_28441,N_28003);
xnor U30696 (N_30696,N_29941,N_28139);
nor U30697 (N_30697,N_28366,N_28705);
nand U30698 (N_30698,N_29764,N_29877);
nor U30699 (N_30699,N_28808,N_29586);
or U30700 (N_30700,N_29958,N_28624);
nand U30701 (N_30701,N_29696,N_28494);
and U30702 (N_30702,N_29030,N_28026);
nand U30703 (N_30703,N_28666,N_29246);
nor U30704 (N_30704,N_28499,N_28392);
or U30705 (N_30705,N_28531,N_29018);
xor U30706 (N_30706,N_29652,N_28419);
nor U30707 (N_30707,N_28742,N_29272);
xnor U30708 (N_30708,N_29402,N_28791);
nor U30709 (N_30709,N_29289,N_29513);
or U30710 (N_30710,N_29538,N_29779);
and U30711 (N_30711,N_28826,N_28720);
xnor U30712 (N_30712,N_28634,N_29333);
and U30713 (N_30713,N_29435,N_28960);
nand U30714 (N_30714,N_29659,N_28498);
nor U30715 (N_30715,N_29765,N_28675);
xor U30716 (N_30716,N_28307,N_29530);
or U30717 (N_30717,N_28617,N_29039);
and U30718 (N_30718,N_28291,N_29218);
nand U30719 (N_30719,N_28079,N_28601);
xnor U30720 (N_30720,N_29033,N_28799);
nor U30721 (N_30721,N_28005,N_29342);
nand U30722 (N_30722,N_29445,N_29541);
and U30723 (N_30723,N_29374,N_29373);
and U30724 (N_30724,N_28284,N_28339);
or U30725 (N_30725,N_29178,N_28031);
nor U30726 (N_30726,N_29575,N_29009);
nor U30727 (N_30727,N_28150,N_29132);
xor U30728 (N_30728,N_28738,N_28912);
nor U30729 (N_30729,N_29181,N_29434);
nor U30730 (N_30730,N_28067,N_28444);
or U30731 (N_30731,N_29507,N_29067);
and U30732 (N_30732,N_29194,N_28133);
or U30733 (N_30733,N_29375,N_29524);
xor U30734 (N_30734,N_29965,N_29052);
xor U30735 (N_30735,N_28070,N_29788);
and U30736 (N_30736,N_29680,N_29353);
xor U30737 (N_30737,N_29479,N_28895);
nand U30738 (N_30738,N_29604,N_29254);
or U30739 (N_30739,N_28804,N_28434);
nand U30740 (N_30740,N_29176,N_29383);
xnor U30741 (N_30741,N_29115,N_28593);
nor U30742 (N_30742,N_28083,N_28245);
nor U30743 (N_30743,N_28215,N_28973);
or U30744 (N_30744,N_29450,N_29539);
nor U30745 (N_30745,N_29572,N_28988);
nor U30746 (N_30746,N_28867,N_29291);
nand U30747 (N_30747,N_28046,N_29872);
xnor U30748 (N_30748,N_29337,N_29408);
and U30749 (N_30749,N_28283,N_29468);
and U30750 (N_30750,N_29088,N_29793);
nor U30751 (N_30751,N_28387,N_29015);
xor U30752 (N_30752,N_28602,N_28632);
and U30753 (N_30753,N_28700,N_28152);
or U30754 (N_30754,N_29858,N_29428);
nor U30755 (N_30755,N_28314,N_29209);
or U30756 (N_30756,N_28349,N_28915);
nand U30757 (N_30757,N_28956,N_29483);
nand U30758 (N_30758,N_29628,N_28935);
xor U30759 (N_30759,N_29276,N_28761);
nor U30760 (N_30760,N_29785,N_28727);
or U30761 (N_30761,N_28414,N_29171);
nand U30762 (N_30762,N_29318,N_29754);
nand U30763 (N_30763,N_28568,N_29833);
and U30764 (N_30764,N_29905,N_29667);
nor U30765 (N_30765,N_28615,N_29578);
and U30766 (N_30766,N_28901,N_28217);
and U30767 (N_30767,N_28971,N_28472);
nand U30768 (N_30768,N_28342,N_29245);
nor U30769 (N_30769,N_28140,N_28119);
or U30770 (N_30770,N_28566,N_29028);
xnor U30771 (N_30771,N_28297,N_29742);
and U30772 (N_30772,N_28145,N_29534);
or U30773 (N_30773,N_28251,N_28709);
xor U30774 (N_30774,N_29642,N_29678);
and U30775 (N_30775,N_29748,N_28739);
nand U30776 (N_30776,N_29114,N_29071);
nand U30777 (N_30777,N_29822,N_28100);
nor U30778 (N_30778,N_29487,N_28591);
nor U30779 (N_30779,N_29596,N_29735);
or U30780 (N_30780,N_28290,N_29564);
or U30781 (N_30781,N_28763,N_28115);
xor U30782 (N_30782,N_28732,N_29255);
nand U30783 (N_30783,N_28101,N_28282);
or U30784 (N_30784,N_28750,N_29376);
nand U30785 (N_30785,N_29149,N_29845);
nand U30786 (N_30786,N_29061,N_28042);
nor U30787 (N_30787,N_28746,N_29000);
or U30788 (N_30788,N_29647,N_29646);
xnor U30789 (N_30789,N_28977,N_29952);
or U30790 (N_30790,N_29938,N_28975);
and U30791 (N_30791,N_29379,N_28747);
nor U30792 (N_30792,N_29955,N_28897);
or U30793 (N_30793,N_28549,N_28928);
and U30794 (N_30794,N_28866,N_29689);
nor U30795 (N_30795,N_28404,N_28500);
or U30796 (N_30796,N_29906,N_29301);
xnor U30797 (N_30797,N_28056,N_28903);
or U30798 (N_30798,N_29990,N_29338);
and U30799 (N_30799,N_28184,N_28830);
and U30800 (N_30800,N_29536,N_29559);
xor U30801 (N_30801,N_29688,N_28018);
or U30802 (N_30802,N_28308,N_29515);
nor U30803 (N_30803,N_29806,N_28663);
nor U30804 (N_30804,N_29908,N_29204);
and U30805 (N_30805,N_28380,N_28969);
and U30806 (N_30806,N_29770,N_29903);
or U30807 (N_30807,N_28117,N_29110);
and U30808 (N_30808,N_29313,N_28881);
and U30809 (N_30809,N_28324,N_28906);
nor U30810 (N_30810,N_28834,N_29810);
nor U30811 (N_30811,N_29285,N_29681);
nand U30812 (N_30812,N_28752,N_29352);
nor U30813 (N_30813,N_29771,N_29606);
nor U30814 (N_30814,N_28431,N_28916);
or U30815 (N_30815,N_28111,N_29839);
or U30816 (N_30816,N_28828,N_29741);
nand U30817 (N_30817,N_28635,N_28898);
xnor U30818 (N_30818,N_28892,N_28475);
and U30819 (N_30819,N_28092,N_28544);
nor U30820 (N_30820,N_29721,N_29282);
or U30821 (N_30821,N_28941,N_29045);
and U30822 (N_30822,N_29610,N_28073);
or U30823 (N_30823,N_28835,N_28124);
and U30824 (N_30824,N_28027,N_29608);
nor U30825 (N_30825,N_29581,N_28200);
or U30826 (N_30826,N_29946,N_28986);
or U30827 (N_30827,N_28418,N_29496);
xnor U30828 (N_30828,N_28193,N_29064);
xor U30829 (N_30829,N_28596,N_29640);
nand U30830 (N_30830,N_28149,N_28760);
nand U30831 (N_30831,N_29709,N_29720);
and U30832 (N_30832,N_28511,N_29056);
nand U30833 (N_30833,N_28611,N_28009);
nor U30834 (N_30834,N_29107,N_29542);
or U30835 (N_30835,N_29821,N_29003);
nor U30836 (N_30836,N_29252,N_28562);
nand U30837 (N_30837,N_29014,N_28861);
nand U30838 (N_30838,N_29177,N_28572);
or U30839 (N_30839,N_29134,N_28530);
xnor U30840 (N_30840,N_29655,N_29320);
or U30841 (N_30841,N_29934,N_29172);
nand U30842 (N_30842,N_28604,N_29244);
nand U30843 (N_30843,N_29164,N_29824);
nand U30844 (N_30844,N_28699,N_29506);
xnor U30845 (N_30845,N_29432,N_29409);
or U30846 (N_30846,N_29274,N_29594);
xnor U30847 (N_30847,N_29654,N_29550);
nor U30848 (N_30848,N_29086,N_28013);
or U30849 (N_30849,N_28902,N_28493);
and U30850 (N_30850,N_29261,N_29311);
nand U30851 (N_30851,N_29008,N_29545);
nor U30852 (N_30852,N_29814,N_29959);
and U30853 (N_30853,N_29713,N_29891);
or U30854 (N_30854,N_29268,N_29059);
nand U30855 (N_30855,N_29104,N_29953);
and U30856 (N_30856,N_28094,N_28476);
nor U30857 (N_30857,N_29570,N_28937);
nand U30858 (N_30858,N_29928,N_29213);
nand U30859 (N_30859,N_28557,N_29523);
and U30860 (N_30860,N_29593,N_29852);
nor U30861 (N_30861,N_29464,N_29371);
nand U30862 (N_30862,N_29792,N_29193);
nand U30863 (N_30863,N_29585,N_28894);
nor U30864 (N_30864,N_29460,N_29591);
xnor U30865 (N_30865,N_29489,N_28123);
xor U30866 (N_30866,N_29238,N_28569);
nor U30867 (N_30867,N_28090,N_29377);
xnor U30868 (N_30868,N_29929,N_28126);
or U30869 (N_30869,N_29695,N_28296);
or U30870 (N_30870,N_29146,N_28506);
nand U30871 (N_30871,N_28240,N_28645);
nor U30872 (N_30872,N_29950,N_29328);
nor U30873 (N_30873,N_29504,N_29312);
or U30874 (N_30874,N_29812,N_29330);
or U30875 (N_30875,N_29119,N_29727);
nor U30876 (N_30876,N_28335,N_28359);
nor U30877 (N_30877,N_29081,N_28972);
or U30878 (N_30878,N_29761,N_28082);
nor U30879 (N_30879,N_29561,N_28024);
nor U30880 (N_30880,N_28260,N_28583);
or U30881 (N_30881,N_29049,N_29349);
xor U30882 (N_30882,N_28468,N_29611);
or U30883 (N_30883,N_28457,N_29766);
and U30884 (N_30884,N_28692,N_28459);
nor U30885 (N_30885,N_28383,N_28166);
xor U30886 (N_30886,N_28248,N_29876);
and U30887 (N_30887,N_28180,N_28657);
nand U30888 (N_30888,N_29174,N_29969);
nor U30889 (N_30889,N_28025,N_29844);
xnor U30890 (N_30890,N_28109,N_29693);
xnor U30891 (N_30891,N_29326,N_28547);
xnor U30892 (N_30892,N_29101,N_29978);
nor U30893 (N_30893,N_29875,N_29102);
xnor U30894 (N_30894,N_29994,N_29942);
nor U30895 (N_30895,N_28650,N_28311);
xor U30896 (N_30896,N_29781,N_29150);
nand U30897 (N_30897,N_29123,N_28756);
nand U30898 (N_30898,N_28438,N_29970);
and U30899 (N_30899,N_29113,N_28030);
nor U30900 (N_30900,N_28777,N_28371);
and U30901 (N_30901,N_29884,N_29500);
xnor U30902 (N_30902,N_28585,N_29414);
nand U30903 (N_30903,N_29520,N_29089);
nor U30904 (N_30904,N_29380,N_29100);
nand U30905 (N_30905,N_29265,N_28702);
or U30906 (N_30906,N_28798,N_28630);
xor U30907 (N_30907,N_28943,N_28931);
nor U30908 (N_30908,N_29022,N_28774);
nand U30909 (N_30909,N_29280,N_29660);
nand U30910 (N_30910,N_28206,N_28685);
or U30911 (N_30911,N_28879,N_29413);
or U30912 (N_30912,N_28991,N_29672);
or U30913 (N_30913,N_29439,N_28770);
and U30914 (N_30914,N_29363,N_28582);
or U30915 (N_30915,N_29264,N_28961);
nor U30916 (N_30916,N_28672,N_29415);
xor U30917 (N_30917,N_28989,N_28347);
xor U30918 (N_30918,N_29579,N_28521);
xnor U30919 (N_30919,N_29615,N_29599);
nand U30920 (N_30920,N_28158,N_29124);
nand U30921 (N_30921,N_28848,N_29573);
or U30922 (N_30922,N_28589,N_28778);
nand U30923 (N_30923,N_29555,N_29871);
nor U30924 (N_30924,N_29354,N_29746);
or U30925 (N_30925,N_28222,N_29921);
and U30926 (N_30926,N_29221,N_28496);
or U30927 (N_30927,N_28393,N_29664);
xnor U30928 (N_30928,N_28886,N_28945);
and U30929 (N_30929,N_28316,N_28226);
nand U30930 (N_30930,N_28823,N_29120);
and U30931 (N_30931,N_28220,N_29188);
xnor U30932 (N_30932,N_28221,N_29456);
or U30933 (N_30933,N_29731,N_28402);
or U30934 (N_30934,N_28529,N_29690);
xor U30935 (N_30935,N_29521,N_29775);
and U30936 (N_30936,N_28388,N_28412);
and U30937 (N_30937,N_28992,N_28536);
xor U30938 (N_30938,N_28563,N_28053);
nor U30939 (N_30939,N_29300,N_28143);
or U30940 (N_30940,N_29577,N_28461);
and U30941 (N_30941,N_29162,N_29492);
or U30942 (N_30942,N_28249,N_29042);
and U30943 (N_30943,N_28071,N_28384);
and U30944 (N_30944,N_29923,N_29035);
nor U30945 (N_30945,N_29710,N_29826);
xnor U30946 (N_30946,N_29662,N_28684);
or U30947 (N_30947,N_29085,N_29079);
or U30948 (N_30948,N_28243,N_28266);
nand U30949 (N_30949,N_28292,N_29926);
nand U30950 (N_30950,N_28427,N_28131);
nor U30951 (N_30951,N_29558,N_28737);
xnor U30952 (N_30952,N_28423,N_28680);
nor U30953 (N_30953,N_28896,N_28689);
nor U30954 (N_30954,N_29911,N_28096);
or U30955 (N_30955,N_28395,N_28656);
nor U30956 (N_30956,N_28618,N_29750);
nand U30957 (N_30957,N_29987,N_29491);
nor U30958 (N_30958,N_29126,N_29525);
nand U30959 (N_30959,N_29183,N_28128);
and U30960 (N_30960,N_29005,N_28279);
xor U30961 (N_30961,N_28889,N_28440);
or U30962 (N_30962,N_28141,N_29616);
nor U30963 (N_30963,N_29046,N_28237);
xor U30964 (N_30964,N_28982,N_29315);
and U30965 (N_30965,N_29029,N_29277);
and U30966 (N_30966,N_29344,N_28033);
and U30967 (N_30967,N_28806,N_29673);
nand U30968 (N_30968,N_29805,N_28164);
or U30969 (N_30969,N_28877,N_28465);
or U30970 (N_30970,N_29986,N_28647);
xnor U30971 (N_30971,N_28186,N_28467);
xor U30972 (N_30972,N_28628,N_28551);
or U30973 (N_30973,N_29856,N_29248);
nand U30974 (N_30974,N_28293,N_28810);
and U30975 (N_30975,N_28087,N_29062);
xnor U30976 (N_30976,N_28102,N_29361);
or U30977 (N_30977,N_28641,N_28662);
nand U30978 (N_30978,N_29691,N_29446);
nand U30979 (N_30979,N_28502,N_28369);
nand U30980 (N_30980,N_28590,N_28398);
nor U30981 (N_30981,N_28010,N_28276);
and U30982 (N_30982,N_28668,N_29778);
nor U30983 (N_30983,N_29198,N_28922);
or U30984 (N_30984,N_29016,N_29230);
xnor U30985 (N_30985,N_28724,N_28032);
and U30986 (N_30986,N_29900,N_28661);
nand U30987 (N_30987,N_28577,N_28614);
nor U30988 (N_30988,N_29816,N_29873);
nand U30989 (N_30989,N_29686,N_28731);
and U30990 (N_30990,N_28396,N_29116);
and U30991 (N_30991,N_29574,N_29977);
xnor U30992 (N_30992,N_28091,N_28978);
nand U30993 (N_30993,N_28512,N_29092);
or U30994 (N_30994,N_28216,N_28406);
nand U30995 (N_30995,N_28085,N_28490);
nand U30996 (N_30996,N_29024,N_29166);
nand U30997 (N_30997,N_29847,N_28045);
and U30998 (N_30998,N_29618,N_28301);
nand U30999 (N_30999,N_29736,N_28766);
xor U31000 (N_31000,N_28069,N_29168);
xnor U31001 (N_31001,N_29770,N_28857);
nor U31002 (N_31002,N_28216,N_28232);
xor U31003 (N_31003,N_28008,N_29680);
and U31004 (N_31004,N_28759,N_28731);
nor U31005 (N_31005,N_28678,N_29250);
xnor U31006 (N_31006,N_28593,N_28583);
and U31007 (N_31007,N_29822,N_28431);
nor U31008 (N_31008,N_29774,N_28593);
nand U31009 (N_31009,N_29168,N_29345);
and U31010 (N_31010,N_28385,N_29570);
nor U31011 (N_31011,N_28354,N_29975);
nor U31012 (N_31012,N_28153,N_28005);
nor U31013 (N_31013,N_28721,N_29145);
or U31014 (N_31014,N_29318,N_28427);
or U31015 (N_31015,N_28009,N_28002);
nand U31016 (N_31016,N_28599,N_28578);
xor U31017 (N_31017,N_29789,N_29036);
and U31018 (N_31018,N_29297,N_29006);
or U31019 (N_31019,N_28450,N_28010);
xor U31020 (N_31020,N_28832,N_28884);
nand U31021 (N_31021,N_28858,N_29291);
nor U31022 (N_31022,N_29442,N_28079);
nor U31023 (N_31023,N_29042,N_29490);
xor U31024 (N_31024,N_29319,N_29763);
or U31025 (N_31025,N_28525,N_28087);
nor U31026 (N_31026,N_28614,N_28313);
nand U31027 (N_31027,N_29444,N_28714);
xor U31028 (N_31028,N_28992,N_29432);
or U31029 (N_31029,N_28919,N_28695);
nor U31030 (N_31030,N_28193,N_28151);
xor U31031 (N_31031,N_29558,N_29565);
nor U31032 (N_31032,N_28078,N_28909);
nand U31033 (N_31033,N_28616,N_28334);
and U31034 (N_31034,N_29343,N_28806);
or U31035 (N_31035,N_29813,N_29256);
xnor U31036 (N_31036,N_29889,N_28443);
xnor U31037 (N_31037,N_28155,N_29284);
and U31038 (N_31038,N_29994,N_29375);
nor U31039 (N_31039,N_28653,N_28976);
xnor U31040 (N_31040,N_29674,N_28552);
xor U31041 (N_31041,N_29906,N_29953);
nand U31042 (N_31042,N_28364,N_28372);
xor U31043 (N_31043,N_28112,N_29208);
or U31044 (N_31044,N_29243,N_28620);
nor U31045 (N_31045,N_29364,N_29348);
nor U31046 (N_31046,N_28171,N_29690);
nand U31047 (N_31047,N_29025,N_29416);
nor U31048 (N_31048,N_29232,N_28688);
nand U31049 (N_31049,N_29624,N_28756);
nand U31050 (N_31050,N_29374,N_29045);
or U31051 (N_31051,N_28993,N_28826);
nand U31052 (N_31052,N_29472,N_28822);
and U31053 (N_31053,N_28515,N_28120);
nor U31054 (N_31054,N_28086,N_29985);
xor U31055 (N_31055,N_28849,N_29757);
nand U31056 (N_31056,N_29963,N_28888);
or U31057 (N_31057,N_29992,N_28652);
nor U31058 (N_31058,N_29441,N_29623);
nor U31059 (N_31059,N_29725,N_29154);
xor U31060 (N_31060,N_29245,N_29899);
nor U31061 (N_31061,N_28989,N_28706);
nor U31062 (N_31062,N_29112,N_28911);
and U31063 (N_31063,N_28247,N_28762);
and U31064 (N_31064,N_28041,N_28357);
xnor U31065 (N_31065,N_29782,N_29082);
or U31066 (N_31066,N_28449,N_29251);
xor U31067 (N_31067,N_28631,N_28177);
nor U31068 (N_31068,N_29619,N_29013);
xnor U31069 (N_31069,N_29172,N_28382);
nand U31070 (N_31070,N_28285,N_29529);
and U31071 (N_31071,N_29997,N_29341);
and U31072 (N_31072,N_29750,N_28739);
nor U31073 (N_31073,N_29757,N_28931);
or U31074 (N_31074,N_28072,N_29789);
or U31075 (N_31075,N_29120,N_28361);
xor U31076 (N_31076,N_28029,N_28255);
and U31077 (N_31077,N_29676,N_29773);
or U31078 (N_31078,N_29087,N_29702);
nor U31079 (N_31079,N_29334,N_28112);
nand U31080 (N_31080,N_29829,N_29460);
nor U31081 (N_31081,N_29161,N_28707);
xor U31082 (N_31082,N_29092,N_29393);
xnor U31083 (N_31083,N_29666,N_28668);
or U31084 (N_31084,N_29472,N_29963);
xor U31085 (N_31085,N_29213,N_29132);
nor U31086 (N_31086,N_28080,N_29258);
nand U31087 (N_31087,N_29607,N_29253);
nor U31088 (N_31088,N_28986,N_29879);
or U31089 (N_31089,N_29072,N_28778);
and U31090 (N_31090,N_28481,N_29692);
or U31091 (N_31091,N_28108,N_28939);
xor U31092 (N_31092,N_28071,N_29661);
or U31093 (N_31093,N_29438,N_29856);
and U31094 (N_31094,N_29668,N_29698);
and U31095 (N_31095,N_29604,N_29119);
nand U31096 (N_31096,N_28340,N_29650);
and U31097 (N_31097,N_29082,N_29747);
nor U31098 (N_31098,N_28707,N_28283);
or U31099 (N_31099,N_28221,N_29270);
nor U31100 (N_31100,N_29819,N_28531);
and U31101 (N_31101,N_29638,N_29417);
nor U31102 (N_31102,N_29848,N_28039);
or U31103 (N_31103,N_29235,N_28269);
nor U31104 (N_31104,N_29192,N_28253);
xnor U31105 (N_31105,N_29116,N_28875);
nor U31106 (N_31106,N_29990,N_28986);
nand U31107 (N_31107,N_29743,N_29299);
nor U31108 (N_31108,N_28690,N_29537);
or U31109 (N_31109,N_28028,N_29944);
or U31110 (N_31110,N_29532,N_28738);
nand U31111 (N_31111,N_29598,N_29041);
nand U31112 (N_31112,N_29692,N_28899);
nand U31113 (N_31113,N_29114,N_28863);
xor U31114 (N_31114,N_28963,N_29959);
xnor U31115 (N_31115,N_29344,N_29854);
xnor U31116 (N_31116,N_29538,N_28844);
and U31117 (N_31117,N_28469,N_29159);
xor U31118 (N_31118,N_28781,N_29025);
nand U31119 (N_31119,N_29157,N_29295);
or U31120 (N_31120,N_29274,N_29995);
xor U31121 (N_31121,N_29131,N_28565);
or U31122 (N_31122,N_28609,N_28404);
or U31123 (N_31123,N_28999,N_29017);
xnor U31124 (N_31124,N_28811,N_28662);
xor U31125 (N_31125,N_29558,N_28386);
or U31126 (N_31126,N_29598,N_28302);
xor U31127 (N_31127,N_28672,N_29866);
nand U31128 (N_31128,N_29799,N_28858);
or U31129 (N_31129,N_28085,N_28022);
nor U31130 (N_31130,N_29852,N_29371);
nor U31131 (N_31131,N_29260,N_29419);
nand U31132 (N_31132,N_29131,N_29539);
xnor U31133 (N_31133,N_28359,N_28237);
nand U31134 (N_31134,N_29425,N_28308);
xor U31135 (N_31135,N_29893,N_29506);
xor U31136 (N_31136,N_28421,N_28471);
and U31137 (N_31137,N_29856,N_28559);
xnor U31138 (N_31138,N_29082,N_29514);
or U31139 (N_31139,N_28473,N_29494);
nand U31140 (N_31140,N_29044,N_29379);
and U31141 (N_31141,N_29374,N_29249);
and U31142 (N_31142,N_29579,N_29853);
nand U31143 (N_31143,N_29469,N_28985);
and U31144 (N_31144,N_29909,N_28384);
or U31145 (N_31145,N_29575,N_28884);
and U31146 (N_31146,N_29714,N_28015);
xnor U31147 (N_31147,N_28906,N_28384);
xor U31148 (N_31148,N_29863,N_28237);
nand U31149 (N_31149,N_28209,N_28164);
nand U31150 (N_31150,N_28222,N_28449);
and U31151 (N_31151,N_28793,N_29323);
nor U31152 (N_31152,N_29655,N_29838);
nor U31153 (N_31153,N_28805,N_29264);
or U31154 (N_31154,N_29180,N_28601);
or U31155 (N_31155,N_29595,N_29868);
nand U31156 (N_31156,N_28659,N_29363);
nand U31157 (N_31157,N_29052,N_28166);
or U31158 (N_31158,N_29171,N_29932);
or U31159 (N_31159,N_29229,N_29748);
nand U31160 (N_31160,N_29755,N_29173);
and U31161 (N_31161,N_29810,N_28926);
nor U31162 (N_31162,N_29398,N_29149);
nand U31163 (N_31163,N_28843,N_28980);
and U31164 (N_31164,N_28145,N_28217);
nand U31165 (N_31165,N_29959,N_28531);
nor U31166 (N_31166,N_29148,N_28372);
or U31167 (N_31167,N_29661,N_29164);
nor U31168 (N_31168,N_29116,N_29409);
nor U31169 (N_31169,N_29868,N_29847);
or U31170 (N_31170,N_29307,N_28746);
nor U31171 (N_31171,N_28782,N_28366);
and U31172 (N_31172,N_29967,N_28997);
nand U31173 (N_31173,N_28315,N_29977);
nor U31174 (N_31174,N_28279,N_28730);
nor U31175 (N_31175,N_29924,N_28968);
xor U31176 (N_31176,N_29569,N_28585);
or U31177 (N_31177,N_28522,N_28471);
or U31178 (N_31178,N_28704,N_29490);
nor U31179 (N_31179,N_29080,N_29965);
or U31180 (N_31180,N_28540,N_29336);
nor U31181 (N_31181,N_29828,N_28680);
nor U31182 (N_31182,N_29286,N_28716);
or U31183 (N_31183,N_28508,N_29382);
xor U31184 (N_31184,N_28027,N_28997);
nor U31185 (N_31185,N_28842,N_28168);
and U31186 (N_31186,N_28370,N_29552);
and U31187 (N_31187,N_29758,N_29610);
nor U31188 (N_31188,N_29424,N_28952);
xnor U31189 (N_31189,N_29391,N_28471);
xor U31190 (N_31190,N_28458,N_29455);
nor U31191 (N_31191,N_28383,N_29535);
and U31192 (N_31192,N_28454,N_29911);
or U31193 (N_31193,N_29290,N_29648);
nor U31194 (N_31194,N_28884,N_28550);
nor U31195 (N_31195,N_29535,N_28563);
nor U31196 (N_31196,N_28682,N_28946);
and U31197 (N_31197,N_29081,N_29999);
xor U31198 (N_31198,N_29944,N_28823);
nor U31199 (N_31199,N_28069,N_29720);
xor U31200 (N_31200,N_29786,N_29973);
or U31201 (N_31201,N_29597,N_28778);
nand U31202 (N_31202,N_28405,N_28594);
nor U31203 (N_31203,N_28945,N_29116);
and U31204 (N_31204,N_29787,N_28450);
xor U31205 (N_31205,N_29387,N_29812);
or U31206 (N_31206,N_29828,N_28109);
nand U31207 (N_31207,N_29949,N_28209);
nor U31208 (N_31208,N_28064,N_29366);
nand U31209 (N_31209,N_29488,N_29583);
nand U31210 (N_31210,N_29275,N_29848);
xnor U31211 (N_31211,N_28249,N_28973);
and U31212 (N_31212,N_28537,N_28736);
nor U31213 (N_31213,N_29153,N_28578);
nand U31214 (N_31214,N_28839,N_28580);
and U31215 (N_31215,N_29828,N_29898);
and U31216 (N_31216,N_28359,N_29780);
nand U31217 (N_31217,N_29247,N_29557);
xnor U31218 (N_31218,N_28463,N_29045);
xor U31219 (N_31219,N_29182,N_28138);
xor U31220 (N_31220,N_28087,N_29424);
nor U31221 (N_31221,N_29757,N_29594);
and U31222 (N_31222,N_28345,N_28386);
nor U31223 (N_31223,N_28560,N_28583);
nand U31224 (N_31224,N_29518,N_28230);
and U31225 (N_31225,N_29962,N_28808);
or U31226 (N_31226,N_28409,N_28208);
xor U31227 (N_31227,N_29596,N_29604);
nor U31228 (N_31228,N_28132,N_28758);
nor U31229 (N_31229,N_29141,N_29872);
xor U31230 (N_31230,N_28321,N_28180);
nand U31231 (N_31231,N_29718,N_29276);
nor U31232 (N_31232,N_29255,N_28129);
nand U31233 (N_31233,N_28796,N_28859);
nor U31234 (N_31234,N_28658,N_28970);
nor U31235 (N_31235,N_29570,N_28471);
xnor U31236 (N_31236,N_29881,N_29246);
xnor U31237 (N_31237,N_28169,N_28179);
xor U31238 (N_31238,N_28995,N_28176);
and U31239 (N_31239,N_28980,N_28587);
and U31240 (N_31240,N_28312,N_28594);
nand U31241 (N_31241,N_29098,N_28835);
xnor U31242 (N_31242,N_28396,N_28306);
xnor U31243 (N_31243,N_28936,N_28536);
and U31244 (N_31244,N_29603,N_28011);
nand U31245 (N_31245,N_29623,N_29956);
xnor U31246 (N_31246,N_29807,N_28888);
xnor U31247 (N_31247,N_28684,N_28189);
nor U31248 (N_31248,N_28666,N_28895);
nand U31249 (N_31249,N_29450,N_28954);
or U31250 (N_31250,N_29654,N_29818);
or U31251 (N_31251,N_29525,N_29992);
nor U31252 (N_31252,N_29364,N_28094);
nand U31253 (N_31253,N_29153,N_29444);
or U31254 (N_31254,N_28895,N_29775);
and U31255 (N_31255,N_28256,N_28440);
nand U31256 (N_31256,N_28223,N_28669);
nand U31257 (N_31257,N_28954,N_28510);
or U31258 (N_31258,N_29276,N_28201);
and U31259 (N_31259,N_28445,N_28361);
xnor U31260 (N_31260,N_28104,N_28319);
or U31261 (N_31261,N_28744,N_28458);
nand U31262 (N_31262,N_29896,N_28264);
xor U31263 (N_31263,N_28806,N_28695);
and U31264 (N_31264,N_29121,N_29359);
nor U31265 (N_31265,N_28675,N_29586);
or U31266 (N_31266,N_29723,N_28272);
and U31267 (N_31267,N_28430,N_29991);
nor U31268 (N_31268,N_28422,N_29426);
and U31269 (N_31269,N_29929,N_29847);
nand U31270 (N_31270,N_29808,N_28685);
or U31271 (N_31271,N_28883,N_28526);
nor U31272 (N_31272,N_29975,N_28248);
xor U31273 (N_31273,N_28467,N_29900);
nor U31274 (N_31274,N_28456,N_29825);
nand U31275 (N_31275,N_28089,N_28323);
and U31276 (N_31276,N_28966,N_29148);
nor U31277 (N_31277,N_28193,N_28307);
nor U31278 (N_31278,N_29686,N_28078);
xnor U31279 (N_31279,N_29618,N_28332);
or U31280 (N_31280,N_28217,N_28048);
and U31281 (N_31281,N_29331,N_28317);
or U31282 (N_31282,N_28438,N_28401);
and U31283 (N_31283,N_28218,N_29269);
and U31284 (N_31284,N_28991,N_29711);
nand U31285 (N_31285,N_29133,N_29934);
xor U31286 (N_31286,N_29417,N_28922);
nor U31287 (N_31287,N_29897,N_29861);
or U31288 (N_31288,N_28117,N_28724);
nor U31289 (N_31289,N_28428,N_29716);
nand U31290 (N_31290,N_28888,N_28498);
xor U31291 (N_31291,N_28948,N_28309);
or U31292 (N_31292,N_28827,N_29272);
xor U31293 (N_31293,N_29131,N_29579);
and U31294 (N_31294,N_28609,N_29317);
and U31295 (N_31295,N_28882,N_29705);
or U31296 (N_31296,N_29948,N_28322);
nand U31297 (N_31297,N_29811,N_29555);
and U31298 (N_31298,N_28561,N_28430);
nand U31299 (N_31299,N_29656,N_28122);
nor U31300 (N_31300,N_29231,N_28794);
xnor U31301 (N_31301,N_29711,N_28474);
xnor U31302 (N_31302,N_28568,N_28958);
and U31303 (N_31303,N_28737,N_28068);
or U31304 (N_31304,N_29941,N_29069);
nor U31305 (N_31305,N_28224,N_29812);
nand U31306 (N_31306,N_29450,N_28812);
nand U31307 (N_31307,N_29567,N_29025);
xor U31308 (N_31308,N_28001,N_29498);
xnor U31309 (N_31309,N_29534,N_29216);
nand U31310 (N_31310,N_28692,N_29149);
or U31311 (N_31311,N_29912,N_28972);
xor U31312 (N_31312,N_28794,N_28606);
or U31313 (N_31313,N_29523,N_29925);
nor U31314 (N_31314,N_28981,N_28872);
nand U31315 (N_31315,N_29112,N_28518);
and U31316 (N_31316,N_29749,N_28975);
or U31317 (N_31317,N_28393,N_28378);
xnor U31318 (N_31318,N_28213,N_28046);
xor U31319 (N_31319,N_28496,N_29628);
and U31320 (N_31320,N_29990,N_28780);
nor U31321 (N_31321,N_28969,N_29314);
and U31322 (N_31322,N_29777,N_28977);
nand U31323 (N_31323,N_28008,N_29138);
or U31324 (N_31324,N_29332,N_29551);
nor U31325 (N_31325,N_29945,N_29332);
nor U31326 (N_31326,N_28340,N_29095);
nand U31327 (N_31327,N_28137,N_28371);
or U31328 (N_31328,N_29147,N_29465);
and U31329 (N_31329,N_28978,N_29826);
xnor U31330 (N_31330,N_28280,N_28176);
or U31331 (N_31331,N_29910,N_28016);
nor U31332 (N_31332,N_28449,N_28358);
xnor U31333 (N_31333,N_28631,N_28889);
nand U31334 (N_31334,N_29471,N_28072);
or U31335 (N_31335,N_28638,N_29577);
nand U31336 (N_31336,N_29284,N_28578);
nor U31337 (N_31337,N_28444,N_29867);
or U31338 (N_31338,N_28416,N_28911);
or U31339 (N_31339,N_28385,N_29777);
nor U31340 (N_31340,N_29988,N_28531);
and U31341 (N_31341,N_28579,N_28245);
or U31342 (N_31342,N_29241,N_29418);
nor U31343 (N_31343,N_28451,N_29610);
nand U31344 (N_31344,N_29200,N_28826);
nor U31345 (N_31345,N_29838,N_29042);
or U31346 (N_31346,N_29683,N_28905);
and U31347 (N_31347,N_29930,N_28242);
nor U31348 (N_31348,N_29129,N_28028);
and U31349 (N_31349,N_28255,N_28200);
and U31350 (N_31350,N_28606,N_28674);
nand U31351 (N_31351,N_29899,N_28303);
and U31352 (N_31352,N_29755,N_29622);
or U31353 (N_31353,N_29502,N_28422);
nor U31354 (N_31354,N_28142,N_28300);
and U31355 (N_31355,N_29447,N_29977);
nor U31356 (N_31356,N_28170,N_29233);
xnor U31357 (N_31357,N_28060,N_28810);
nor U31358 (N_31358,N_29521,N_28005);
nand U31359 (N_31359,N_29210,N_28824);
nand U31360 (N_31360,N_29101,N_29259);
and U31361 (N_31361,N_29318,N_29889);
and U31362 (N_31362,N_28065,N_29074);
nor U31363 (N_31363,N_28389,N_29948);
or U31364 (N_31364,N_28567,N_29992);
xnor U31365 (N_31365,N_29352,N_28861);
and U31366 (N_31366,N_29756,N_29716);
nand U31367 (N_31367,N_29180,N_28855);
nand U31368 (N_31368,N_29695,N_28819);
nor U31369 (N_31369,N_28909,N_28686);
nand U31370 (N_31370,N_28882,N_28184);
nand U31371 (N_31371,N_29861,N_28656);
nand U31372 (N_31372,N_28667,N_28782);
xor U31373 (N_31373,N_29008,N_29795);
nand U31374 (N_31374,N_28921,N_29766);
nand U31375 (N_31375,N_29823,N_28131);
nor U31376 (N_31376,N_29888,N_28845);
nand U31377 (N_31377,N_28889,N_28399);
xnor U31378 (N_31378,N_29219,N_29082);
or U31379 (N_31379,N_28629,N_29426);
and U31380 (N_31380,N_29228,N_28129);
nand U31381 (N_31381,N_29087,N_28709);
xnor U31382 (N_31382,N_29853,N_28991);
and U31383 (N_31383,N_28563,N_29635);
and U31384 (N_31384,N_29736,N_28082);
xnor U31385 (N_31385,N_29912,N_29252);
nor U31386 (N_31386,N_29175,N_28639);
xor U31387 (N_31387,N_28394,N_29292);
xor U31388 (N_31388,N_29401,N_28267);
nand U31389 (N_31389,N_29417,N_29835);
nor U31390 (N_31390,N_29816,N_28044);
nand U31391 (N_31391,N_29618,N_28850);
and U31392 (N_31392,N_28396,N_29045);
nand U31393 (N_31393,N_28959,N_28468);
xor U31394 (N_31394,N_29663,N_28296);
nor U31395 (N_31395,N_28825,N_28995);
nor U31396 (N_31396,N_29985,N_28593);
xor U31397 (N_31397,N_28327,N_29960);
or U31398 (N_31398,N_29860,N_28982);
nand U31399 (N_31399,N_28534,N_28586);
or U31400 (N_31400,N_28428,N_29002);
nor U31401 (N_31401,N_28099,N_28840);
or U31402 (N_31402,N_29216,N_29413);
nand U31403 (N_31403,N_29335,N_29476);
and U31404 (N_31404,N_29745,N_29332);
nor U31405 (N_31405,N_29336,N_29050);
nand U31406 (N_31406,N_28839,N_29607);
or U31407 (N_31407,N_28053,N_28963);
nand U31408 (N_31408,N_28403,N_29399);
and U31409 (N_31409,N_28897,N_28153);
xor U31410 (N_31410,N_29548,N_29411);
and U31411 (N_31411,N_28348,N_29972);
nor U31412 (N_31412,N_28260,N_29951);
and U31413 (N_31413,N_28251,N_28961);
nor U31414 (N_31414,N_29689,N_29302);
xnor U31415 (N_31415,N_28497,N_29445);
and U31416 (N_31416,N_29979,N_29080);
nor U31417 (N_31417,N_29306,N_28142);
nor U31418 (N_31418,N_29049,N_28028);
xnor U31419 (N_31419,N_29987,N_28188);
or U31420 (N_31420,N_28051,N_28257);
or U31421 (N_31421,N_28175,N_29072);
nand U31422 (N_31422,N_28958,N_29664);
nand U31423 (N_31423,N_29071,N_29283);
or U31424 (N_31424,N_29446,N_29612);
or U31425 (N_31425,N_28686,N_28816);
nand U31426 (N_31426,N_28248,N_29789);
nand U31427 (N_31427,N_29549,N_29849);
nor U31428 (N_31428,N_29450,N_28213);
xnor U31429 (N_31429,N_28739,N_29610);
and U31430 (N_31430,N_28115,N_29049);
and U31431 (N_31431,N_28808,N_29883);
or U31432 (N_31432,N_29417,N_28411);
nor U31433 (N_31433,N_29393,N_28863);
xnor U31434 (N_31434,N_28431,N_28451);
nor U31435 (N_31435,N_28606,N_28642);
nor U31436 (N_31436,N_28637,N_29733);
and U31437 (N_31437,N_28893,N_28730);
and U31438 (N_31438,N_29746,N_29691);
and U31439 (N_31439,N_28195,N_29257);
nor U31440 (N_31440,N_28166,N_29034);
xor U31441 (N_31441,N_28011,N_28741);
nor U31442 (N_31442,N_28178,N_28126);
nand U31443 (N_31443,N_28009,N_29966);
nor U31444 (N_31444,N_28249,N_28047);
nor U31445 (N_31445,N_28280,N_29240);
nand U31446 (N_31446,N_28215,N_29850);
xnor U31447 (N_31447,N_28250,N_29777);
nor U31448 (N_31448,N_29711,N_28322);
nor U31449 (N_31449,N_29023,N_28198);
and U31450 (N_31450,N_28021,N_29865);
xor U31451 (N_31451,N_28399,N_29049);
xnor U31452 (N_31452,N_29048,N_29069);
nand U31453 (N_31453,N_29546,N_29380);
or U31454 (N_31454,N_28494,N_28282);
nor U31455 (N_31455,N_28573,N_28344);
or U31456 (N_31456,N_29351,N_29257);
and U31457 (N_31457,N_29340,N_29598);
nand U31458 (N_31458,N_28339,N_29642);
nand U31459 (N_31459,N_28430,N_29194);
and U31460 (N_31460,N_28368,N_28048);
or U31461 (N_31461,N_28361,N_28487);
and U31462 (N_31462,N_29645,N_28698);
and U31463 (N_31463,N_28847,N_28778);
or U31464 (N_31464,N_29461,N_28873);
xor U31465 (N_31465,N_28641,N_29598);
or U31466 (N_31466,N_29873,N_29292);
nor U31467 (N_31467,N_29271,N_28965);
xor U31468 (N_31468,N_29758,N_29911);
xor U31469 (N_31469,N_28770,N_28466);
nor U31470 (N_31470,N_29055,N_28774);
and U31471 (N_31471,N_29126,N_28799);
nand U31472 (N_31472,N_28675,N_28877);
and U31473 (N_31473,N_29540,N_28672);
nand U31474 (N_31474,N_28179,N_29231);
nor U31475 (N_31475,N_29380,N_29932);
nor U31476 (N_31476,N_28983,N_28802);
and U31477 (N_31477,N_28314,N_28986);
nand U31478 (N_31478,N_28531,N_28046);
nor U31479 (N_31479,N_28748,N_29626);
nand U31480 (N_31480,N_28517,N_29707);
or U31481 (N_31481,N_29638,N_28528);
xor U31482 (N_31482,N_29562,N_29479);
xor U31483 (N_31483,N_29651,N_28925);
nand U31484 (N_31484,N_28631,N_28112);
and U31485 (N_31485,N_28076,N_29264);
nor U31486 (N_31486,N_28669,N_29995);
and U31487 (N_31487,N_29286,N_28223);
nor U31488 (N_31488,N_29660,N_28549);
xnor U31489 (N_31489,N_29089,N_29461);
or U31490 (N_31490,N_29763,N_28750);
nand U31491 (N_31491,N_28014,N_29965);
nor U31492 (N_31492,N_29354,N_28433);
or U31493 (N_31493,N_29316,N_28645);
or U31494 (N_31494,N_29848,N_28001);
or U31495 (N_31495,N_29521,N_29271);
or U31496 (N_31496,N_28820,N_29542);
and U31497 (N_31497,N_29961,N_28717);
xnor U31498 (N_31498,N_28795,N_28389);
nand U31499 (N_31499,N_28386,N_28806);
or U31500 (N_31500,N_29765,N_29688);
nand U31501 (N_31501,N_28049,N_29238);
nor U31502 (N_31502,N_28791,N_29702);
or U31503 (N_31503,N_28701,N_29588);
nor U31504 (N_31504,N_28549,N_29786);
nand U31505 (N_31505,N_29078,N_28198);
nand U31506 (N_31506,N_29442,N_28404);
and U31507 (N_31507,N_29254,N_28498);
nand U31508 (N_31508,N_28925,N_29824);
and U31509 (N_31509,N_29003,N_29016);
and U31510 (N_31510,N_29554,N_29701);
or U31511 (N_31511,N_28719,N_28587);
and U31512 (N_31512,N_28848,N_29702);
and U31513 (N_31513,N_29722,N_28831);
xnor U31514 (N_31514,N_29439,N_29446);
or U31515 (N_31515,N_29569,N_28052);
nand U31516 (N_31516,N_29350,N_28014);
nand U31517 (N_31517,N_28377,N_28256);
nand U31518 (N_31518,N_29060,N_29479);
nor U31519 (N_31519,N_28690,N_28179);
nor U31520 (N_31520,N_29792,N_28516);
xor U31521 (N_31521,N_28519,N_29059);
nor U31522 (N_31522,N_29748,N_29260);
or U31523 (N_31523,N_28328,N_28038);
xnor U31524 (N_31524,N_28219,N_28943);
nor U31525 (N_31525,N_29074,N_29838);
nand U31526 (N_31526,N_28672,N_28025);
xnor U31527 (N_31527,N_28147,N_28078);
nand U31528 (N_31528,N_29777,N_29329);
nand U31529 (N_31529,N_29554,N_29306);
nor U31530 (N_31530,N_29852,N_29205);
and U31531 (N_31531,N_28993,N_29721);
nor U31532 (N_31532,N_28120,N_28020);
or U31533 (N_31533,N_29512,N_28913);
and U31534 (N_31534,N_28598,N_28611);
or U31535 (N_31535,N_29635,N_28014);
and U31536 (N_31536,N_29184,N_29432);
nor U31537 (N_31537,N_29577,N_28227);
nand U31538 (N_31538,N_28957,N_28035);
or U31539 (N_31539,N_29518,N_29889);
nand U31540 (N_31540,N_29213,N_29950);
xnor U31541 (N_31541,N_29651,N_29429);
xnor U31542 (N_31542,N_29685,N_28834);
or U31543 (N_31543,N_29435,N_28046);
nand U31544 (N_31544,N_29647,N_28990);
and U31545 (N_31545,N_29990,N_28646);
nor U31546 (N_31546,N_28691,N_28459);
nor U31547 (N_31547,N_29279,N_28372);
nand U31548 (N_31548,N_28516,N_29348);
nand U31549 (N_31549,N_29745,N_28460);
and U31550 (N_31550,N_29162,N_29663);
xnor U31551 (N_31551,N_28040,N_28221);
and U31552 (N_31552,N_29277,N_28976);
nand U31553 (N_31553,N_28452,N_29496);
nand U31554 (N_31554,N_29217,N_28185);
nand U31555 (N_31555,N_28880,N_28570);
xor U31556 (N_31556,N_29405,N_28769);
nor U31557 (N_31557,N_28871,N_29503);
and U31558 (N_31558,N_29781,N_29529);
and U31559 (N_31559,N_29257,N_29534);
nor U31560 (N_31560,N_29726,N_28068);
or U31561 (N_31561,N_28314,N_29119);
or U31562 (N_31562,N_28423,N_28313);
nand U31563 (N_31563,N_29971,N_29562);
nor U31564 (N_31564,N_29334,N_28130);
nor U31565 (N_31565,N_28428,N_29465);
and U31566 (N_31566,N_29249,N_29719);
or U31567 (N_31567,N_28054,N_29208);
xnor U31568 (N_31568,N_28905,N_28780);
and U31569 (N_31569,N_28045,N_29396);
xnor U31570 (N_31570,N_29707,N_28230);
or U31571 (N_31571,N_28283,N_29571);
and U31572 (N_31572,N_28094,N_29375);
xor U31573 (N_31573,N_29678,N_28925);
and U31574 (N_31574,N_28569,N_29113);
nor U31575 (N_31575,N_29426,N_29849);
nor U31576 (N_31576,N_29188,N_28736);
and U31577 (N_31577,N_28291,N_29578);
xnor U31578 (N_31578,N_29334,N_29719);
or U31579 (N_31579,N_28588,N_28228);
nand U31580 (N_31580,N_28623,N_28022);
nand U31581 (N_31581,N_28041,N_29519);
and U31582 (N_31582,N_29217,N_28313);
or U31583 (N_31583,N_29687,N_28383);
nand U31584 (N_31584,N_29455,N_28327);
or U31585 (N_31585,N_29759,N_28451);
nor U31586 (N_31586,N_28277,N_28845);
nand U31587 (N_31587,N_29745,N_28445);
and U31588 (N_31588,N_29384,N_29329);
xnor U31589 (N_31589,N_29866,N_28881);
and U31590 (N_31590,N_28950,N_28526);
nor U31591 (N_31591,N_28290,N_28817);
xor U31592 (N_31592,N_29988,N_29515);
and U31593 (N_31593,N_28764,N_28323);
nor U31594 (N_31594,N_29159,N_28385);
and U31595 (N_31595,N_28747,N_29524);
or U31596 (N_31596,N_29100,N_29962);
xor U31597 (N_31597,N_29239,N_29898);
and U31598 (N_31598,N_29354,N_29449);
nand U31599 (N_31599,N_28312,N_29125);
and U31600 (N_31600,N_28892,N_28331);
xnor U31601 (N_31601,N_28921,N_29380);
xor U31602 (N_31602,N_28069,N_29612);
nand U31603 (N_31603,N_29149,N_28728);
or U31604 (N_31604,N_29440,N_28635);
or U31605 (N_31605,N_29672,N_29927);
nor U31606 (N_31606,N_29322,N_28076);
xor U31607 (N_31607,N_28050,N_29665);
xor U31608 (N_31608,N_28867,N_28327);
nor U31609 (N_31609,N_28508,N_29581);
nor U31610 (N_31610,N_29941,N_28521);
nor U31611 (N_31611,N_29105,N_29758);
xor U31612 (N_31612,N_28366,N_29794);
nand U31613 (N_31613,N_29664,N_29589);
or U31614 (N_31614,N_28468,N_28008);
or U31615 (N_31615,N_28469,N_29069);
xnor U31616 (N_31616,N_29631,N_28062);
or U31617 (N_31617,N_29887,N_29496);
and U31618 (N_31618,N_28001,N_29363);
xnor U31619 (N_31619,N_28198,N_28510);
or U31620 (N_31620,N_28919,N_29746);
nor U31621 (N_31621,N_29692,N_29064);
nor U31622 (N_31622,N_28902,N_29239);
or U31623 (N_31623,N_29190,N_28794);
nand U31624 (N_31624,N_29134,N_29665);
and U31625 (N_31625,N_28070,N_28937);
nor U31626 (N_31626,N_28929,N_28550);
nand U31627 (N_31627,N_29579,N_29448);
nor U31628 (N_31628,N_28010,N_29136);
xor U31629 (N_31629,N_28445,N_29011);
nand U31630 (N_31630,N_28240,N_29383);
nand U31631 (N_31631,N_28303,N_28455);
nor U31632 (N_31632,N_29030,N_29759);
or U31633 (N_31633,N_28963,N_29718);
and U31634 (N_31634,N_29691,N_29283);
nor U31635 (N_31635,N_28836,N_29568);
nor U31636 (N_31636,N_29108,N_28327);
nand U31637 (N_31637,N_29448,N_28068);
nor U31638 (N_31638,N_28562,N_28546);
or U31639 (N_31639,N_29942,N_28402);
or U31640 (N_31640,N_28563,N_29594);
or U31641 (N_31641,N_28268,N_28290);
or U31642 (N_31642,N_28977,N_28537);
nand U31643 (N_31643,N_29533,N_28780);
xnor U31644 (N_31644,N_28424,N_28559);
or U31645 (N_31645,N_29368,N_28803);
xnor U31646 (N_31646,N_29350,N_29825);
xnor U31647 (N_31647,N_28279,N_29756);
nand U31648 (N_31648,N_29733,N_28226);
nand U31649 (N_31649,N_28619,N_29781);
nor U31650 (N_31650,N_28093,N_29728);
xnor U31651 (N_31651,N_28641,N_28755);
nand U31652 (N_31652,N_28512,N_29525);
and U31653 (N_31653,N_29654,N_28976);
or U31654 (N_31654,N_28498,N_29989);
or U31655 (N_31655,N_28560,N_29435);
nand U31656 (N_31656,N_29293,N_28041);
nor U31657 (N_31657,N_29444,N_28648);
nand U31658 (N_31658,N_28766,N_29648);
xnor U31659 (N_31659,N_29654,N_28467);
or U31660 (N_31660,N_28658,N_28193);
nand U31661 (N_31661,N_28947,N_29571);
or U31662 (N_31662,N_28149,N_28180);
or U31663 (N_31663,N_29308,N_29196);
nand U31664 (N_31664,N_28933,N_29452);
and U31665 (N_31665,N_29374,N_28991);
nand U31666 (N_31666,N_29360,N_28224);
xnor U31667 (N_31667,N_28783,N_28124);
xor U31668 (N_31668,N_28138,N_28825);
nor U31669 (N_31669,N_29630,N_29414);
nand U31670 (N_31670,N_28137,N_29173);
nand U31671 (N_31671,N_28493,N_28752);
or U31672 (N_31672,N_28081,N_28443);
xor U31673 (N_31673,N_28574,N_29062);
and U31674 (N_31674,N_28950,N_28573);
nand U31675 (N_31675,N_28318,N_29801);
or U31676 (N_31676,N_28299,N_28102);
or U31677 (N_31677,N_28449,N_28684);
xor U31678 (N_31678,N_28160,N_29260);
or U31679 (N_31679,N_29912,N_28420);
nor U31680 (N_31680,N_29716,N_29616);
xor U31681 (N_31681,N_29403,N_28485);
nand U31682 (N_31682,N_29115,N_28877);
nor U31683 (N_31683,N_29593,N_28698);
xnor U31684 (N_31684,N_28959,N_28511);
nor U31685 (N_31685,N_28946,N_29286);
or U31686 (N_31686,N_29657,N_29323);
or U31687 (N_31687,N_29012,N_29638);
and U31688 (N_31688,N_29706,N_29836);
and U31689 (N_31689,N_29660,N_28282);
xor U31690 (N_31690,N_28894,N_28416);
nor U31691 (N_31691,N_28735,N_29613);
nor U31692 (N_31692,N_29069,N_28181);
nand U31693 (N_31693,N_29147,N_29579);
xnor U31694 (N_31694,N_29169,N_28865);
nor U31695 (N_31695,N_28851,N_29197);
xnor U31696 (N_31696,N_28403,N_28750);
xor U31697 (N_31697,N_28426,N_29214);
or U31698 (N_31698,N_29575,N_28197);
or U31699 (N_31699,N_29493,N_28372);
xor U31700 (N_31700,N_28646,N_28780);
nand U31701 (N_31701,N_28103,N_28436);
xnor U31702 (N_31702,N_28163,N_28800);
xor U31703 (N_31703,N_29205,N_29389);
nand U31704 (N_31704,N_29406,N_29091);
and U31705 (N_31705,N_29648,N_28414);
xnor U31706 (N_31706,N_28460,N_29590);
nor U31707 (N_31707,N_29239,N_29166);
and U31708 (N_31708,N_29287,N_29912);
nor U31709 (N_31709,N_28811,N_28145);
nor U31710 (N_31710,N_28951,N_28911);
or U31711 (N_31711,N_29593,N_28131);
nand U31712 (N_31712,N_28071,N_28580);
and U31713 (N_31713,N_29007,N_29126);
nand U31714 (N_31714,N_29873,N_28582);
xor U31715 (N_31715,N_29386,N_28835);
and U31716 (N_31716,N_29704,N_28609);
or U31717 (N_31717,N_29041,N_29369);
nor U31718 (N_31718,N_28962,N_28891);
xor U31719 (N_31719,N_29879,N_29514);
nand U31720 (N_31720,N_28022,N_29274);
and U31721 (N_31721,N_28616,N_28582);
nor U31722 (N_31722,N_28487,N_28329);
or U31723 (N_31723,N_28495,N_29421);
or U31724 (N_31724,N_29061,N_29771);
and U31725 (N_31725,N_29506,N_29778);
xnor U31726 (N_31726,N_28893,N_28482);
or U31727 (N_31727,N_28730,N_28377);
xor U31728 (N_31728,N_28545,N_29291);
nand U31729 (N_31729,N_28696,N_29439);
nor U31730 (N_31730,N_29892,N_28279);
nor U31731 (N_31731,N_29919,N_29333);
and U31732 (N_31732,N_29712,N_29846);
nand U31733 (N_31733,N_28057,N_29042);
nor U31734 (N_31734,N_29959,N_28256);
nand U31735 (N_31735,N_28187,N_28616);
and U31736 (N_31736,N_28708,N_28528);
and U31737 (N_31737,N_29907,N_28165);
nor U31738 (N_31738,N_29476,N_28983);
nor U31739 (N_31739,N_28085,N_29792);
and U31740 (N_31740,N_29191,N_28947);
xor U31741 (N_31741,N_28356,N_28199);
nor U31742 (N_31742,N_29128,N_28621);
nor U31743 (N_31743,N_29372,N_29728);
nand U31744 (N_31744,N_28883,N_29242);
nand U31745 (N_31745,N_29673,N_28440);
nor U31746 (N_31746,N_29111,N_28786);
and U31747 (N_31747,N_29197,N_28087);
nand U31748 (N_31748,N_29357,N_29843);
and U31749 (N_31749,N_29878,N_29494);
and U31750 (N_31750,N_28208,N_28136);
and U31751 (N_31751,N_28969,N_28876);
or U31752 (N_31752,N_28657,N_28422);
xnor U31753 (N_31753,N_29579,N_29398);
and U31754 (N_31754,N_29275,N_28215);
and U31755 (N_31755,N_29709,N_29126);
nand U31756 (N_31756,N_28460,N_28147);
nand U31757 (N_31757,N_28071,N_29082);
xnor U31758 (N_31758,N_28148,N_28297);
xor U31759 (N_31759,N_29074,N_29756);
xnor U31760 (N_31760,N_28615,N_28898);
and U31761 (N_31761,N_28786,N_28987);
xnor U31762 (N_31762,N_28971,N_29122);
and U31763 (N_31763,N_28181,N_28688);
or U31764 (N_31764,N_29465,N_29606);
nor U31765 (N_31765,N_29835,N_29777);
nand U31766 (N_31766,N_28265,N_28814);
nor U31767 (N_31767,N_29474,N_28896);
nand U31768 (N_31768,N_28606,N_28263);
nand U31769 (N_31769,N_28567,N_29375);
or U31770 (N_31770,N_29247,N_29497);
nor U31771 (N_31771,N_29979,N_28348);
xor U31772 (N_31772,N_29644,N_29273);
or U31773 (N_31773,N_29183,N_28272);
nand U31774 (N_31774,N_29391,N_29736);
nor U31775 (N_31775,N_29776,N_28038);
nor U31776 (N_31776,N_28147,N_28621);
nor U31777 (N_31777,N_29174,N_28867);
nand U31778 (N_31778,N_29348,N_28480);
nor U31779 (N_31779,N_28721,N_28411);
nor U31780 (N_31780,N_29865,N_29627);
xor U31781 (N_31781,N_28137,N_28684);
and U31782 (N_31782,N_29075,N_29134);
or U31783 (N_31783,N_28952,N_29867);
nor U31784 (N_31784,N_28820,N_29252);
nor U31785 (N_31785,N_28551,N_28160);
xor U31786 (N_31786,N_29852,N_29846);
or U31787 (N_31787,N_28182,N_28341);
or U31788 (N_31788,N_29515,N_28898);
xor U31789 (N_31789,N_29595,N_29894);
or U31790 (N_31790,N_28961,N_28165);
or U31791 (N_31791,N_28467,N_29660);
and U31792 (N_31792,N_29765,N_29114);
xor U31793 (N_31793,N_29811,N_28113);
nand U31794 (N_31794,N_28387,N_28996);
xor U31795 (N_31795,N_28351,N_28603);
nand U31796 (N_31796,N_28798,N_28816);
or U31797 (N_31797,N_29385,N_28490);
or U31798 (N_31798,N_28241,N_28350);
nor U31799 (N_31799,N_28688,N_28785);
xnor U31800 (N_31800,N_28675,N_29564);
and U31801 (N_31801,N_28995,N_28965);
xor U31802 (N_31802,N_28665,N_28526);
and U31803 (N_31803,N_29177,N_29135);
or U31804 (N_31804,N_28877,N_29092);
or U31805 (N_31805,N_28881,N_28641);
nor U31806 (N_31806,N_28693,N_29459);
nor U31807 (N_31807,N_28436,N_28466);
xor U31808 (N_31808,N_29365,N_28336);
nand U31809 (N_31809,N_28049,N_28973);
and U31810 (N_31810,N_29319,N_29502);
xor U31811 (N_31811,N_28713,N_29507);
nor U31812 (N_31812,N_28872,N_29019);
nand U31813 (N_31813,N_28657,N_28053);
nor U31814 (N_31814,N_29068,N_29806);
and U31815 (N_31815,N_29427,N_28997);
nand U31816 (N_31816,N_29048,N_29800);
xor U31817 (N_31817,N_29324,N_29797);
or U31818 (N_31818,N_29300,N_28083);
xor U31819 (N_31819,N_28723,N_29832);
nor U31820 (N_31820,N_28465,N_28918);
nor U31821 (N_31821,N_29411,N_29696);
nand U31822 (N_31822,N_29216,N_28186);
nor U31823 (N_31823,N_28718,N_28665);
nor U31824 (N_31824,N_29949,N_29063);
xor U31825 (N_31825,N_28380,N_29164);
or U31826 (N_31826,N_28555,N_28409);
and U31827 (N_31827,N_28243,N_28163);
xor U31828 (N_31828,N_28518,N_28950);
or U31829 (N_31829,N_29945,N_28130);
xnor U31830 (N_31830,N_28338,N_28359);
and U31831 (N_31831,N_28524,N_28765);
nand U31832 (N_31832,N_29713,N_29489);
nor U31833 (N_31833,N_28928,N_28769);
xor U31834 (N_31834,N_28058,N_29619);
or U31835 (N_31835,N_29194,N_28833);
xnor U31836 (N_31836,N_29333,N_29810);
nor U31837 (N_31837,N_29878,N_29686);
or U31838 (N_31838,N_29320,N_28769);
nor U31839 (N_31839,N_29400,N_28536);
or U31840 (N_31840,N_29599,N_29296);
nand U31841 (N_31841,N_28647,N_29467);
nand U31842 (N_31842,N_28113,N_29063);
xor U31843 (N_31843,N_28393,N_29827);
or U31844 (N_31844,N_28113,N_28579);
or U31845 (N_31845,N_28410,N_28832);
nand U31846 (N_31846,N_29217,N_28897);
and U31847 (N_31847,N_28570,N_29223);
nor U31848 (N_31848,N_28408,N_28452);
nand U31849 (N_31849,N_29554,N_28225);
nand U31850 (N_31850,N_28332,N_29959);
or U31851 (N_31851,N_29979,N_29543);
nand U31852 (N_31852,N_28366,N_29337);
or U31853 (N_31853,N_29334,N_28206);
or U31854 (N_31854,N_28132,N_28750);
and U31855 (N_31855,N_28578,N_28311);
xor U31856 (N_31856,N_29373,N_28748);
xnor U31857 (N_31857,N_28668,N_29847);
xnor U31858 (N_31858,N_28288,N_29163);
nand U31859 (N_31859,N_28192,N_29334);
nand U31860 (N_31860,N_28345,N_28634);
or U31861 (N_31861,N_29414,N_28364);
and U31862 (N_31862,N_28371,N_28321);
or U31863 (N_31863,N_28074,N_28424);
xnor U31864 (N_31864,N_28430,N_29110);
nor U31865 (N_31865,N_29683,N_29179);
or U31866 (N_31866,N_29536,N_28962);
xor U31867 (N_31867,N_29373,N_28916);
or U31868 (N_31868,N_29745,N_29147);
xnor U31869 (N_31869,N_29151,N_29861);
and U31870 (N_31870,N_28269,N_28506);
nor U31871 (N_31871,N_29105,N_29434);
nand U31872 (N_31872,N_28023,N_29951);
nand U31873 (N_31873,N_28706,N_29760);
or U31874 (N_31874,N_28170,N_28581);
nor U31875 (N_31875,N_29952,N_28956);
or U31876 (N_31876,N_28359,N_28057);
nor U31877 (N_31877,N_29320,N_29355);
nor U31878 (N_31878,N_28407,N_28992);
and U31879 (N_31879,N_28766,N_29552);
or U31880 (N_31880,N_28769,N_29752);
xnor U31881 (N_31881,N_28954,N_29372);
xnor U31882 (N_31882,N_28113,N_29373);
nor U31883 (N_31883,N_29244,N_28247);
and U31884 (N_31884,N_28170,N_29043);
nand U31885 (N_31885,N_28188,N_29814);
or U31886 (N_31886,N_28621,N_29307);
nand U31887 (N_31887,N_28486,N_28896);
nand U31888 (N_31888,N_29443,N_29418);
nand U31889 (N_31889,N_28921,N_28422);
or U31890 (N_31890,N_29384,N_28579);
xnor U31891 (N_31891,N_29206,N_28822);
or U31892 (N_31892,N_29471,N_28936);
xnor U31893 (N_31893,N_28646,N_29372);
and U31894 (N_31894,N_28584,N_28231);
nor U31895 (N_31895,N_28707,N_28563);
and U31896 (N_31896,N_29051,N_28509);
and U31897 (N_31897,N_28396,N_29741);
xnor U31898 (N_31898,N_28002,N_28102);
nor U31899 (N_31899,N_29567,N_29012);
or U31900 (N_31900,N_29392,N_28884);
or U31901 (N_31901,N_28214,N_29778);
xor U31902 (N_31902,N_29107,N_29580);
and U31903 (N_31903,N_29430,N_28935);
xor U31904 (N_31904,N_29792,N_28244);
and U31905 (N_31905,N_28303,N_28916);
and U31906 (N_31906,N_29746,N_29748);
nor U31907 (N_31907,N_29374,N_29520);
nor U31908 (N_31908,N_29256,N_29769);
xor U31909 (N_31909,N_28322,N_29273);
or U31910 (N_31910,N_28727,N_28739);
nand U31911 (N_31911,N_28930,N_29742);
and U31912 (N_31912,N_28744,N_29316);
or U31913 (N_31913,N_28723,N_29875);
xnor U31914 (N_31914,N_28376,N_28454);
xnor U31915 (N_31915,N_28557,N_28446);
or U31916 (N_31916,N_28966,N_29439);
and U31917 (N_31917,N_28801,N_29541);
xnor U31918 (N_31918,N_29211,N_29224);
nand U31919 (N_31919,N_29870,N_28113);
nor U31920 (N_31920,N_28613,N_28904);
and U31921 (N_31921,N_29183,N_28668);
nor U31922 (N_31922,N_29319,N_29328);
nand U31923 (N_31923,N_28603,N_29927);
nor U31924 (N_31924,N_29492,N_28808);
nor U31925 (N_31925,N_28585,N_28868);
and U31926 (N_31926,N_28444,N_28114);
nor U31927 (N_31927,N_29934,N_28572);
nor U31928 (N_31928,N_29678,N_29163);
nand U31929 (N_31929,N_28615,N_29944);
nand U31930 (N_31930,N_29125,N_28545);
nand U31931 (N_31931,N_29015,N_28231);
nor U31932 (N_31932,N_29052,N_29031);
and U31933 (N_31933,N_29030,N_29331);
nand U31934 (N_31934,N_29698,N_28374);
xnor U31935 (N_31935,N_29651,N_29951);
xnor U31936 (N_31936,N_29571,N_29209);
nor U31937 (N_31937,N_28105,N_29666);
xor U31938 (N_31938,N_29940,N_28489);
xnor U31939 (N_31939,N_29234,N_29945);
and U31940 (N_31940,N_29377,N_29328);
and U31941 (N_31941,N_28565,N_28555);
and U31942 (N_31942,N_28335,N_28544);
nor U31943 (N_31943,N_28022,N_28689);
xor U31944 (N_31944,N_28423,N_29251);
nand U31945 (N_31945,N_29326,N_29138);
nand U31946 (N_31946,N_29197,N_28618);
xor U31947 (N_31947,N_29395,N_29455);
or U31948 (N_31948,N_28029,N_29898);
and U31949 (N_31949,N_28333,N_29444);
xor U31950 (N_31950,N_28328,N_29531);
or U31951 (N_31951,N_29823,N_28922);
or U31952 (N_31952,N_28782,N_29482);
xnor U31953 (N_31953,N_28053,N_29465);
and U31954 (N_31954,N_29582,N_29600);
nand U31955 (N_31955,N_28542,N_29662);
and U31956 (N_31956,N_28065,N_29598);
nand U31957 (N_31957,N_28273,N_29405);
nor U31958 (N_31958,N_28593,N_29321);
xnor U31959 (N_31959,N_29855,N_28312);
xnor U31960 (N_31960,N_29167,N_29075);
or U31961 (N_31961,N_28058,N_28325);
nor U31962 (N_31962,N_29024,N_29267);
and U31963 (N_31963,N_29004,N_28175);
nor U31964 (N_31964,N_29330,N_29672);
nor U31965 (N_31965,N_28438,N_29126);
nor U31966 (N_31966,N_29408,N_29788);
or U31967 (N_31967,N_29389,N_28876);
and U31968 (N_31968,N_29766,N_29524);
nor U31969 (N_31969,N_28976,N_28335);
and U31970 (N_31970,N_29981,N_29402);
and U31971 (N_31971,N_29537,N_28637);
and U31972 (N_31972,N_29704,N_29947);
and U31973 (N_31973,N_29910,N_29659);
xnor U31974 (N_31974,N_29227,N_28960);
or U31975 (N_31975,N_28986,N_29283);
and U31976 (N_31976,N_29756,N_28861);
or U31977 (N_31977,N_29192,N_28274);
and U31978 (N_31978,N_29380,N_28845);
and U31979 (N_31979,N_29080,N_28732);
xnor U31980 (N_31980,N_29184,N_28286);
and U31981 (N_31981,N_28858,N_29232);
nand U31982 (N_31982,N_28241,N_29352);
nor U31983 (N_31983,N_29807,N_29266);
nor U31984 (N_31984,N_29257,N_29932);
xor U31985 (N_31985,N_29143,N_28196);
nand U31986 (N_31986,N_29944,N_28617);
nor U31987 (N_31987,N_28270,N_29568);
nand U31988 (N_31988,N_29383,N_29339);
or U31989 (N_31989,N_28583,N_29608);
xnor U31990 (N_31990,N_28291,N_29680);
nor U31991 (N_31991,N_29450,N_28094);
and U31992 (N_31992,N_29409,N_28695);
or U31993 (N_31993,N_28007,N_29053);
and U31994 (N_31994,N_29482,N_28709);
nand U31995 (N_31995,N_28840,N_29428);
or U31996 (N_31996,N_29785,N_29478);
xnor U31997 (N_31997,N_29714,N_29465);
nand U31998 (N_31998,N_28221,N_29327);
nand U31999 (N_31999,N_29006,N_29109);
nand U32000 (N_32000,N_31030,N_30451);
nand U32001 (N_32001,N_31162,N_31277);
or U32002 (N_32002,N_31955,N_30119);
or U32003 (N_32003,N_31238,N_30516);
or U32004 (N_32004,N_30917,N_31788);
and U32005 (N_32005,N_31660,N_31027);
nand U32006 (N_32006,N_31863,N_31598);
nand U32007 (N_32007,N_30342,N_30739);
nor U32008 (N_32008,N_30117,N_30840);
and U32009 (N_32009,N_30462,N_31237);
nand U32010 (N_32010,N_31946,N_31632);
and U32011 (N_32011,N_30711,N_30726);
nor U32012 (N_32012,N_31222,N_31518);
or U32013 (N_32013,N_31704,N_31415);
or U32014 (N_32014,N_31752,N_31491);
xnor U32015 (N_32015,N_31777,N_31144);
nand U32016 (N_32016,N_30386,N_30586);
nor U32017 (N_32017,N_31726,N_30373);
nor U32018 (N_32018,N_30653,N_31104);
or U32019 (N_32019,N_30245,N_31380);
nand U32020 (N_32020,N_31792,N_30659);
xor U32021 (N_32021,N_30897,N_31472);
xnor U32022 (N_32022,N_31166,N_31947);
nand U32023 (N_32023,N_31125,N_31705);
xor U32024 (N_32024,N_30389,N_30454);
or U32025 (N_32025,N_30699,N_30460);
nand U32026 (N_32026,N_31119,N_30062);
or U32027 (N_32027,N_30965,N_30625);
and U32028 (N_32028,N_31572,N_31213);
and U32029 (N_32029,N_30508,N_31248);
nor U32030 (N_32030,N_31790,N_30555);
nand U32031 (N_32031,N_31844,N_30996);
or U32032 (N_32032,N_30227,N_30091);
nand U32033 (N_32033,N_30667,N_31379);
nor U32034 (N_32034,N_30989,N_31061);
or U32035 (N_32035,N_31188,N_30638);
and U32036 (N_32036,N_31214,N_31171);
nand U32037 (N_32037,N_30219,N_31991);
nand U32038 (N_32038,N_31130,N_31732);
or U32039 (N_32039,N_31000,N_30866);
or U32040 (N_32040,N_31892,N_30115);
nand U32041 (N_32041,N_30490,N_31891);
and U32042 (N_32042,N_30118,N_31227);
xnor U32043 (N_32043,N_31658,N_31260);
nor U32044 (N_32044,N_30352,N_30515);
nor U32045 (N_32045,N_30283,N_31908);
and U32046 (N_32046,N_30400,N_30693);
and U32047 (N_32047,N_31833,N_31668);
xnor U32048 (N_32048,N_31507,N_30871);
xnor U32049 (N_32049,N_31387,N_30754);
xor U32050 (N_32050,N_30941,N_30177);
xnor U32051 (N_32051,N_30150,N_31490);
nor U32052 (N_32052,N_30253,N_30856);
nor U32053 (N_32053,N_30341,N_30696);
nor U32054 (N_32054,N_30790,N_30632);
nor U32055 (N_32055,N_30345,N_31739);
nand U32056 (N_32056,N_31943,N_30873);
or U32057 (N_32057,N_31841,N_31635);
and U32058 (N_32058,N_30438,N_30288);
or U32059 (N_32059,N_30361,N_30616);
nor U32060 (N_32060,N_30331,N_31604);
nor U32061 (N_32061,N_31366,N_30461);
and U32062 (N_32062,N_30836,N_30011);
nor U32063 (N_32063,N_31583,N_31143);
nor U32064 (N_32064,N_31595,N_30466);
nand U32065 (N_32065,N_30885,N_31318);
and U32066 (N_32066,N_30683,N_31981);
xor U32067 (N_32067,N_30966,N_30259);
or U32068 (N_32068,N_31519,N_31483);
nand U32069 (N_32069,N_30000,N_30909);
nor U32070 (N_32070,N_31120,N_30041);
nand U32071 (N_32071,N_30145,N_31454);
nor U32072 (N_32072,N_30872,N_31703);
and U32073 (N_32073,N_31170,N_30380);
xnor U32074 (N_32074,N_30825,N_31858);
nor U32075 (N_32075,N_30070,N_30753);
xnor U32076 (N_32076,N_30126,N_31763);
or U32077 (N_32077,N_31046,N_30995);
nor U32078 (N_32078,N_30561,N_30621);
and U32079 (N_32079,N_31169,N_30196);
or U32080 (N_32080,N_30901,N_30709);
and U32081 (N_32081,N_30633,N_30073);
and U32082 (N_32082,N_30808,N_31330);
or U32083 (N_32083,N_31830,N_30647);
nand U32084 (N_32084,N_31573,N_31346);
xnor U32085 (N_32085,N_30101,N_30988);
nor U32086 (N_32086,N_31612,N_31811);
and U32087 (N_32087,N_30583,N_31857);
and U32088 (N_32088,N_31562,N_31839);
xnor U32089 (N_32089,N_30356,N_31862);
xor U32090 (N_32090,N_30278,N_31345);
nand U32091 (N_32091,N_30784,N_31702);
and U32092 (N_32092,N_31296,N_30521);
nand U32093 (N_32093,N_31544,N_30025);
xor U32094 (N_32094,N_30804,N_30611);
nand U32095 (N_32095,N_30795,N_30176);
nand U32096 (N_32096,N_31771,N_30534);
nor U32097 (N_32097,N_31650,N_30172);
nand U32098 (N_32098,N_30056,N_31560);
xnor U32099 (N_32099,N_31968,N_30701);
nor U32100 (N_32100,N_30147,N_30817);
nor U32101 (N_32101,N_30299,N_30982);
nand U32102 (N_32102,N_30890,N_30854);
nand U32103 (N_32103,N_31928,N_30525);
or U32104 (N_32104,N_30788,N_31556);
nand U32105 (N_32105,N_30628,N_31075);
and U32106 (N_32106,N_31499,N_31493);
and U32107 (N_32107,N_31189,N_30455);
nand U32108 (N_32108,N_31740,N_31090);
xor U32109 (N_32109,N_30403,N_31459);
nand U32110 (N_32110,N_30927,N_30411);
or U32111 (N_32111,N_31682,N_30751);
nand U32112 (N_32112,N_31087,N_30656);
nor U32113 (N_32113,N_31926,N_31288);
and U32114 (N_32114,N_31464,N_31698);
nand U32115 (N_32115,N_31787,N_31023);
or U32116 (N_32116,N_30363,N_31010);
nor U32117 (N_32117,N_30435,N_30348);
nor U32118 (N_32118,N_30410,N_31450);
or U32119 (N_32119,N_31411,N_31951);
nand U32120 (N_32120,N_31097,N_31205);
and U32121 (N_32121,N_30421,N_30758);
xor U32122 (N_32122,N_30413,N_30522);
xnor U32123 (N_32123,N_30047,N_31901);
and U32124 (N_32124,N_30406,N_30979);
or U32125 (N_32125,N_31550,N_30067);
and U32126 (N_32126,N_30669,N_30578);
nand U32127 (N_32127,N_30963,N_31389);
and U32128 (N_32128,N_30130,N_31314);
or U32129 (N_32129,N_31184,N_31385);
and U32130 (N_32130,N_30512,N_31948);
xor U32131 (N_32131,N_30530,N_31126);
nor U32132 (N_32132,N_31983,N_30194);
or U32133 (N_32133,N_31079,N_31223);
and U32134 (N_32134,N_30477,N_30900);
xor U32135 (N_32135,N_30506,N_31909);
or U32136 (N_32136,N_31799,N_31683);
or U32137 (N_32137,N_30549,N_31744);
nand U32138 (N_32138,N_31128,N_30376);
nor U32139 (N_32139,N_31866,N_30293);
and U32140 (N_32140,N_31358,N_30281);
and U32141 (N_32141,N_31502,N_31225);
xor U32142 (N_32142,N_30390,N_30449);
xnor U32143 (N_32143,N_31462,N_30811);
and U32144 (N_32144,N_31309,N_31714);
or U32145 (N_32145,N_30095,N_30159);
xor U32146 (N_32146,N_31673,N_31504);
or U32147 (N_32147,N_30504,N_31655);
or U32148 (N_32148,N_31966,N_31069);
or U32149 (N_32149,N_30407,N_31390);
and U32150 (N_32150,N_31378,N_31074);
nor U32151 (N_32151,N_30307,N_30318);
and U32152 (N_32152,N_30317,N_31108);
nor U32153 (N_32153,N_31717,N_31640);
nand U32154 (N_32154,N_31369,N_31756);
xor U32155 (N_32155,N_30241,N_30644);
and U32156 (N_32156,N_31755,N_31810);
and U32157 (N_32157,N_31876,N_31797);
nor U32158 (N_32158,N_30960,N_31293);
or U32159 (N_32159,N_31012,N_31172);
and U32160 (N_32160,N_31896,N_30173);
xor U32161 (N_32161,N_31158,N_30572);
nand U32162 (N_32162,N_31581,N_31988);
xor U32163 (N_32163,N_30843,N_30266);
nor U32164 (N_32164,N_31233,N_30916);
xnor U32165 (N_32165,N_31461,N_30268);
or U32166 (N_32166,N_30273,N_31699);
nor U32167 (N_32167,N_30886,N_31035);
or U32168 (N_32168,N_30735,N_30167);
and U32169 (N_32169,N_31443,N_31394);
nand U32170 (N_32170,N_30304,N_30322);
or U32171 (N_32171,N_30676,N_30598);
and U32172 (N_32172,N_30985,N_30132);
nand U32173 (N_32173,N_31528,N_31460);
nor U32174 (N_32174,N_30412,N_31515);
xnor U32175 (N_32175,N_31364,N_30509);
nand U32176 (N_32176,N_30626,N_30657);
xnor U32177 (N_32177,N_30102,N_30548);
xnor U32178 (N_32178,N_31984,N_30113);
xnor U32179 (N_32179,N_30500,N_30848);
and U32180 (N_32180,N_31999,N_30655);
and U32181 (N_32181,N_31545,N_31949);
nor U32182 (N_32182,N_31342,N_30404);
nand U32183 (N_32183,N_30128,N_30265);
or U32184 (N_32184,N_31548,N_30929);
or U32185 (N_32185,N_31816,N_31791);
or U32186 (N_32186,N_31430,N_30813);
xnor U32187 (N_32187,N_31818,N_31589);
xnor U32188 (N_32188,N_31445,N_30577);
or U32189 (N_32189,N_30715,N_31956);
nor U32190 (N_32190,N_30296,N_31016);
and U32191 (N_32191,N_30685,N_30141);
or U32192 (N_32192,N_31840,N_30098);
nand U32193 (N_32193,N_30756,N_30546);
xnor U32194 (N_32194,N_31398,N_30272);
xor U32195 (N_32195,N_30684,N_31256);
xor U32196 (N_32196,N_30202,N_30816);
and U32197 (N_32197,N_30153,N_31219);
xnor U32198 (N_32198,N_31925,N_31247);
or U32199 (N_32199,N_30999,N_30243);
nor U32200 (N_32200,N_31310,N_30465);
xnor U32201 (N_32201,N_30215,N_30923);
xnor U32202 (N_32202,N_30239,N_30297);
and U32203 (N_32203,N_30742,N_30086);
nand U32204 (N_32204,N_30275,N_30183);
or U32205 (N_32205,N_31147,N_30221);
and U32206 (N_32206,N_31643,N_31940);
nand U32207 (N_32207,N_30907,N_30977);
or U32208 (N_32208,N_30928,N_30889);
or U32209 (N_32209,N_31820,N_30639);
xnor U32210 (N_32210,N_31480,N_31628);
or U32211 (N_32211,N_30133,N_30827);
or U32212 (N_32212,N_30671,N_30946);
nor U32213 (N_32213,N_30589,N_31465);
xor U32214 (N_32214,N_31105,N_30094);
nor U32215 (N_32215,N_30605,N_30984);
and U32216 (N_32216,N_31880,N_31979);
and U32217 (N_32217,N_31985,N_31442);
nor U32218 (N_32218,N_31588,N_31639);
nand U32219 (N_32219,N_31989,N_31211);
and U32220 (N_32220,N_31152,N_31760);
and U32221 (N_32221,N_31495,N_30016);
nor U32222 (N_32222,N_31533,N_31031);
nor U32223 (N_32223,N_30280,N_31070);
or U32224 (N_32224,N_30012,N_31438);
xnor U32225 (N_32225,N_30953,N_30303);
or U32226 (N_32226,N_30931,N_30838);
nor U32227 (N_32227,N_30485,N_30142);
xor U32228 (N_32228,N_31451,N_30707);
nand U32229 (N_32229,N_30483,N_31789);
nor U32230 (N_32230,N_31769,N_31334);
nor U32231 (N_32231,N_30203,N_30375);
and U32232 (N_32232,N_31902,N_31403);
nor U32233 (N_32233,N_30229,N_30934);
or U32234 (N_32234,N_30591,N_30416);
nand U32235 (N_32235,N_30064,N_30498);
nand U32236 (N_32236,N_31974,N_30374);
nor U32237 (N_32237,N_31043,N_31384);
and U32238 (N_32238,N_30986,N_31585);
nor U32239 (N_32239,N_30261,N_30351);
and U32240 (N_32240,N_30563,N_30046);
nor U32241 (N_32241,N_30759,N_31522);
nor U32242 (N_32242,N_30765,N_31295);
nor U32243 (N_32243,N_30214,N_30733);
or U32244 (N_32244,N_31854,N_30803);
nand U32245 (N_32245,N_31764,N_31933);
nand U32246 (N_32246,N_30396,N_30855);
nand U32247 (N_32247,N_31142,N_31889);
and U32248 (N_32248,N_30913,N_30370);
nand U32249 (N_32249,N_31540,N_30039);
nand U32250 (N_32250,N_30852,N_30295);
xnor U32251 (N_32251,N_31441,N_30391);
nor U32252 (N_32252,N_30526,N_31374);
xnor U32253 (N_32253,N_30007,N_31412);
and U32254 (N_32254,N_31496,N_30550);
xnor U32255 (N_32255,N_30335,N_31750);
nand U32256 (N_32256,N_31199,N_31065);
nor U32257 (N_32257,N_30689,N_30874);
xor U32258 (N_32258,N_30725,N_30010);
nor U32259 (N_32259,N_30722,N_30734);
or U32260 (N_32260,N_31605,N_30088);
nor U32261 (N_32261,N_30264,N_30514);
and U32262 (N_32262,N_30328,N_30161);
nand U32263 (N_32263,N_30542,N_30660);
and U32264 (N_32264,N_31049,N_30154);
xor U32265 (N_32265,N_31823,N_31821);
or U32266 (N_32266,N_31831,N_31303);
and U32267 (N_32267,N_31838,N_30812);
nor U32268 (N_32268,N_30155,N_31530);
and U32269 (N_32269,N_30355,N_30998);
xor U32270 (N_32270,N_31526,N_31102);
or U32271 (N_32271,N_30031,N_31014);
or U32272 (N_32272,N_30573,N_31709);
and U32273 (N_32273,N_31196,N_30450);
nand U32274 (N_32274,N_30912,N_30581);
xor U32275 (N_32275,N_30131,N_30895);
or U32276 (N_32276,N_31264,N_30877);
nor U32277 (N_32277,N_31032,N_30805);
nand U32278 (N_32278,N_30997,N_30050);
nor U32279 (N_32279,N_30973,N_31922);
xor U32280 (N_32280,N_31843,N_31052);
nor U32281 (N_32281,N_31853,N_30978);
xor U32282 (N_32282,N_31961,N_31718);
nand U32283 (N_32283,N_31837,N_31145);
xor U32284 (N_32284,N_30782,N_31748);
and U32285 (N_32285,N_30298,N_31117);
xnor U32286 (N_32286,N_31054,N_31186);
and U32287 (N_32287,N_31878,N_31575);
or U32288 (N_32288,N_31910,N_30301);
nor U32289 (N_32289,N_30736,N_30747);
nor U32290 (N_32290,N_31067,N_31363);
or U32291 (N_32291,N_31351,N_30059);
nor U32292 (N_32292,N_30242,N_30922);
and U32293 (N_32293,N_31611,N_31313);
and U32294 (N_32294,N_31352,N_30821);
and U32295 (N_32295,N_31060,N_30137);
xor U32296 (N_32296,N_30664,N_30030);
or U32297 (N_32297,N_30743,N_31904);
nor U32298 (N_32298,N_30994,N_31886);
nand U32299 (N_32299,N_30648,N_30008);
and U32300 (N_32300,N_31906,N_30652);
xnor U32301 (N_32301,N_30513,N_31934);
xor U32302 (N_32302,N_31558,N_31630);
nand U32303 (N_32303,N_30938,N_30990);
or U32304 (N_32304,N_30096,N_30034);
or U32305 (N_32305,N_30206,N_31554);
nor U32306 (N_32306,N_30192,N_30472);
nor U32307 (N_32307,N_31805,N_30106);
nor U32308 (N_32308,N_31423,N_31336);
nand U32309 (N_32309,N_31399,N_31393);
nand U32310 (N_32310,N_31834,N_31557);
or U32311 (N_32311,N_30104,N_30255);
nand U32312 (N_32312,N_30346,N_30222);
xor U32313 (N_32313,N_30055,N_30860);
nor U32314 (N_32314,N_30910,N_30232);
and U32315 (N_32315,N_31681,N_30402);
and U32316 (N_32316,N_31218,N_30085);
nand U32317 (N_32317,N_31111,N_30859);
or U32318 (N_32318,N_30405,N_31191);
nor U32319 (N_32319,N_30190,N_30427);
nand U32320 (N_32320,N_30392,N_31871);
or U32321 (N_32321,N_30875,N_31765);
and U32322 (N_32322,N_31970,N_31672);
nor U32323 (N_32323,N_30757,N_30467);
and U32324 (N_32324,N_31254,N_30839);
nand U32325 (N_32325,N_30724,N_30475);
nand U32326 (N_32326,N_30114,N_31872);
nand U32327 (N_32327,N_31089,N_30809);
or U32328 (N_32328,N_31576,N_30970);
or U32329 (N_32329,N_30668,N_31965);
xor U32330 (N_32330,N_31440,N_31665);
nand U32331 (N_32331,N_30179,N_30246);
or U32332 (N_32332,N_30425,N_31424);
or U32333 (N_32333,N_31996,N_30893);
or U32334 (N_32334,N_30920,N_30325);
or U32335 (N_32335,N_30395,N_30672);
xnor U32336 (N_32336,N_31347,N_31680);
nand U32337 (N_32337,N_31915,N_30223);
or U32338 (N_32338,N_30310,N_30112);
or U32339 (N_32339,N_30925,N_31221);
xor U32340 (N_32340,N_31053,N_31239);
nor U32341 (N_32341,N_30276,N_31669);
xnor U32342 (N_32342,N_31794,N_30491);
nand U32343 (N_32343,N_31434,N_30021);
or U32344 (N_32344,N_31874,N_31124);
or U32345 (N_32345,N_30957,N_30072);
and U32346 (N_32346,N_30362,N_30005);
nor U32347 (N_32347,N_30774,N_31969);
nor U32348 (N_32348,N_31729,N_31944);
nor U32349 (N_32349,N_30603,N_31259);
and U32350 (N_32350,N_31435,N_30123);
nor U32351 (N_32351,N_30712,N_31500);
xor U32352 (N_32352,N_31931,N_30623);
xor U32353 (N_32353,N_30732,N_31649);
and U32354 (N_32354,N_31180,N_30252);
nor U32355 (N_32355,N_30705,N_31082);
nor U32356 (N_32356,N_31381,N_31092);
xor U32357 (N_32357,N_31177,N_31918);
and U32358 (N_32358,N_31255,N_30908);
nor U32359 (N_32359,N_31410,N_31973);
and U32360 (N_32360,N_31676,N_31618);
nor U32361 (N_32361,N_31859,N_30251);
and U32362 (N_32362,N_30204,N_30409);
and U32363 (N_32363,N_31281,N_30612);
nand U32364 (N_32364,N_30778,N_30936);
and U32365 (N_32365,N_31916,N_30051);
nor U32366 (N_32366,N_30480,N_30650);
nor U32367 (N_32367,N_31975,N_31482);
xor U32368 (N_32368,N_31447,N_30903);
and U32369 (N_32369,N_31139,N_31463);
nor U32370 (N_32370,N_30093,N_30146);
or U32371 (N_32371,N_31062,N_30822);
or U32372 (N_32372,N_30954,N_31229);
xnor U32373 (N_32373,N_31994,N_30339);
nand U32374 (N_32374,N_30919,N_31924);
nor U32375 (N_32375,N_30902,N_30023);
xnor U32376 (N_32376,N_30151,N_30422);
nand U32377 (N_32377,N_30748,N_31962);
nand U32378 (N_32378,N_30697,N_30330);
or U32379 (N_32379,N_31091,N_31539);
xor U32380 (N_32380,N_30593,N_31429);
nor U32381 (N_32381,N_30823,N_30143);
nor U32382 (N_32382,N_31116,N_31813);
nor U32383 (N_32383,N_30474,N_31311);
nand U32384 (N_32384,N_31800,N_30810);
or U32385 (N_32385,N_31865,N_31768);
nor U32386 (N_32386,N_30718,N_31426);
or U32387 (N_32387,N_31298,N_30198);
or U32388 (N_32388,N_31037,N_30887);
nand U32389 (N_32389,N_30270,N_31603);
nor U32390 (N_32390,N_30899,N_31449);
and U32391 (N_32391,N_31127,N_30388);
and U32392 (N_32392,N_31033,N_31409);
nand U32393 (N_32393,N_31098,N_31825);
and U32394 (N_32394,N_30429,N_30230);
or U32395 (N_32395,N_31722,N_31942);
nor U32396 (N_32396,N_30746,N_31072);
nor U32397 (N_32397,N_31025,N_31802);
nand U32398 (N_32398,N_30289,N_31829);
nor U32399 (N_32399,N_31354,N_31088);
and U32400 (N_32400,N_31324,N_30048);
or U32401 (N_32401,N_30596,N_31814);
xnor U32402 (N_32402,N_31512,N_31761);
xnor U32403 (N_32403,N_31776,N_31028);
nand U32404 (N_32404,N_30499,N_31505);
or U32405 (N_32405,N_30829,N_30529);
or U32406 (N_32406,N_31101,N_30698);
nand U32407 (N_32407,N_30993,N_31206);
and U32408 (N_32408,N_30158,N_31847);
xor U32409 (N_32409,N_31633,N_31690);
and U32410 (N_32410,N_30523,N_31738);
xor U32411 (N_32411,N_30584,N_31960);
nand U32412 (N_32412,N_31086,N_31574);
xor U32413 (N_32413,N_30505,N_31634);
and U32414 (N_32414,N_31867,N_31316);
nor U32415 (N_32415,N_31846,N_30456);
and U32416 (N_32416,N_31757,N_31967);
and U32417 (N_32417,N_31836,N_31479);
and U32418 (N_32418,N_30134,N_30641);
or U32419 (N_32419,N_30801,N_30643);
or U32420 (N_32420,N_31596,N_31484);
nand U32421 (N_32421,N_31289,N_31064);
and U32422 (N_32422,N_30930,N_31671);
or U32423 (N_32423,N_30002,N_30020);
or U32424 (N_32424,N_30367,N_31011);
or U32425 (N_32425,N_30939,N_31686);
xor U32426 (N_32426,N_31921,N_31520);
xnor U32427 (N_32427,N_30567,N_31341);
and U32428 (N_32428,N_31263,N_31822);
or U32429 (N_32429,N_31852,N_30981);
and U32430 (N_32430,N_31536,N_31236);
and U32431 (N_32431,N_30217,N_30369);
xor U32432 (N_32432,N_31276,N_30068);
nor U32433 (N_32433,N_30675,N_30862);
or U32434 (N_32434,N_31266,N_31273);
xnor U32435 (N_32435,N_31093,N_31995);
and U32436 (N_32436,N_31448,N_30831);
or U32437 (N_32437,N_31506,N_30849);
xnor U32438 (N_32438,N_30181,N_31715);
nor U32439 (N_32439,N_31096,N_30590);
nand U32440 (N_32440,N_31428,N_30687);
nand U32441 (N_32441,N_31468,N_31785);
and U32442 (N_32442,N_30481,N_31657);
and U32443 (N_32443,N_30017,N_30263);
nand U32444 (N_32444,N_31712,N_31986);
nor U32445 (N_32445,N_31489,N_30383);
and U32446 (N_32446,N_30798,N_30891);
nor U32447 (N_32447,N_30964,N_30600);
or U32448 (N_32448,N_31741,N_31308);
and U32449 (N_32449,N_31856,N_31244);
nor U32450 (N_32450,N_30894,N_31485);
xor U32451 (N_32451,N_30360,N_30597);
and U32452 (N_32452,N_31267,N_30807);
or U32453 (N_32453,N_31272,N_31231);
nor U32454 (N_32454,N_31458,N_30863);
nor U32455 (N_32455,N_31514,N_30914);
nand U32456 (N_32456,N_31624,N_31240);
xnor U32457 (N_32457,N_30719,N_31486);
or U32458 (N_32458,N_31401,N_30287);
xor U32459 (N_32459,N_31007,N_30384);
and U32460 (N_32460,N_31181,N_30089);
xor U32461 (N_32461,N_30975,N_30492);
and U32462 (N_32462,N_31537,N_30237);
and U32463 (N_32463,N_30527,N_30180);
and U32464 (N_32464,N_30174,N_31224);
nand U32465 (N_32465,N_31020,N_30184);
nor U32466 (N_32466,N_31553,N_30967);
nand U32467 (N_32467,N_30018,N_30976);
or U32468 (N_32468,N_30501,N_30607);
and U32469 (N_32469,N_30524,N_30164);
nand U32470 (N_32470,N_30285,N_30741);
or U32471 (N_32471,N_30015,N_31466);
xnor U32472 (N_32472,N_30710,N_30442);
nor U32473 (N_32473,N_31076,N_31534);
xor U32474 (N_32474,N_30200,N_31809);
or U32475 (N_32475,N_30444,N_30175);
nand U32476 (N_32476,N_30845,N_31746);
nand U32477 (N_32477,N_30552,N_30453);
and U32478 (N_32478,N_31622,N_31066);
and U32479 (N_32479,N_31971,N_31201);
or U32480 (N_32480,N_30762,N_31297);
or U32481 (N_32481,N_31779,N_30703);
and U32482 (N_32482,N_31579,N_30775);
and U32483 (N_32483,N_31099,N_30320);
and U32484 (N_32484,N_30528,N_30169);
or U32485 (N_32485,N_30940,N_30764);
xor U32486 (N_32486,N_30961,N_30436);
nor U32487 (N_32487,N_30418,N_30447);
and U32488 (N_32488,N_31707,N_31652);
nand U32489 (N_32489,N_31470,N_30654);
and U32490 (N_32490,N_30614,N_31135);
and U32491 (N_32491,N_30543,N_31662);
xnor U32492 (N_32492,N_30945,N_30063);
nand U32493 (N_32493,N_31675,N_31724);
and U32494 (N_32494,N_31864,N_30099);
and U32495 (N_32495,N_30446,N_30915);
nand U32496 (N_32496,N_30306,N_30588);
or U32497 (N_32497,N_31780,N_30417);
and U32498 (N_32498,N_31348,N_31538);
and U32499 (N_32499,N_31938,N_31762);
xnor U32500 (N_32500,N_30918,N_31727);
nand U32501 (N_32501,N_30236,N_31121);
nor U32502 (N_32502,N_30437,N_30448);
nor U32503 (N_32503,N_31736,N_30334);
and U32504 (N_32504,N_30044,N_31359);
xnor U32505 (N_32505,N_31932,N_31895);
nand U32506 (N_32506,N_31408,N_30212);
and U32507 (N_32507,N_31375,N_30789);
or U32508 (N_32508,N_30076,N_30359);
or U32509 (N_32509,N_30924,N_31026);
nor U32510 (N_32510,N_31807,N_31344);
nor U32511 (N_32511,N_31929,N_31160);
or U32512 (N_32512,N_31647,N_30079);
nand U32513 (N_32513,N_31663,N_31559);
or U32514 (N_32514,N_31317,N_30308);
nand U32515 (N_32515,N_31029,N_31642);
or U32516 (N_32516,N_30933,N_30081);
or U32517 (N_32517,N_30559,N_31356);
and U32518 (N_32518,N_30001,N_30111);
nand U32519 (N_32519,N_31391,N_31148);
or U32520 (N_32520,N_31587,N_31701);
nor U32521 (N_32521,N_31508,N_30533);
nor U32522 (N_32522,N_31950,N_30329);
xor U32523 (N_32523,N_31436,N_30032);
or U32524 (N_32524,N_30116,N_30983);
nand U32525 (N_32525,N_30019,N_31850);
nand U32526 (N_32526,N_30470,N_31275);
or U32527 (N_32527,N_30148,N_31728);
nor U32528 (N_32528,N_30870,N_30309);
xor U32529 (N_32529,N_31209,N_31377);
xnor U32530 (N_32530,N_31936,N_30054);
nand U32531 (N_32531,N_30424,N_30868);
nand U32532 (N_32532,N_31163,N_31455);
or U32533 (N_32533,N_30692,N_31306);
and U32534 (N_32534,N_31417,N_30952);
xnor U32535 (N_32535,N_31107,N_31165);
nand U32536 (N_32536,N_30898,N_31555);
nand U32537 (N_32537,N_30408,N_30932);
nor U32538 (N_32538,N_31656,N_30974);
nand U32539 (N_32539,N_30841,N_31582);
nor U32540 (N_32540,N_30835,N_30440);
xnor U32541 (N_32541,N_31469,N_30959);
nor U32542 (N_32542,N_31751,N_31110);
nor U32543 (N_32543,N_30233,N_30152);
nor U32544 (N_32544,N_31242,N_30187);
nand U32545 (N_32545,N_30646,N_30228);
nand U32546 (N_32546,N_30368,N_30881);
and U32547 (N_32547,N_31040,N_31427);
and U32548 (N_32548,N_31195,N_31137);
and U32549 (N_32549,N_30551,N_31939);
xor U32550 (N_32550,N_30888,N_31868);
nand U32551 (N_32551,N_31319,N_30794);
or U32552 (N_32552,N_31759,N_31888);
nand U32553 (N_32553,N_31246,N_30084);
or U32554 (N_32554,N_30028,N_31235);
xnor U32555 (N_32555,N_30702,N_30262);
or U32556 (N_32556,N_30987,N_30796);
or U32557 (N_32557,N_30162,N_30224);
or U32558 (N_32558,N_31198,N_30120);
nand U32559 (N_32559,N_30730,N_31659);
xnor U32560 (N_32560,N_30629,N_30014);
xnor U32561 (N_32561,N_31106,N_30721);
or U32562 (N_32562,N_30791,N_31339);
xor U32563 (N_32563,N_30171,N_30880);
and U32564 (N_32564,N_31400,N_30122);
and U32565 (N_32565,N_31179,N_30968);
xnor U32566 (N_32566,N_30502,N_30980);
and U32567 (N_32567,N_31613,N_30087);
or U32568 (N_32568,N_30785,N_30185);
or U32569 (N_32569,N_31362,N_30029);
nor U32570 (N_32570,N_31963,N_30053);
nor U32571 (N_32571,N_31685,N_31190);
xnor U32572 (N_32572,N_30282,N_31457);
nor U32573 (N_32573,N_31623,N_31848);
and U32574 (N_32574,N_30457,N_30714);
nand U32575 (N_32575,N_30950,N_31568);
nand U32576 (N_32576,N_30832,N_30770);
nor U32577 (N_32577,N_30136,N_30992);
or U32578 (N_32578,N_30844,N_30344);
or U32579 (N_32579,N_31591,N_31332);
or U32580 (N_32580,N_30826,N_30319);
or U32581 (N_32581,N_31100,N_31903);
or U32582 (N_32582,N_30750,N_30324);
xor U32583 (N_32583,N_31719,N_31274);
nor U32584 (N_32584,N_30249,N_31808);
xnor U32585 (N_32585,N_30878,N_30149);
or U32586 (N_32586,N_30824,N_30833);
nor U32587 (N_32587,N_30210,N_30225);
nor U32588 (N_32588,N_30484,N_31475);
and U32589 (N_32589,N_30956,N_30302);
and U32590 (N_32590,N_30949,N_31115);
or U32591 (N_32591,N_30830,N_30350);
or U32592 (N_32592,N_31648,N_30565);
xnor U32593 (N_32593,N_30323,N_31042);
nor U32594 (N_32594,N_30582,N_30060);
nand U32595 (N_32595,N_31775,N_31290);
nor U32596 (N_32596,N_30627,N_31887);
and U32597 (N_32597,N_30165,N_30497);
xnor U32598 (N_32598,N_30495,N_31057);
xnor U32599 (N_32599,N_31284,N_31019);
and U32600 (N_32600,N_31959,N_31433);
and U32601 (N_32601,N_31592,N_30414);
nor U32602 (N_32602,N_30846,N_30315);
nand U32603 (N_32603,N_31419,N_31812);
nand U32604 (N_32604,N_31370,N_31118);
nand U32605 (N_32605,N_30250,N_31159);
and U32606 (N_32606,N_31045,N_31047);
or U32607 (N_32607,N_31329,N_30071);
nor U32608 (N_32608,N_30544,N_31149);
xor U32609 (N_32609,N_30381,N_31621);
and U32610 (N_32610,N_31826,N_31210);
xnor U32611 (N_32611,N_30459,N_30205);
or U32612 (N_32612,N_31899,N_30858);
and U32613 (N_32613,N_30077,N_30615);
xnor U32614 (N_32614,N_30479,N_31208);
or U32615 (N_32615,N_30662,N_30574);
nor U32616 (N_32616,N_30160,N_31133);
nor U32617 (N_32617,N_30037,N_31516);
xor U32618 (N_32618,N_30135,N_31280);
xnor U32619 (N_32619,N_31474,N_31795);
xor U32620 (N_32620,N_31845,N_30943);
xor U32621 (N_32621,N_31140,N_31476);
xor U32622 (N_32622,N_30393,N_30906);
or U32623 (N_32623,N_30078,N_31571);
nand U32624 (N_32624,N_31781,N_31954);
xnor U32625 (N_32625,N_31155,N_30622);
xor U32626 (N_32626,N_30353,N_30004);
nand U32627 (N_32627,N_31747,N_31883);
nor U32628 (N_32628,N_31957,N_30896);
nand U32629 (N_32629,N_30690,N_30636);
and U32630 (N_32630,N_31262,N_31194);
xor U32631 (N_32631,N_31422,N_31234);
xnor U32632 (N_32632,N_31285,N_30942);
nor U32633 (N_32633,N_30478,N_31667);
and U32634 (N_32634,N_30024,N_30640);
or U32635 (N_32635,N_30052,N_30378);
nand U32636 (N_32636,N_30300,N_30321);
xor U32637 (N_32637,N_30314,N_31200);
nand U32638 (N_32638,N_30663,N_31644);
nand U32639 (N_32639,N_30686,N_31692);
or U32640 (N_32640,N_30489,N_30536);
xor U32641 (N_32641,N_30178,N_31215);
or U32642 (N_32642,N_30882,N_31203);
or U32643 (N_32643,N_31299,N_30163);
xor U32644 (N_32644,N_31625,N_31881);
nor U32645 (N_32645,N_30673,N_30948);
and U32646 (N_32646,N_31212,N_30487);
nor U32647 (N_32647,N_31723,N_30058);
or U32648 (N_32648,N_31232,N_31230);
xnor U32649 (N_32649,N_31315,N_30608);
xnor U32650 (N_32650,N_30631,N_31251);
and U32651 (N_32651,N_31292,N_31168);
nand U32652 (N_32652,N_30554,N_30911);
and U32653 (N_32653,N_31349,N_31395);
nor U32654 (N_32654,N_30464,N_30792);
xor U32655 (N_32655,N_30651,N_30129);
nand U32656 (N_32656,N_30797,N_31404);
and U32657 (N_32657,N_31183,N_31529);
and U32658 (N_32658,N_31733,N_31081);
nor U32659 (N_32659,N_30026,N_30027);
and U32660 (N_32660,N_30556,N_31982);
nor U32661 (N_32661,N_31123,N_31245);
nor U32662 (N_32662,N_31627,N_30090);
nand U32663 (N_32663,N_31202,N_30138);
nor U32664 (N_32664,N_31036,N_31626);
or U32665 (N_32665,N_31094,N_30763);
nor U32666 (N_32666,N_31471,N_31584);
and U32667 (N_32667,N_30166,N_31980);
nand U32668 (N_32668,N_31873,N_30354);
or U32669 (N_32669,N_31013,N_30327);
or U32670 (N_32670,N_31523,N_31002);
xor U32671 (N_32671,N_31610,N_30517);
nor U32672 (N_32672,N_30040,N_31446);
or U32673 (N_32673,N_30951,N_30947);
xor U32674 (N_32674,N_31564,N_30100);
nor U32675 (N_32675,N_30793,N_31498);
nor U32676 (N_32676,N_31481,N_31693);
or U32677 (N_32677,N_31197,N_31801);
nor U32678 (N_32678,N_30290,N_31269);
nand U32679 (N_32679,N_30476,N_30486);
or U32680 (N_32680,N_31753,N_30080);
nand U32681 (N_32681,N_30364,N_30431);
nand U32682 (N_32682,N_31713,N_30731);
or U32683 (N_32683,N_30274,N_31919);
and U32684 (N_32684,N_30575,N_30433);
nand U32685 (N_32685,N_30110,N_31321);
nand U32686 (N_32686,N_30806,N_30022);
or U32687 (N_32687,N_31397,N_30065);
nor U32688 (N_32688,N_31376,N_30197);
and U32689 (N_32689,N_30884,N_31048);
xor U32690 (N_32690,N_31882,N_31804);
nor U32691 (N_32691,N_30679,N_30170);
nor U32692 (N_32692,N_30082,N_31382);
or U32693 (N_32693,N_30038,N_30208);
or U32694 (N_32694,N_30876,N_30316);
and U32695 (N_32695,N_30540,N_30248);
or U32696 (N_32696,N_30347,N_31488);
or U32697 (N_32697,N_31608,N_31945);
xnor U32698 (N_32698,N_31827,N_30760);
and U32699 (N_32699,N_30857,N_31937);
nand U32700 (N_32700,N_31594,N_30420);
or U32701 (N_32701,N_31414,N_31793);
or U32702 (N_32702,N_31770,N_31542);
nand U32703 (N_32703,N_31294,N_31337);
nor U32704 (N_32704,N_31270,N_30292);
nand U32705 (N_32705,N_30771,N_31917);
and U32706 (N_32706,N_31521,N_31073);
xnor U32707 (N_32707,N_30235,N_30247);
and U32708 (N_32708,N_30372,N_31510);
nand U32709 (N_32709,N_30538,N_31257);
xor U32710 (N_32710,N_31367,N_30043);
nand U32711 (N_32711,N_30695,N_30820);
and U32712 (N_32712,N_31085,N_31103);
nand U32713 (N_32713,N_31607,N_31952);
and U32714 (N_32714,N_31661,N_31372);
xor U32715 (N_32715,N_30193,N_31637);
xor U32716 (N_32716,N_31720,N_30510);
or U32717 (N_32717,N_31786,N_30861);
and U32718 (N_32718,N_31055,N_31861);
and U32719 (N_32719,N_30665,N_30682);
or U32720 (N_32720,N_30366,N_30610);
nand U32721 (N_32721,N_30568,N_31599);
nand U32722 (N_32722,N_30207,N_30260);
nand U32723 (N_32723,N_31645,N_31425);
or U32724 (N_32724,N_30604,N_30592);
xnor U32725 (N_32725,N_31977,N_31532);
nor U32726 (N_32726,N_30969,N_31687);
and U32727 (N_32727,N_31879,N_31478);
xnor U32728 (N_32728,N_31405,N_30313);
or U32729 (N_32729,N_30269,N_31877);
or U32730 (N_32730,N_30777,N_31629);
nor U32731 (N_32731,N_30426,N_31905);
nand U32732 (N_32732,N_30564,N_31580);
and U32733 (N_32733,N_31900,N_30704);
xnor U32734 (N_32734,N_30258,N_30333);
and U32735 (N_32735,N_30006,N_30780);
or U32736 (N_32736,N_30140,N_30365);
nand U32737 (N_32737,N_30294,N_30057);
xnor U32738 (N_32738,N_31819,N_30620);
and U32739 (N_32739,N_31041,N_30452);
xnor U32740 (N_32740,N_31051,N_31511);
xor U32741 (N_32741,N_31972,N_31122);
nor U32742 (N_32742,N_30769,N_31708);
nand U32743 (N_32743,N_31009,N_31978);
nand U32744 (N_32744,N_31546,N_30828);
nor U32745 (N_32745,N_30286,N_31824);
and U32746 (N_32746,N_31323,N_30853);
or U32747 (N_32747,N_31001,N_31456);
or U32748 (N_32748,N_30291,N_30594);
nand U32749 (N_32749,N_30921,N_31694);
xnor U32750 (N_32750,N_30061,N_31509);
and U32751 (N_32751,N_31935,N_30767);
and U32752 (N_32752,N_30772,N_30441);
xor U32753 (N_32753,N_30199,N_31320);
and U32754 (N_32754,N_31386,N_30571);
or U32755 (N_32755,N_31586,N_31525);
or U32756 (N_32756,N_31563,N_31678);
nand U32757 (N_32757,N_31444,N_30851);
xnor U32758 (N_32758,N_31742,N_30944);
xnor U32759 (N_32759,N_30188,N_31340);
nand U32760 (N_32760,N_31735,N_30209);
and U32761 (N_32761,N_30864,N_30271);
or U32762 (N_32762,N_31174,N_31305);
or U32763 (N_32763,N_30469,N_30991);
and U32764 (N_32764,N_31930,N_31015);
and U32765 (N_32765,N_31396,N_31796);
nor U32766 (N_32766,N_31371,N_30482);
and U32767 (N_32767,N_31920,N_30326);
xnor U32768 (N_32768,N_30800,N_31684);
and U32769 (N_32769,N_31907,N_31268);
and U32770 (N_32770,N_31279,N_30541);
nand U32771 (N_32771,N_30531,N_31439);
nand U32772 (N_32772,N_30557,N_31361);
or U32773 (N_32773,N_31431,N_31646);
and U32774 (N_32774,N_30520,N_30737);
or U32775 (N_32775,N_31497,N_31651);
xnor U32776 (N_32776,N_30972,N_30905);
nor U32777 (N_32777,N_30398,N_30720);
nor U32778 (N_32778,N_30189,N_30637);
nand U32779 (N_32779,N_30926,N_31250);
xor U32780 (N_32780,N_31192,N_30439);
nor U32781 (N_32781,N_31849,N_31129);
nor U32782 (N_32782,N_31368,N_31283);
nand U32783 (N_32783,N_31653,N_30428);
xor U32784 (N_32784,N_31688,N_30691);
or U32785 (N_32785,N_31593,N_31253);
or U32786 (N_32786,N_31156,N_31737);
nand U32787 (N_32787,N_30749,N_30045);
and U32788 (N_32788,N_31700,N_31291);
nor U32789 (N_32789,N_31893,N_31549);
xor U32790 (N_32790,N_30267,N_31870);
nand U32791 (N_32791,N_30401,N_31696);
nand U32792 (N_32792,N_30847,N_31601);
and U32793 (N_32793,N_30445,N_30867);
nand U32794 (N_32794,N_31437,N_31416);
nor U32795 (N_32795,N_31413,N_30745);
or U32796 (N_32796,N_31730,N_30680);
or U32797 (N_32797,N_30545,N_31182);
nand U32798 (N_32798,N_30256,N_30535);
nand U32799 (N_32799,N_31561,N_31338);
nor U32800 (N_32800,N_30240,N_30075);
or U32801 (N_32801,N_30013,N_30168);
xor U32802 (N_32802,N_30624,N_31531);
xor U32803 (N_32803,N_31402,N_30674);
nand U32804 (N_32804,N_30139,N_30432);
nor U32805 (N_32805,N_30602,N_31654);
or U32806 (N_32806,N_30511,N_30083);
xnor U32807 (N_32807,N_31706,N_31252);
or U32808 (N_32808,N_31567,N_30182);
nand U32809 (N_32809,N_30216,N_31617);
nand U32810 (N_32810,N_30716,N_30234);
and U32811 (N_32811,N_31913,N_30092);
nand U32812 (N_32812,N_30103,N_31132);
xnor U32813 (N_32813,N_31597,N_31039);
xor U32814 (N_32814,N_31590,N_31569);
nor U32815 (N_32815,N_31923,N_30587);
nand U32816 (N_32816,N_31038,N_31835);
nor U32817 (N_32817,N_31220,N_31998);
nand U32818 (N_32818,N_30773,N_31078);
nand U32819 (N_32819,N_31421,N_30678);
nor U32820 (N_32820,N_30312,N_31691);
and U32821 (N_32821,N_30708,N_31958);
xnor U32822 (N_32822,N_30609,N_30599);
or U32823 (N_32823,N_31578,N_31373);
and U32824 (N_32824,N_31674,N_31494);
xnor U32825 (N_32825,N_31745,N_30618);
nand U32826 (N_32826,N_30787,N_30560);
and U32827 (N_32827,N_31734,N_31501);
nand U32828 (N_32828,N_31150,N_31616);
nand U32829 (N_32829,N_31355,N_31914);
and U32830 (N_32830,N_31327,N_30144);
nand U32831 (N_32831,N_31987,N_31365);
and U32832 (N_32832,N_30727,N_30358);
nor U32833 (N_32833,N_30254,N_31912);
nand U32834 (N_32834,N_31541,N_31050);
or U32835 (N_32835,N_31524,N_31547);
and U32836 (N_32836,N_30332,N_31249);
or U32837 (N_32837,N_30471,N_30033);
nor U32838 (N_32838,N_31803,N_31084);
and U32839 (N_32839,N_31207,N_31021);
and U32840 (N_32840,N_30869,N_31911);
nor U32841 (N_32841,N_31187,N_31302);
nand U32842 (N_32842,N_31024,N_31614);
xnor U32843 (N_32843,N_30488,N_30645);
and U32844 (N_32844,N_31452,N_30336);
nor U32845 (N_32845,N_31286,N_31976);
nor U32846 (N_32846,N_31301,N_30186);
or U32847 (N_32847,N_30815,N_30415);
xnor U32848 (N_32848,N_30430,N_31095);
nor U32849 (N_32849,N_31503,N_30097);
nand U32850 (N_32850,N_30971,N_31175);
or U32851 (N_32851,N_30661,N_31226);
and U32852 (N_32852,N_31551,N_31216);
nand U32853 (N_32853,N_30157,N_31134);
or U32854 (N_32854,N_30958,N_31897);
xor U32855 (N_32855,N_30766,N_31300);
or U32856 (N_32856,N_30562,N_31157);
and U32857 (N_32857,N_31034,N_30201);
and U32858 (N_32858,N_31725,N_30700);
or U32859 (N_32859,N_30728,N_31204);
and U32860 (N_32860,N_30337,N_30569);
nand U32861 (N_32861,N_30738,N_31059);
xnor U32862 (N_32862,N_31953,N_30619);
nand U32863 (N_32863,N_30883,N_31068);
nor U32864 (N_32864,N_31282,N_31842);
and U32865 (N_32865,N_30681,N_30387);
nand U32866 (N_32866,N_30677,N_30494);
or U32867 (N_32867,N_30009,N_31278);
nor U32868 (N_32868,N_30752,N_31261);
and U32869 (N_32869,N_30419,N_30580);
xnor U32870 (N_32870,N_30109,N_31056);
and U32871 (N_32871,N_30496,N_30379);
nand U32872 (N_32872,N_30305,N_31477);
and U32873 (N_32873,N_30507,N_31328);
xor U32874 (N_32874,N_31772,N_30226);
nor U32875 (N_32875,N_30107,N_31333);
xnor U32876 (N_32876,N_30503,N_31018);
and U32877 (N_32877,N_31176,N_30311);
and U32878 (N_32878,N_30779,N_31265);
xor U32879 (N_32879,N_31602,N_31326);
or U32880 (N_32880,N_31392,N_31992);
xnor U32881 (N_32881,N_31606,N_30613);
or U32882 (N_32882,N_31335,N_31631);
or U32883 (N_32883,N_31828,N_31941);
nand U32884 (N_32884,N_30213,N_30191);
nand U32885 (N_32885,N_30642,N_31406);
and U32886 (N_32886,N_30850,N_31679);
and U32887 (N_32887,N_31322,N_30035);
or U32888 (N_32888,N_31570,N_31193);
or U32889 (N_32889,N_30127,N_30658);
and U32890 (N_32890,N_30717,N_31875);
or U32891 (N_32891,N_30399,N_31527);
or U32892 (N_32892,N_30105,N_30049);
or U32893 (N_32893,N_31312,N_30340);
nor U32894 (N_32894,N_30036,N_30519);
and U32895 (N_32895,N_31766,N_31894);
nor U32896 (N_32896,N_31161,N_31141);
and U32897 (N_32897,N_30688,N_30397);
nor U32898 (N_32898,N_31005,N_31331);
and U32899 (N_32899,N_31990,N_30744);
nand U32900 (N_32900,N_30601,N_30904);
nor U32901 (N_32901,N_30108,N_31615);
or U32902 (N_32902,N_30570,N_31178);
or U32903 (N_32903,N_30357,N_31418);
or U32904 (N_32904,N_31185,N_30786);
nor U32905 (N_32905,N_31666,N_31885);
or U32906 (N_32906,N_31860,N_31407);
or U32907 (N_32907,N_30566,N_31600);
xor U32908 (N_32908,N_31778,N_31711);
xor U32909 (N_32909,N_30124,N_31151);
xnor U32910 (N_32910,N_31003,N_31044);
nor U32911 (N_32911,N_30579,N_30649);
nor U32912 (N_32912,N_30121,N_31077);
nor U32913 (N_32913,N_30394,N_30635);
nor U32914 (N_32914,N_31492,N_31927);
nor U32915 (N_32915,N_30617,N_31287);
nor U32916 (N_32916,N_30865,N_30585);
nor U32917 (N_32917,N_31513,N_31173);
nand U32918 (N_32918,N_31517,N_30238);
nand U32919 (N_32919,N_30837,N_31721);
xnor U32920 (N_32920,N_30694,N_30799);
xnor U32921 (N_32921,N_30069,N_31716);
or U32922 (N_32922,N_31304,N_30231);
and U32923 (N_32923,N_30761,N_31432);
or U32924 (N_32924,N_31784,N_30783);
nand U32925 (N_32925,N_31664,N_31350);
nand U32926 (N_32926,N_30218,N_31677);
nor U32927 (N_32927,N_30935,N_31782);
nor U32928 (N_32928,N_31535,N_31058);
nand U32929 (N_32929,N_30723,N_31697);
xnor U32930 (N_32930,N_31487,N_30125);
or U32931 (N_32931,N_31063,N_31343);
nor U32932 (N_32932,N_31758,N_31353);
or U32933 (N_32933,N_30074,N_31638);
nand U32934 (N_32934,N_30729,N_30003);
xor U32935 (N_32935,N_30937,N_31153);
nand U32936 (N_32936,N_31243,N_31228);
nand U32937 (N_32937,N_31217,N_31817);
nor U32938 (N_32938,N_30343,N_30670);
nor U32939 (N_32939,N_31783,N_31743);
xnor U32940 (N_32940,N_31552,N_30814);
xor U32941 (N_32941,N_31006,N_31258);
and U32942 (N_32942,N_30634,N_31307);
or U32943 (N_32943,N_31388,N_30532);
or U32944 (N_32944,N_30537,N_30156);
or U32945 (N_32945,N_31898,N_31473);
nand U32946 (N_32946,N_31083,N_30434);
nand U32947 (N_32947,N_30338,N_31731);
or U32948 (N_32948,N_31131,N_30195);
and U32949 (N_32949,N_31884,N_31004);
nor U32950 (N_32950,N_30558,N_30818);
and U32951 (N_32951,N_31806,N_30834);
nor U32952 (N_32952,N_30802,N_31855);
or U32953 (N_32953,N_30666,N_31167);
nor U32954 (N_32954,N_30955,N_30066);
nor U32955 (N_32955,N_30706,N_30042);
nor U32956 (N_32956,N_31851,N_30423);
nand U32957 (N_32957,N_31997,N_30371);
nand U32958 (N_32958,N_31577,N_31113);
and U32959 (N_32959,N_31271,N_30740);
or U32960 (N_32960,N_31114,N_31383);
xnor U32961 (N_32961,N_30220,N_31670);
and U32962 (N_32962,N_31754,N_31453);
xor U32963 (N_32963,N_31774,N_30377);
and U32964 (N_32964,N_30349,N_31008);
nand U32965 (N_32965,N_30277,N_30776);
and U32966 (N_32966,N_30382,N_30755);
nor U32967 (N_32967,N_31609,N_31749);
nor U32968 (N_32968,N_31565,N_31798);
xor U32969 (N_32969,N_31112,N_30879);
and U32970 (N_32970,N_30284,N_30768);
nand U32971 (N_32971,N_31071,N_30630);
and U32972 (N_32972,N_31109,N_31964);
nand U32973 (N_32973,N_31815,N_31832);
or U32974 (N_32974,N_31164,N_30576);
and U32975 (N_32975,N_31146,N_31543);
xor U32976 (N_32976,N_31993,N_30892);
nand U32977 (N_32977,N_31710,N_30713);
xor U32978 (N_32978,N_30385,N_30819);
or U32979 (N_32979,N_31641,N_31420);
xnor U32980 (N_32980,N_31467,N_31360);
nand U32981 (N_32981,N_31022,N_31773);
nor U32982 (N_32982,N_30443,N_31566);
or U32983 (N_32983,N_30595,N_31325);
or U32984 (N_32984,N_31890,N_30606);
xnor U32985 (N_32985,N_30473,N_31619);
and U32986 (N_32986,N_31620,N_30257);
or U32987 (N_32987,N_31357,N_31869);
and U32988 (N_32988,N_31241,N_30781);
or U32989 (N_32989,N_31689,N_30553);
and U32990 (N_32990,N_31136,N_30547);
nor U32991 (N_32991,N_31017,N_31695);
nor U32992 (N_32992,N_30279,N_31767);
nor U32993 (N_32993,N_30518,N_30539);
or U32994 (N_32994,N_30244,N_31080);
or U32995 (N_32995,N_31636,N_30463);
nor U32996 (N_32996,N_30842,N_31154);
or U32997 (N_32997,N_30962,N_30468);
or U32998 (N_32998,N_31138,N_30493);
and U32999 (N_32999,N_30458,N_30211);
xor U33000 (N_33000,N_30357,N_31512);
nand U33001 (N_33001,N_31637,N_31793);
and U33002 (N_33002,N_30139,N_30413);
nand U33003 (N_33003,N_30746,N_31130);
and U33004 (N_33004,N_31606,N_30731);
and U33005 (N_33005,N_31406,N_30921);
or U33006 (N_33006,N_31779,N_31067);
and U33007 (N_33007,N_30840,N_30518);
and U33008 (N_33008,N_30375,N_30968);
nand U33009 (N_33009,N_31563,N_30728);
and U33010 (N_33010,N_30872,N_31945);
and U33011 (N_33011,N_30499,N_31656);
nor U33012 (N_33012,N_30154,N_30518);
xnor U33013 (N_33013,N_31896,N_30145);
and U33014 (N_33014,N_31958,N_31372);
and U33015 (N_33015,N_30212,N_31457);
nor U33016 (N_33016,N_30281,N_30298);
nand U33017 (N_33017,N_31554,N_31926);
and U33018 (N_33018,N_30436,N_30439);
nor U33019 (N_33019,N_30649,N_31354);
nor U33020 (N_33020,N_31467,N_30563);
nor U33021 (N_33021,N_31687,N_30018);
or U33022 (N_33022,N_31592,N_31151);
xor U33023 (N_33023,N_31864,N_30733);
and U33024 (N_33024,N_31200,N_30543);
xor U33025 (N_33025,N_31819,N_31202);
xnor U33026 (N_33026,N_30018,N_31547);
or U33027 (N_33027,N_31171,N_31873);
nor U33028 (N_33028,N_30875,N_31399);
or U33029 (N_33029,N_30331,N_30074);
nor U33030 (N_33030,N_31069,N_31887);
or U33031 (N_33031,N_31071,N_30003);
nand U33032 (N_33032,N_30358,N_31530);
nand U33033 (N_33033,N_30248,N_31820);
and U33034 (N_33034,N_30525,N_30125);
nand U33035 (N_33035,N_30274,N_30786);
or U33036 (N_33036,N_31483,N_31738);
xor U33037 (N_33037,N_31926,N_31937);
nor U33038 (N_33038,N_30166,N_31134);
and U33039 (N_33039,N_30143,N_30945);
nor U33040 (N_33040,N_31995,N_30411);
xnor U33041 (N_33041,N_30253,N_30125);
nand U33042 (N_33042,N_31405,N_31104);
xnor U33043 (N_33043,N_31192,N_30273);
and U33044 (N_33044,N_31710,N_30219);
nand U33045 (N_33045,N_31657,N_31550);
and U33046 (N_33046,N_30217,N_30146);
xnor U33047 (N_33047,N_31002,N_31439);
xor U33048 (N_33048,N_30340,N_30982);
or U33049 (N_33049,N_31664,N_31939);
nor U33050 (N_33050,N_30737,N_31130);
or U33051 (N_33051,N_30416,N_30248);
nor U33052 (N_33052,N_30640,N_31932);
or U33053 (N_33053,N_31006,N_30733);
nor U33054 (N_33054,N_31349,N_30955);
and U33055 (N_33055,N_31699,N_31641);
nand U33056 (N_33056,N_31866,N_30383);
xor U33057 (N_33057,N_30024,N_30250);
nor U33058 (N_33058,N_30503,N_30788);
xor U33059 (N_33059,N_30619,N_30260);
xor U33060 (N_33060,N_30536,N_30788);
and U33061 (N_33061,N_30390,N_31411);
and U33062 (N_33062,N_31581,N_30557);
or U33063 (N_33063,N_30718,N_30781);
or U33064 (N_33064,N_30929,N_30049);
xor U33065 (N_33065,N_31818,N_30812);
nand U33066 (N_33066,N_30270,N_30959);
and U33067 (N_33067,N_31997,N_31078);
nor U33068 (N_33068,N_30433,N_30579);
or U33069 (N_33069,N_30021,N_31412);
xnor U33070 (N_33070,N_30331,N_31852);
or U33071 (N_33071,N_30971,N_31879);
nor U33072 (N_33072,N_31010,N_30305);
nand U33073 (N_33073,N_31388,N_31532);
or U33074 (N_33074,N_31637,N_30271);
or U33075 (N_33075,N_31735,N_31219);
and U33076 (N_33076,N_31625,N_31882);
or U33077 (N_33077,N_30759,N_31936);
xor U33078 (N_33078,N_31853,N_30819);
or U33079 (N_33079,N_31257,N_31946);
xnor U33080 (N_33080,N_30363,N_31490);
or U33081 (N_33081,N_31267,N_31983);
xnor U33082 (N_33082,N_31056,N_31896);
or U33083 (N_33083,N_30404,N_30234);
nor U33084 (N_33084,N_30975,N_31966);
xnor U33085 (N_33085,N_31330,N_30098);
nand U33086 (N_33086,N_30764,N_31074);
xnor U33087 (N_33087,N_30709,N_30950);
nand U33088 (N_33088,N_30940,N_30539);
nand U33089 (N_33089,N_31068,N_31991);
xnor U33090 (N_33090,N_31366,N_30510);
or U33091 (N_33091,N_31845,N_31366);
or U33092 (N_33092,N_30249,N_31822);
nor U33093 (N_33093,N_31499,N_30975);
xor U33094 (N_33094,N_31707,N_31275);
nor U33095 (N_33095,N_31890,N_30505);
nor U33096 (N_33096,N_30070,N_31434);
xnor U33097 (N_33097,N_31673,N_31159);
nand U33098 (N_33098,N_31833,N_31757);
nor U33099 (N_33099,N_31647,N_30462);
or U33100 (N_33100,N_30913,N_30015);
nor U33101 (N_33101,N_31514,N_31155);
nor U33102 (N_33102,N_31493,N_31813);
nand U33103 (N_33103,N_30180,N_30979);
nor U33104 (N_33104,N_30495,N_30651);
and U33105 (N_33105,N_31127,N_31564);
and U33106 (N_33106,N_31417,N_31957);
or U33107 (N_33107,N_30704,N_30743);
and U33108 (N_33108,N_30040,N_31038);
and U33109 (N_33109,N_31955,N_31416);
or U33110 (N_33110,N_31467,N_30998);
and U33111 (N_33111,N_31348,N_31861);
and U33112 (N_33112,N_30770,N_30424);
and U33113 (N_33113,N_31438,N_30536);
or U33114 (N_33114,N_30854,N_31560);
xnor U33115 (N_33115,N_30566,N_31755);
xnor U33116 (N_33116,N_30683,N_31785);
and U33117 (N_33117,N_30956,N_30414);
and U33118 (N_33118,N_31836,N_31379);
or U33119 (N_33119,N_31626,N_31375);
nand U33120 (N_33120,N_31348,N_31727);
nand U33121 (N_33121,N_30519,N_31866);
xor U33122 (N_33122,N_31203,N_30196);
and U33123 (N_33123,N_30061,N_30611);
nand U33124 (N_33124,N_30981,N_30447);
or U33125 (N_33125,N_31897,N_31484);
nor U33126 (N_33126,N_31876,N_31764);
or U33127 (N_33127,N_30273,N_30214);
nor U33128 (N_33128,N_31912,N_30902);
nand U33129 (N_33129,N_30614,N_31526);
nand U33130 (N_33130,N_30851,N_31986);
or U33131 (N_33131,N_31171,N_31448);
nand U33132 (N_33132,N_30701,N_30385);
or U33133 (N_33133,N_31626,N_30969);
nor U33134 (N_33134,N_31903,N_30134);
xor U33135 (N_33135,N_30144,N_30735);
nor U33136 (N_33136,N_30303,N_30863);
and U33137 (N_33137,N_31724,N_30627);
xnor U33138 (N_33138,N_31089,N_30687);
or U33139 (N_33139,N_30804,N_30597);
xor U33140 (N_33140,N_30367,N_31834);
xnor U33141 (N_33141,N_31900,N_30883);
nand U33142 (N_33142,N_31445,N_30410);
and U33143 (N_33143,N_30217,N_31977);
or U33144 (N_33144,N_30526,N_31653);
xor U33145 (N_33145,N_30777,N_30513);
nor U33146 (N_33146,N_30202,N_30758);
nand U33147 (N_33147,N_30701,N_31887);
nor U33148 (N_33148,N_30364,N_31032);
or U33149 (N_33149,N_30959,N_30140);
and U33150 (N_33150,N_31858,N_30949);
nand U33151 (N_33151,N_31444,N_31744);
and U33152 (N_33152,N_31437,N_31973);
or U33153 (N_33153,N_30606,N_30921);
xnor U33154 (N_33154,N_31536,N_31307);
xnor U33155 (N_33155,N_31325,N_30357);
xnor U33156 (N_33156,N_30463,N_30947);
and U33157 (N_33157,N_30753,N_31543);
nand U33158 (N_33158,N_30118,N_30796);
or U33159 (N_33159,N_31278,N_31580);
xor U33160 (N_33160,N_30887,N_30014);
nand U33161 (N_33161,N_31386,N_31145);
and U33162 (N_33162,N_30702,N_31213);
and U33163 (N_33163,N_31685,N_30109);
nand U33164 (N_33164,N_31006,N_31595);
nand U33165 (N_33165,N_31607,N_31089);
xor U33166 (N_33166,N_31074,N_30811);
nor U33167 (N_33167,N_31649,N_30349);
nor U33168 (N_33168,N_31100,N_31055);
and U33169 (N_33169,N_31517,N_30646);
nor U33170 (N_33170,N_30967,N_31654);
or U33171 (N_33171,N_31009,N_30770);
and U33172 (N_33172,N_31107,N_30569);
xnor U33173 (N_33173,N_30977,N_31207);
nand U33174 (N_33174,N_31713,N_31411);
or U33175 (N_33175,N_30003,N_31842);
nor U33176 (N_33176,N_31183,N_30377);
nand U33177 (N_33177,N_30010,N_30004);
or U33178 (N_33178,N_31456,N_31393);
and U33179 (N_33179,N_30128,N_30924);
nand U33180 (N_33180,N_30338,N_30373);
and U33181 (N_33181,N_31677,N_31948);
xor U33182 (N_33182,N_31449,N_31030);
nor U33183 (N_33183,N_30262,N_30000);
or U33184 (N_33184,N_31243,N_30605);
nand U33185 (N_33185,N_31628,N_31168);
xor U33186 (N_33186,N_30723,N_30169);
nor U33187 (N_33187,N_30723,N_31392);
and U33188 (N_33188,N_31414,N_31574);
and U33189 (N_33189,N_30745,N_30813);
nor U33190 (N_33190,N_31892,N_31960);
xor U33191 (N_33191,N_30754,N_30203);
nor U33192 (N_33192,N_31400,N_30710);
or U33193 (N_33193,N_30297,N_31622);
or U33194 (N_33194,N_30121,N_30879);
and U33195 (N_33195,N_30092,N_30036);
nor U33196 (N_33196,N_30313,N_31415);
or U33197 (N_33197,N_31784,N_30994);
nor U33198 (N_33198,N_31575,N_30262);
nor U33199 (N_33199,N_30721,N_31669);
xor U33200 (N_33200,N_30967,N_31011);
nand U33201 (N_33201,N_30600,N_30089);
nor U33202 (N_33202,N_30365,N_30195);
or U33203 (N_33203,N_30459,N_31443);
and U33204 (N_33204,N_30886,N_31857);
or U33205 (N_33205,N_30524,N_30669);
nand U33206 (N_33206,N_30634,N_31093);
and U33207 (N_33207,N_31188,N_30757);
or U33208 (N_33208,N_31729,N_30580);
nor U33209 (N_33209,N_31880,N_30077);
nand U33210 (N_33210,N_31408,N_31223);
nand U33211 (N_33211,N_31972,N_31055);
nor U33212 (N_33212,N_31707,N_31272);
nor U33213 (N_33213,N_30147,N_31531);
or U33214 (N_33214,N_30074,N_31799);
nand U33215 (N_33215,N_30342,N_31852);
nor U33216 (N_33216,N_30949,N_30521);
or U33217 (N_33217,N_31962,N_30488);
or U33218 (N_33218,N_30694,N_31923);
nor U33219 (N_33219,N_31677,N_31333);
xnor U33220 (N_33220,N_30810,N_31254);
xnor U33221 (N_33221,N_30166,N_30812);
or U33222 (N_33222,N_30660,N_30865);
nand U33223 (N_33223,N_30708,N_30866);
nor U33224 (N_33224,N_30319,N_30196);
or U33225 (N_33225,N_31399,N_31287);
and U33226 (N_33226,N_31850,N_30271);
xnor U33227 (N_33227,N_30095,N_30662);
nor U33228 (N_33228,N_31381,N_31911);
or U33229 (N_33229,N_30350,N_30037);
nand U33230 (N_33230,N_31249,N_31594);
and U33231 (N_33231,N_31566,N_30535);
and U33232 (N_33232,N_30020,N_31617);
nor U33233 (N_33233,N_30421,N_31430);
or U33234 (N_33234,N_31801,N_30797);
nor U33235 (N_33235,N_30189,N_30164);
or U33236 (N_33236,N_31420,N_30974);
nand U33237 (N_33237,N_31887,N_31399);
nor U33238 (N_33238,N_30929,N_31818);
or U33239 (N_33239,N_30227,N_30083);
or U33240 (N_33240,N_31549,N_30888);
and U33241 (N_33241,N_31593,N_31553);
nand U33242 (N_33242,N_30237,N_30783);
or U33243 (N_33243,N_31182,N_30057);
nand U33244 (N_33244,N_30610,N_30155);
nor U33245 (N_33245,N_31203,N_31602);
or U33246 (N_33246,N_31493,N_30311);
nor U33247 (N_33247,N_30997,N_31594);
nand U33248 (N_33248,N_30989,N_31169);
and U33249 (N_33249,N_30653,N_30009);
and U33250 (N_33250,N_30918,N_30950);
nand U33251 (N_33251,N_30115,N_30375);
xnor U33252 (N_33252,N_31488,N_31419);
and U33253 (N_33253,N_31685,N_31645);
nand U33254 (N_33254,N_30824,N_30543);
and U33255 (N_33255,N_31875,N_31306);
and U33256 (N_33256,N_30673,N_31906);
and U33257 (N_33257,N_31672,N_30996);
or U33258 (N_33258,N_31694,N_31246);
xor U33259 (N_33259,N_31830,N_30682);
or U33260 (N_33260,N_31930,N_31024);
xor U33261 (N_33261,N_30164,N_30204);
nand U33262 (N_33262,N_30390,N_30546);
xor U33263 (N_33263,N_30884,N_30171);
and U33264 (N_33264,N_31526,N_31832);
and U33265 (N_33265,N_30471,N_30734);
nor U33266 (N_33266,N_30344,N_31237);
nor U33267 (N_33267,N_30550,N_30912);
or U33268 (N_33268,N_31049,N_30179);
nor U33269 (N_33269,N_30246,N_30747);
xor U33270 (N_33270,N_30747,N_31517);
nor U33271 (N_33271,N_30891,N_30914);
and U33272 (N_33272,N_31784,N_30558);
and U33273 (N_33273,N_31108,N_30072);
nand U33274 (N_33274,N_30782,N_30288);
xor U33275 (N_33275,N_31146,N_31539);
nor U33276 (N_33276,N_30180,N_30310);
nand U33277 (N_33277,N_31431,N_30265);
or U33278 (N_33278,N_31096,N_30786);
nand U33279 (N_33279,N_30644,N_30050);
or U33280 (N_33280,N_30814,N_30499);
or U33281 (N_33281,N_30614,N_31358);
xor U33282 (N_33282,N_30020,N_31078);
xor U33283 (N_33283,N_30269,N_31741);
xnor U33284 (N_33284,N_30133,N_31140);
nand U33285 (N_33285,N_30575,N_30309);
nand U33286 (N_33286,N_31703,N_30891);
and U33287 (N_33287,N_30309,N_31159);
nand U33288 (N_33288,N_30175,N_31820);
or U33289 (N_33289,N_31775,N_31042);
nor U33290 (N_33290,N_30587,N_30056);
nor U33291 (N_33291,N_31179,N_31950);
and U33292 (N_33292,N_30143,N_31335);
or U33293 (N_33293,N_30104,N_30574);
xor U33294 (N_33294,N_31541,N_30679);
xnor U33295 (N_33295,N_31877,N_31750);
xor U33296 (N_33296,N_30935,N_31624);
and U33297 (N_33297,N_31973,N_31591);
nor U33298 (N_33298,N_31371,N_31443);
nand U33299 (N_33299,N_31992,N_31441);
xnor U33300 (N_33300,N_30616,N_31724);
nand U33301 (N_33301,N_30512,N_31883);
xnor U33302 (N_33302,N_30049,N_30252);
nand U33303 (N_33303,N_30007,N_31832);
nand U33304 (N_33304,N_31123,N_31920);
nor U33305 (N_33305,N_31233,N_30273);
xnor U33306 (N_33306,N_30971,N_30748);
and U33307 (N_33307,N_31352,N_31780);
nor U33308 (N_33308,N_30970,N_30385);
and U33309 (N_33309,N_31602,N_31475);
or U33310 (N_33310,N_31453,N_30146);
nand U33311 (N_33311,N_31481,N_30476);
nand U33312 (N_33312,N_31898,N_30984);
nor U33313 (N_33313,N_31072,N_31966);
nand U33314 (N_33314,N_30491,N_30729);
and U33315 (N_33315,N_31668,N_31866);
nor U33316 (N_33316,N_30790,N_31863);
xor U33317 (N_33317,N_30333,N_30723);
nor U33318 (N_33318,N_31208,N_31413);
or U33319 (N_33319,N_31928,N_31337);
xor U33320 (N_33320,N_30175,N_30763);
xnor U33321 (N_33321,N_30767,N_30397);
nand U33322 (N_33322,N_31614,N_30851);
and U33323 (N_33323,N_30468,N_31918);
nand U33324 (N_33324,N_31570,N_30780);
nand U33325 (N_33325,N_31773,N_30323);
xor U33326 (N_33326,N_31092,N_31936);
or U33327 (N_33327,N_31384,N_30966);
xnor U33328 (N_33328,N_31422,N_30224);
and U33329 (N_33329,N_30177,N_30602);
and U33330 (N_33330,N_31075,N_30441);
nor U33331 (N_33331,N_31523,N_30929);
xnor U33332 (N_33332,N_30269,N_30117);
xnor U33333 (N_33333,N_31259,N_31274);
or U33334 (N_33334,N_30902,N_30263);
xor U33335 (N_33335,N_31195,N_31872);
nor U33336 (N_33336,N_30894,N_30079);
xnor U33337 (N_33337,N_31840,N_30946);
xor U33338 (N_33338,N_30764,N_31257);
nor U33339 (N_33339,N_31574,N_30203);
xor U33340 (N_33340,N_31866,N_31985);
and U33341 (N_33341,N_31856,N_31059);
nand U33342 (N_33342,N_30823,N_31153);
nand U33343 (N_33343,N_30120,N_30123);
and U33344 (N_33344,N_30066,N_31360);
nand U33345 (N_33345,N_30727,N_31329);
xor U33346 (N_33346,N_31210,N_30725);
or U33347 (N_33347,N_31651,N_30351);
and U33348 (N_33348,N_31073,N_31319);
and U33349 (N_33349,N_30274,N_30788);
xor U33350 (N_33350,N_30769,N_30690);
and U33351 (N_33351,N_31732,N_30728);
or U33352 (N_33352,N_31556,N_31648);
nand U33353 (N_33353,N_30744,N_30720);
xnor U33354 (N_33354,N_31122,N_30348);
or U33355 (N_33355,N_31204,N_31120);
nor U33356 (N_33356,N_30571,N_30230);
or U33357 (N_33357,N_30192,N_31538);
or U33358 (N_33358,N_31051,N_30595);
nand U33359 (N_33359,N_31050,N_30361);
nand U33360 (N_33360,N_31836,N_30503);
nor U33361 (N_33361,N_31839,N_30735);
nor U33362 (N_33362,N_31257,N_30045);
and U33363 (N_33363,N_30689,N_31100);
nand U33364 (N_33364,N_31739,N_30505);
nor U33365 (N_33365,N_30443,N_30296);
or U33366 (N_33366,N_30054,N_30253);
xor U33367 (N_33367,N_30824,N_31535);
xor U33368 (N_33368,N_31772,N_31023);
xor U33369 (N_33369,N_31774,N_30745);
and U33370 (N_33370,N_31591,N_31835);
xor U33371 (N_33371,N_30514,N_31072);
and U33372 (N_33372,N_31658,N_30663);
xnor U33373 (N_33373,N_30314,N_30758);
and U33374 (N_33374,N_31850,N_30201);
or U33375 (N_33375,N_30082,N_30386);
nor U33376 (N_33376,N_30503,N_30904);
nand U33377 (N_33377,N_31760,N_31977);
nand U33378 (N_33378,N_30783,N_30914);
nor U33379 (N_33379,N_30196,N_31572);
nand U33380 (N_33380,N_31154,N_31204);
and U33381 (N_33381,N_30926,N_30156);
nand U33382 (N_33382,N_30571,N_31655);
xnor U33383 (N_33383,N_30528,N_30818);
xnor U33384 (N_33384,N_31016,N_31655);
nor U33385 (N_33385,N_31698,N_31445);
or U33386 (N_33386,N_30710,N_30040);
xnor U33387 (N_33387,N_30555,N_31171);
nand U33388 (N_33388,N_31940,N_31784);
xnor U33389 (N_33389,N_31259,N_31075);
nand U33390 (N_33390,N_31119,N_30683);
nand U33391 (N_33391,N_30568,N_31047);
and U33392 (N_33392,N_31082,N_31940);
or U33393 (N_33393,N_30906,N_31721);
and U33394 (N_33394,N_30082,N_31515);
or U33395 (N_33395,N_30300,N_31982);
xor U33396 (N_33396,N_31219,N_30086);
nor U33397 (N_33397,N_31818,N_31791);
nand U33398 (N_33398,N_31513,N_30564);
and U33399 (N_33399,N_31703,N_30320);
and U33400 (N_33400,N_30588,N_30484);
and U33401 (N_33401,N_30799,N_31990);
or U33402 (N_33402,N_31568,N_31903);
and U33403 (N_33403,N_30404,N_30033);
or U33404 (N_33404,N_30441,N_31277);
and U33405 (N_33405,N_30063,N_31528);
nor U33406 (N_33406,N_31808,N_31735);
nand U33407 (N_33407,N_30490,N_30794);
xor U33408 (N_33408,N_31030,N_31256);
and U33409 (N_33409,N_30233,N_30936);
xnor U33410 (N_33410,N_31356,N_30865);
nor U33411 (N_33411,N_30008,N_31300);
or U33412 (N_33412,N_31872,N_31450);
or U33413 (N_33413,N_31631,N_31903);
and U33414 (N_33414,N_30416,N_30216);
nor U33415 (N_33415,N_31937,N_30828);
and U33416 (N_33416,N_30485,N_31259);
or U33417 (N_33417,N_30719,N_30342);
nand U33418 (N_33418,N_31942,N_30693);
xor U33419 (N_33419,N_30929,N_30297);
nor U33420 (N_33420,N_30602,N_31052);
xor U33421 (N_33421,N_30816,N_31620);
xnor U33422 (N_33422,N_31582,N_30755);
or U33423 (N_33423,N_30942,N_30871);
or U33424 (N_33424,N_30119,N_30983);
or U33425 (N_33425,N_31451,N_30971);
nor U33426 (N_33426,N_31946,N_30300);
and U33427 (N_33427,N_30583,N_31680);
nand U33428 (N_33428,N_31371,N_30646);
or U33429 (N_33429,N_30372,N_30875);
and U33430 (N_33430,N_31393,N_31413);
and U33431 (N_33431,N_31889,N_30608);
nand U33432 (N_33432,N_31553,N_30600);
xnor U33433 (N_33433,N_30099,N_31645);
or U33434 (N_33434,N_30309,N_31047);
nand U33435 (N_33435,N_30787,N_30031);
nor U33436 (N_33436,N_30282,N_31899);
nor U33437 (N_33437,N_31512,N_30966);
nor U33438 (N_33438,N_31709,N_31377);
and U33439 (N_33439,N_30875,N_30907);
or U33440 (N_33440,N_31499,N_31304);
and U33441 (N_33441,N_30684,N_31986);
xnor U33442 (N_33442,N_31915,N_31679);
or U33443 (N_33443,N_30787,N_30433);
and U33444 (N_33444,N_31993,N_30867);
or U33445 (N_33445,N_30439,N_31521);
or U33446 (N_33446,N_31316,N_31701);
and U33447 (N_33447,N_31163,N_30058);
and U33448 (N_33448,N_31845,N_31675);
xor U33449 (N_33449,N_30410,N_31841);
or U33450 (N_33450,N_31788,N_30299);
and U33451 (N_33451,N_31862,N_30260);
and U33452 (N_33452,N_30875,N_31588);
and U33453 (N_33453,N_31462,N_30598);
xor U33454 (N_33454,N_30977,N_31345);
or U33455 (N_33455,N_31011,N_30954);
xnor U33456 (N_33456,N_31435,N_31323);
and U33457 (N_33457,N_31854,N_30190);
or U33458 (N_33458,N_31560,N_30778);
and U33459 (N_33459,N_31047,N_30234);
and U33460 (N_33460,N_30496,N_30564);
and U33461 (N_33461,N_30470,N_31388);
nor U33462 (N_33462,N_30878,N_31720);
nor U33463 (N_33463,N_30611,N_30984);
nand U33464 (N_33464,N_31996,N_31968);
or U33465 (N_33465,N_30162,N_30134);
or U33466 (N_33466,N_31539,N_31516);
nand U33467 (N_33467,N_31512,N_31200);
nand U33468 (N_33468,N_31352,N_31235);
or U33469 (N_33469,N_30381,N_31972);
or U33470 (N_33470,N_30814,N_31233);
or U33471 (N_33471,N_31598,N_30667);
nand U33472 (N_33472,N_31499,N_30595);
nand U33473 (N_33473,N_30179,N_31622);
nor U33474 (N_33474,N_31376,N_30395);
nand U33475 (N_33475,N_30386,N_31490);
nor U33476 (N_33476,N_31039,N_31398);
and U33477 (N_33477,N_30380,N_30839);
xnor U33478 (N_33478,N_31927,N_30076);
nand U33479 (N_33479,N_31130,N_30145);
and U33480 (N_33480,N_31408,N_30256);
and U33481 (N_33481,N_30818,N_30542);
nor U33482 (N_33482,N_30468,N_31563);
or U33483 (N_33483,N_30745,N_30259);
nor U33484 (N_33484,N_30610,N_31435);
nand U33485 (N_33485,N_30532,N_30828);
and U33486 (N_33486,N_31238,N_31566);
nor U33487 (N_33487,N_30045,N_30911);
or U33488 (N_33488,N_31091,N_31233);
xnor U33489 (N_33489,N_30668,N_31364);
or U33490 (N_33490,N_30171,N_31957);
xnor U33491 (N_33491,N_31073,N_31530);
nor U33492 (N_33492,N_31164,N_30036);
and U33493 (N_33493,N_31050,N_31011);
xor U33494 (N_33494,N_30940,N_30469);
nand U33495 (N_33495,N_30828,N_30470);
nor U33496 (N_33496,N_31928,N_31894);
or U33497 (N_33497,N_31734,N_31304);
or U33498 (N_33498,N_30780,N_31048);
xnor U33499 (N_33499,N_31130,N_30005);
nand U33500 (N_33500,N_30413,N_31342);
and U33501 (N_33501,N_31274,N_30731);
xor U33502 (N_33502,N_30159,N_31739);
and U33503 (N_33503,N_30192,N_30833);
or U33504 (N_33504,N_31787,N_31355);
nand U33505 (N_33505,N_30577,N_30516);
and U33506 (N_33506,N_31704,N_31609);
or U33507 (N_33507,N_30876,N_30487);
nand U33508 (N_33508,N_30579,N_30693);
and U33509 (N_33509,N_31132,N_31342);
or U33510 (N_33510,N_30151,N_30704);
nor U33511 (N_33511,N_30113,N_30102);
xnor U33512 (N_33512,N_31835,N_30018);
nor U33513 (N_33513,N_31483,N_30358);
nor U33514 (N_33514,N_30603,N_30801);
or U33515 (N_33515,N_31376,N_30700);
nor U33516 (N_33516,N_31952,N_31439);
xnor U33517 (N_33517,N_30512,N_30346);
nor U33518 (N_33518,N_30064,N_30188);
or U33519 (N_33519,N_30298,N_31718);
or U33520 (N_33520,N_30024,N_31104);
nand U33521 (N_33521,N_30263,N_31502);
nand U33522 (N_33522,N_30524,N_31771);
nand U33523 (N_33523,N_31059,N_31880);
and U33524 (N_33524,N_30113,N_31019);
or U33525 (N_33525,N_31763,N_31548);
xor U33526 (N_33526,N_31762,N_31713);
nor U33527 (N_33527,N_30075,N_30472);
xor U33528 (N_33528,N_31403,N_31707);
or U33529 (N_33529,N_30817,N_31816);
xor U33530 (N_33530,N_31955,N_31968);
or U33531 (N_33531,N_30140,N_31380);
nor U33532 (N_33532,N_31688,N_31171);
or U33533 (N_33533,N_30934,N_31103);
nand U33534 (N_33534,N_30453,N_30567);
and U33535 (N_33535,N_31809,N_30978);
or U33536 (N_33536,N_31612,N_31680);
and U33537 (N_33537,N_31423,N_31611);
nor U33538 (N_33538,N_31291,N_31979);
and U33539 (N_33539,N_31178,N_31597);
or U33540 (N_33540,N_30900,N_31191);
or U33541 (N_33541,N_30256,N_30438);
nor U33542 (N_33542,N_31335,N_31862);
nor U33543 (N_33543,N_31206,N_30553);
xnor U33544 (N_33544,N_30815,N_31413);
nor U33545 (N_33545,N_31626,N_31462);
or U33546 (N_33546,N_30203,N_30417);
and U33547 (N_33547,N_30831,N_31415);
nand U33548 (N_33548,N_31243,N_30186);
nand U33549 (N_33549,N_31039,N_30078);
nor U33550 (N_33550,N_30543,N_31773);
or U33551 (N_33551,N_31352,N_30842);
nand U33552 (N_33552,N_30696,N_31106);
nand U33553 (N_33553,N_31606,N_31533);
nand U33554 (N_33554,N_30837,N_31172);
or U33555 (N_33555,N_31722,N_31067);
and U33556 (N_33556,N_31380,N_31845);
xnor U33557 (N_33557,N_31438,N_30527);
and U33558 (N_33558,N_30821,N_30063);
nand U33559 (N_33559,N_31404,N_31658);
xnor U33560 (N_33560,N_31655,N_30103);
nor U33561 (N_33561,N_30350,N_31621);
nor U33562 (N_33562,N_30898,N_30144);
nand U33563 (N_33563,N_31902,N_31571);
xnor U33564 (N_33564,N_30586,N_30868);
nand U33565 (N_33565,N_30436,N_31211);
and U33566 (N_33566,N_31369,N_30917);
nand U33567 (N_33567,N_30914,N_30341);
and U33568 (N_33568,N_31922,N_30244);
xnor U33569 (N_33569,N_30177,N_30760);
and U33570 (N_33570,N_30400,N_30450);
and U33571 (N_33571,N_30775,N_31687);
nand U33572 (N_33572,N_30709,N_30107);
xnor U33573 (N_33573,N_31959,N_31418);
nor U33574 (N_33574,N_31789,N_31087);
or U33575 (N_33575,N_31765,N_30733);
xnor U33576 (N_33576,N_30248,N_31172);
or U33577 (N_33577,N_31638,N_31567);
xnor U33578 (N_33578,N_31056,N_30195);
nor U33579 (N_33579,N_30220,N_30279);
or U33580 (N_33580,N_30153,N_30082);
and U33581 (N_33581,N_31699,N_31311);
or U33582 (N_33582,N_30642,N_31755);
nand U33583 (N_33583,N_31304,N_30907);
nand U33584 (N_33584,N_30920,N_31058);
and U33585 (N_33585,N_31011,N_30467);
xnor U33586 (N_33586,N_30068,N_30621);
xnor U33587 (N_33587,N_30176,N_30808);
nor U33588 (N_33588,N_30971,N_30072);
and U33589 (N_33589,N_30188,N_30207);
nor U33590 (N_33590,N_30455,N_31944);
nand U33591 (N_33591,N_31316,N_31501);
nor U33592 (N_33592,N_31490,N_30077);
xor U33593 (N_33593,N_31993,N_30298);
and U33594 (N_33594,N_30098,N_31039);
xor U33595 (N_33595,N_30676,N_30997);
or U33596 (N_33596,N_31154,N_30902);
or U33597 (N_33597,N_31468,N_30244);
nand U33598 (N_33598,N_30512,N_30422);
nand U33599 (N_33599,N_31277,N_31651);
xnor U33600 (N_33600,N_31332,N_31211);
nor U33601 (N_33601,N_30626,N_30740);
or U33602 (N_33602,N_31270,N_31902);
and U33603 (N_33603,N_31940,N_30635);
or U33604 (N_33604,N_30822,N_30330);
nor U33605 (N_33605,N_31875,N_30093);
and U33606 (N_33606,N_31286,N_30663);
nor U33607 (N_33607,N_30464,N_31370);
nor U33608 (N_33608,N_30482,N_30056);
or U33609 (N_33609,N_31651,N_30379);
xor U33610 (N_33610,N_30733,N_30890);
nand U33611 (N_33611,N_30592,N_31959);
xor U33612 (N_33612,N_31570,N_30238);
or U33613 (N_33613,N_31686,N_31987);
and U33614 (N_33614,N_30196,N_31088);
xnor U33615 (N_33615,N_30254,N_31596);
nand U33616 (N_33616,N_30779,N_30880);
nor U33617 (N_33617,N_31250,N_31199);
nand U33618 (N_33618,N_30822,N_30657);
nor U33619 (N_33619,N_31391,N_30085);
nand U33620 (N_33620,N_30596,N_30619);
and U33621 (N_33621,N_31107,N_31565);
and U33622 (N_33622,N_30907,N_30590);
xnor U33623 (N_33623,N_30225,N_30735);
or U33624 (N_33624,N_30688,N_30693);
nor U33625 (N_33625,N_31496,N_31455);
nor U33626 (N_33626,N_31586,N_31330);
nand U33627 (N_33627,N_30206,N_31541);
or U33628 (N_33628,N_31067,N_31256);
xor U33629 (N_33629,N_30711,N_31819);
or U33630 (N_33630,N_31914,N_30646);
or U33631 (N_33631,N_30673,N_30237);
or U33632 (N_33632,N_31365,N_30665);
or U33633 (N_33633,N_30633,N_30903);
and U33634 (N_33634,N_31353,N_31393);
or U33635 (N_33635,N_30073,N_31468);
nor U33636 (N_33636,N_31269,N_30452);
nor U33637 (N_33637,N_30923,N_30435);
nand U33638 (N_33638,N_31561,N_30553);
nor U33639 (N_33639,N_31915,N_31319);
or U33640 (N_33640,N_30799,N_30374);
nand U33641 (N_33641,N_30437,N_30967);
nand U33642 (N_33642,N_30439,N_31489);
xor U33643 (N_33643,N_30821,N_30025);
nand U33644 (N_33644,N_30290,N_31263);
and U33645 (N_33645,N_31016,N_31918);
or U33646 (N_33646,N_31764,N_30602);
and U33647 (N_33647,N_30235,N_30628);
nand U33648 (N_33648,N_30293,N_31395);
nand U33649 (N_33649,N_31687,N_30899);
and U33650 (N_33650,N_30662,N_30800);
nor U33651 (N_33651,N_31320,N_31799);
nor U33652 (N_33652,N_31268,N_30322);
nand U33653 (N_33653,N_31947,N_30405);
nor U33654 (N_33654,N_30197,N_30125);
and U33655 (N_33655,N_30816,N_30226);
nand U33656 (N_33656,N_31352,N_31351);
xor U33657 (N_33657,N_31653,N_30286);
and U33658 (N_33658,N_30926,N_31856);
nor U33659 (N_33659,N_30246,N_30231);
xnor U33660 (N_33660,N_30552,N_30468);
and U33661 (N_33661,N_30661,N_30909);
xor U33662 (N_33662,N_31688,N_30983);
xor U33663 (N_33663,N_30552,N_31376);
nand U33664 (N_33664,N_31247,N_31294);
nand U33665 (N_33665,N_31648,N_31849);
nor U33666 (N_33666,N_31394,N_30365);
and U33667 (N_33667,N_31833,N_31518);
nand U33668 (N_33668,N_30873,N_31717);
and U33669 (N_33669,N_31845,N_30057);
and U33670 (N_33670,N_31427,N_30599);
nand U33671 (N_33671,N_31940,N_30191);
and U33672 (N_33672,N_31872,N_31953);
nor U33673 (N_33673,N_31072,N_30980);
and U33674 (N_33674,N_30510,N_30943);
or U33675 (N_33675,N_31633,N_31515);
nor U33676 (N_33676,N_30285,N_31176);
or U33677 (N_33677,N_30885,N_31652);
nor U33678 (N_33678,N_30449,N_31775);
and U33679 (N_33679,N_30480,N_30987);
nand U33680 (N_33680,N_30548,N_31548);
nor U33681 (N_33681,N_30445,N_30915);
xor U33682 (N_33682,N_31399,N_31628);
and U33683 (N_33683,N_30098,N_31100);
nor U33684 (N_33684,N_31857,N_31422);
and U33685 (N_33685,N_31717,N_30915);
or U33686 (N_33686,N_30513,N_31439);
nor U33687 (N_33687,N_31909,N_31337);
xnor U33688 (N_33688,N_31219,N_31124);
or U33689 (N_33689,N_30579,N_30786);
xnor U33690 (N_33690,N_31808,N_30578);
xnor U33691 (N_33691,N_31690,N_30978);
nand U33692 (N_33692,N_30344,N_31629);
nor U33693 (N_33693,N_31709,N_31352);
nand U33694 (N_33694,N_31825,N_30023);
xor U33695 (N_33695,N_30250,N_31922);
nor U33696 (N_33696,N_30919,N_31513);
nand U33697 (N_33697,N_30070,N_31226);
nor U33698 (N_33698,N_31951,N_31993);
xnor U33699 (N_33699,N_30792,N_30225);
nor U33700 (N_33700,N_30457,N_30216);
nor U33701 (N_33701,N_30196,N_31292);
nand U33702 (N_33702,N_31447,N_31697);
nand U33703 (N_33703,N_31773,N_30793);
or U33704 (N_33704,N_31268,N_31059);
nand U33705 (N_33705,N_30439,N_30551);
nand U33706 (N_33706,N_31179,N_31267);
and U33707 (N_33707,N_31595,N_31517);
xor U33708 (N_33708,N_31661,N_31921);
nand U33709 (N_33709,N_31454,N_30987);
nor U33710 (N_33710,N_30733,N_31668);
xnor U33711 (N_33711,N_31764,N_31453);
and U33712 (N_33712,N_30510,N_30620);
xnor U33713 (N_33713,N_31841,N_30417);
nand U33714 (N_33714,N_31055,N_30804);
nand U33715 (N_33715,N_31138,N_31350);
xnor U33716 (N_33716,N_30764,N_31442);
or U33717 (N_33717,N_31330,N_31149);
and U33718 (N_33718,N_31803,N_30820);
nand U33719 (N_33719,N_30076,N_30060);
nand U33720 (N_33720,N_31917,N_31443);
nor U33721 (N_33721,N_31824,N_31871);
or U33722 (N_33722,N_31093,N_31070);
nand U33723 (N_33723,N_31266,N_31684);
or U33724 (N_33724,N_30883,N_31698);
and U33725 (N_33725,N_30279,N_31130);
nand U33726 (N_33726,N_30012,N_30177);
or U33727 (N_33727,N_31002,N_30399);
xnor U33728 (N_33728,N_30032,N_30016);
xor U33729 (N_33729,N_31410,N_30468);
nand U33730 (N_33730,N_30941,N_31786);
nor U33731 (N_33731,N_31319,N_30020);
or U33732 (N_33732,N_30224,N_31116);
or U33733 (N_33733,N_30206,N_30484);
xnor U33734 (N_33734,N_31138,N_31840);
nor U33735 (N_33735,N_30835,N_30973);
and U33736 (N_33736,N_31843,N_30174);
nand U33737 (N_33737,N_30060,N_31368);
nor U33738 (N_33738,N_31428,N_30468);
or U33739 (N_33739,N_30132,N_30564);
and U33740 (N_33740,N_31069,N_31348);
nand U33741 (N_33741,N_31249,N_30494);
or U33742 (N_33742,N_31996,N_30989);
nor U33743 (N_33743,N_31257,N_30098);
nand U33744 (N_33744,N_31641,N_31560);
nand U33745 (N_33745,N_30564,N_30457);
xnor U33746 (N_33746,N_30244,N_30165);
xor U33747 (N_33747,N_30397,N_31822);
and U33748 (N_33748,N_30450,N_30436);
nand U33749 (N_33749,N_30062,N_31283);
or U33750 (N_33750,N_30211,N_31702);
or U33751 (N_33751,N_30296,N_30957);
and U33752 (N_33752,N_30890,N_31859);
nand U33753 (N_33753,N_30302,N_31213);
or U33754 (N_33754,N_30339,N_30606);
xnor U33755 (N_33755,N_31276,N_31949);
nor U33756 (N_33756,N_31059,N_30162);
nand U33757 (N_33757,N_31953,N_30951);
nor U33758 (N_33758,N_30062,N_30146);
and U33759 (N_33759,N_31578,N_30524);
nand U33760 (N_33760,N_30040,N_31030);
nand U33761 (N_33761,N_31150,N_30180);
nor U33762 (N_33762,N_31294,N_31848);
nor U33763 (N_33763,N_31234,N_31949);
nand U33764 (N_33764,N_30842,N_31647);
nand U33765 (N_33765,N_31970,N_30601);
nor U33766 (N_33766,N_31949,N_31547);
xnor U33767 (N_33767,N_30637,N_30141);
or U33768 (N_33768,N_30279,N_31710);
and U33769 (N_33769,N_31067,N_30962);
nand U33770 (N_33770,N_31490,N_30103);
xnor U33771 (N_33771,N_31183,N_30424);
nand U33772 (N_33772,N_30081,N_30540);
and U33773 (N_33773,N_31955,N_30375);
and U33774 (N_33774,N_31693,N_31364);
xnor U33775 (N_33775,N_31023,N_30287);
and U33776 (N_33776,N_31071,N_31113);
nand U33777 (N_33777,N_30381,N_30250);
or U33778 (N_33778,N_30477,N_31042);
xnor U33779 (N_33779,N_31221,N_31897);
nand U33780 (N_33780,N_30330,N_31825);
and U33781 (N_33781,N_30815,N_31727);
xnor U33782 (N_33782,N_31727,N_30317);
and U33783 (N_33783,N_31270,N_30565);
and U33784 (N_33784,N_31510,N_31601);
and U33785 (N_33785,N_30411,N_31836);
and U33786 (N_33786,N_31045,N_30788);
or U33787 (N_33787,N_31816,N_30843);
and U33788 (N_33788,N_30373,N_31324);
or U33789 (N_33789,N_30950,N_31641);
nor U33790 (N_33790,N_31050,N_31748);
nand U33791 (N_33791,N_30903,N_31924);
nand U33792 (N_33792,N_31493,N_30568);
nor U33793 (N_33793,N_30027,N_31380);
xor U33794 (N_33794,N_31715,N_30947);
and U33795 (N_33795,N_30334,N_31794);
or U33796 (N_33796,N_31678,N_31319);
xor U33797 (N_33797,N_31283,N_30924);
nor U33798 (N_33798,N_31494,N_30624);
or U33799 (N_33799,N_31136,N_30754);
or U33800 (N_33800,N_31103,N_30526);
nor U33801 (N_33801,N_30647,N_31231);
and U33802 (N_33802,N_31313,N_30021);
or U33803 (N_33803,N_30465,N_30973);
and U33804 (N_33804,N_31378,N_31942);
or U33805 (N_33805,N_31052,N_30396);
nor U33806 (N_33806,N_31556,N_30614);
xnor U33807 (N_33807,N_30661,N_31280);
and U33808 (N_33808,N_31731,N_30460);
and U33809 (N_33809,N_31876,N_30350);
nand U33810 (N_33810,N_30001,N_30176);
xor U33811 (N_33811,N_30795,N_30491);
xor U33812 (N_33812,N_30573,N_31741);
nand U33813 (N_33813,N_30893,N_31960);
nand U33814 (N_33814,N_31593,N_30718);
or U33815 (N_33815,N_31014,N_31040);
or U33816 (N_33816,N_31871,N_30630);
xnor U33817 (N_33817,N_31042,N_30082);
or U33818 (N_33818,N_31075,N_31693);
nand U33819 (N_33819,N_30554,N_31896);
or U33820 (N_33820,N_30474,N_31216);
nand U33821 (N_33821,N_31649,N_30081);
or U33822 (N_33822,N_31438,N_31486);
nand U33823 (N_33823,N_30327,N_31298);
nand U33824 (N_33824,N_31127,N_31658);
and U33825 (N_33825,N_30916,N_30381);
nand U33826 (N_33826,N_30694,N_31059);
nand U33827 (N_33827,N_30805,N_30094);
and U33828 (N_33828,N_31285,N_30040);
and U33829 (N_33829,N_31929,N_31895);
and U33830 (N_33830,N_30881,N_30311);
nor U33831 (N_33831,N_30508,N_31653);
xor U33832 (N_33832,N_30302,N_31400);
xor U33833 (N_33833,N_31138,N_31333);
and U33834 (N_33834,N_30180,N_31336);
nand U33835 (N_33835,N_31048,N_31315);
nor U33836 (N_33836,N_31080,N_30438);
nor U33837 (N_33837,N_31736,N_30315);
or U33838 (N_33838,N_31826,N_31098);
and U33839 (N_33839,N_30166,N_30831);
nand U33840 (N_33840,N_30116,N_31944);
and U33841 (N_33841,N_31287,N_30635);
xnor U33842 (N_33842,N_30951,N_31260);
nand U33843 (N_33843,N_31807,N_30319);
nor U33844 (N_33844,N_30954,N_30433);
nand U33845 (N_33845,N_31836,N_30452);
or U33846 (N_33846,N_30891,N_31874);
nor U33847 (N_33847,N_31515,N_31010);
nor U33848 (N_33848,N_31560,N_31427);
and U33849 (N_33849,N_30663,N_30789);
nand U33850 (N_33850,N_30420,N_30104);
nand U33851 (N_33851,N_30517,N_31345);
nor U33852 (N_33852,N_31621,N_30376);
xor U33853 (N_33853,N_31908,N_30954);
nand U33854 (N_33854,N_31183,N_30982);
nand U33855 (N_33855,N_31739,N_30476);
xnor U33856 (N_33856,N_30731,N_31351);
nor U33857 (N_33857,N_30335,N_31074);
or U33858 (N_33858,N_31579,N_30434);
nor U33859 (N_33859,N_30402,N_30078);
xor U33860 (N_33860,N_31371,N_31479);
xnor U33861 (N_33861,N_31068,N_31207);
and U33862 (N_33862,N_30157,N_31702);
or U33863 (N_33863,N_31685,N_30165);
nor U33864 (N_33864,N_31298,N_30316);
or U33865 (N_33865,N_30100,N_30399);
and U33866 (N_33866,N_30295,N_31126);
nor U33867 (N_33867,N_31456,N_31138);
or U33868 (N_33868,N_30018,N_31499);
and U33869 (N_33869,N_31148,N_30473);
xor U33870 (N_33870,N_31074,N_30178);
or U33871 (N_33871,N_31346,N_31791);
and U33872 (N_33872,N_31340,N_30487);
xnor U33873 (N_33873,N_31542,N_31035);
xnor U33874 (N_33874,N_30105,N_31892);
and U33875 (N_33875,N_30078,N_31669);
and U33876 (N_33876,N_30608,N_30689);
and U33877 (N_33877,N_30782,N_30801);
nor U33878 (N_33878,N_30317,N_31868);
nor U33879 (N_33879,N_30360,N_31588);
or U33880 (N_33880,N_31830,N_30730);
nor U33881 (N_33881,N_30603,N_30506);
nor U33882 (N_33882,N_30380,N_31635);
nand U33883 (N_33883,N_31597,N_30797);
and U33884 (N_33884,N_30789,N_31439);
nand U33885 (N_33885,N_31266,N_30575);
nor U33886 (N_33886,N_31825,N_30943);
or U33887 (N_33887,N_31667,N_30614);
nor U33888 (N_33888,N_31157,N_31415);
nand U33889 (N_33889,N_31533,N_30184);
xor U33890 (N_33890,N_31885,N_30215);
xnor U33891 (N_33891,N_31978,N_31408);
nor U33892 (N_33892,N_31557,N_31836);
nand U33893 (N_33893,N_31664,N_31701);
xnor U33894 (N_33894,N_30312,N_31486);
and U33895 (N_33895,N_30224,N_30844);
xnor U33896 (N_33896,N_30893,N_31762);
nand U33897 (N_33897,N_31789,N_30737);
nand U33898 (N_33898,N_30463,N_30438);
or U33899 (N_33899,N_30359,N_31300);
or U33900 (N_33900,N_30124,N_31238);
and U33901 (N_33901,N_30049,N_30640);
nor U33902 (N_33902,N_31356,N_31167);
and U33903 (N_33903,N_31529,N_31119);
or U33904 (N_33904,N_31759,N_31321);
xnor U33905 (N_33905,N_30419,N_30131);
xor U33906 (N_33906,N_31195,N_30102);
nand U33907 (N_33907,N_31488,N_31745);
and U33908 (N_33908,N_30441,N_31535);
or U33909 (N_33909,N_31895,N_31196);
and U33910 (N_33910,N_30538,N_30514);
or U33911 (N_33911,N_31867,N_31728);
nand U33912 (N_33912,N_31260,N_31624);
nor U33913 (N_33913,N_30125,N_30607);
xor U33914 (N_33914,N_30280,N_31813);
or U33915 (N_33915,N_31355,N_31025);
nand U33916 (N_33916,N_30579,N_31969);
xnor U33917 (N_33917,N_31205,N_30845);
or U33918 (N_33918,N_30814,N_30001);
nor U33919 (N_33919,N_31086,N_31492);
nor U33920 (N_33920,N_30165,N_30333);
nor U33921 (N_33921,N_31152,N_30545);
or U33922 (N_33922,N_31895,N_30331);
nand U33923 (N_33923,N_30526,N_30449);
and U33924 (N_33924,N_30933,N_31563);
or U33925 (N_33925,N_31753,N_30686);
nor U33926 (N_33926,N_30997,N_30557);
nor U33927 (N_33927,N_30931,N_30932);
nand U33928 (N_33928,N_31406,N_30617);
nand U33929 (N_33929,N_31574,N_31028);
nor U33930 (N_33930,N_31134,N_30225);
and U33931 (N_33931,N_30219,N_31364);
nand U33932 (N_33932,N_30158,N_30785);
and U33933 (N_33933,N_31208,N_30561);
or U33934 (N_33934,N_30654,N_31088);
or U33935 (N_33935,N_30552,N_30776);
xnor U33936 (N_33936,N_31904,N_31758);
or U33937 (N_33937,N_31767,N_30338);
xnor U33938 (N_33938,N_31066,N_31966);
and U33939 (N_33939,N_30107,N_31140);
nand U33940 (N_33940,N_30184,N_31145);
and U33941 (N_33941,N_30962,N_31267);
or U33942 (N_33942,N_31748,N_30979);
nand U33943 (N_33943,N_30144,N_30969);
nor U33944 (N_33944,N_31822,N_30546);
nand U33945 (N_33945,N_30800,N_31593);
or U33946 (N_33946,N_31452,N_30940);
or U33947 (N_33947,N_31020,N_30202);
and U33948 (N_33948,N_31050,N_31524);
xor U33949 (N_33949,N_30632,N_30579);
nor U33950 (N_33950,N_31738,N_30069);
and U33951 (N_33951,N_30057,N_30936);
nand U33952 (N_33952,N_31862,N_30878);
or U33953 (N_33953,N_30393,N_31635);
nand U33954 (N_33954,N_31258,N_31672);
nand U33955 (N_33955,N_31979,N_30184);
and U33956 (N_33956,N_30882,N_30096);
and U33957 (N_33957,N_30799,N_30854);
xor U33958 (N_33958,N_31804,N_30498);
nand U33959 (N_33959,N_30552,N_30687);
nor U33960 (N_33960,N_30975,N_30655);
xnor U33961 (N_33961,N_30038,N_30817);
or U33962 (N_33962,N_30447,N_30148);
and U33963 (N_33963,N_31208,N_30771);
nand U33964 (N_33964,N_30020,N_30077);
xor U33965 (N_33965,N_31967,N_31656);
or U33966 (N_33966,N_30102,N_31177);
nor U33967 (N_33967,N_31843,N_30461);
xor U33968 (N_33968,N_30366,N_31030);
xnor U33969 (N_33969,N_31811,N_30473);
nor U33970 (N_33970,N_31096,N_31792);
or U33971 (N_33971,N_30834,N_31448);
nand U33972 (N_33972,N_31922,N_31269);
nand U33973 (N_33973,N_30756,N_30077);
or U33974 (N_33974,N_31736,N_31083);
xnor U33975 (N_33975,N_30343,N_31125);
and U33976 (N_33976,N_31419,N_31576);
xor U33977 (N_33977,N_31638,N_31816);
nand U33978 (N_33978,N_31622,N_30724);
xnor U33979 (N_33979,N_30066,N_31403);
nand U33980 (N_33980,N_30585,N_30980);
xnor U33981 (N_33981,N_31578,N_30365);
xor U33982 (N_33982,N_31670,N_31660);
nand U33983 (N_33983,N_31670,N_30177);
nand U33984 (N_33984,N_30097,N_30769);
xnor U33985 (N_33985,N_31581,N_30141);
nor U33986 (N_33986,N_31814,N_30256);
and U33987 (N_33987,N_31478,N_30498);
and U33988 (N_33988,N_31460,N_31533);
xnor U33989 (N_33989,N_30843,N_31132);
or U33990 (N_33990,N_31028,N_30326);
xor U33991 (N_33991,N_30782,N_31708);
nand U33992 (N_33992,N_30099,N_30635);
nor U33993 (N_33993,N_31303,N_30047);
xor U33994 (N_33994,N_30131,N_30182);
xnor U33995 (N_33995,N_30647,N_31621);
and U33996 (N_33996,N_30584,N_31837);
nor U33997 (N_33997,N_30252,N_31980);
nand U33998 (N_33998,N_31791,N_30289);
nand U33999 (N_33999,N_30807,N_30470);
xnor U34000 (N_34000,N_33473,N_33478);
nand U34001 (N_34001,N_32207,N_33755);
and U34002 (N_34002,N_33687,N_32203);
nand U34003 (N_34003,N_33309,N_32667);
or U34004 (N_34004,N_33583,N_33059);
nand U34005 (N_34005,N_32285,N_33470);
nand U34006 (N_34006,N_32430,N_33963);
xnor U34007 (N_34007,N_32149,N_32323);
or U34008 (N_34008,N_32061,N_33632);
nor U34009 (N_34009,N_32234,N_32373);
xnor U34010 (N_34010,N_32941,N_33357);
nor U34011 (N_34011,N_33346,N_33715);
nand U34012 (N_34012,N_33073,N_32568);
or U34013 (N_34013,N_33783,N_33421);
or U34014 (N_34014,N_32503,N_33328);
and U34015 (N_34015,N_33873,N_32458);
nor U34016 (N_34016,N_33926,N_33941);
or U34017 (N_34017,N_33829,N_32728);
xnor U34018 (N_34018,N_32489,N_33146);
nor U34019 (N_34019,N_33033,N_32699);
nand U34020 (N_34020,N_32355,N_33114);
nor U34021 (N_34021,N_32339,N_32624);
and U34022 (N_34022,N_32960,N_32722);
or U34023 (N_34023,N_33965,N_33657);
and U34024 (N_34024,N_33377,N_32327);
or U34025 (N_34025,N_32215,N_33789);
or U34026 (N_34026,N_32438,N_33944);
and U34027 (N_34027,N_32023,N_33369);
or U34028 (N_34028,N_33663,N_32427);
nor U34029 (N_34029,N_32603,N_33525);
nand U34030 (N_34030,N_33822,N_33919);
nand U34031 (N_34031,N_33824,N_32771);
nor U34032 (N_34032,N_32409,N_32147);
and U34033 (N_34033,N_32175,N_32093);
nor U34034 (N_34034,N_33600,N_33008);
nor U34035 (N_34035,N_32530,N_33801);
nor U34036 (N_34036,N_33752,N_33484);
nand U34037 (N_34037,N_33539,N_33215);
nor U34038 (N_34038,N_33007,N_33798);
nor U34039 (N_34039,N_33452,N_32273);
and U34040 (N_34040,N_33474,N_32159);
nand U34041 (N_34041,N_32414,N_33904);
xnor U34042 (N_34042,N_32721,N_33046);
nand U34043 (N_34043,N_33998,N_33709);
xor U34044 (N_34044,N_33440,N_33994);
or U34045 (N_34045,N_33052,N_33287);
and U34046 (N_34046,N_33678,N_32270);
and U34047 (N_34047,N_32152,N_33480);
nor U34048 (N_34048,N_32027,N_33603);
nor U34049 (N_34049,N_33067,N_32357);
or U34050 (N_34050,N_32957,N_33886);
and U34051 (N_34051,N_32112,N_33285);
and U34052 (N_34052,N_32221,N_33284);
and U34053 (N_34053,N_32882,N_33496);
xor U34054 (N_34054,N_33292,N_33895);
or U34055 (N_34055,N_33934,N_32782);
nand U34056 (N_34056,N_32440,N_32294);
xnor U34057 (N_34057,N_33051,N_33072);
and U34058 (N_34058,N_32878,N_33320);
xor U34059 (N_34059,N_32226,N_32080);
xnor U34060 (N_34060,N_33802,N_33071);
and U34061 (N_34061,N_32311,N_33862);
nor U34062 (N_34062,N_32309,N_32401);
nand U34063 (N_34063,N_33395,N_32816);
nand U34064 (N_34064,N_33710,N_33265);
and U34065 (N_34065,N_33524,N_33240);
or U34066 (N_34066,N_33701,N_32094);
and U34067 (N_34067,N_33803,N_32527);
nor U34068 (N_34068,N_33355,N_33411);
or U34069 (N_34069,N_32399,N_32677);
and U34070 (N_34070,N_33375,N_33262);
and U34071 (N_34071,N_33960,N_32165);
or U34072 (N_34072,N_32714,N_32923);
nor U34073 (N_34073,N_32451,N_33549);
or U34074 (N_34074,N_33273,N_32808);
and U34075 (N_34075,N_32161,N_32640);
and U34076 (N_34076,N_32108,N_33201);
or U34077 (N_34077,N_32184,N_32884);
or U34078 (N_34078,N_32491,N_33612);
xnor U34079 (N_34079,N_32068,N_32111);
nor U34080 (N_34080,N_32597,N_32452);
nand U34081 (N_34081,N_33106,N_32576);
nand U34082 (N_34082,N_32509,N_32439);
nand U34083 (N_34083,N_33171,N_32420);
xnor U34084 (N_34084,N_32138,N_32158);
xnor U34085 (N_34085,N_33724,N_32441);
xor U34086 (N_34086,N_32672,N_33365);
or U34087 (N_34087,N_33719,N_33380);
or U34088 (N_34088,N_32818,N_33143);
or U34089 (N_34089,N_33630,N_32856);
nand U34090 (N_34090,N_32828,N_33455);
or U34091 (N_34091,N_32510,N_32867);
and U34092 (N_34092,N_33676,N_33510);
xnor U34093 (N_34093,N_33604,N_32933);
nor U34094 (N_34094,N_33808,N_33288);
xor U34095 (N_34095,N_32873,N_33069);
nor U34096 (N_34096,N_33775,N_32574);
xor U34097 (N_34097,N_33209,N_32251);
nand U34098 (N_34098,N_32666,N_33537);
or U34099 (N_34099,N_32442,N_32349);
xor U34100 (N_34100,N_33990,N_33207);
nand U34101 (N_34101,N_33551,N_32620);
nand U34102 (N_34102,N_33232,N_32935);
and U34103 (N_34103,N_33279,N_32275);
nand U34104 (N_34104,N_33139,N_33823);
and U34105 (N_34105,N_33268,N_33979);
nand U34106 (N_34106,N_32801,N_32484);
nand U34107 (N_34107,N_33386,N_32186);
xor U34108 (N_34108,N_32348,N_33521);
and U34109 (N_34109,N_32747,N_33160);
or U34110 (N_34110,N_33336,N_33693);
xor U34111 (N_34111,N_33836,N_32696);
or U34112 (N_34112,N_32182,N_33865);
xnor U34113 (N_34113,N_33057,N_32318);
nor U34114 (N_34114,N_33573,N_33690);
nand U34115 (N_34115,N_32560,N_32085);
nand U34116 (N_34116,N_33408,N_32483);
xor U34117 (N_34117,N_32997,N_32836);
and U34118 (N_34118,N_32717,N_33857);
xor U34119 (N_34119,N_33061,N_32287);
xor U34120 (N_34120,N_33419,N_32129);
or U34121 (N_34121,N_33140,N_33195);
nand U34122 (N_34122,N_32268,N_33964);
xnor U34123 (N_34123,N_32972,N_32209);
or U34124 (N_34124,N_32245,N_33736);
and U34125 (N_34125,N_33000,N_32352);
and U34126 (N_34126,N_32598,N_32365);
or U34127 (N_34127,N_33515,N_32211);
or U34128 (N_34128,N_33306,N_33432);
and U34129 (N_34129,N_33435,N_33954);
and U34130 (N_34130,N_32927,N_33307);
or U34131 (N_34131,N_32999,N_32661);
and U34132 (N_34132,N_32858,N_33368);
xor U34133 (N_34133,N_33290,N_33298);
xnor U34134 (N_34134,N_32854,N_33224);
nor U34135 (N_34135,N_33413,N_32086);
nand U34136 (N_34136,N_32631,N_33325);
nand U34137 (N_34137,N_32437,N_33389);
and U34138 (N_34138,N_32014,N_32976);
xor U34139 (N_34139,N_33397,N_33312);
nand U34140 (N_34140,N_33592,N_32306);
and U34141 (N_34141,N_33134,N_33472);
and U34142 (N_34142,N_32272,N_32101);
or U34143 (N_34143,N_32859,N_33983);
nand U34144 (N_34144,N_32267,N_32792);
and U34145 (N_34145,N_33444,N_32787);
and U34146 (N_34146,N_33210,N_33782);
nand U34147 (N_34147,N_33514,N_33576);
xor U34148 (N_34148,N_33556,N_33247);
nand U34149 (N_34149,N_33070,N_33703);
nand U34150 (N_34150,N_33508,N_32024);
nor U34151 (N_34151,N_33550,N_32403);
xor U34152 (N_34152,N_32778,N_33436);
xor U34153 (N_34153,N_33850,N_32394);
xnor U34154 (N_34154,N_32644,N_32555);
or U34155 (N_34155,N_33372,N_33216);
xor U34156 (N_34156,N_32536,N_32078);
nor U34157 (N_34157,N_33929,N_33644);
or U34158 (N_34158,N_32166,N_32404);
and U34159 (N_34159,N_32632,N_33077);
or U34160 (N_34160,N_33342,N_32822);
xor U34161 (N_34161,N_32300,N_33699);
nand U34162 (N_34162,N_32075,N_33203);
or U34163 (N_34163,N_32682,N_33655);
or U34164 (N_34164,N_32838,N_32673);
nand U34165 (N_34165,N_32379,N_33396);
or U34166 (N_34166,N_32235,N_33907);
nand U34167 (N_34167,N_32876,N_32942);
and U34168 (N_34168,N_33962,N_33161);
nand U34169 (N_34169,N_33781,N_32140);
and U34170 (N_34170,N_32196,N_33691);
nand U34171 (N_34171,N_32614,N_33560);
nor U34172 (N_34172,N_32160,N_32225);
xor U34173 (N_34173,N_33037,N_32383);
nor U34174 (N_34174,N_32797,N_32183);
nand U34175 (N_34175,N_32350,N_33731);
or U34176 (N_34176,N_33587,N_32675);
or U34177 (N_34177,N_33433,N_33289);
nand U34178 (N_34178,N_32082,N_32072);
xnor U34179 (N_34179,N_32926,N_32587);
and U34180 (N_34180,N_33011,N_32843);
or U34181 (N_34181,N_33658,N_32331);
xor U34182 (N_34182,N_33733,N_32304);
xnor U34183 (N_34183,N_33950,N_32125);
nand U34184 (N_34184,N_33916,N_32839);
nor U34185 (N_34185,N_33887,N_33559);
nand U34186 (N_34186,N_33189,N_33393);
nand U34187 (N_34187,N_33429,N_32146);
nand U34188 (N_34188,N_32040,N_32793);
or U34189 (N_34189,N_32929,N_32353);
nand U34190 (N_34190,N_32260,N_32993);
and U34191 (N_34191,N_33115,N_32518);
or U34192 (N_34192,N_32475,N_33107);
xnor U34193 (N_34193,N_32756,N_33304);
xor U34194 (N_34194,N_32232,N_33953);
xor U34195 (N_34195,N_33347,N_32141);
xor U34196 (N_34196,N_33099,N_33980);
nor U34197 (N_34197,N_32594,N_33184);
and U34198 (N_34198,N_32785,N_32638);
and U34199 (N_34199,N_32174,N_33152);
nor U34200 (N_34200,N_33669,N_33374);
or U34201 (N_34201,N_32837,N_33970);
nand U34202 (N_34202,N_33238,N_32951);
or U34203 (N_34203,N_32692,N_33523);
nor U34204 (N_34204,N_33625,N_32637);
or U34205 (N_34205,N_33384,N_33038);
nor U34206 (N_34206,N_32197,N_32849);
or U34207 (N_34207,N_32916,N_32543);
and U34208 (N_34208,N_32513,N_33925);
nand U34209 (N_34209,N_32768,N_33951);
nand U34210 (N_34210,N_33827,N_32986);
or U34211 (N_34211,N_33972,N_32761);
nor U34212 (N_34212,N_32004,N_32307);
or U34213 (N_34213,N_33391,N_32554);
or U34214 (N_34214,N_32522,N_33302);
nor U34215 (N_34215,N_32487,N_32636);
and U34216 (N_34216,N_32443,N_33494);
or U34217 (N_34217,N_32319,N_32674);
or U34218 (N_34218,N_33686,N_33150);
nor U34219 (N_34219,N_32264,N_32544);
or U34220 (N_34220,N_33588,N_33174);
nor U34221 (N_34221,N_33349,N_33175);
and U34222 (N_34222,N_33404,N_33042);
nor U34223 (N_34223,N_32000,N_32959);
nor U34224 (N_34224,N_32780,N_32378);
xnor U34225 (N_34225,N_32851,N_32120);
or U34226 (N_34226,N_32700,N_32609);
and U34227 (N_34227,N_33414,N_33572);
nor U34228 (N_34228,N_32137,N_33029);
or U34229 (N_34229,N_33405,N_32645);
and U34230 (N_34230,N_33875,N_33027);
and U34231 (N_34231,N_32312,N_33351);
nand U34232 (N_34232,N_33567,N_32848);
nor U34233 (N_34233,N_32062,N_32930);
or U34234 (N_34234,N_32978,N_32833);
xnor U34235 (N_34235,N_32217,N_32759);
and U34236 (N_34236,N_32727,N_32514);
nand U34237 (N_34237,N_33527,N_32054);
or U34238 (N_34238,N_32222,N_32563);
or U34239 (N_34239,N_33729,N_33622);
and U34240 (N_34240,N_33677,N_33235);
or U34241 (N_34241,N_32936,N_33424);
and U34242 (N_34242,N_32177,N_33698);
nor U34243 (N_34243,N_33859,N_33271);
nand U34244 (N_34244,N_33503,N_33125);
nor U34245 (N_34245,N_33529,N_33996);
nor U34246 (N_34246,N_33048,N_32567);
xnor U34247 (N_34247,N_32920,N_32725);
and U34248 (N_34248,N_32372,N_33236);
xor U34249 (N_34249,N_33502,N_33530);
nand U34250 (N_34250,N_33640,N_32476);
nor U34251 (N_34251,N_32965,N_32382);
and U34252 (N_34252,N_32366,N_33229);
xnor U34253 (N_34253,N_32444,N_32336);
and U34254 (N_34254,N_32810,N_32283);
nor U34255 (N_34255,N_32893,N_32201);
or U34256 (N_34256,N_33138,N_33773);
nor U34257 (N_34257,N_32391,N_32777);
or U34258 (N_34258,N_33155,N_33939);
or U34259 (N_34259,N_32274,N_32504);
or U34260 (N_34260,N_33096,N_33418);
and U34261 (N_34261,N_32477,N_33400);
nor U34262 (N_34262,N_33804,N_33810);
and U34263 (N_34263,N_33330,N_33725);
xnor U34264 (N_34264,N_33883,N_33322);
nand U34265 (N_34265,N_32398,N_33518);
xor U34266 (N_34266,N_32332,N_33423);
or U34267 (N_34267,N_32124,N_32607);
or U34268 (N_34268,N_33874,N_33467);
nand U34269 (N_34269,N_33516,N_33682);
and U34270 (N_34270,N_33860,N_33075);
nand U34271 (N_34271,N_32055,N_32255);
or U34272 (N_34272,N_32938,N_32694);
nor U34273 (N_34273,N_33674,N_33517);
or U34274 (N_34274,N_33915,N_33564);
nand U34275 (N_34275,N_32626,N_33280);
nor U34276 (N_34276,N_32465,N_33596);
nand U34277 (N_34277,N_33259,N_33745);
or U34278 (N_34278,N_33202,N_33017);
or U34279 (N_34279,N_33512,N_33332);
nand U34280 (N_34280,N_32259,N_33797);
nor U34281 (N_34281,N_32962,N_33590);
nand U34282 (N_34282,N_32276,N_33722);
nand U34283 (N_34283,N_32831,N_33899);
nand U34284 (N_34284,N_33918,N_32749);
nand U34285 (N_34285,N_32032,N_32115);
or U34286 (N_34286,N_32605,N_33794);
nand U34287 (N_34287,N_33519,N_33233);
nand U34288 (N_34288,N_32776,N_32257);
and U34289 (N_34289,N_33645,N_32971);
nor U34290 (N_34290,N_33402,N_33947);
or U34291 (N_34291,N_32531,N_33805);
nor U34292 (N_34292,N_33465,N_33911);
xnor U34293 (N_34293,N_32190,N_33853);
or U34294 (N_34294,N_33989,N_32669);
or U34295 (N_34295,N_33049,N_32116);
and U34296 (N_34296,N_33345,N_32153);
or U34297 (N_34297,N_32520,N_32416);
nor U34298 (N_34298,N_32515,N_32407);
or U34299 (N_34299,N_33392,N_33685);
nand U34300 (N_34300,N_33754,N_32301);
nand U34301 (N_34301,N_33593,N_33006);
xnor U34302 (N_34302,N_33252,N_32067);
or U34303 (N_34303,N_33969,N_32150);
nand U34304 (N_34304,N_33806,N_33223);
xor U34305 (N_34305,N_32195,N_32846);
xor U34306 (N_34306,N_33132,N_32519);
and U34307 (N_34307,N_32627,N_33881);
nor U34308 (N_34308,N_32013,N_33277);
or U34309 (N_34309,N_32244,N_32271);
nor U34310 (N_34310,N_33013,N_32719);
or U34311 (N_34311,N_33153,N_33777);
xor U34312 (N_34312,N_33430,N_33296);
nand U34313 (N_34313,N_32910,N_32526);
or U34314 (N_34314,N_33167,N_33591);
nor U34315 (N_34315,N_32584,N_33780);
nand U34316 (N_34316,N_33667,N_33364);
xor U34317 (N_34317,N_33741,N_32709);
nor U34318 (N_34318,N_33636,N_33065);
nand U34319 (N_34319,N_32381,N_33927);
and U34320 (N_34320,N_32964,N_33986);
and U34321 (N_34321,N_32208,N_33565);
nor U34322 (N_34322,N_32090,N_33659);
nand U34323 (N_34323,N_33917,N_33680);
or U34324 (N_34324,N_33906,N_33876);
and U34325 (N_34325,N_33879,N_32252);
or U34326 (N_34326,N_32593,N_32046);
xnor U34327 (N_34327,N_32303,N_33270);
nand U34328 (N_34328,N_33118,N_33100);
or U34329 (N_34329,N_33102,N_33267);
nor U34330 (N_34330,N_32900,N_32875);
xnor U34331 (N_34331,N_33749,N_32180);
xor U34332 (N_34332,N_33889,N_32652);
nor U34333 (N_34333,N_33513,N_33818);
and U34334 (N_34334,N_33620,N_33053);
and U34335 (N_34335,N_32360,N_32803);
or U34336 (N_34336,N_33942,N_33714);
nand U34337 (N_34337,N_32523,N_33083);
or U34338 (N_34338,N_33757,N_33028);
nand U34339 (N_34339,N_33828,N_33727);
and U34340 (N_34340,N_33205,N_33766);
or U34341 (N_34341,N_33263,N_32495);
xor U34342 (N_34342,N_32230,N_32281);
nor U34343 (N_34343,N_33373,N_33973);
or U34344 (N_34344,N_32337,N_33842);
xor U34345 (N_34345,N_33089,N_33511);
nand U34346 (N_34346,N_33534,N_32114);
nand U34347 (N_34347,N_33054,N_33326);
nand U34348 (N_34348,N_32676,N_32421);
nor U34349 (N_34349,N_32755,N_32043);
nand U34350 (N_34350,N_33156,N_32500);
nand U34351 (N_34351,N_33605,N_32585);
and U34352 (N_34352,N_32842,N_32928);
nor U34353 (N_34353,N_33087,N_33159);
nand U34354 (N_34354,N_33169,N_32826);
or U34355 (N_34355,N_33643,N_32733);
nand U34356 (N_34356,N_32660,N_32254);
nor U34357 (N_34357,N_33381,N_33213);
nand U34358 (N_34358,N_32422,N_33335);
nand U34359 (N_34359,N_32871,N_32293);
or U34360 (N_34360,N_32435,N_33334);
and U34361 (N_34361,N_33490,N_32074);
nand U34362 (N_34362,N_33219,N_32047);
xor U34363 (N_34363,N_33713,N_33097);
and U34364 (N_34364,N_33191,N_33062);
and U34365 (N_34365,N_33726,N_32497);
xnor U34366 (N_34366,N_33343,N_33275);
nor U34367 (N_34367,N_32739,N_32091);
or U34368 (N_34368,N_32097,N_33554);
and U34369 (N_34369,N_32498,N_33449);
nor U34370 (N_34370,N_33743,N_32821);
and U34371 (N_34371,N_33672,N_33291);
and U34372 (N_34372,N_33226,N_32912);
nor U34373 (N_34373,N_32118,N_33858);
nor U34374 (N_34374,N_32006,N_32214);
nor U34375 (N_34375,N_32646,N_32892);
xnor U34376 (N_34376,N_33193,N_33647);
nor U34377 (N_34377,N_33378,N_33997);
or U34378 (N_34378,N_33767,N_33788);
or U34379 (N_34379,N_32814,N_32123);
or U34380 (N_34380,N_33181,N_32164);
and U34381 (N_34381,N_33297,N_32246);
nand U34382 (N_34382,N_32872,N_33208);
nor U34383 (N_34383,N_32983,N_33589);
nor U34384 (N_34384,N_33353,N_32376);
nand U34385 (N_34385,N_32695,N_32885);
xnor U34386 (N_34386,N_32918,N_32501);
and U34387 (N_34387,N_33183,N_32641);
or U34388 (N_34388,N_32480,N_32305);
nor U34389 (N_34389,N_33464,N_32291);
nor U34390 (N_34390,N_33885,N_33579);
or U34391 (N_34391,N_32809,N_33661);
xor U34392 (N_34392,N_32764,N_32098);
xnor U34393 (N_34393,N_32107,N_32359);
xor U34394 (N_34394,N_33570,N_33383);
and U34395 (N_34395,N_32173,N_33370);
and U34396 (N_34396,N_33629,N_33103);
or U34397 (N_34397,N_32845,N_32994);
and U34398 (N_34398,N_33833,N_33684);
and U34399 (N_34399,N_32426,N_32343);
xor U34400 (N_34400,N_32070,N_33656);
and U34401 (N_34401,N_32945,N_32529);
or U34402 (N_34402,N_33366,N_32857);
or U34403 (N_34403,N_32686,N_33136);
nand U34404 (N_34404,N_32693,N_33064);
and U34405 (N_34405,N_33618,N_32711);
or U34406 (N_34406,N_32237,N_32344);
nor U34407 (N_34407,N_33759,N_33555);
nand U34408 (N_34408,N_33166,N_33839);
or U34409 (N_34409,N_32330,N_32862);
nand U34410 (N_34410,N_32369,N_32290);
or U34411 (N_34411,N_32664,N_33142);
or U34412 (N_34412,N_33675,N_33617);
xor U34413 (N_34413,N_33420,N_33966);
or U34414 (N_34414,N_33900,N_33540);
xnor U34415 (N_34415,N_33938,N_32135);
or U34416 (N_34416,N_33108,N_33552);
nor U34417 (N_34417,N_32807,N_32987);
xnor U34418 (N_34418,N_33192,N_32657);
or U34419 (N_34419,N_32580,N_33212);
and U34420 (N_34420,N_32741,N_33720);
nor U34421 (N_34421,N_33882,N_33748);
nor U34422 (N_34422,N_33324,N_32413);
and U34423 (N_34423,N_32868,N_32528);
or U34424 (N_34424,N_33295,N_33946);
nor U34425 (N_34425,N_32316,N_32705);
and U34426 (N_34426,N_33756,N_32202);
and U34427 (N_34427,N_32653,N_32418);
and U34428 (N_34428,N_33303,N_32760);
nand U34429 (N_34429,N_32618,N_32685);
and U34430 (N_34430,N_32703,N_32975);
or U34431 (N_34431,N_33878,N_33081);
xnor U34432 (N_34432,N_32619,N_33739);
and U34433 (N_34433,N_32089,N_32581);
nor U34434 (N_34434,N_32017,N_33563);
nand U34435 (N_34435,N_33761,N_33485);
and U34436 (N_34436,N_33975,N_33457);
nor U34437 (N_34437,N_32015,N_33388);
xnor U34438 (N_34438,N_32397,N_33182);
xor U34439 (N_34439,N_33113,N_33646);
or U34440 (N_34440,N_33410,N_33492);
nand U34441 (N_34441,N_32967,N_32710);
xnor U34442 (N_34442,N_32284,N_33261);
xnor U34443 (N_34443,N_32461,N_32315);
or U34444 (N_34444,N_32852,N_32434);
xor U34445 (N_34445,N_32151,N_33225);
or U34446 (N_34446,N_33427,N_33045);
xnor U34447 (N_34447,N_33104,N_33660);
xnor U34448 (N_34448,N_32813,N_32772);
and U34449 (N_34449,N_33574,N_32371);
xor U34450 (N_34450,N_32362,N_33673);
and U34451 (N_34451,N_32718,N_32865);
and U34452 (N_34452,N_32448,N_32651);
or U34453 (N_34453,N_33471,N_33004);
nor U34454 (N_34454,N_32163,N_33039);
xnor U34455 (N_34455,N_33451,N_33015);
and U34456 (N_34456,N_33456,N_32402);
nand U34457 (N_34457,N_32248,N_32634);
or U34458 (N_34458,N_33854,N_32263);
nand U34459 (N_34459,N_33498,N_32410);
and U34460 (N_34460,N_33041,N_32600);
and U34461 (N_34461,N_32026,N_32313);
xor U34462 (N_34462,N_32494,N_33935);
and U34463 (N_34463,N_33122,N_33584);
nor U34464 (N_34464,N_33095,N_32570);
or U34465 (N_34465,N_32170,N_33744);
or U34466 (N_34466,N_33269,N_33704);
xor U34467 (N_34467,N_33621,N_32083);
nor U34468 (N_34468,N_32454,N_33415);
nor U34469 (N_34469,N_32322,N_32016);
nor U34470 (N_34470,N_33123,N_32079);
and U34471 (N_34471,N_32431,N_33441);
nor U34472 (N_34472,N_32968,N_32656);
xor U34473 (N_34473,N_33601,N_33896);
and U34474 (N_34474,N_33825,N_33250);
and U34475 (N_34475,N_33256,N_33448);
and U34476 (N_34476,N_33898,N_33982);
nand U34477 (N_34477,N_33931,N_33790);
nor U34478 (N_34478,N_33785,N_33412);
xnor U34479 (N_34479,N_32577,N_33598);
or U34480 (N_34480,N_32535,N_33683);
and U34481 (N_34481,N_32025,N_33901);
nor U34482 (N_34482,N_33043,N_32770);
and U34483 (N_34483,N_33910,N_33024);
and U34484 (N_34484,N_32623,N_33079);
nor U34485 (N_34485,N_33428,N_32297);
nand U34486 (N_34486,N_32850,N_33650);
nand U34487 (N_34487,N_32866,N_33821);
nor U34488 (N_34488,N_33034,N_33361);
and U34489 (N_34489,N_32335,N_32466);
or U34490 (N_34490,N_33458,N_32888);
nand U34491 (N_34491,N_32233,N_33746);
nor U34492 (N_34492,N_32474,N_32648);
or U34493 (N_34493,N_32156,N_32406);
nand U34494 (N_34494,N_32552,N_32549);
and U34495 (N_34495,N_33016,N_33179);
nand U34496 (N_34496,N_33085,N_33023);
or U34497 (N_34497,N_33194,N_32102);
nor U34498 (N_34498,N_33945,N_33877);
nor U34499 (N_34499,N_32388,N_33119);
nor U34500 (N_34500,N_33407,N_32035);
and U34501 (N_34501,N_32385,N_33249);
nand U34502 (N_34502,N_33417,N_32613);
and U34503 (N_34503,N_33692,N_32277);
xor U34504 (N_34504,N_33974,N_33301);
xor U34505 (N_34505,N_32745,N_33522);
nor U34506 (N_34506,N_33545,N_33120);
xor U34507 (N_34507,N_33316,N_32204);
or U34508 (N_34508,N_32553,N_33770);
nor U34509 (N_34509,N_32502,N_32996);
nand U34510 (N_34510,N_32469,N_32056);
nand U34511 (N_34511,N_32393,N_32713);
nand U34512 (N_34512,N_33282,N_32049);
nor U34513 (N_34513,N_33792,N_33491);
xnor U34514 (N_34514,N_32969,N_32429);
xor U34515 (N_34515,N_33864,N_32973);
and U34516 (N_34516,N_33126,N_32701);
or U34517 (N_34517,N_32425,N_33558);
or U34518 (N_34518,N_33594,N_33735);
nand U34519 (N_34519,N_33553,N_32286);
nand U34520 (N_34520,N_33466,N_32172);
nor U34521 (N_34521,N_32187,N_33264);
xor U34522 (N_34522,N_33211,N_33716);
nand U34523 (N_34523,N_32625,N_32148);
xor U34524 (N_34524,N_33718,N_32863);
nand U34525 (N_34525,N_32485,N_32559);
or U34526 (N_34526,N_33813,N_32053);
and U34527 (N_34527,N_32988,N_32302);
xnor U34528 (N_34528,N_32145,N_32939);
xnor U34529 (N_34529,N_33036,N_32805);
nand U34530 (N_34530,N_32189,N_33535);
and U34531 (N_34531,N_32065,N_32881);
xor U34532 (N_34532,N_32341,N_33568);
or U34533 (N_34533,N_33493,N_33765);
nor U34534 (N_34534,N_32925,N_32524);
nor U34535 (N_34535,N_32869,N_32687);
and U34536 (N_34536,N_33406,N_33241);
xor U34537 (N_34537,N_32508,N_32752);
nor U34538 (N_34538,N_33454,N_33932);
nor U34539 (N_34539,N_33231,N_33019);
xor U34540 (N_34540,N_32649,N_33164);
xnor U34541 (N_34541,N_32110,N_32179);
or U34542 (N_34542,N_33838,N_33403);
and U34543 (N_34543,N_33832,N_32931);
or U34544 (N_34544,N_33178,N_33367);
or U34545 (N_34545,N_32671,N_32130);
and U34546 (N_34546,N_32706,N_33300);
xor U34547 (N_34547,N_32169,N_33504);
nand U34548 (N_34548,N_33543,N_33967);
xor U34549 (N_34549,N_32540,N_32966);
nand U34550 (N_34550,N_32105,N_32030);
and U34551 (N_34551,N_33921,N_33751);
or U34552 (N_34552,N_32462,N_33486);
nor U34553 (N_34553,N_33255,N_32762);
nor U34554 (N_34554,N_32569,N_33796);
and U34555 (N_34555,N_33637,N_33442);
and U34556 (N_34556,N_33246,N_33317);
and U34557 (N_34557,N_32142,N_32561);
or U34558 (N_34558,N_33010,N_33483);
xnor U34559 (N_34559,N_32773,N_32157);
xnor U34560 (N_34560,N_33278,N_33337);
xor U34561 (N_34561,N_33350,N_32578);
and U34562 (N_34562,N_32117,N_33538);
xor U34563 (N_34563,N_32363,N_32847);
xnor U34564 (N_34564,N_32310,N_32827);
xnor U34565 (N_34565,N_32901,N_32299);
nor U34566 (N_34566,N_33830,N_32723);
xor U34567 (N_34567,N_32880,N_33602);
or U34568 (N_34568,N_33666,N_33641);
or U34569 (N_34569,N_32533,N_33708);
nand U34570 (N_34570,N_33871,N_33848);
nor U34571 (N_34571,N_33460,N_32539);
or U34572 (N_34572,N_33443,N_33826);
and U34573 (N_34573,N_33670,N_33068);
nor U34574 (N_34574,N_32704,N_32039);
and U34575 (N_34575,N_33109,N_33482);
nor U34576 (N_34576,N_32953,N_32617);
and U34577 (N_34577,N_32450,N_32269);
and U34578 (N_34578,N_32481,N_32546);
or U34579 (N_34579,N_33628,N_32591);
nor U34580 (N_34580,N_33999,N_33204);
nand U34581 (N_34581,N_32021,N_32218);
nand U34582 (N_34582,N_32775,N_32432);
nor U34583 (N_34583,N_33190,N_32800);
and U34584 (N_34584,N_33799,N_32794);
and U34585 (N_34585,N_33323,N_32952);
xnor U34586 (N_34586,N_32358,N_32396);
xnor U34587 (N_34587,N_32734,N_32943);
and U34588 (N_34588,N_33541,N_33141);
nor U34589 (N_34589,N_32368,N_32899);
or U34590 (N_34590,N_33144,N_33679);
or U34591 (N_34591,N_32282,N_33131);
nand U34592 (N_34592,N_33501,N_32817);
xnor U34593 (N_34593,N_33258,N_32288);
nand U34594 (N_34594,N_32127,N_33002);
xor U34595 (N_34595,N_33499,N_32735);
xor U34596 (N_34596,N_32011,N_33327);
xor U34597 (N_34597,N_32832,N_32730);
xnor U34598 (N_34598,N_32512,N_32538);
or U34599 (N_34599,N_33705,N_33253);
and U34600 (N_34600,N_32904,N_32903);
nor U34601 (N_34601,N_33091,N_32034);
and U34602 (N_34602,N_33923,N_32915);
or U34603 (N_34603,N_32921,N_32162);
nor U34604 (N_34604,N_32781,N_32192);
and U34605 (N_34605,N_32961,N_32963);
and U34606 (N_34606,N_32970,N_32855);
and U34607 (N_34607,N_32799,N_33385);
or U34608 (N_34608,N_33993,N_32236);
nand U34609 (N_34609,N_32223,N_33148);
nand U34610 (N_34610,N_33198,N_33940);
nor U34611 (N_34611,N_32377,N_32937);
nand U34612 (N_34612,N_32076,N_33738);
nor U34613 (N_34613,N_32629,N_32550);
nor U34614 (N_34614,N_33121,N_32956);
xnor U34615 (N_34615,N_33807,N_33607);
and U34616 (N_34616,N_33771,N_33446);
xor U34617 (N_34617,N_32909,N_33768);
nand U34618 (N_34618,N_32732,N_33283);
nor U34619 (N_34619,N_33800,N_32100);
nor U34620 (N_34620,N_32408,N_32642);
nor U34621 (N_34621,N_32798,N_32249);
nor U34622 (N_34622,N_32493,N_33450);
nand U34623 (N_34623,N_32499,N_32212);
nor U34624 (N_34624,N_33248,N_33050);
nor U34625 (N_34625,N_32680,N_32630);
nor U34626 (N_34626,N_32171,N_33093);
or U34627 (N_34627,N_32314,N_32911);
nor U34628 (N_34628,N_33154,N_32806);
and U34629 (N_34629,N_33462,N_33913);
nand U34630 (N_34630,N_32354,N_33943);
nand U34631 (N_34631,N_33218,N_33394);
or U34632 (N_34632,N_32517,N_33651);
nor U34633 (N_34633,N_32947,N_32003);
nand U34634 (N_34634,N_33197,N_33723);
and U34635 (N_34635,N_32840,N_33787);
and U34636 (N_34636,N_32906,N_32690);
or U34637 (N_34637,N_32333,N_33489);
xnor U34638 (N_34638,N_33333,N_32726);
or U34639 (N_34639,N_33852,N_32940);
or U34640 (N_34640,N_32573,N_32445);
nor U34641 (N_34641,N_33681,N_33884);
nand U34642 (N_34642,N_32824,N_32562);
or U34643 (N_34643,N_32586,N_33129);
nand U34644 (N_34644,N_32134,N_33903);
or U34645 (N_34645,N_33098,N_32841);
xnor U34646 (N_34646,N_32823,N_33112);
xnor U34647 (N_34647,N_32886,N_33058);
and U34648 (N_34648,N_33030,N_33784);
or U34649 (N_34649,N_32018,N_33055);
and U34650 (N_34650,N_33005,N_33294);
nand U34651 (N_34651,N_33763,N_32473);
and U34652 (N_34652,N_32932,N_32889);
nor U34653 (N_34653,N_32606,N_32796);
nand U34654 (N_34654,N_33653,N_32883);
xnor U34655 (N_34655,N_33338,N_33076);
xnor U34656 (N_34656,N_33868,N_32922);
nor U34657 (N_34657,N_33870,N_33151);
and U34658 (N_34658,N_33426,N_32122);
nand U34659 (N_34659,N_33227,N_32596);
xor U34660 (N_34660,N_32985,N_33992);
xor U34661 (N_34661,N_32662,N_33634);
nand U34662 (N_34662,N_32007,N_33831);
nor U34663 (N_34663,N_32488,N_33595);
xor U34664 (N_34664,N_33459,N_32989);
xnor U34665 (N_34665,N_33642,N_33340);
nor U34666 (N_34666,N_33044,N_33506);
and U34667 (N_34667,N_32433,N_32521);
nor U34668 (N_34668,N_33398,N_32659);
and U34669 (N_34669,N_32505,N_33528);
nand U34670 (N_34670,N_33185,N_32329);
or U34671 (N_34671,N_32069,N_32811);
nand U34672 (N_34672,N_33176,N_33671);
and U34673 (N_34673,N_33665,N_33902);
or U34674 (N_34674,N_32712,N_32386);
and U34675 (N_34675,N_33243,N_32374);
nand U34676 (N_34676,N_32325,N_32320);
xnor U34677 (N_34677,N_33707,N_33863);
nand U34678 (N_34678,N_33124,N_32265);
xnor U34679 (N_34679,N_32317,N_33308);
and U34680 (N_34680,N_33128,N_32051);
xnor U34681 (N_34681,N_33758,N_33180);
nand U34682 (N_34682,N_33082,N_32820);
nor U34683 (N_34683,N_33170,N_33186);
xor U34684 (N_34684,N_33688,N_33157);
nand U34685 (N_34685,N_33111,N_32608);
nor U34686 (N_34686,N_33257,N_32788);
or U34687 (N_34687,N_33562,N_32575);
xor U34688 (N_34688,N_32126,N_32389);
nand U34689 (N_34689,N_32042,N_33214);
or U34690 (N_34690,N_33696,N_33276);
and U34691 (N_34691,N_33497,N_32470);
and U34692 (N_34692,N_32144,N_32572);
and U34693 (N_34693,N_32496,N_33611);
or U34694 (N_34694,N_32022,N_33845);
nand U34695 (N_34695,N_32219,N_33623);
nor U34696 (N_34696,N_32001,N_32698);
or U34697 (N_34697,N_32804,N_32955);
and U34698 (N_34698,N_32417,N_32944);
or U34699 (N_34699,N_33984,N_33117);
and U34700 (N_34700,N_33409,N_32557);
xor U34701 (N_34701,N_33200,N_32834);
xnor U34702 (N_34702,N_33893,N_32790);
nor U34703 (N_34703,N_32380,N_32063);
xor U34704 (N_34704,N_32551,N_33228);
nand U34705 (N_34705,N_32340,N_33321);
xor U34706 (N_34706,N_32099,N_33387);
nor U34707 (N_34707,N_33585,N_32191);
or U34708 (N_34708,N_32342,N_32482);
xnor U34709 (N_34709,N_33507,N_33837);
nand U34710 (N_34710,N_33487,N_33379);
or U34711 (N_34711,N_32279,N_33237);
xor U34712 (N_34712,N_33786,N_33626);
and U34713 (N_34713,N_32511,N_32891);
and U34714 (N_34714,N_32471,N_33542);
nand U34715 (N_34715,N_32104,N_33905);
nand U34716 (N_34716,N_32029,N_33137);
nor U34717 (N_34717,N_32456,N_32870);
or U34718 (N_34718,N_32890,N_33872);
or U34719 (N_34719,N_33090,N_32009);
nor U34720 (N_34720,N_32128,N_33371);
nand U34721 (N_34721,N_33614,N_32984);
nand U34722 (N_34722,N_33425,N_32280);
xnor U34723 (N_34723,N_33732,N_33274);
and U34724 (N_34724,N_32532,N_32250);
and U34725 (N_34725,N_32036,N_33382);
and U34726 (N_34726,N_33834,N_33221);
nor U34727 (N_34727,N_33581,N_32981);
and U34728 (N_34728,N_32213,N_32742);
xor U34729 (N_34729,N_33234,N_32261);
nand U34730 (N_34730,N_32789,N_33074);
and U34731 (N_34731,N_33447,N_33001);
nand U34732 (N_34732,N_33509,N_32479);
nor U34733 (N_34733,N_32507,N_33488);
nor U34734 (N_34734,N_32347,N_32419);
xnor U34735 (N_34735,N_32020,N_33286);
xnor U34736 (N_34736,N_33933,N_33217);
or U34737 (N_34737,N_33866,N_32242);
nor U34738 (N_34738,N_33110,N_32253);
or U34739 (N_34739,N_33697,N_32113);
and U34740 (N_34740,N_32905,N_32744);
nor U34741 (N_34741,N_32423,N_32949);
or U34742 (N_34742,N_32542,N_33762);
nand U34743 (N_34743,N_33840,N_32057);
nor U34744 (N_34744,N_33376,N_32058);
nor U34745 (N_34745,N_33694,N_33662);
or U34746 (N_34746,N_32556,N_32908);
nor U34747 (N_34747,N_32459,N_32689);
nand U34748 (N_34748,N_33897,N_32031);
and U34749 (N_34749,N_33668,N_33463);
or U34750 (N_34750,N_32784,N_33158);
nand U34751 (N_34751,N_32492,N_32033);
and U34752 (N_34752,N_32181,N_33242);
nor U34753 (N_34753,N_33165,N_32008);
and U34754 (N_34754,N_33314,N_32467);
nor U34755 (N_34755,N_33299,N_32103);
nor U34756 (N_34756,N_33056,N_33025);
nand U34757 (N_34757,N_32589,N_33546);
or U34758 (N_34758,N_33843,N_32564);
or U34759 (N_34759,N_32326,N_33500);
xor U34760 (N_34760,N_33955,N_33244);
and U34761 (N_34761,N_33084,N_32464);
nand U34762 (N_34762,N_33481,N_32610);
nand U34763 (N_34763,N_32795,N_33088);
nand U34764 (N_34764,N_32205,N_32375);
nand U34765 (N_34765,N_32622,N_33101);
nor U34766 (N_34766,N_32980,N_32240);
xor U34767 (N_34767,N_33772,N_33706);
and U34768 (N_34768,N_33520,N_33461);
or U34769 (N_34769,N_32861,N_33561);
nor U34770 (N_34770,N_32829,N_32655);
and U34771 (N_34771,N_32289,N_33260);
nor U34772 (N_34772,N_32753,N_33608);
nor U34773 (N_34773,N_33092,N_32715);
xor U34774 (N_34774,N_33020,N_32411);
nor U34775 (N_34775,N_33914,N_33846);
or U34776 (N_34776,N_32954,N_33548);
xnor U34777 (N_34777,N_33855,N_32835);
and U34778 (N_34778,N_32193,N_32478);
xnor U34779 (N_34779,N_33847,N_32256);
or U34780 (N_34780,N_32119,N_33615);
xnor U34781 (N_34781,N_33695,N_33116);
or U34782 (N_34782,N_33894,N_33348);
and U34783 (N_34783,N_32229,N_33740);
nand U34784 (N_34784,N_33835,N_32298);
or U34785 (N_34785,N_32059,N_32131);
nor U34786 (N_34786,N_33390,N_32825);
or U34787 (N_34787,N_33578,N_33779);
xnor U34788 (N_34788,N_33976,N_33254);
xor U34789 (N_34789,N_32948,N_32616);
xor U34790 (N_34790,N_32974,N_32992);
nand U34791 (N_34791,N_33434,N_32545);
and U34792 (N_34792,N_33168,N_32633);
nand U34793 (N_34793,N_32449,N_33819);
or U34794 (N_34794,N_33445,N_33479);
nand U34795 (N_34795,N_32864,N_32628);
xnor U34796 (N_34796,N_32356,N_33750);
nand U34797 (N_34797,N_33599,N_32751);
or U34798 (N_34798,N_33776,N_33401);
nand U34799 (N_34799,N_33577,N_33721);
nor U34800 (N_34800,N_32802,N_33012);
and U34801 (N_34801,N_33547,N_32109);
nor U34802 (N_34802,N_33616,N_33293);
nor U34803 (N_34803,N_32198,N_32950);
nor U34804 (N_34804,N_33851,N_32194);
nand U34805 (N_34805,N_33961,N_33689);
xor U34806 (N_34806,N_32262,N_32769);
nand U34807 (N_34807,N_32132,N_32447);
nand U34808 (N_34808,N_33431,N_33957);
or U34809 (N_34809,N_32334,N_32238);
nand U34810 (N_34810,N_33968,N_33639);
or U34811 (N_34811,N_32351,N_33891);
and U34812 (N_34812,N_32604,N_33145);
and U34813 (N_34813,N_32812,N_33035);
xnor U34814 (N_34814,N_32005,N_33469);
xor U34815 (N_34815,N_32748,N_33610);
nor U34816 (N_34816,N_33439,N_33022);
nor U34817 (N_34817,N_32977,N_33026);
nor U34818 (N_34818,N_33888,N_32924);
and U34819 (N_34819,N_32258,N_32045);
nor U34820 (N_34820,N_32227,N_33815);
or U34821 (N_34821,N_33606,N_32220);
and U34822 (N_34822,N_32590,N_32081);
nand U34823 (N_34823,N_33222,N_32914);
nor U34824 (N_34824,N_33795,N_33654);
nand U34825 (N_34825,N_32092,N_32472);
or U34826 (N_34826,N_32178,N_32844);
nand U34827 (N_34827,N_33638,N_32716);
xor U34828 (N_34828,N_32037,N_32185);
nand U34829 (N_34829,N_33717,N_33339);
and U34830 (N_34830,N_33649,N_33760);
and U34831 (N_34831,N_32670,N_33571);
xor U34832 (N_34832,N_32424,N_32830);
and U34833 (N_34833,N_33437,N_33149);
nor U34834 (N_34834,N_32278,N_33196);
and U34835 (N_34835,N_33251,N_33014);
and U34836 (N_34836,N_32763,N_33924);
or U34837 (N_34837,N_33536,N_32541);
nor U34838 (N_34838,N_33040,N_32247);
xnor U34839 (N_34839,N_32815,N_32757);
or U34840 (N_34840,N_33861,N_32077);
nand U34841 (N_34841,N_33597,N_33816);
xnor U34842 (N_34842,N_32002,N_32758);
xnor U34843 (N_34843,N_33199,N_33477);
xor U34844 (N_34844,N_33206,N_33526);
and U34845 (N_34845,N_32579,N_33354);
and U34846 (N_34846,N_33018,N_33930);
or U34847 (N_34847,N_33438,N_33468);
nor U34848 (N_34848,N_32525,N_33609);
nor U34849 (N_34849,N_32583,N_32879);
nor U34850 (N_34850,N_33817,N_33566);
xnor U34851 (N_34851,N_33147,N_33952);
nand U34852 (N_34852,N_33769,N_32460);
nand U34853 (N_34853,N_33532,N_33814);
nand U34854 (N_34854,N_33230,N_33912);
xor U34855 (N_34855,N_33909,N_33753);
and U34856 (N_34856,N_33172,N_32995);
and U34857 (N_34857,N_32958,N_33310);
and U34858 (N_34858,N_32765,N_32064);
nor U34859 (N_34859,N_32746,N_33245);
and U34860 (N_34860,N_32681,N_32990);
nand U34861 (N_34861,N_32041,N_32346);
or U34862 (N_34862,N_32946,N_33774);
nor U34863 (N_34863,N_33711,N_33177);
nand U34864 (N_34864,N_33987,N_32463);
and U34865 (N_34865,N_33495,N_32658);
xnor U34866 (N_34866,N_32010,N_32917);
and U34867 (N_34867,N_33892,N_33331);
or U34868 (N_34868,N_33003,N_32361);
xnor U34869 (N_34869,N_33356,N_33032);
xnor U34870 (N_34870,N_32907,N_32683);
or U34871 (N_34871,N_33991,N_32457);
nor U34872 (N_34872,N_32654,N_32691);
or U34873 (N_34873,N_32860,N_32621);
and U34874 (N_34874,N_32877,N_33313);
and U34875 (N_34875,N_33582,N_32324);
nand U34876 (N_34876,N_32436,N_32121);
xnor U34877 (N_34877,N_32743,N_32206);
nand U34878 (N_34878,N_33948,N_33127);
or U34879 (N_34879,N_32665,N_32766);
nor U34880 (N_34880,N_33981,N_32679);
nor U34881 (N_34881,N_33311,N_33187);
nor U34882 (N_34882,N_33880,N_32643);
nand U34883 (N_34883,N_32668,N_32897);
nand U34884 (N_34884,N_32143,N_32702);
xor U34885 (N_34885,N_32663,N_33531);
and U34886 (N_34886,N_32345,N_32200);
or U34887 (N_34887,N_32453,N_32216);
xor U34888 (N_34888,N_32754,N_32446);
xor U34889 (N_34889,N_33856,N_33569);
nand U34890 (N_34890,N_32095,N_32096);
and U34891 (N_34891,N_32534,N_33633);
xor U34892 (N_34892,N_33047,N_33133);
and U34893 (N_34893,N_32228,N_32736);
nand U34894 (N_34894,N_33737,N_32729);
nand U34895 (N_34895,N_33958,N_33820);
or U34896 (N_34896,N_32592,N_33844);
nor U34897 (N_34897,N_32139,N_32052);
nor U34898 (N_34898,N_33778,N_32737);
or U34899 (N_34899,N_33580,N_33031);
nand U34900 (N_34900,N_32601,N_32210);
nand U34901 (N_34901,N_32913,N_32919);
or U34902 (N_34902,N_32073,N_32239);
xor U34903 (N_34903,N_33239,N_32328);
and U34904 (N_34904,N_33978,N_33809);
nor U34905 (N_34905,N_32615,N_33476);
or U34906 (N_34906,N_33742,N_33890);
and U34907 (N_34907,N_33533,N_33700);
and U34908 (N_34908,N_32998,N_32635);
nor U34909 (N_34909,N_32566,N_33937);
nand U34910 (N_34910,N_32338,N_33747);
or U34911 (N_34911,N_33624,N_33163);
nand U34912 (N_34912,N_32243,N_33977);
xor U34913 (N_34913,N_33173,N_32548);
and U34914 (N_34914,N_33360,N_33764);
and U34915 (N_34915,N_32087,N_33712);
xnor U34916 (N_34916,N_32395,N_33575);
and U34917 (N_34917,N_33220,N_32367);
nor U34918 (N_34918,N_33627,N_33869);
xnor U34919 (N_34919,N_32364,N_32647);
nand U34920 (N_34920,N_32292,N_32415);
nor U34921 (N_34921,N_33130,N_32688);
and U34922 (N_34922,N_33908,N_32547);
and U34923 (N_34923,N_32894,N_32106);
nand U34924 (N_34924,N_32786,N_33094);
xnor U34925 (N_34925,N_32168,N_32896);
and U34926 (N_34926,N_32791,N_32708);
nand U34927 (N_34927,N_33922,N_32038);
xor U34928 (N_34928,N_32571,N_32991);
xor U34929 (N_34929,N_32199,N_32516);
and U34930 (N_34930,N_32012,N_32819);
or U34931 (N_34931,N_33453,N_33730);
nand U34932 (N_34932,N_32241,N_33849);
or U34933 (N_34933,N_33631,N_32071);
nand U34934 (N_34934,N_32537,N_33272);
nor U34935 (N_34935,N_33359,N_32612);
nand U34936 (N_34936,N_32066,N_32979);
nor U34937 (N_34937,N_33949,N_32599);
nand U34938 (N_34938,N_33793,N_33341);
or U34939 (N_34939,N_33080,N_33063);
or U34940 (N_34940,N_33009,N_33652);
and U34941 (N_34941,N_32084,N_33988);
and U34942 (N_34942,N_32028,N_32588);
xnor U34943 (N_34943,N_32296,N_32188);
or U34944 (N_34944,N_32740,N_33305);
nand U34945 (N_34945,N_32176,N_33956);
or U34946 (N_34946,N_33021,N_32155);
nor U34947 (N_34947,N_32611,N_32490);
or U34948 (N_34948,N_33505,N_33920);
nor U34949 (N_34949,N_32684,N_32088);
and U34950 (N_34950,N_33329,N_33078);
and U34951 (N_34951,N_32384,N_33086);
nor U34952 (N_34952,N_33812,N_32874);
and U34953 (N_34953,N_32898,N_32295);
or U34954 (N_34954,N_32400,N_32390);
nand U34955 (N_34955,N_33619,N_33702);
nor U34956 (N_34956,N_32231,N_33664);
nand U34957 (N_34957,N_32738,N_33867);
xnor U34958 (N_34958,N_33358,N_33648);
and U34959 (N_34959,N_33416,N_32678);
or U34960 (N_34960,N_32224,N_32582);
and U34961 (N_34961,N_32895,N_32468);
nor U34962 (N_34962,N_32308,N_32783);
xnor U34963 (N_34963,N_33734,N_32019);
or U34964 (N_34964,N_33728,N_33060);
nand U34965 (N_34965,N_32154,N_32602);
and U34966 (N_34966,N_32266,N_33586);
nand U34967 (N_34967,N_32720,N_33399);
nand U34968 (N_34968,N_32767,N_33162);
nand U34969 (N_34969,N_32558,N_32392);
and U34970 (N_34970,N_33344,N_32731);
or U34971 (N_34971,N_32412,N_33557);
or U34972 (N_34972,N_32853,N_32387);
xnor U34973 (N_34973,N_33422,N_32486);
nor U34974 (N_34974,N_32506,N_33936);
xnor U34975 (N_34975,N_33971,N_32902);
and U34976 (N_34976,N_33995,N_32779);
or U34977 (N_34977,N_33841,N_33352);
xor U34978 (N_34978,N_32934,N_32060);
and U34979 (N_34979,N_33266,N_33475);
xnor U34980 (N_34980,N_32774,N_33135);
nand U34981 (N_34981,N_33928,N_32050);
xor U34982 (N_34982,N_33635,N_32697);
xor U34983 (N_34983,N_33959,N_32565);
nor U34984 (N_34984,N_33066,N_33188);
or U34985 (N_34985,N_32750,N_32639);
nor U34986 (N_34986,N_32321,N_32428);
or U34987 (N_34987,N_33281,N_32136);
xor U34988 (N_34988,N_33363,N_32887);
xor U34989 (N_34989,N_32707,N_33318);
nand U34990 (N_34990,N_33791,N_33105);
or U34991 (N_34991,N_33613,N_33544);
xor U34992 (N_34992,N_33811,N_32370);
or U34993 (N_34993,N_33319,N_33985);
nand U34994 (N_34994,N_32982,N_32167);
and U34995 (N_34995,N_32650,N_33315);
nor U34996 (N_34996,N_32595,N_32455);
and U34997 (N_34997,N_32044,N_33362);
or U34998 (N_34998,N_32405,N_32724);
nand U34999 (N_34999,N_32133,N_32048);
nor U35000 (N_35000,N_32772,N_32814);
nand U35001 (N_35001,N_32284,N_33052);
or U35002 (N_35002,N_32472,N_32775);
and U35003 (N_35003,N_32492,N_33941);
nor U35004 (N_35004,N_33701,N_32923);
nand U35005 (N_35005,N_32638,N_32233);
xnor U35006 (N_35006,N_33321,N_32864);
and U35007 (N_35007,N_33958,N_33239);
xnor U35008 (N_35008,N_32908,N_32724);
or U35009 (N_35009,N_32059,N_33800);
xor U35010 (N_35010,N_33740,N_32453);
nand U35011 (N_35011,N_32660,N_32862);
xor U35012 (N_35012,N_32766,N_32564);
and U35013 (N_35013,N_32726,N_32691);
and U35014 (N_35014,N_32011,N_33577);
xnor U35015 (N_35015,N_33210,N_33536);
xnor U35016 (N_35016,N_33752,N_33142);
nor U35017 (N_35017,N_32325,N_32149);
and U35018 (N_35018,N_32520,N_32101);
and U35019 (N_35019,N_33880,N_32665);
nand U35020 (N_35020,N_32290,N_33770);
and U35021 (N_35021,N_33248,N_33241);
nor U35022 (N_35022,N_32384,N_33792);
and U35023 (N_35023,N_32800,N_32646);
and U35024 (N_35024,N_32403,N_32457);
nand U35025 (N_35025,N_32186,N_32555);
nor U35026 (N_35026,N_32666,N_33149);
or U35027 (N_35027,N_33863,N_33519);
nor U35028 (N_35028,N_33298,N_32202);
nand U35029 (N_35029,N_32370,N_32186);
nand U35030 (N_35030,N_33944,N_32391);
nor U35031 (N_35031,N_32746,N_32908);
or U35032 (N_35032,N_33832,N_33523);
nor U35033 (N_35033,N_33017,N_33041);
and U35034 (N_35034,N_33541,N_33456);
and U35035 (N_35035,N_33993,N_32393);
or U35036 (N_35036,N_32791,N_32768);
or U35037 (N_35037,N_32794,N_33124);
and U35038 (N_35038,N_33295,N_33518);
nor U35039 (N_35039,N_32834,N_33895);
nand U35040 (N_35040,N_33415,N_33975);
xor U35041 (N_35041,N_32540,N_33353);
nor U35042 (N_35042,N_32137,N_33751);
or U35043 (N_35043,N_32405,N_32296);
nor U35044 (N_35044,N_33788,N_32888);
or U35045 (N_35045,N_32847,N_32493);
xnor U35046 (N_35046,N_33117,N_33628);
and U35047 (N_35047,N_32191,N_32337);
nand U35048 (N_35048,N_33589,N_33804);
nor U35049 (N_35049,N_32742,N_32402);
or U35050 (N_35050,N_32980,N_32158);
xor U35051 (N_35051,N_32273,N_32175);
and U35052 (N_35052,N_33084,N_32191);
xor U35053 (N_35053,N_32792,N_32298);
xor U35054 (N_35054,N_33866,N_32364);
nor U35055 (N_35055,N_32525,N_32821);
xnor U35056 (N_35056,N_33958,N_33879);
nor U35057 (N_35057,N_33577,N_32775);
and U35058 (N_35058,N_32115,N_32722);
or U35059 (N_35059,N_33768,N_32916);
nor U35060 (N_35060,N_33215,N_32664);
and U35061 (N_35061,N_32353,N_33054);
xnor U35062 (N_35062,N_32397,N_32136);
or U35063 (N_35063,N_32933,N_33482);
and U35064 (N_35064,N_33419,N_32425);
nand U35065 (N_35065,N_32941,N_33703);
nor U35066 (N_35066,N_33413,N_33330);
nor U35067 (N_35067,N_32915,N_32199);
xor U35068 (N_35068,N_33508,N_32888);
nor U35069 (N_35069,N_32861,N_32687);
nand U35070 (N_35070,N_32072,N_32561);
xnor U35071 (N_35071,N_32825,N_33577);
and U35072 (N_35072,N_32616,N_32831);
nand U35073 (N_35073,N_32200,N_32322);
xnor U35074 (N_35074,N_32749,N_33409);
and U35075 (N_35075,N_33064,N_33560);
and U35076 (N_35076,N_33672,N_32600);
nand U35077 (N_35077,N_33335,N_33778);
or U35078 (N_35078,N_33059,N_33604);
and U35079 (N_35079,N_33784,N_32262);
nor U35080 (N_35080,N_32681,N_32502);
or U35081 (N_35081,N_32299,N_32872);
or U35082 (N_35082,N_33774,N_33150);
and U35083 (N_35083,N_33524,N_32911);
nor U35084 (N_35084,N_33313,N_33600);
nand U35085 (N_35085,N_32249,N_33803);
and U35086 (N_35086,N_32457,N_32058);
nand U35087 (N_35087,N_32934,N_32008);
xnor U35088 (N_35088,N_32740,N_32952);
xnor U35089 (N_35089,N_32061,N_33113);
nand U35090 (N_35090,N_33112,N_33730);
nor U35091 (N_35091,N_33453,N_33411);
and U35092 (N_35092,N_33056,N_33694);
nor U35093 (N_35093,N_33170,N_33124);
nand U35094 (N_35094,N_33891,N_33506);
and U35095 (N_35095,N_32868,N_33401);
or U35096 (N_35096,N_32963,N_32587);
xor U35097 (N_35097,N_32940,N_33940);
or U35098 (N_35098,N_32581,N_32969);
or U35099 (N_35099,N_32931,N_33693);
xor U35100 (N_35100,N_32191,N_33671);
or U35101 (N_35101,N_32729,N_32028);
or U35102 (N_35102,N_33450,N_32141);
xor U35103 (N_35103,N_32189,N_33855);
or U35104 (N_35104,N_32398,N_33203);
nor U35105 (N_35105,N_32738,N_32260);
nand U35106 (N_35106,N_32284,N_32247);
xnor U35107 (N_35107,N_32542,N_32807);
xnor U35108 (N_35108,N_32807,N_32918);
xnor U35109 (N_35109,N_33095,N_33050);
and U35110 (N_35110,N_33767,N_32339);
nand U35111 (N_35111,N_32879,N_32420);
or U35112 (N_35112,N_32366,N_33230);
or U35113 (N_35113,N_33882,N_32116);
and U35114 (N_35114,N_32892,N_33810);
nor U35115 (N_35115,N_33346,N_33508);
nor U35116 (N_35116,N_33195,N_32716);
and U35117 (N_35117,N_33011,N_32997);
or U35118 (N_35118,N_33327,N_32253);
xnor U35119 (N_35119,N_33020,N_32333);
nor U35120 (N_35120,N_32850,N_32039);
nor U35121 (N_35121,N_33858,N_32379);
or U35122 (N_35122,N_32455,N_32859);
nor U35123 (N_35123,N_33730,N_33530);
nor U35124 (N_35124,N_32344,N_32572);
and U35125 (N_35125,N_33775,N_32557);
or U35126 (N_35126,N_32167,N_33202);
xor U35127 (N_35127,N_33950,N_32861);
and U35128 (N_35128,N_32591,N_33511);
and U35129 (N_35129,N_33403,N_32140);
xor U35130 (N_35130,N_32443,N_32958);
nor U35131 (N_35131,N_33793,N_33589);
nand U35132 (N_35132,N_33809,N_32690);
nor U35133 (N_35133,N_32415,N_33871);
nor U35134 (N_35134,N_32140,N_32514);
nand U35135 (N_35135,N_32004,N_32501);
xor U35136 (N_35136,N_33366,N_32105);
and U35137 (N_35137,N_32327,N_32466);
or U35138 (N_35138,N_32093,N_32704);
or U35139 (N_35139,N_33847,N_33831);
or U35140 (N_35140,N_33649,N_32141);
nand U35141 (N_35141,N_32694,N_33428);
nor U35142 (N_35142,N_32588,N_32030);
nand U35143 (N_35143,N_33478,N_33489);
nor U35144 (N_35144,N_32989,N_33828);
nand U35145 (N_35145,N_32367,N_32253);
nor U35146 (N_35146,N_32818,N_32333);
and U35147 (N_35147,N_32725,N_32703);
and U35148 (N_35148,N_32354,N_32913);
nand U35149 (N_35149,N_33720,N_32991);
and U35150 (N_35150,N_33239,N_33675);
nand U35151 (N_35151,N_33395,N_33833);
or U35152 (N_35152,N_32937,N_33018);
xnor U35153 (N_35153,N_32670,N_32895);
and U35154 (N_35154,N_32397,N_33653);
or U35155 (N_35155,N_33811,N_33908);
and U35156 (N_35156,N_32795,N_32003);
nand U35157 (N_35157,N_33825,N_33339);
and U35158 (N_35158,N_32253,N_32209);
and U35159 (N_35159,N_33911,N_32965);
nand U35160 (N_35160,N_32352,N_33475);
xor U35161 (N_35161,N_33242,N_33275);
nor U35162 (N_35162,N_33807,N_32212);
xnor U35163 (N_35163,N_33600,N_33283);
and U35164 (N_35164,N_32365,N_33646);
or U35165 (N_35165,N_33715,N_33940);
nand U35166 (N_35166,N_32799,N_33526);
and U35167 (N_35167,N_33375,N_32432);
xnor U35168 (N_35168,N_33829,N_33737);
nand U35169 (N_35169,N_32925,N_33221);
nand U35170 (N_35170,N_33871,N_32412);
xor U35171 (N_35171,N_32359,N_33644);
or U35172 (N_35172,N_32468,N_32781);
and U35173 (N_35173,N_33436,N_33854);
xnor U35174 (N_35174,N_32207,N_33735);
xor U35175 (N_35175,N_33484,N_33357);
nor U35176 (N_35176,N_33825,N_32784);
nor U35177 (N_35177,N_33451,N_32905);
and U35178 (N_35178,N_33361,N_33853);
or U35179 (N_35179,N_33261,N_33897);
nand U35180 (N_35180,N_33383,N_33632);
nor U35181 (N_35181,N_32537,N_32996);
and U35182 (N_35182,N_32299,N_33019);
nand U35183 (N_35183,N_32587,N_33302);
nand U35184 (N_35184,N_32870,N_33796);
nor U35185 (N_35185,N_32262,N_32695);
nor U35186 (N_35186,N_33980,N_32672);
xnor U35187 (N_35187,N_33475,N_33510);
nor U35188 (N_35188,N_33822,N_33145);
and U35189 (N_35189,N_33525,N_33954);
or U35190 (N_35190,N_33652,N_33644);
and U35191 (N_35191,N_32830,N_32892);
or U35192 (N_35192,N_33182,N_32671);
xor U35193 (N_35193,N_32086,N_32974);
nand U35194 (N_35194,N_33583,N_32533);
nand U35195 (N_35195,N_33831,N_32824);
nand U35196 (N_35196,N_32355,N_33438);
and U35197 (N_35197,N_32935,N_33286);
nor U35198 (N_35198,N_32490,N_32226);
and U35199 (N_35199,N_33146,N_33700);
nand U35200 (N_35200,N_32543,N_33136);
nand U35201 (N_35201,N_32437,N_32813);
xnor U35202 (N_35202,N_32422,N_32636);
or U35203 (N_35203,N_33709,N_32652);
or U35204 (N_35204,N_33296,N_33966);
nand U35205 (N_35205,N_32668,N_33992);
xnor U35206 (N_35206,N_33883,N_33642);
xor U35207 (N_35207,N_32915,N_32023);
or U35208 (N_35208,N_33139,N_33793);
and U35209 (N_35209,N_32667,N_33174);
xnor U35210 (N_35210,N_33852,N_33891);
xnor U35211 (N_35211,N_33510,N_32510);
nor U35212 (N_35212,N_33560,N_33031);
nor U35213 (N_35213,N_33842,N_33962);
or U35214 (N_35214,N_33467,N_33801);
nand U35215 (N_35215,N_33047,N_33306);
nor U35216 (N_35216,N_33886,N_32802);
xnor U35217 (N_35217,N_33898,N_32161);
nand U35218 (N_35218,N_33379,N_33277);
xnor U35219 (N_35219,N_33661,N_32974);
and U35220 (N_35220,N_32201,N_32510);
nor U35221 (N_35221,N_32053,N_32523);
xor U35222 (N_35222,N_33779,N_33522);
or U35223 (N_35223,N_32382,N_32869);
or U35224 (N_35224,N_33191,N_32589);
or U35225 (N_35225,N_32600,N_32835);
and U35226 (N_35226,N_32438,N_33420);
and U35227 (N_35227,N_32183,N_32546);
and U35228 (N_35228,N_33810,N_32438);
xor U35229 (N_35229,N_32396,N_32083);
nand U35230 (N_35230,N_33550,N_32885);
xor U35231 (N_35231,N_32923,N_32384);
or U35232 (N_35232,N_32376,N_32756);
and U35233 (N_35233,N_32286,N_32540);
nand U35234 (N_35234,N_33148,N_33103);
and U35235 (N_35235,N_33950,N_32586);
or U35236 (N_35236,N_32875,N_32884);
and U35237 (N_35237,N_32346,N_32668);
nor U35238 (N_35238,N_32185,N_32253);
or U35239 (N_35239,N_32500,N_32818);
and U35240 (N_35240,N_33646,N_33266);
nor U35241 (N_35241,N_32436,N_32913);
xor U35242 (N_35242,N_32764,N_32193);
nand U35243 (N_35243,N_33362,N_32724);
or U35244 (N_35244,N_32447,N_33031);
or U35245 (N_35245,N_32581,N_32905);
nand U35246 (N_35246,N_32325,N_32078);
or U35247 (N_35247,N_33980,N_32405);
xnor U35248 (N_35248,N_32329,N_33788);
nor U35249 (N_35249,N_32566,N_33396);
and U35250 (N_35250,N_33942,N_32217);
xor U35251 (N_35251,N_32520,N_32519);
nor U35252 (N_35252,N_33021,N_32825);
or U35253 (N_35253,N_32285,N_32731);
nand U35254 (N_35254,N_33677,N_32374);
xor U35255 (N_35255,N_33747,N_32603);
and U35256 (N_35256,N_32381,N_33297);
or U35257 (N_35257,N_32368,N_32457);
xor U35258 (N_35258,N_32407,N_33143);
and U35259 (N_35259,N_33876,N_33774);
or U35260 (N_35260,N_33276,N_33216);
xor U35261 (N_35261,N_33999,N_33147);
and U35262 (N_35262,N_32583,N_32890);
xnor U35263 (N_35263,N_33576,N_32989);
xor U35264 (N_35264,N_32132,N_32053);
and U35265 (N_35265,N_32109,N_32853);
nand U35266 (N_35266,N_32368,N_32117);
nor U35267 (N_35267,N_32980,N_33589);
nand U35268 (N_35268,N_33225,N_32632);
xor U35269 (N_35269,N_33939,N_32318);
and U35270 (N_35270,N_33558,N_32763);
nor U35271 (N_35271,N_33506,N_32035);
and U35272 (N_35272,N_33816,N_32453);
and U35273 (N_35273,N_32706,N_33272);
and U35274 (N_35274,N_33458,N_32829);
xnor U35275 (N_35275,N_32522,N_32793);
or U35276 (N_35276,N_33011,N_32055);
and U35277 (N_35277,N_32243,N_33566);
and U35278 (N_35278,N_32651,N_33854);
or U35279 (N_35279,N_32928,N_32975);
nor U35280 (N_35280,N_32469,N_33703);
or U35281 (N_35281,N_32293,N_33613);
nor U35282 (N_35282,N_33982,N_32386);
nor U35283 (N_35283,N_33349,N_33335);
or U35284 (N_35284,N_33022,N_33154);
nand U35285 (N_35285,N_33001,N_33410);
and U35286 (N_35286,N_33673,N_33105);
xor U35287 (N_35287,N_32850,N_33945);
xor U35288 (N_35288,N_32879,N_33454);
or U35289 (N_35289,N_33893,N_32202);
nor U35290 (N_35290,N_33722,N_32480);
xnor U35291 (N_35291,N_33437,N_33755);
or U35292 (N_35292,N_33566,N_33329);
nand U35293 (N_35293,N_33917,N_32526);
nor U35294 (N_35294,N_33670,N_32327);
nor U35295 (N_35295,N_33952,N_33417);
xnor U35296 (N_35296,N_33031,N_33720);
nand U35297 (N_35297,N_33892,N_32122);
or U35298 (N_35298,N_33889,N_33332);
xor U35299 (N_35299,N_32250,N_32457);
and U35300 (N_35300,N_33590,N_32035);
nand U35301 (N_35301,N_32166,N_32656);
and U35302 (N_35302,N_32351,N_32903);
nand U35303 (N_35303,N_32214,N_33627);
and U35304 (N_35304,N_33429,N_33582);
nand U35305 (N_35305,N_33508,N_33409);
nand U35306 (N_35306,N_32246,N_33214);
and U35307 (N_35307,N_32290,N_32714);
nor U35308 (N_35308,N_32734,N_32222);
xor U35309 (N_35309,N_32497,N_32169);
or U35310 (N_35310,N_33224,N_33764);
xor U35311 (N_35311,N_33593,N_32053);
xnor U35312 (N_35312,N_32644,N_33117);
and U35313 (N_35313,N_32666,N_33861);
nor U35314 (N_35314,N_33071,N_32421);
nor U35315 (N_35315,N_32967,N_33900);
and U35316 (N_35316,N_33425,N_32782);
or U35317 (N_35317,N_32706,N_32759);
and U35318 (N_35318,N_32309,N_32098);
xnor U35319 (N_35319,N_32751,N_33243);
and U35320 (N_35320,N_32437,N_33532);
xnor U35321 (N_35321,N_32372,N_32788);
and U35322 (N_35322,N_33173,N_32402);
xnor U35323 (N_35323,N_32845,N_32367);
or U35324 (N_35324,N_33903,N_33933);
nand U35325 (N_35325,N_32743,N_33809);
and U35326 (N_35326,N_32825,N_33353);
nor U35327 (N_35327,N_32907,N_32381);
or U35328 (N_35328,N_33410,N_33997);
nand U35329 (N_35329,N_33202,N_33114);
nand U35330 (N_35330,N_33507,N_33252);
and U35331 (N_35331,N_32546,N_32728);
xor U35332 (N_35332,N_32351,N_32630);
and U35333 (N_35333,N_32756,N_33025);
or U35334 (N_35334,N_32728,N_33171);
nand U35335 (N_35335,N_32156,N_33747);
and U35336 (N_35336,N_32812,N_33385);
or U35337 (N_35337,N_32449,N_32789);
nand U35338 (N_35338,N_32717,N_32216);
nand U35339 (N_35339,N_33703,N_33653);
xor U35340 (N_35340,N_32037,N_33723);
nand U35341 (N_35341,N_33599,N_33846);
nor U35342 (N_35342,N_32732,N_33358);
or U35343 (N_35343,N_33708,N_32825);
and U35344 (N_35344,N_33664,N_32445);
xor U35345 (N_35345,N_33720,N_33704);
nand U35346 (N_35346,N_32497,N_33446);
or U35347 (N_35347,N_32357,N_33846);
xor U35348 (N_35348,N_33462,N_33216);
or U35349 (N_35349,N_33442,N_32423);
and U35350 (N_35350,N_33510,N_32066);
or U35351 (N_35351,N_33431,N_32663);
and U35352 (N_35352,N_32303,N_32895);
nand U35353 (N_35353,N_33136,N_32629);
and U35354 (N_35354,N_33706,N_33911);
nand U35355 (N_35355,N_32595,N_32705);
nand U35356 (N_35356,N_33295,N_33948);
or U35357 (N_35357,N_32162,N_33127);
or U35358 (N_35358,N_32416,N_33484);
nand U35359 (N_35359,N_33816,N_32804);
nor U35360 (N_35360,N_32763,N_33046);
nand U35361 (N_35361,N_32947,N_32956);
nor U35362 (N_35362,N_32475,N_32309);
nor U35363 (N_35363,N_33249,N_33930);
nand U35364 (N_35364,N_32507,N_32253);
xnor U35365 (N_35365,N_32962,N_33830);
xor U35366 (N_35366,N_32377,N_33616);
and U35367 (N_35367,N_33913,N_32300);
or U35368 (N_35368,N_32195,N_33037);
nor U35369 (N_35369,N_32516,N_32935);
nand U35370 (N_35370,N_32141,N_32483);
or U35371 (N_35371,N_32311,N_33205);
and U35372 (N_35372,N_32238,N_33850);
xor U35373 (N_35373,N_33331,N_32499);
and U35374 (N_35374,N_32823,N_33196);
xor U35375 (N_35375,N_33167,N_33673);
xnor U35376 (N_35376,N_33153,N_32262);
xor U35377 (N_35377,N_33066,N_32108);
nand U35378 (N_35378,N_32936,N_32861);
and U35379 (N_35379,N_32571,N_32763);
or U35380 (N_35380,N_33168,N_32728);
or U35381 (N_35381,N_32238,N_33733);
nor U35382 (N_35382,N_33652,N_32236);
nand U35383 (N_35383,N_33660,N_33885);
or U35384 (N_35384,N_33925,N_32515);
or U35385 (N_35385,N_32438,N_32916);
or U35386 (N_35386,N_33305,N_32552);
nor U35387 (N_35387,N_32994,N_33403);
nor U35388 (N_35388,N_33426,N_32270);
nand U35389 (N_35389,N_33348,N_33808);
or U35390 (N_35390,N_33704,N_33475);
xnor U35391 (N_35391,N_33848,N_33635);
xnor U35392 (N_35392,N_33052,N_32544);
nand U35393 (N_35393,N_33903,N_32343);
or U35394 (N_35394,N_33194,N_33570);
nor U35395 (N_35395,N_33022,N_33554);
and U35396 (N_35396,N_32288,N_32950);
xor U35397 (N_35397,N_33937,N_33796);
xor U35398 (N_35398,N_32451,N_33193);
or U35399 (N_35399,N_32094,N_33076);
and U35400 (N_35400,N_32931,N_32272);
nor U35401 (N_35401,N_33038,N_32502);
nand U35402 (N_35402,N_33387,N_33936);
or U35403 (N_35403,N_32720,N_33953);
xor U35404 (N_35404,N_32260,N_32783);
nand U35405 (N_35405,N_32028,N_33839);
or U35406 (N_35406,N_33630,N_33731);
nor U35407 (N_35407,N_32124,N_33225);
or U35408 (N_35408,N_32466,N_33605);
nand U35409 (N_35409,N_32467,N_33317);
and U35410 (N_35410,N_33024,N_33774);
or U35411 (N_35411,N_32329,N_33826);
and U35412 (N_35412,N_32180,N_32132);
nor U35413 (N_35413,N_33647,N_33887);
nor U35414 (N_35414,N_33301,N_33401);
and U35415 (N_35415,N_33540,N_32954);
xor U35416 (N_35416,N_33133,N_32358);
nand U35417 (N_35417,N_32452,N_33148);
and U35418 (N_35418,N_32816,N_33940);
nor U35419 (N_35419,N_32095,N_33068);
or U35420 (N_35420,N_32351,N_33794);
xnor U35421 (N_35421,N_32981,N_32396);
and U35422 (N_35422,N_33704,N_32196);
and U35423 (N_35423,N_33838,N_33441);
nor U35424 (N_35424,N_33197,N_32730);
xnor U35425 (N_35425,N_32726,N_32887);
nand U35426 (N_35426,N_33890,N_33579);
xor U35427 (N_35427,N_32363,N_32576);
nand U35428 (N_35428,N_32722,N_33558);
or U35429 (N_35429,N_32997,N_33334);
nor U35430 (N_35430,N_33159,N_32484);
nand U35431 (N_35431,N_32785,N_33092);
nand U35432 (N_35432,N_33045,N_32719);
nor U35433 (N_35433,N_33290,N_32048);
xnor U35434 (N_35434,N_33589,N_33408);
or U35435 (N_35435,N_32976,N_33757);
and U35436 (N_35436,N_33329,N_32866);
nor U35437 (N_35437,N_33657,N_32307);
xnor U35438 (N_35438,N_32380,N_32217);
and U35439 (N_35439,N_33279,N_32551);
and U35440 (N_35440,N_33211,N_33082);
nor U35441 (N_35441,N_33661,N_32194);
and U35442 (N_35442,N_32826,N_32572);
or U35443 (N_35443,N_33607,N_32741);
and U35444 (N_35444,N_32793,N_33624);
nand U35445 (N_35445,N_33944,N_32911);
or U35446 (N_35446,N_33849,N_33161);
xnor U35447 (N_35447,N_32017,N_32828);
or U35448 (N_35448,N_32543,N_32142);
nand U35449 (N_35449,N_33161,N_32655);
nand U35450 (N_35450,N_32251,N_32909);
and U35451 (N_35451,N_32105,N_32945);
nor U35452 (N_35452,N_33803,N_33563);
nand U35453 (N_35453,N_33625,N_32821);
nor U35454 (N_35454,N_32131,N_33563);
xor U35455 (N_35455,N_32613,N_32216);
or U35456 (N_35456,N_32254,N_33763);
nor U35457 (N_35457,N_33530,N_32804);
or U35458 (N_35458,N_33437,N_33853);
nand U35459 (N_35459,N_32212,N_33370);
or U35460 (N_35460,N_33878,N_33438);
xnor U35461 (N_35461,N_33168,N_32323);
and U35462 (N_35462,N_32139,N_32434);
and U35463 (N_35463,N_32351,N_33118);
nor U35464 (N_35464,N_33061,N_33191);
and U35465 (N_35465,N_33017,N_32320);
nand U35466 (N_35466,N_32057,N_32823);
or U35467 (N_35467,N_32935,N_32214);
and U35468 (N_35468,N_33868,N_32568);
nor U35469 (N_35469,N_32173,N_33105);
xor U35470 (N_35470,N_32693,N_33436);
xnor U35471 (N_35471,N_32149,N_32007);
nand U35472 (N_35472,N_33817,N_32093);
xor U35473 (N_35473,N_33514,N_33941);
nand U35474 (N_35474,N_33648,N_33413);
nand U35475 (N_35475,N_32421,N_32662);
nor U35476 (N_35476,N_33898,N_33498);
nand U35477 (N_35477,N_32696,N_33209);
nor U35478 (N_35478,N_33991,N_33077);
nand U35479 (N_35479,N_33498,N_33082);
or U35480 (N_35480,N_32900,N_33212);
xor U35481 (N_35481,N_33531,N_33282);
nor U35482 (N_35482,N_33493,N_33411);
nor U35483 (N_35483,N_32137,N_32552);
or U35484 (N_35484,N_32675,N_32008);
nand U35485 (N_35485,N_33509,N_32518);
xor U35486 (N_35486,N_33833,N_32133);
and U35487 (N_35487,N_32532,N_33074);
and U35488 (N_35488,N_33469,N_33097);
and U35489 (N_35489,N_32458,N_33268);
xor U35490 (N_35490,N_33333,N_33052);
nand U35491 (N_35491,N_32944,N_32229);
nor U35492 (N_35492,N_33085,N_32927);
xnor U35493 (N_35493,N_33110,N_33823);
nor U35494 (N_35494,N_32065,N_32240);
nand U35495 (N_35495,N_32085,N_32058);
and U35496 (N_35496,N_33683,N_32901);
and U35497 (N_35497,N_32451,N_33901);
nand U35498 (N_35498,N_32288,N_32409);
or U35499 (N_35499,N_32391,N_33060);
xnor U35500 (N_35500,N_32284,N_33102);
xnor U35501 (N_35501,N_33479,N_32030);
or U35502 (N_35502,N_33016,N_32222);
xnor U35503 (N_35503,N_33142,N_33466);
xor U35504 (N_35504,N_33864,N_32322);
nand U35505 (N_35505,N_33353,N_33515);
nor U35506 (N_35506,N_32641,N_33269);
xor U35507 (N_35507,N_32624,N_32395);
or U35508 (N_35508,N_32247,N_33023);
or U35509 (N_35509,N_32190,N_33770);
nor U35510 (N_35510,N_32398,N_33916);
nand U35511 (N_35511,N_33854,N_33814);
xor U35512 (N_35512,N_33094,N_32178);
and U35513 (N_35513,N_33233,N_32959);
and U35514 (N_35514,N_32522,N_32325);
xor U35515 (N_35515,N_32021,N_32393);
or U35516 (N_35516,N_33279,N_33780);
xnor U35517 (N_35517,N_33877,N_33750);
xnor U35518 (N_35518,N_33234,N_32488);
or U35519 (N_35519,N_32282,N_33953);
or U35520 (N_35520,N_33790,N_32346);
xnor U35521 (N_35521,N_33456,N_32471);
and U35522 (N_35522,N_32232,N_33420);
and U35523 (N_35523,N_33960,N_33812);
and U35524 (N_35524,N_32104,N_33393);
nor U35525 (N_35525,N_32655,N_33315);
nor U35526 (N_35526,N_33417,N_32964);
nor U35527 (N_35527,N_33120,N_33691);
nand U35528 (N_35528,N_32460,N_32472);
xor U35529 (N_35529,N_33042,N_32624);
xnor U35530 (N_35530,N_32159,N_32736);
and U35531 (N_35531,N_33604,N_32278);
nor U35532 (N_35532,N_32650,N_32501);
and U35533 (N_35533,N_33837,N_32437);
or U35534 (N_35534,N_32465,N_32701);
or U35535 (N_35535,N_33700,N_33322);
xor U35536 (N_35536,N_32711,N_33730);
nor U35537 (N_35537,N_32218,N_33262);
nand U35538 (N_35538,N_33392,N_32694);
nand U35539 (N_35539,N_33214,N_33269);
or U35540 (N_35540,N_33848,N_32574);
xor U35541 (N_35541,N_32356,N_32028);
xnor U35542 (N_35542,N_32460,N_33056);
and U35543 (N_35543,N_33153,N_33850);
and U35544 (N_35544,N_33792,N_32478);
and U35545 (N_35545,N_32592,N_33010);
and U35546 (N_35546,N_32176,N_33769);
nor U35547 (N_35547,N_32143,N_32730);
and U35548 (N_35548,N_32947,N_32070);
xor U35549 (N_35549,N_33375,N_32158);
or U35550 (N_35550,N_33852,N_32472);
or U35551 (N_35551,N_33680,N_33078);
nand U35552 (N_35552,N_32480,N_33129);
nor U35553 (N_35553,N_32538,N_32258);
nand U35554 (N_35554,N_33518,N_32051);
nand U35555 (N_35555,N_32543,N_33327);
and U35556 (N_35556,N_33229,N_32018);
or U35557 (N_35557,N_33762,N_32502);
nor U35558 (N_35558,N_32691,N_32737);
or U35559 (N_35559,N_33519,N_32576);
nand U35560 (N_35560,N_33394,N_33112);
nand U35561 (N_35561,N_32469,N_32783);
nor U35562 (N_35562,N_32618,N_32078);
xor U35563 (N_35563,N_33477,N_33731);
xnor U35564 (N_35564,N_32307,N_32354);
or U35565 (N_35565,N_33429,N_33672);
nor U35566 (N_35566,N_32794,N_32010);
or U35567 (N_35567,N_32433,N_33118);
nand U35568 (N_35568,N_32699,N_32058);
nor U35569 (N_35569,N_33326,N_33804);
xnor U35570 (N_35570,N_33186,N_33487);
xor U35571 (N_35571,N_33341,N_33162);
nor U35572 (N_35572,N_32914,N_33541);
xor U35573 (N_35573,N_32873,N_32855);
nand U35574 (N_35574,N_33489,N_33572);
and U35575 (N_35575,N_32640,N_33961);
or U35576 (N_35576,N_32516,N_32030);
or U35577 (N_35577,N_32135,N_33162);
or U35578 (N_35578,N_32308,N_33590);
xor U35579 (N_35579,N_32625,N_32429);
or U35580 (N_35580,N_32806,N_33230);
nand U35581 (N_35581,N_32064,N_33514);
nor U35582 (N_35582,N_33259,N_32799);
nor U35583 (N_35583,N_33621,N_33708);
and U35584 (N_35584,N_32315,N_32517);
and U35585 (N_35585,N_32044,N_33241);
and U35586 (N_35586,N_32680,N_32359);
and U35587 (N_35587,N_32750,N_33876);
nor U35588 (N_35588,N_33745,N_33823);
xor U35589 (N_35589,N_33618,N_33638);
nor U35590 (N_35590,N_32006,N_33872);
nand U35591 (N_35591,N_33367,N_32176);
xor U35592 (N_35592,N_33027,N_32998);
and U35593 (N_35593,N_33598,N_33044);
nand U35594 (N_35594,N_32238,N_33372);
nor U35595 (N_35595,N_33214,N_33809);
and U35596 (N_35596,N_33006,N_32822);
nand U35597 (N_35597,N_33802,N_32384);
nor U35598 (N_35598,N_32806,N_32125);
nor U35599 (N_35599,N_33294,N_32640);
nand U35600 (N_35600,N_33448,N_33928);
and U35601 (N_35601,N_33662,N_33197);
and U35602 (N_35602,N_33126,N_33723);
nor U35603 (N_35603,N_33841,N_33033);
or U35604 (N_35604,N_33136,N_33125);
and U35605 (N_35605,N_32977,N_32853);
nor U35606 (N_35606,N_32855,N_32281);
nor U35607 (N_35607,N_33612,N_32335);
xor U35608 (N_35608,N_32152,N_33209);
nor U35609 (N_35609,N_32386,N_32150);
nand U35610 (N_35610,N_32630,N_32622);
nand U35611 (N_35611,N_33078,N_33819);
or U35612 (N_35612,N_32258,N_32920);
nor U35613 (N_35613,N_33857,N_33715);
nand U35614 (N_35614,N_33537,N_33526);
nor U35615 (N_35615,N_33698,N_33161);
or U35616 (N_35616,N_32230,N_32321);
or U35617 (N_35617,N_32193,N_32717);
nor U35618 (N_35618,N_33112,N_33212);
nand U35619 (N_35619,N_32742,N_32639);
xor U35620 (N_35620,N_33123,N_32847);
nor U35621 (N_35621,N_32707,N_33394);
or U35622 (N_35622,N_32156,N_32982);
and U35623 (N_35623,N_33690,N_33851);
or U35624 (N_35624,N_32859,N_32254);
xor U35625 (N_35625,N_33525,N_33834);
nand U35626 (N_35626,N_32853,N_33782);
xnor U35627 (N_35627,N_33600,N_33409);
xor U35628 (N_35628,N_32727,N_32443);
nand U35629 (N_35629,N_32963,N_33843);
and U35630 (N_35630,N_32099,N_32675);
xnor U35631 (N_35631,N_32961,N_33555);
xor U35632 (N_35632,N_33804,N_33541);
nor U35633 (N_35633,N_32167,N_33966);
or U35634 (N_35634,N_33732,N_33840);
nor U35635 (N_35635,N_33387,N_32891);
or U35636 (N_35636,N_32858,N_32557);
and U35637 (N_35637,N_32490,N_33194);
or U35638 (N_35638,N_32004,N_32449);
and U35639 (N_35639,N_32593,N_32378);
nand U35640 (N_35640,N_33908,N_32923);
and U35641 (N_35641,N_33126,N_32706);
nor U35642 (N_35642,N_32312,N_33344);
and U35643 (N_35643,N_32597,N_32804);
or U35644 (N_35644,N_33879,N_32209);
nand U35645 (N_35645,N_32289,N_32977);
nand U35646 (N_35646,N_33440,N_33149);
nand U35647 (N_35647,N_32051,N_33653);
or U35648 (N_35648,N_33214,N_33226);
nor U35649 (N_35649,N_32280,N_32641);
or U35650 (N_35650,N_33691,N_33860);
xnor U35651 (N_35651,N_33375,N_32337);
nor U35652 (N_35652,N_32193,N_33042);
or U35653 (N_35653,N_32578,N_32503);
and U35654 (N_35654,N_33361,N_33267);
nand U35655 (N_35655,N_33062,N_33615);
nor U35656 (N_35656,N_32034,N_33844);
xor U35657 (N_35657,N_32737,N_32035);
xnor U35658 (N_35658,N_33611,N_32920);
nand U35659 (N_35659,N_32720,N_32920);
and U35660 (N_35660,N_33225,N_32995);
nand U35661 (N_35661,N_33513,N_32589);
and U35662 (N_35662,N_33637,N_32179);
and U35663 (N_35663,N_33401,N_33811);
nor U35664 (N_35664,N_33574,N_32958);
or U35665 (N_35665,N_32988,N_32541);
xor U35666 (N_35666,N_33632,N_32865);
nor U35667 (N_35667,N_32324,N_33248);
and U35668 (N_35668,N_33287,N_32307);
nand U35669 (N_35669,N_33345,N_33101);
nand U35670 (N_35670,N_33431,N_32023);
or U35671 (N_35671,N_33875,N_32204);
or U35672 (N_35672,N_33117,N_33199);
nor U35673 (N_35673,N_33437,N_32301);
or U35674 (N_35674,N_33936,N_33071);
xnor U35675 (N_35675,N_33743,N_32929);
and U35676 (N_35676,N_33590,N_32275);
nand U35677 (N_35677,N_33849,N_32142);
nor U35678 (N_35678,N_32130,N_32748);
nor U35679 (N_35679,N_32690,N_32762);
xor U35680 (N_35680,N_33181,N_33627);
nand U35681 (N_35681,N_33191,N_32223);
xnor U35682 (N_35682,N_33004,N_32564);
and U35683 (N_35683,N_32153,N_33107);
or U35684 (N_35684,N_32023,N_32578);
xnor U35685 (N_35685,N_32069,N_33926);
xor U35686 (N_35686,N_33595,N_33316);
xnor U35687 (N_35687,N_32908,N_32487);
xnor U35688 (N_35688,N_32877,N_33204);
and U35689 (N_35689,N_33966,N_32317);
or U35690 (N_35690,N_33499,N_32298);
and U35691 (N_35691,N_32765,N_32061);
nor U35692 (N_35692,N_33379,N_33292);
or U35693 (N_35693,N_32502,N_33287);
nand U35694 (N_35694,N_32398,N_33469);
xor U35695 (N_35695,N_32445,N_32792);
and U35696 (N_35696,N_33672,N_32943);
xnor U35697 (N_35697,N_32219,N_33920);
nand U35698 (N_35698,N_32181,N_32581);
and U35699 (N_35699,N_33841,N_33798);
nand U35700 (N_35700,N_32901,N_32215);
xor U35701 (N_35701,N_32554,N_32052);
and U35702 (N_35702,N_33877,N_32547);
xor U35703 (N_35703,N_33240,N_32745);
nand U35704 (N_35704,N_33323,N_33769);
nand U35705 (N_35705,N_32147,N_33502);
nor U35706 (N_35706,N_33291,N_33812);
nor U35707 (N_35707,N_33786,N_32849);
nor U35708 (N_35708,N_33272,N_33455);
nand U35709 (N_35709,N_32639,N_32158);
nand U35710 (N_35710,N_32570,N_33127);
nor U35711 (N_35711,N_32068,N_33308);
and U35712 (N_35712,N_33893,N_33634);
xor U35713 (N_35713,N_32290,N_32028);
nor U35714 (N_35714,N_33901,N_33586);
xor U35715 (N_35715,N_33374,N_32035);
xnor U35716 (N_35716,N_33277,N_32565);
nand U35717 (N_35717,N_33372,N_32357);
and U35718 (N_35718,N_32753,N_33051);
nor U35719 (N_35719,N_33501,N_32306);
nand U35720 (N_35720,N_33406,N_32338);
or U35721 (N_35721,N_32907,N_33197);
or U35722 (N_35722,N_32209,N_33668);
nand U35723 (N_35723,N_32361,N_33202);
and U35724 (N_35724,N_32941,N_32436);
xnor U35725 (N_35725,N_32038,N_32275);
and U35726 (N_35726,N_32525,N_33096);
xor U35727 (N_35727,N_32185,N_33685);
or U35728 (N_35728,N_32481,N_32119);
xnor U35729 (N_35729,N_32335,N_32272);
nor U35730 (N_35730,N_32069,N_32301);
nor U35731 (N_35731,N_33416,N_32677);
xor U35732 (N_35732,N_33284,N_32699);
nor U35733 (N_35733,N_32576,N_33722);
nor U35734 (N_35734,N_33953,N_33820);
or U35735 (N_35735,N_33533,N_32519);
nor U35736 (N_35736,N_32735,N_32588);
xnor U35737 (N_35737,N_33486,N_33039);
or U35738 (N_35738,N_32948,N_33893);
or U35739 (N_35739,N_33325,N_33125);
nand U35740 (N_35740,N_32209,N_32214);
xor U35741 (N_35741,N_33812,N_33757);
nand U35742 (N_35742,N_32194,N_32008);
nand U35743 (N_35743,N_33515,N_33172);
nor U35744 (N_35744,N_32049,N_33241);
nand U35745 (N_35745,N_33875,N_33536);
or U35746 (N_35746,N_33283,N_32598);
nand U35747 (N_35747,N_32032,N_32133);
nor U35748 (N_35748,N_32425,N_32862);
nor U35749 (N_35749,N_33974,N_33223);
and U35750 (N_35750,N_32635,N_33118);
or U35751 (N_35751,N_32875,N_33733);
or U35752 (N_35752,N_33627,N_32846);
or U35753 (N_35753,N_32237,N_32783);
and U35754 (N_35754,N_33418,N_32841);
xor U35755 (N_35755,N_33071,N_33897);
nor U35756 (N_35756,N_32315,N_33337);
xnor U35757 (N_35757,N_32515,N_33661);
or U35758 (N_35758,N_33747,N_32439);
or U35759 (N_35759,N_32899,N_32589);
nor U35760 (N_35760,N_33820,N_33322);
xnor U35761 (N_35761,N_32166,N_33548);
nor U35762 (N_35762,N_33487,N_32537);
and U35763 (N_35763,N_33196,N_32980);
or U35764 (N_35764,N_33580,N_32489);
and U35765 (N_35765,N_32121,N_32084);
xor U35766 (N_35766,N_33768,N_32466);
xor U35767 (N_35767,N_32118,N_32517);
and U35768 (N_35768,N_32606,N_33386);
nand U35769 (N_35769,N_32214,N_33097);
nand U35770 (N_35770,N_32503,N_32790);
nor U35771 (N_35771,N_33047,N_32696);
nand U35772 (N_35772,N_33516,N_33574);
nand U35773 (N_35773,N_33230,N_32471);
xnor U35774 (N_35774,N_32574,N_32250);
and U35775 (N_35775,N_32994,N_33660);
nor U35776 (N_35776,N_32430,N_32137);
and U35777 (N_35777,N_32225,N_32596);
nand U35778 (N_35778,N_33187,N_32363);
xor U35779 (N_35779,N_33609,N_33843);
or U35780 (N_35780,N_32656,N_33025);
xor U35781 (N_35781,N_32213,N_33991);
xnor U35782 (N_35782,N_33949,N_33772);
and U35783 (N_35783,N_32461,N_32000);
nor U35784 (N_35784,N_32463,N_33930);
xor U35785 (N_35785,N_33763,N_33884);
xor U35786 (N_35786,N_32543,N_33640);
nor U35787 (N_35787,N_33650,N_32341);
nand U35788 (N_35788,N_32981,N_32012);
or U35789 (N_35789,N_33766,N_33393);
and U35790 (N_35790,N_33785,N_33131);
xnor U35791 (N_35791,N_32915,N_32940);
nand U35792 (N_35792,N_32730,N_32843);
or U35793 (N_35793,N_33913,N_32172);
nand U35794 (N_35794,N_33425,N_33941);
xnor U35795 (N_35795,N_32684,N_33572);
or U35796 (N_35796,N_32909,N_32437);
and U35797 (N_35797,N_32373,N_32109);
or U35798 (N_35798,N_33787,N_32608);
nand U35799 (N_35799,N_32358,N_32012);
or U35800 (N_35800,N_33664,N_32905);
or U35801 (N_35801,N_33414,N_32237);
and U35802 (N_35802,N_32206,N_33382);
or U35803 (N_35803,N_32922,N_32906);
nand U35804 (N_35804,N_32026,N_33555);
or U35805 (N_35805,N_32301,N_32035);
nand U35806 (N_35806,N_33969,N_33372);
and U35807 (N_35807,N_32342,N_33590);
nor U35808 (N_35808,N_33298,N_33800);
or U35809 (N_35809,N_32087,N_33228);
and U35810 (N_35810,N_32856,N_32731);
nand U35811 (N_35811,N_32550,N_32784);
or U35812 (N_35812,N_33531,N_32756);
nand U35813 (N_35813,N_33189,N_32129);
nor U35814 (N_35814,N_33684,N_33577);
nor U35815 (N_35815,N_33110,N_33670);
nor U35816 (N_35816,N_33682,N_33100);
nand U35817 (N_35817,N_33177,N_32794);
and U35818 (N_35818,N_32686,N_33279);
or U35819 (N_35819,N_33415,N_33284);
nor U35820 (N_35820,N_32328,N_32907);
nand U35821 (N_35821,N_33760,N_33821);
and U35822 (N_35822,N_33545,N_33359);
and U35823 (N_35823,N_32750,N_32312);
and U35824 (N_35824,N_33964,N_33823);
or U35825 (N_35825,N_32461,N_33511);
nand U35826 (N_35826,N_33959,N_33938);
or U35827 (N_35827,N_32116,N_33643);
nor U35828 (N_35828,N_32695,N_32138);
nor U35829 (N_35829,N_32746,N_32625);
nor U35830 (N_35830,N_32372,N_33712);
nand U35831 (N_35831,N_33116,N_33018);
or U35832 (N_35832,N_33851,N_32738);
nor U35833 (N_35833,N_33891,N_33853);
or U35834 (N_35834,N_32795,N_32895);
nand U35835 (N_35835,N_32484,N_32921);
and U35836 (N_35836,N_32802,N_33362);
and U35837 (N_35837,N_33036,N_33072);
nand U35838 (N_35838,N_33858,N_33474);
or U35839 (N_35839,N_33667,N_32098);
xnor U35840 (N_35840,N_32859,N_32771);
nand U35841 (N_35841,N_33938,N_33275);
nor U35842 (N_35842,N_32530,N_33579);
nand U35843 (N_35843,N_32667,N_33564);
and U35844 (N_35844,N_33982,N_33029);
xor U35845 (N_35845,N_32542,N_32938);
nor U35846 (N_35846,N_32749,N_32358);
nand U35847 (N_35847,N_33249,N_32672);
and U35848 (N_35848,N_32242,N_33192);
nor U35849 (N_35849,N_33259,N_32152);
xnor U35850 (N_35850,N_32048,N_33967);
nor U35851 (N_35851,N_33532,N_32436);
nand U35852 (N_35852,N_32860,N_33126);
nand U35853 (N_35853,N_33497,N_33336);
nand U35854 (N_35854,N_33433,N_32729);
nor U35855 (N_35855,N_32245,N_32150);
nand U35856 (N_35856,N_32827,N_33545);
nor U35857 (N_35857,N_33455,N_33341);
or U35858 (N_35858,N_33563,N_32204);
xnor U35859 (N_35859,N_32145,N_32997);
and U35860 (N_35860,N_33021,N_33407);
xnor U35861 (N_35861,N_32212,N_32181);
nand U35862 (N_35862,N_33432,N_33888);
nand U35863 (N_35863,N_32339,N_32836);
xnor U35864 (N_35864,N_32327,N_33869);
nand U35865 (N_35865,N_33255,N_33221);
nand U35866 (N_35866,N_32301,N_33649);
nor U35867 (N_35867,N_32893,N_32905);
or U35868 (N_35868,N_33779,N_32836);
nand U35869 (N_35869,N_32467,N_33531);
nand U35870 (N_35870,N_33998,N_32894);
or U35871 (N_35871,N_32176,N_33309);
nand U35872 (N_35872,N_33253,N_32867);
and U35873 (N_35873,N_32321,N_33422);
nor U35874 (N_35874,N_32782,N_32795);
or U35875 (N_35875,N_32936,N_33236);
nand U35876 (N_35876,N_33663,N_33376);
and U35877 (N_35877,N_32127,N_32930);
nor U35878 (N_35878,N_33119,N_32944);
nand U35879 (N_35879,N_32050,N_33570);
nor U35880 (N_35880,N_33250,N_33243);
nand U35881 (N_35881,N_32653,N_33581);
nor U35882 (N_35882,N_33141,N_33490);
or U35883 (N_35883,N_32867,N_33887);
nand U35884 (N_35884,N_32404,N_32890);
and U35885 (N_35885,N_32007,N_32968);
nor U35886 (N_35886,N_32557,N_33538);
xnor U35887 (N_35887,N_33520,N_32213);
nand U35888 (N_35888,N_33131,N_32685);
and U35889 (N_35889,N_33581,N_32410);
or U35890 (N_35890,N_32937,N_33641);
xor U35891 (N_35891,N_32979,N_33727);
nor U35892 (N_35892,N_32759,N_32185);
xnor U35893 (N_35893,N_33498,N_32690);
nand U35894 (N_35894,N_33056,N_32613);
xnor U35895 (N_35895,N_32305,N_33198);
or U35896 (N_35896,N_32968,N_33275);
nor U35897 (N_35897,N_32322,N_32239);
xnor U35898 (N_35898,N_33586,N_33391);
nand U35899 (N_35899,N_32334,N_33936);
nand U35900 (N_35900,N_33728,N_32886);
or U35901 (N_35901,N_33629,N_32220);
nor U35902 (N_35902,N_33312,N_32464);
nand U35903 (N_35903,N_32577,N_32049);
or U35904 (N_35904,N_33066,N_32856);
nand U35905 (N_35905,N_32238,N_32889);
and U35906 (N_35906,N_32752,N_33639);
or U35907 (N_35907,N_32795,N_32055);
or U35908 (N_35908,N_32089,N_33301);
and U35909 (N_35909,N_33645,N_32671);
nand U35910 (N_35910,N_33298,N_33649);
or U35911 (N_35911,N_33159,N_32962);
nor U35912 (N_35912,N_33899,N_32947);
or U35913 (N_35913,N_32205,N_33720);
xor U35914 (N_35914,N_32799,N_32047);
or U35915 (N_35915,N_32968,N_33843);
nand U35916 (N_35916,N_32913,N_32294);
and U35917 (N_35917,N_33194,N_33380);
nand U35918 (N_35918,N_33417,N_32325);
xor U35919 (N_35919,N_32845,N_32590);
nand U35920 (N_35920,N_33559,N_32395);
nor U35921 (N_35921,N_33311,N_33504);
nor U35922 (N_35922,N_32304,N_32580);
nand U35923 (N_35923,N_32219,N_32892);
nand U35924 (N_35924,N_33566,N_33004);
or U35925 (N_35925,N_32709,N_33063);
xor U35926 (N_35926,N_32661,N_33085);
nor U35927 (N_35927,N_33834,N_33562);
and U35928 (N_35928,N_32259,N_33014);
nor U35929 (N_35929,N_33947,N_32516);
nand U35930 (N_35930,N_33948,N_33868);
nand U35931 (N_35931,N_33267,N_32008);
xnor U35932 (N_35932,N_32957,N_33563);
xor U35933 (N_35933,N_33664,N_33131);
nor U35934 (N_35934,N_33209,N_32494);
xnor U35935 (N_35935,N_33234,N_33578);
xor U35936 (N_35936,N_32887,N_32472);
and U35937 (N_35937,N_32785,N_33296);
nor U35938 (N_35938,N_33191,N_32999);
xnor U35939 (N_35939,N_32955,N_33337);
nor U35940 (N_35940,N_32002,N_33013);
xor U35941 (N_35941,N_33745,N_33117);
or U35942 (N_35942,N_33666,N_32958);
nand U35943 (N_35943,N_33655,N_33699);
and U35944 (N_35944,N_32662,N_32631);
nand U35945 (N_35945,N_32244,N_33204);
and U35946 (N_35946,N_32253,N_33333);
nand U35947 (N_35947,N_33954,N_33761);
nand U35948 (N_35948,N_33713,N_33804);
nand U35949 (N_35949,N_33102,N_33837);
nand U35950 (N_35950,N_33625,N_33087);
nor U35951 (N_35951,N_33401,N_33416);
or U35952 (N_35952,N_33527,N_33595);
nand U35953 (N_35953,N_32153,N_32037);
nand U35954 (N_35954,N_32354,N_33407);
nor U35955 (N_35955,N_32432,N_32893);
nand U35956 (N_35956,N_33613,N_32893);
nor U35957 (N_35957,N_33595,N_33716);
and U35958 (N_35958,N_33193,N_33879);
or U35959 (N_35959,N_32445,N_33063);
and U35960 (N_35960,N_33673,N_32065);
and U35961 (N_35961,N_32966,N_33319);
or U35962 (N_35962,N_32097,N_32699);
nand U35963 (N_35963,N_33303,N_33720);
xnor U35964 (N_35964,N_32754,N_33516);
nand U35965 (N_35965,N_32339,N_33594);
xor U35966 (N_35966,N_33100,N_33899);
xnor U35967 (N_35967,N_32323,N_32577);
xnor U35968 (N_35968,N_33317,N_32212);
or U35969 (N_35969,N_33657,N_32130);
nor U35970 (N_35970,N_32382,N_32520);
xnor U35971 (N_35971,N_33734,N_33678);
or U35972 (N_35972,N_33041,N_33950);
xnor U35973 (N_35973,N_33579,N_32086);
nor U35974 (N_35974,N_33084,N_33384);
nand U35975 (N_35975,N_33341,N_33070);
nor U35976 (N_35976,N_33419,N_32908);
nor U35977 (N_35977,N_33195,N_32158);
and U35978 (N_35978,N_33375,N_32125);
nand U35979 (N_35979,N_32292,N_32548);
nand U35980 (N_35980,N_32238,N_33727);
nor U35981 (N_35981,N_33555,N_33755);
nor U35982 (N_35982,N_32893,N_33085);
xnor U35983 (N_35983,N_32623,N_32862);
nor U35984 (N_35984,N_32731,N_33913);
nand U35985 (N_35985,N_33870,N_33600);
nand U35986 (N_35986,N_32857,N_32769);
nand U35987 (N_35987,N_33732,N_33700);
and U35988 (N_35988,N_33794,N_33852);
or U35989 (N_35989,N_33557,N_32697);
nand U35990 (N_35990,N_33992,N_33975);
or U35991 (N_35991,N_33030,N_32481);
or U35992 (N_35992,N_32837,N_33548);
nand U35993 (N_35993,N_32034,N_33258);
or U35994 (N_35994,N_33814,N_32285);
and U35995 (N_35995,N_33579,N_33175);
and U35996 (N_35996,N_33666,N_33591);
nand U35997 (N_35997,N_32641,N_32843);
and U35998 (N_35998,N_33062,N_32288);
xnor U35999 (N_35999,N_33313,N_32933);
nand U36000 (N_36000,N_35898,N_35467);
and U36001 (N_36001,N_35570,N_34251);
xor U36002 (N_36002,N_34472,N_34287);
xnor U36003 (N_36003,N_35262,N_35210);
or U36004 (N_36004,N_35515,N_35571);
or U36005 (N_36005,N_35585,N_34324);
or U36006 (N_36006,N_34598,N_34098);
or U36007 (N_36007,N_35400,N_35142);
or U36008 (N_36008,N_35138,N_35963);
or U36009 (N_36009,N_34206,N_34089);
nand U36010 (N_36010,N_34395,N_35477);
nor U36011 (N_36011,N_34981,N_34175);
and U36012 (N_36012,N_34360,N_35633);
or U36013 (N_36013,N_35954,N_34152);
and U36014 (N_36014,N_34694,N_35098);
nor U36015 (N_36015,N_34257,N_34496);
nand U36016 (N_36016,N_34773,N_34457);
and U36017 (N_36017,N_34831,N_34374);
nand U36018 (N_36018,N_34302,N_34428);
nor U36019 (N_36019,N_34872,N_34873);
xnor U36020 (N_36020,N_35893,N_34580);
xnor U36021 (N_36021,N_35705,N_34477);
or U36022 (N_36022,N_35785,N_34433);
and U36023 (N_36023,N_35835,N_34401);
nand U36024 (N_36024,N_34862,N_34029);
and U36025 (N_36025,N_34241,N_35036);
nor U36026 (N_36026,N_34057,N_34337);
nor U36027 (N_36027,N_35843,N_35830);
nand U36028 (N_36028,N_34413,N_34420);
or U36029 (N_36029,N_34454,N_35704);
or U36030 (N_36030,N_34312,N_35975);
xnor U36031 (N_36031,N_35317,N_34161);
nor U36032 (N_36032,N_34054,N_34533);
xnor U36033 (N_36033,N_34438,N_34279);
and U36034 (N_36034,N_35209,N_34855);
xor U36035 (N_36035,N_34995,N_34227);
nand U36036 (N_36036,N_35584,N_34911);
nor U36037 (N_36037,N_34667,N_34844);
nand U36038 (N_36038,N_35120,N_35780);
and U36039 (N_36039,N_35324,N_35225);
nor U36040 (N_36040,N_35053,N_34609);
or U36041 (N_36041,N_35792,N_34572);
or U36042 (N_36042,N_34463,N_34311);
nand U36043 (N_36043,N_34197,N_34107);
nand U36044 (N_36044,N_35701,N_34789);
xnor U36045 (N_36045,N_35831,N_35154);
nand U36046 (N_36046,N_34895,N_34309);
nand U36047 (N_36047,N_34822,N_34385);
xor U36048 (N_36048,N_34129,N_34881);
xor U36049 (N_36049,N_34756,N_34845);
nand U36050 (N_36050,N_35685,N_35594);
and U36051 (N_36051,N_34444,N_35998);
nand U36052 (N_36052,N_34173,N_35493);
xor U36053 (N_36053,N_34458,N_35109);
xnor U36054 (N_36054,N_34787,N_35474);
xnor U36055 (N_36055,N_34733,N_34735);
nor U36056 (N_36056,N_35124,N_34514);
and U36057 (N_36057,N_35667,N_34292);
or U36058 (N_36058,N_35414,N_35356);
and U36059 (N_36059,N_34544,N_35728);
xnor U36060 (N_36060,N_35659,N_35466);
nor U36061 (N_36061,N_34488,N_35838);
nand U36062 (N_36062,N_34059,N_35741);
xnor U36063 (N_36063,N_34531,N_34585);
xnor U36064 (N_36064,N_34936,N_34908);
nor U36065 (N_36065,N_35945,N_35265);
nand U36066 (N_36066,N_35921,N_35086);
and U36067 (N_36067,N_35037,N_35385);
xor U36068 (N_36068,N_35894,N_35828);
nand U36069 (N_36069,N_35146,N_35745);
and U36070 (N_36070,N_34866,N_35191);
nand U36071 (N_36071,N_35253,N_34269);
and U36072 (N_36072,N_34763,N_35343);
xor U36073 (N_36073,N_35798,N_34080);
nand U36074 (N_36074,N_35079,N_35607);
and U36075 (N_36075,N_34655,N_34856);
nor U36076 (N_36076,N_35510,N_34805);
or U36077 (N_36077,N_34320,N_35471);
xnor U36078 (N_36078,N_35600,N_35361);
nor U36079 (N_36079,N_35230,N_34613);
and U36080 (N_36080,N_34846,N_35379);
nor U36081 (N_36081,N_34048,N_35605);
or U36082 (N_36082,N_35276,N_35058);
and U36083 (N_36083,N_34941,N_34732);
and U36084 (N_36084,N_35853,N_34754);
and U36085 (N_36085,N_34299,N_34145);
nand U36086 (N_36086,N_34939,N_35689);
xor U36087 (N_36087,N_35617,N_34335);
and U36088 (N_36088,N_35820,N_35383);
or U36089 (N_36089,N_34124,N_35782);
nand U36090 (N_36090,N_34310,N_35115);
nand U36091 (N_36091,N_34712,N_35775);
or U36092 (N_36092,N_35270,N_34677);
nor U36093 (N_36093,N_35983,N_35074);
xor U36094 (N_36094,N_35604,N_35358);
xor U36095 (N_36095,N_35917,N_34923);
nor U36096 (N_36096,N_35874,N_34875);
or U36097 (N_36097,N_34199,N_35248);
xnor U36098 (N_36098,N_35234,N_34614);
xnor U36099 (N_36099,N_35955,N_34952);
and U36100 (N_36100,N_34709,N_35478);
and U36101 (N_36101,N_35402,N_35895);
xnor U36102 (N_36102,N_34705,N_35596);
and U36103 (N_36103,N_34737,N_35988);
xor U36104 (N_36104,N_34326,N_35006);
and U36105 (N_36105,N_34110,N_34740);
xor U36106 (N_36106,N_35991,N_34810);
or U36107 (N_36107,N_35871,N_35004);
xnor U36108 (N_36108,N_34800,N_34077);
nand U36109 (N_36109,N_34377,N_34935);
or U36110 (N_36110,N_34209,N_35390);
nand U36111 (N_36111,N_34903,N_35859);
and U36112 (N_36112,N_34180,N_34745);
nand U36113 (N_36113,N_34041,N_34512);
nand U36114 (N_36114,N_35176,N_35735);
or U36115 (N_36115,N_34524,N_35307);
or U36116 (N_36116,N_34548,N_35677);
nor U36117 (N_36117,N_34529,N_34725);
or U36118 (N_36118,N_34301,N_35612);
xnor U36119 (N_36119,N_35919,N_34564);
nand U36120 (N_36120,N_34039,N_34502);
xor U36121 (N_36121,N_35540,N_34461);
and U36122 (N_36122,N_35511,N_35198);
and U36123 (N_36123,N_34654,N_34834);
nand U36124 (N_36124,N_34357,N_34925);
nand U36125 (N_36125,N_35531,N_34644);
or U36126 (N_36126,N_35359,N_35099);
or U36127 (N_36127,N_35372,N_34499);
and U36128 (N_36128,N_34042,N_35536);
nor U36129 (N_36129,N_35131,N_35501);
nor U36130 (N_36130,N_34347,N_35756);
and U36131 (N_36131,N_34992,N_35714);
xor U36132 (N_36132,N_34121,N_34298);
and U36133 (N_36133,N_34096,N_35371);
xnor U36134 (N_36134,N_34031,N_35772);
nor U36135 (N_36135,N_34777,N_34661);
and U36136 (N_36136,N_34552,N_34393);
and U36137 (N_36137,N_34523,N_35936);
or U36138 (N_36138,N_34711,N_35937);
xor U36139 (N_36139,N_34703,N_34730);
nor U36140 (N_36140,N_35156,N_35715);
nor U36141 (N_36141,N_35241,N_35100);
or U36142 (N_36142,N_35311,N_35473);
and U36143 (N_36143,N_35942,N_35207);
nand U36144 (N_36144,N_35212,N_34052);
nor U36145 (N_36145,N_34081,N_35444);
nor U36146 (N_36146,N_35171,N_35861);
nand U36147 (N_36147,N_34728,N_35533);
nand U36148 (N_36148,N_34863,N_35255);
nor U36149 (N_36149,N_35578,N_34134);
nand U36150 (N_36150,N_34827,N_34859);
and U36151 (N_36151,N_35681,N_35630);
xnor U36152 (N_36152,N_35970,N_35783);
xor U36153 (N_36153,N_34007,N_34790);
and U36154 (N_36154,N_34664,N_35545);
or U36155 (N_36155,N_34507,N_34118);
nor U36156 (N_36156,N_35899,N_35136);
nand U36157 (N_36157,N_34250,N_35579);
nor U36158 (N_36158,N_35308,N_35202);
and U36159 (N_36159,N_34044,N_35513);
xor U36160 (N_36160,N_34813,N_34683);
and U36161 (N_36161,N_34045,N_34541);
xnor U36162 (N_36162,N_34394,N_35934);
nand U36163 (N_36163,N_35427,N_35254);
and U36164 (N_36164,N_35418,N_35470);
or U36165 (N_36165,N_34167,N_35897);
nor U36166 (N_36166,N_34253,N_34435);
xnor U36167 (N_36167,N_35818,N_35774);
or U36168 (N_36168,N_35521,N_35071);
and U36169 (N_36169,N_35344,N_35232);
nand U36170 (N_36170,N_35304,N_35526);
nand U36171 (N_36171,N_35683,N_35182);
xnor U36172 (N_36172,N_34976,N_35117);
nor U36173 (N_36173,N_34753,N_35582);
nor U36174 (N_36174,N_34806,N_35297);
or U36175 (N_36175,N_34877,N_35087);
nand U36176 (N_36176,N_34874,N_35137);
xor U36177 (N_36177,N_35047,N_34914);
and U36178 (N_36178,N_34088,N_35193);
and U36179 (N_36179,N_35490,N_34238);
nand U36180 (N_36180,N_34318,N_34485);
nor U36181 (N_36181,N_35802,N_35291);
or U36182 (N_36182,N_35458,N_34473);
or U36183 (N_36183,N_34097,N_35694);
nor U36184 (N_36184,N_34761,N_34469);
xor U36185 (N_36185,N_35797,N_35550);
nor U36186 (N_36186,N_35215,N_34876);
or U36187 (N_36187,N_34932,N_35038);
and U36188 (N_36188,N_34902,N_35111);
and U36189 (N_36189,N_35391,N_34517);
and U36190 (N_36190,N_34672,N_34071);
or U36191 (N_36191,N_35589,N_34108);
nand U36192 (N_36192,N_35731,N_35882);
nor U36193 (N_36193,N_35488,N_35077);
or U36194 (N_36194,N_34565,N_34092);
and U36195 (N_36195,N_34372,N_35247);
and U36196 (N_36196,N_34074,N_35367);
nor U36197 (N_36197,N_34078,N_35849);
nor U36198 (N_36198,N_35009,N_34616);
nor U36199 (N_36199,N_34601,N_34645);
and U36200 (N_36200,N_35776,N_34102);
nand U36201 (N_36201,N_35483,N_34781);
or U36202 (N_36202,N_34604,N_34901);
xor U36203 (N_36203,N_35051,N_34228);
xor U36204 (N_36204,N_34772,N_34766);
nor U36205 (N_36205,N_34525,N_35025);
nor U36206 (N_36206,N_35816,N_34618);
and U36207 (N_36207,N_34303,N_35267);
nor U36208 (N_36208,N_34245,N_35869);
and U36209 (N_36209,N_34406,N_34638);
and U36210 (N_36210,N_34530,N_34949);
and U36211 (N_36211,N_34398,N_34599);
or U36212 (N_36212,N_35627,N_34095);
nand U36213 (N_36213,N_34704,N_35128);
xor U36214 (N_36214,N_35479,N_35014);
and U36215 (N_36215,N_34261,N_35147);
and U36216 (N_36216,N_35887,N_35145);
and U36217 (N_36217,N_34955,N_35903);
xnor U36218 (N_36218,N_35445,N_34422);
xnor U36219 (N_36219,N_35794,N_34101);
nand U36220 (N_36220,N_34627,N_34893);
xnor U36221 (N_36221,N_34757,N_35836);
or U36222 (N_36222,N_35964,N_34028);
nor U36223 (N_36223,N_35277,N_34346);
or U36224 (N_36224,N_35839,N_35539);
xor U36225 (N_36225,N_34837,N_34194);
and U36226 (N_36226,N_35956,N_34380);
and U36227 (N_36227,N_35151,N_35054);
nor U36228 (N_36228,N_34629,N_35016);
nand U36229 (N_36229,N_35494,N_35177);
and U36230 (N_36230,N_35012,N_35181);
or U36231 (N_36231,N_35387,N_34315);
and U36232 (N_36232,N_34000,N_35727);
nand U36233 (N_36233,N_35810,N_34069);
and U36234 (N_36234,N_35765,N_34437);
nand U36235 (N_36235,N_35746,N_34578);
nand U36236 (N_36236,N_34662,N_35425);
or U36237 (N_36237,N_35879,N_34807);
or U36238 (N_36238,N_35654,N_34626);
nand U36239 (N_36239,N_35590,N_35468);
nor U36240 (N_36240,N_35841,N_35434);
or U36241 (N_36241,N_35781,N_35906);
and U36242 (N_36242,N_35586,N_35748);
nor U36243 (N_36243,N_35062,N_34275);
or U36244 (N_36244,N_34900,N_35965);
nand U36245 (N_36245,N_34791,N_34288);
or U36246 (N_36246,N_35985,N_34587);
nor U36247 (N_36247,N_34091,N_35236);
xnor U36248 (N_36248,N_35284,N_34693);
and U36249 (N_36249,N_34624,N_35522);
or U36250 (N_36250,N_35668,N_35365);
nor U36251 (N_36251,N_35368,N_35346);
nor U36252 (N_36252,N_34792,N_35646);
nand U36253 (N_36253,N_35085,N_35024);
nor U36254 (N_36254,N_34033,N_34389);
or U36255 (N_36255,N_34522,N_35377);
nor U36256 (N_36256,N_34963,N_34202);
or U36257 (N_36257,N_35339,N_35670);
nor U36258 (N_36258,N_35327,N_34242);
xnor U36259 (N_36259,N_34159,N_35263);
nand U36260 (N_36260,N_35624,N_34894);
and U36261 (N_36261,N_35423,N_34285);
and U36262 (N_36262,N_35846,N_35747);
and U36263 (N_36263,N_34073,N_34594);
xor U36264 (N_36264,N_35245,N_35957);
nand U36265 (N_36265,N_35930,N_34714);
nand U36266 (N_36266,N_34403,N_34224);
xnor U36267 (N_36267,N_34615,N_34960);
xor U36268 (N_36268,N_35873,N_34852);
xnor U36269 (N_36269,N_35194,N_34668);
and U36270 (N_36270,N_35966,N_35000);
nand U36271 (N_36271,N_34741,N_35103);
nor U36272 (N_36272,N_34980,N_34602);
and U36273 (N_36273,N_35121,N_34946);
nand U36274 (N_36274,N_34723,N_34188);
or U36275 (N_36275,N_34414,N_34650);
nor U36276 (N_36276,N_34294,N_34503);
nor U36277 (N_36277,N_35105,N_34688);
xor U36278 (N_36278,N_34133,N_34775);
xor U36279 (N_36279,N_34400,N_35457);
or U36280 (N_36280,N_34550,N_34127);
nor U36281 (N_36281,N_34481,N_35002);
nor U36282 (N_36282,N_34061,N_35082);
nor U36283 (N_36283,N_34112,N_34090);
or U36284 (N_36284,N_34256,N_34451);
or U36285 (N_36285,N_34370,N_34486);
xor U36286 (N_36286,N_34783,N_34579);
or U36287 (N_36287,N_34561,N_34453);
and U36288 (N_36288,N_35360,N_34853);
xnor U36289 (N_36289,N_34718,N_35127);
nor U36290 (N_36290,N_35565,N_35272);
nor U36291 (N_36291,N_35489,N_34833);
nor U36292 (N_36292,N_34079,N_35114);
and U36293 (N_36293,N_34971,N_34483);
nor U36294 (N_36294,N_34032,N_34888);
nand U36295 (N_36295,N_35953,N_35227);
or U36296 (N_36296,N_35443,N_34828);
and U36297 (N_36297,N_34402,N_35939);
nor U36298 (N_36298,N_34396,N_35560);
nand U36299 (N_36299,N_34633,N_35003);
xor U36300 (N_36300,N_35635,N_35028);
nand U36301 (N_36301,N_34919,N_35070);
xnor U36302 (N_36302,N_35821,N_35113);
and U36303 (N_36303,N_35150,N_35048);
nor U36304 (N_36304,N_35091,N_34291);
nand U36305 (N_36305,N_34429,N_35692);
or U36306 (N_36306,N_35461,N_35996);
nor U36307 (N_36307,N_35132,N_35433);
and U36308 (N_36308,N_34043,N_34518);
nor U36309 (N_36309,N_35938,N_35329);
xnor U36310 (N_36310,N_35732,N_34751);
xnor U36311 (N_36311,N_35296,N_34412);
nor U36312 (N_36312,N_34493,N_35250);
and U36313 (N_36313,N_34538,N_34917);
nand U36314 (N_36314,N_34012,N_34839);
and U36315 (N_36315,N_34549,N_35858);
nand U36316 (N_36316,N_34177,N_35349);
nand U36317 (N_36317,N_35569,N_34094);
xnor U36318 (N_36318,N_35703,N_34912);
nand U36319 (N_36319,N_35602,N_35905);
or U36320 (N_36320,N_34008,N_34479);
nor U36321 (N_36321,N_34314,N_35357);
nor U36322 (N_36322,N_34722,N_35778);
nand U36323 (N_36323,N_34205,N_34086);
or U36324 (N_36324,N_34968,N_35352);
nand U36325 (N_36325,N_34082,N_34904);
nor U36326 (N_36326,N_34116,N_35476);
nor U36327 (N_36327,N_34267,N_35110);
or U36328 (N_36328,N_35010,N_35971);
nand U36329 (N_36329,N_34390,N_34213);
nor U36330 (N_36330,N_35753,N_35574);
xor U36331 (N_36331,N_34063,N_35926);
nand U36332 (N_36332,N_34055,N_34018);
xor U36333 (N_36333,N_35106,N_34427);
nand U36334 (N_36334,N_34560,N_34141);
nand U36335 (N_36335,N_35279,N_34219);
nand U36336 (N_36336,N_34996,N_34411);
nand U36337 (N_36337,N_35647,N_34821);
nand U36338 (N_36338,N_35382,N_35200);
nand U36339 (N_36339,N_35587,N_35711);
nand U36340 (N_36340,N_34038,N_34710);
or U36341 (N_36341,N_34641,N_34210);
nor U36342 (N_36342,N_35626,N_34870);
or U36343 (N_36343,N_34836,N_34913);
nand U36344 (N_36344,N_35686,N_34563);
and U36345 (N_36345,N_34047,N_35164);
nor U36346 (N_36346,N_34474,N_35969);
nand U36347 (N_36347,N_35076,N_34305);
or U36348 (N_36348,N_35561,N_35097);
or U36349 (N_36349,N_34956,N_34924);
nand U36350 (N_36350,N_34617,N_35287);
and U36351 (N_36351,N_35655,N_35240);
nand U36352 (N_36352,N_34640,N_35682);
and U36353 (N_36353,N_35381,N_35422);
and U36354 (N_36354,N_35543,N_35648);
nand U36355 (N_36355,N_35914,N_34665);
nor U36356 (N_36356,N_34378,N_35631);
or U36357 (N_36357,N_35410,N_35322);
or U36358 (N_36358,N_34966,N_34099);
and U36359 (N_36359,N_34931,N_34929);
and U36360 (N_36360,N_35237,N_34017);
or U36361 (N_36361,N_34409,N_35834);
nor U36362 (N_36362,N_35595,N_34537);
nand U36363 (N_36363,N_34154,N_34252);
nand U36364 (N_36364,N_35021,N_34573);
nand U36365 (N_36365,N_35052,N_35736);
xnor U36366 (N_36366,N_35657,N_35761);
and U36367 (N_36367,N_34439,N_35502);
nand U36368 (N_36368,N_34114,N_35231);
xor U36369 (N_36369,N_34105,N_34068);
or U36370 (N_36370,N_35651,N_34804);
and U36371 (N_36371,N_34520,N_35188);
or U36372 (N_36372,N_35043,N_35300);
and U36373 (N_36373,N_34359,N_35876);
xor U36374 (N_36374,N_35395,N_35354);
and U36375 (N_36375,N_35321,N_35323);
xor U36376 (N_36376,N_35397,N_35661);
and U36377 (N_36377,N_35454,N_34184);
nor U36378 (N_36378,N_35049,N_34132);
xor U36379 (N_36379,N_35497,N_34690);
or U36380 (N_36380,N_35573,N_34636);
xnor U36381 (N_36381,N_35057,N_35216);
nor U36382 (N_36382,N_35598,N_35301);
xor U36383 (N_36383,N_34799,N_34660);
and U36384 (N_36384,N_34570,N_34339);
nor U36385 (N_36385,N_35447,N_34014);
or U36386 (N_36386,N_35503,N_34947);
nand U36387 (N_36387,N_35716,N_34990);
nor U36388 (N_36388,N_35822,N_35973);
or U36389 (N_36389,N_35591,N_35481);
nor U36390 (N_36390,N_35165,N_35817);
or U36391 (N_36391,N_34967,N_34084);
or U36392 (N_36392,N_34826,N_34679);
xnor U36393 (N_36393,N_34340,N_35157);
and U36394 (N_36394,N_35017,N_34490);
nor U36395 (N_36395,N_35168,N_35409);
nor U36396 (N_36396,N_34172,N_35396);
nand U36397 (N_36397,N_34752,N_35325);
and U36398 (N_36398,N_34700,N_35777);
and U36399 (N_36399,N_34207,N_35636);
xor U36400 (N_36400,N_35644,N_34943);
nand U36401 (N_36401,N_34215,N_35228);
and U36402 (N_36402,N_35941,N_34953);
and U36403 (N_36403,N_35528,N_34345);
or U36404 (N_36404,N_35482,N_35266);
nand U36405 (N_36405,N_34200,N_34854);
and U36406 (N_36406,N_35465,N_34268);
or U36407 (N_36407,N_34743,N_35239);
and U36408 (N_36408,N_35485,N_34801);
nor U36409 (N_36409,N_35886,N_35653);
nor U36410 (N_36410,N_34191,N_35226);
or U36411 (N_36411,N_35555,N_35195);
xnor U36412 (N_36412,N_35345,N_35787);
xor U36413 (N_36413,N_34659,N_35450);
and U36414 (N_36414,N_34060,N_35880);
xnor U36415 (N_36415,N_35336,N_34696);
nor U36416 (N_36416,N_35441,N_35637);
xnor U36417 (N_36417,N_35740,N_34443);
nand U36418 (N_36418,N_34596,N_34729);
or U36419 (N_36419,N_34386,N_34779);
nand U36420 (N_36420,N_35011,N_35394);
or U36421 (N_36421,N_34687,N_35238);
xor U36422 (N_36422,N_35133,N_35069);
nor U36423 (N_36423,N_34897,N_34482);
xnor U36424 (N_36424,N_34366,N_34630);
xnor U36425 (N_36425,N_35684,N_34764);
and U36426 (N_36426,N_35527,N_35439);
xor U36427 (N_36427,N_35650,N_34109);
and U36428 (N_36428,N_34449,N_34150);
or U36429 (N_36429,N_35388,N_35178);
nor U36430 (N_36430,N_34887,N_35722);
nand U36431 (N_36431,N_35122,N_35404);
and U36432 (N_36432,N_34658,N_34379);
nor U36433 (N_36433,N_35842,N_35083);
nor U36434 (N_36434,N_35924,N_34815);
or U36435 (N_36435,N_35629,N_34126);
nand U36436 (N_36436,N_35155,N_34260);
and U36437 (N_36437,N_35860,N_35107);
nand U36438 (N_36438,N_34566,N_34915);
nand U36439 (N_36439,N_34719,N_34405);
and U36440 (N_36440,N_35658,N_34500);
and U36441 (N_36441,N_34222,N_34878);
or U36442 (N_36442,N_35826,N_35205);
xnor U36443 (N_36443,N_34162,N_35623);
or U36444 (N_36444,N_35912,N_34610);
and U36445 (N_36445,N_34882,N_34857);
and U36446 (N_36446,N_35334,N_34509);
and U36447 (N_36447,N_35980,N_35348);
xnor U36448 (N_36448,N_34954,N_34111);
nor U36449 (N_36449,N_35801,N_35370);
nand U36450 (N_36450,N_34982,N_35932);
xor U36451 (N_36451,N_34365,N_35743);
nand U36452 (N_36452,N_35328,N_34323);
and U36453 (N_36453,N_35034,N_35326);
nor U36454 (N_36454,N_35663,N_35197);
nor U36455 (N_36455,N_34342,N_35749);
and U36456 (N_36456,N_34006,N_35015);
or U36457 (N_36457,N_35420,N_35362);
or U36458 (N_36458,N_34138,N_35175);
xor U36459 (N_36459,N_35729,N_34391);
xor U36460 (N_36460,N_35518,N_35019);
xor U36461 (N_36461,N_35438,N_35844);
or U36462 (N_36462,N_34113,N_35744);
xor U36463 (N_36463,N_34249,N_35866);
nand U36464 (N_36464,N_34495,N_35073);
nand U36465 (N_36465,N_35752,N_34803);
nor U36466 (N_36466,N_35862,N_34861);
nand U36467 (N_36467,N_34717,N_35910);
nand U36468 (N_36468,N_34065,N_35351);
nand U36469 (N_36469,N_34684,N_35916);
nor U36470 (N_36470,N_34284,N_35718);
xnor U36471 (N_36471,N_34183,N_35529);
nand U36472 (N_36472,N_35104,N_35101);
xnor U36473 (N_36473,N_34234,N_34583);
nand U36474 (N_36474,N_35733,N_35833);
nand U36475 (N_36475,N_35896,N_35314);
nand U36476 (N_36476,N_35976,N_35763);
nand U36477 (N_36477,N_34363,N_34950);
nor U36478 (N_36478,N_35566,N_34369);
nor U36479 (N_36479,N_35755,N_35620);
or U36480 (N_36480,N_35641,N_34991);
nor U36481 (N_36481,N_35773,N_35261);
or U36482 (N_36482,N_35562,N_34848);
or U36483 (N_36483,N_35995,N_35577);
nand U36484 (N_36484,N_35621,N_34958);
nand U36485 (N_36485,N_35224,N_35319);
nand U36486 (N_36486,N_35639,N_35556);
or U36487 (N_36487,N_34588,N_35166);
nand U36488 (N_36488,N_35614,N_35676);
xnor U36489 (N_36489,N_35405,N_35152);
or U36490 (N_36490,N_35134,N_35870);
or U36491 (N_36491,N_35472,N_35213);
xor U36492 (N_36492,N_35567,N_35417);
and U36493 (N_36493,N_34970,N_34144);
nand U36494 (N_36494,N_34179,N_35649);
nand U36495 (N_36495,N_35616,N_34584);
and U36496 (N_36496,N_34930,N_34013);
xor U36497 (N_36497,N_35524,N_34170);
and U36498 (N_36498,N_35688,N_34721);
nand U36499 (N_36499,N_34623,N_34759);
xnor U36500 (N_36500,N_35597,N_34621);
and U36501 (N_36501,N_34731,N_34064);
or U36502 (N_36502,N_35534,N_34166);
nand U36503 (N_36503,N_34460,N_34383);
nor U36504 (N_36504,N_35519,N_34168);
and U36505 (N_36505,N_34104,N_35112);
and U36506 (N_36506,N_34217,N_34446);
and U36507 (N_36507,N_34993,N_34050);
nor U36508 (N_36508,N_34122,N_34015);
nor U36509 (N_36509,N_34332,N_34760);
and U36510 (N_36510,N_35159,N_34281);
and U36511 (N_36511,N_35712,N_34497);
and U36512 (N_36512,N_35544,N_35719);
nand U36513 (N_36513,N_34997,N_34160);
nand U36514 (N_36514,N_35935,N_34663);
or U36515 (N_36515,N_34201,N_35353);
nand U36516 (N_36516,N_35889,N_34973);
nor U36517 (N_36517,N_34333,N_35143);
or U36518 (N_36518,N_34328,N_35538);
xor U36519 (N_36519,N_35766,N_35446);
nor U36520 (N_36520,N_35455,N_35271);
xor U36521 (N_36521,N_34325,N_35373);
nor U36522 (N_36522,N_35599,N_34466);
nand U36523 (N_36523,N_35153,N_35603);
and U36524 (N_36524,N_35552,N_35979);
nor U36525 (N_36525,N_35007,N_35464);
xnor U36526 (N_36526,N_34130,N_35967);
nand U36527 (N_36527,N_34592,N_34825);
or U36528 (N_36528,N_35229,N_34832);
and U36529 (N_36529,N_34478,N_34851);
nor U36530 (N_36530,N_34922,N_35340);
and U36531 (N_36531,N_34796,N_34646);
and U36532 (N_36532,N_35710,N_34539);
xnor U36533 (N_36533,N_35699,N_34891);
nand U36534 (N_36534,N_34504,N_34410);
xnor U36535 (N_36535,N_35305,N_34998);
and U36536 (N_36536,N_34536,N_35811);
xor U36537 (N_36537,N_34978,N_34909);
nor U36538 (N_36538,N_35815,N_35827);
and U36539 (N_36539,N_34979,N_35135);
and U36540 (N_36540,N_35666,N_34083);
nand U36541 (N_36541,N_35848,N_35242);
or U36542 (N_36542,N_35299,N_34336);
xnor U36543 (N_36543,N_34841,N_35280);
xnor U36544 (N_36544,N_35078,N_34480);
xnor U36545 (N_36545,N_35588,N_35642);
or U36546 (N_36546,N_35302,N_35804);
or U36547 (N_36547,N_34830,N_35974);
xnor U36548 (N_36548,N_35431,N_34304);
nand U36549 (N_36549,N_34415,N_35056);
nor U36550 (N_36550,N_34498,N_35116);
or U36551 (N_36551,N_34066,N_34785);
nand U36552 (N_36552,N_34678,N_35695);
nand U36553 (N_36553,N_34475,N_34755);
or U36554 (N_36554,N_34046,N_34569);
and U36555 (N_36555,N_34484,N_35063);
xnor U36556 (N_36556,N_34165,N_35259);
and U36557 (N_36557,N_34426,N_35211);
and U36558 (N_36558,N_35293,N_35295);
or U36559 (N_36559,N_34212,N_35440);
and U36560 (N_36560,N_35790,N_35881);
nand U36561 (N_36561,N_34534,N_35281);
or U36562 (N_36562,N_35192,N_35480);
nand U36563 (N_36563,N_34231,N_34697);
or U36564 (N_36564,N_35851,N_35864);
and U36565 (N_36565,N_35369,N_34959);
xor U36566 (N_36566,N_34270,N_35179);
nand U36567 (N_36567,N_34628,N_34140);
and U36568 (N_36568,N_34421,N_34809);
nand U36569 (N_36569,N_34739,N_34467);
nand U36570 (N_36570,N_34771,N_34300);
nand U36571 (N_36571,N_35350,N_35093);
and U36572 (N_36572,N_35313,N_35809);
and U36573 (N_36573,N_34748,N_34576);
nand U36574 (N_36574,N_35907,N_35032);
xor U36575 (N_36575,N_34164,N_35981);
nor U36576 (N_36576,N_34178,N_35316);
xnor U36577 (N_36577,N_34715,N_34049);
and U36578 (N_36578,N_34948,N_34643);
xor U36579 (N_36579,N_34375,N_35274);
xor U36580 (N_36580,N_34035,N_35918);
and U36581 (N_36581,N_34965,N_35257);
and U36582 (N_36582,N_34648,N_34425);
or U36583 (N_36583,N_34158,N_35947);
xnor U36584 (N_36584,N_35987,N_35581);
or U36585 (N_36585,N_35922,N_34277);
nand U36586 (N_36586,N_34797,N_34196);
nor U36587 (N_36587,N_35506,N_35413);
xor U36588 (N_36588,N_34487,N_35931);
and U36589 (N_36589,N_34037,N_34254);
xnor U36590 (N_36590,N_34169,N_34330);
or U36591 (N_36591,N_35608,N_34637);
nand U36592 (N_36592,N_35542,N_34937);
nor U36593 (N_36593,N_35268,N_34392);
nor U36594 (N_36594,N_35872,N_35392);
nor U36595 (N_36595,N_35315,N_35429);
nand U36596 (N_36596,N_34788,N_35913);
nand U36597 (N_36597,N_34009,N_34543);
xnor U36598 (N_36598,N_35726,N_35335);
xor U36599 (N_36599,N_34961,N_34174);
nand U36600 (N_36600,N_34899,N_35702);
or U36601 (N_36601,N_34026,N_35788);
nor U36602 (N_36602,N_35499,N_34442);
nand U36603 (N_36603,N_35278,N_35144);
nor U36604 (N_36604,N_35375,N_35096);
or U36605 (N_36605,N_35977,N_35282);
nor U36606 (N_36606,N_34258,N_35094);
or U36607 (N_36607,N_34575,N_35199);
and U36608 (N_36608,N_34100,N_35487);
nand U36609 (N_36609,N_35338,N_34554);
or U36610 (N_36610,N_34376,N_35514);
nor U36611 (N_36611,N_34259,N_34351);
xnor U36612 (N_36612,N_35767,N_34526);
xor U36613 (N_36613,N_35026,N_35366);
nand U36614 (N_36614,N_34293,N_35123);
nor U36615 (N_36615,N_35671,N_35800);
or U36616 (N_36616,N_35771,N_34508);
and U36617 (N_36617,N_34972,N_34273);
nor U36618 (N_36618,N_35796,N_35374);
xnor U36619 (N_36619,N_35784,N_34190);
nor U36620 (N_36620,N_34634,N_34556);
and U36621 (N_36621,N_34087,N_35084);
nand U36622 (N_36622,N_34384,N_35050);
xor U36623 (N_36623,N_35709,N_35678);
xnor U36624 (N_36624,N_34255,N_35532);
xor U36625 (N_36625,N_35416,N_35244);
or U36626 (N_36626,N_35865,N_34148);
and U36627 (N_36627,N_34235,N_35005);
xor U36628 (N_36628,N_35525,N_35419);
and U36629 (N_36629,N_34942,N_35553);
nand U36630 (N_36630,N_34767,N_34053);
nor U36631 (N_36631,N_35795,N_34984);
and U36632 (N_36632,N_35341,N_35462);
nand U36633 (N_36633,N_35915,N_34265);
nor U36634 (N_36634,N_35535,N_35972);
nand U36635 (N_36635,N_35061,N_34135);
xor U36636 (N_36636,N_34321,N_35952);
nor U36637 (N_36637,N_35332,N_34156);
and U36638 (N_36638,N_35246,N_35713);
nor U36639 (N_36639,N_34289,N_34608);
nand U36640 (N_36640,N_35475,N_34501);
nor U36641 (N_36641,N_34653,N_35029);
and U36642 (N_36642,N_34746,N_34944);
xor U36643 (N_36643,N_35496,N_34417);
xnor U36644 (N_36644,N_34176,N_35610);
xor U36645 (N_36645,N_35593,N_34632);
nand U36646 (N_36646,N_35060,N_35500);
or U36647 (N_36647,N_35769,N_35331);
nor U36648 (N_36648,N_35933,N_34577);
nand U36649 (N_36649,N_35723,N_35436);
nor U36650 (N_36650,N_35508,N_35923);
and U36651 (N_36651,N_35885,N_35551);
and U36652 (N_36652,N_34515,N_35807);
nor U36653 (N_36653,N_35102,N_35852);
nand U36654 (N_36654,N_34812,N_34910);
nand U36655 (N_36655,N_34666,N_34155);
xor U36656 (N_36656,N_35492,N_35559);
or U36657 (N_36657,N_34720,N_34491);
and U36658 (N_36658,N_34203,N_35611);
and U36659 (N_36659,N_35814,N_34142);
nor U36660 (N_36660,N_35068,N_35946);
or U36661 (N_36661,N_35576,N_35813);
or U36662 (N_36662,N_35090,N_35857);
and U36663 (N_36663,N_34244,N_34692);
or U36664 (N_36664,N_35920,N_34353);
or U36665 (N_36665,N_35613,N_35721);
nor U36666 (N_36666,N_35812,N_35298);
nand U36667 (N_36667,N_35994,N_35355);
nand U36668 (N_36668,N_34016,N_35672);
nand U36669 (N_36669,N_34838,N_34186);
xor U36670 (N_36670,N_35498,N_34597);
or U36671 (N_36671,N_34708,N_34171);
and U36672 (N_36672,N_34713,N_34620);
or U36673 (N_36673,N_34331,N_35386);
xnor U36674 (N_36674,N_34371,N_34283);
and U36675 (N_36675,N_34456,N_35186);
and U36676 (N_36676,N_35258,N_35805);
xor U36677 (N_36677,N_34595,N_35690);
nor U36678 (N_36678,N_34001,N_35950);
or U36679 (N_36679,N_34407,N_34139);
and U36680 (N_36680,N_35495,N_35799);
nor U36681 (N_36681,N_34975,N_35260);
and U36682 (N_36682,N_34886,N_34865);
nor U36683 (N_36683,N_35027,N_35592);
nor U36684 (N_36684,N_34682,N_34770);
or U36685 (N_36685,N_35606,N_35252);
xor U36686 (N_36686,N_34387,N_35185);
and U36687 (N_36687,N_35888,N_34286);
nand U36688 (N_36688,N_35214,N_34675);
nand U36689 (N_36689,N_35163,N_35758);
or U36690 (N_36690,N_34204,N_35033);
or U36691 (N_36691,N_34674,N_34418);
nand U36692 (N_36692,N_35825,N_35768);
nor U36693 (N_36693,N_35218,N_35958);
xor U36694 (N_36694,N_34793,N_35982);
nor U36695 (N_36695,N_34698,N_35541);
and U36696 (N_36696,N_34811,N_34471);
and U36697 (N_36697,N_34974,N_35660);
or U36698 (N_36698,N_34987,N_34419);
or U36699 (N_36699,N_34408,N_34798);
nand U36700 (N_36700,N_34892,N_34535);
and U36701 (N_36701,N_34056,N_35537);
and U36702 (N_36702,N_35680,N_35558);
or U36703 (N_36703,N_34808,N_35824);
xor U36704 (N_36704,N_35364,N_35092);
or U36705 (N_36705,N_35789,N_35220);
and U36706 (N_36706,N_34225,N_35868);
xnor U36707 (N_36707,N_35160,N_34600);
nand U36708 (N_36708,N_34274,N_35845);
or U36709 (N_36709,N_35643,N_35949);
or U36710 (N_36710,N_34605,N_35294);
nor U36711 (N_36711,N_35530,N_35256);
nand U36712 (N_36712,N_34358,N_35734);
and U36713 (N_36713,N_34440,N_35453);
xnor U36714 (N_36714,N_34233,N_35679);
nand U36715 (N_36715,N_34510,N_34896);
or U36716 (N_36716,N_34562,N_35285);
nor U36717 (N_36717,N_35398,N_35548);
or U36718 (N_36718,N_34404,N_35564);
and U36719 (N_36719,N_34858,N_35306);
nand U36720 (N_36720,N_34143,N_34706);
nor U36721 (N_36721,N_34557,N_35928);
or U36722 (N_36722,N_34680,N_34308);
and U36723 (N_36723,N_35554,N_35180);
nor U36724 (N_36724,N_34747,N_35459);
nor U36725 (N_36725,N_34117,N_35040);
nand U36726 (N_36726,N_35618,N_34367);
xnor U36727 (N_36727,N_35696,N_34794);
nor U36728 (N_36728,N_35437,N_34424);
nor U36729 (N_36729,N_34527,N_34867);
nor U36730 (N_36730,N_34181,N_34603);
nand U36731 (N_36731,N_35632,N_35042);
nor U36732 (N_36732,N_34847,N_34373);
nand U36733 (N_36733,N_35243,N_34040);
and U36734 (N_36734,N_35878,N_34727);
or U36735 (N_36735,N_34356,N_34452);
nand U36736 (N_36736,N_35992,N_35547);
nor U36737 (N_36737,N_35962,N_35832);
or U36738 (N_36738,N_34010,N_35219);
xor U36739 (N_36739,N_34067,N_34307);
nand U36740 (N_36740,N_34749,N_35900);
nor U36741 (N_36741,N_34296,N_35619);
nand U36742 (N_36742,N_35129,N_34591);
or U36743 (N_36743,N_34334,N_35925);
or U36744 (N_36744,N_34671,N_34951);
nor U36745 (N_36745,N_35075,N_35999);
and U36746 (N_36746,N_34983,N_35803);
nand U36747 (N_36747,N_34670,N_35516);
and U36748 (N_36748,N_35172,N_34651);
and U36749 (N_36749,N_34631,N_34208);
and U36750 (N_36750,N_34780,N_35850);
and U36751 (N_36751,N_34860,N_34187);
or U36752 (N_36752,N_34136,N_35189);
xor U36753 (N_36753,N_35430,N_34151);
or U36754 (N_36754,N_35856,N_35867);
nor U36755 (N_36755,N_35786,N_35568);
nand U36756 (N_36756,N_35310,N_35233);
or U36757 (N_36757,N_35884,N_34619);
xnor U36758 (N_36758,N_35406,N_34574);
nand U36759 (N_36759,N_34989,N_35108);
nand U36760 (N_36760,N_34450,N_35819);
nand U36761 (N_36761,N_34957,N_35162);
and U36762 (N_36762,N_34232,N_35309);
nor U36763 (N_36763,N_34239,N_35095);
nand U36764 (N_36764,N_35421,N_34316);
or U36765 (N_36765,N_34297,N_34189);
xor U36766 (N_36766,N_35855,N_34945);
or U36767 (N_36767,N_35717,N_35424);
or U36768 (N_36768,N_34229,N_35908);
nand U36769 (N_36769,N_35615,N_34364);
nor U36770 (N_36770,N_35628,N_34985);
nor U36771 (N_36771,N_35426,N_34004);
and U36772 (N_36772,N_35407,N_34445);
nand U36773 (N_36773,N_34938,N_34243);
xnor U36774 (N_36774,N_35401,N_34221);
or U36775 (N_36775,N_35389,N_35520);
xnor U36776 (N_36776,N_35442,N_35669);
nand U36777 (N_36777,N_34062,N_35173);
nand U36778 (N_36778,N_34784,N_34149);
xnor U36779 (N_36779,N_34927,N_34625);
nor U36780 (N_36780,N_35697,N_34934);
and U36781 (N_36781,N_35890,N_35484);
nand U36782 (N_36782,N_35428,N_34817);
or U36783 (N_36783,N_35303,N_34476);
or U36784 (N_36784,N_34519,N_35720);
nand U36785 (N_36785,N_34553,N_34397);
and U36786 (N_36786,N_35959,N_34317);
or U36787 (N_36787,N_35235,N_35762);
xnor U36788 (N_36788,N_34468,N_35055);
nand U36789 (N_36789,N_35290,N_35877);
or U36790 (N_36790,N_35563,N_35580);
xor U36791 (N_36791,N_34218,N_35640);
and U36792 (N_36792,N_34214,N_34350);
or U36793 (N_36793,N_34622,N_35652);
nand U36794 (N_36794,N_35609,N_34685);
nand U36795 (N_36795,N_34220,N_34890);
and U36796 (N_36796,N_34933,N_35288);
nand U36797 (N_36797,N_35549,N_35901);
and U36798 (N_36798,N_35840,N_34920);
and U36799 (N_36799,N_35759,N_34494);
nor U36800 (N_36800,N_35902,N_35013);
nor U36801 (N_36801,N_35645,N_34532);
nand U36802 (N_36802,N_34020,N_35403);
nand U36803 (N_36803,N_35089,N_34612);
xor U36804 (N_36804,N_34319,N_34230);
xor U36805 (N_36805,N_34195,N_35854);
xnor U36806 (N_36806,N_35708,N_34883);
xor U36807 (N_36807,N_34586,N_34348);
or U36808 (N_36808,N_34030,N_34738);
nand U36809 (N_36809,N_34926,N_35863);
or U36810 (N_36810,N_35039,N_35673);
and U36811 (N_36811,N_34464,N_34216);
xor U36812 (N_36812,N_35273,N_34362);
xnor U36813 (N_36813,N_35251,N_35337);
xor U36814 (N_36814,N_35312,N_34076);
and U36815 (N_36815,N_35754,N_34673);
xor U36816 (N_36816,N_35512,N_34907);
or U36817 (N_36817,N_35738,N_34123);
nand U36818 (N_36818,N_34119,N_34051);
or U36819 (N_36819,N_35960,N_35023);
or U36820 (N_36820,N_35691,N_34416);
nand U36821 (N_36821,N_34147,N_34448);
nor U36822 (N_36822,N_35384,N_34432);
nor U36823 (N_36823,N_34656,N_35546);
and U36824 (N_36824,N_35411,N_35432);
nand U36825 (N_36825,N_35206,N_35140);
and U36826 (N_36826,N_34115,N_34816);
nand U36827 (N_36827,N_35978,N_34768);
nor U36828 (N_36828,N_34511,N_35875);
and U36829 (N_36829,N_34106,N_35190);
nand U36830 (N_36830,N_34248,N_35045);
nor U36831 (N_36831,N_34582,N_35739);
or U36832 (N_36832,N_34840,N_35700);
and U36833 (N_36833,N_35041,N_34226);
or U36834 (N_36834,N_34782,N_34681);
xnor U36835 (N_36835,N_35779,N_34567);
and U36836 (N_36836,N_35320,N_34036);
nor U36837 (N_36837,N_34880,N_35662);
nand U36838 (N_36838,N_34824,N_34676);
and U36839 (N_36839,N_34551,N_34581);
xor U36840 (N_36840,N_35764,N_34354);
nor U36841 (N_36841,N_34399,N_34750);
and U36842 (N_36842,N_35951,N_34898);
or U36843 (N_36843,N_35141,N_34322);
or U36844 (N_36844,N_35183,N_35601);
nor U36845 (N_36845,N_34223,N_35196);
and U36846 (N_36846,N_34075,N_34829);
xnor U36847 (N_36847,N_34264,N_35126);
nand U36848 (N_36848,N_35001,N_35031);
nor U36849 (N_36849,N_34262,N_34423);
nand U36850 (N_36850,N_34338,N_34528);
and U36851 (N_36851,N_35161,N_34192);
nor U36852 (N_36852,N_35289,N_34327);
xor U36853 (N_36853,N_35412,N_35064);
and U36854 (N_36854,N_34885,N_35363);
nor U36855 (N_36855,N_34125,N_34736);
nor U36856 (N_36856,N_35080,N_34611);
xor U36857 (N_36857,N_35904,N_35557);
nand U36858 (N_36858,N_34352,N_34879);
or U36859 (N_36859,N_34999,N_35008);
or U36860 (N_36860,N_35059,N_34093);
or U36861 (N_36861,N_35275,N_35249);
and U36862 (N_36862,N_34814,N_34128);
xnor U36863 (N_36863,N_34916,N_34868);
xnor U36864 (N_36864,N_34278,N_35724);
nor U36865 (N_36865,N_35793,N_35943);
nor U36866 (N_36866,N_34388,N_34027);
xor U36867 (N_36867,N_34185,N_35463);
and U36868 (N_36868,N_35393,N_34237);
xor U36869 (N_36869,N_35698,N_34470);
xor U36870 (N_36870,N_34988,N_34702);
nand U36871 (N_36871,N_35330,N_35823);
nor U36872 (N_36872,N_34489,N_35469);
nand U36873 (N_36873,N_35158,N_35847);
and U36874 (N_36874,N_35507,N_35449);
nor U36875 (N_36875,N_35452,N_35118);
and U36876 (N_36876,N_34969,N_34003);
nand U36877 (N_36877,N_34034,N_35687);
nor U36878 (N_36878,N_34021,N_35169);
xnor U36879 (N_36879,N_34559,N_34590);
xor U36880 (N_36880,N_34441,N_35378);
nor U36881 (N_36881,N_35451,N_34306);
and U36882 (N_36882,N_34647,N_34381);
or U36883 (N_36883,N_35737,N_35707);
nor U36884 (N_36884,N_34236,N_35829);
or U36885 (N_36885,N_34246,N_34940);
nor U36886 (N_36886,N_34329,N_34313);
or U36887 (N_36887,N_34349,N_34850);
and U36888 (N_36888,N_34455,N_35020);
nand U36889 (N_36889,N_34540,N_34744);
or U36890 (N_36890,N_35583,N_34689);
nand U36891 (N_36891,N_34994,N_35760);
nand U36892 (N_36892,N_34153,N_34607);
or U36893 (N_36893,N_34011,N_34157);
and U36894 (N_36894,N_35929,N_34819);
or U36895 (N_36895,N_35342,N_34716);
xnor U36896 (N_36896,N_35993,N_35292);
nor U36897 (N_36897,N_35380,N_35486);
and U36898 (N_36898,N_35656,N_35415);
nor U36899 (N_36899,N_35035,N_34843);
or U36900 (N_36900,N_35204,N_35791);
nand U36901 (N_36901,N_35170,N_34431);
or U36902 (N_36902,N_35523,N_35022);
nor U36903 (N_36903,N_34542,N_35675);
nand U36904 (N_36904,N_34382,N_35961);
xnor U36905 (N_36905,N_34669,N_35944);
or U36906 (N_36906,N_34657,N_35167);
xor U36907 (N_36907,N_34778,N_34505);
and U36908 (N_36908,N_35725,N_34884);
and U36909 (N_36909,N_35030,N_34002);
and U36910 (N_36910,N_34025,N_35505);
and U36911 (N_36911,N_34459,N_35770);
and U36912 (N_36912,N_34103,N_34465);
or U36913 (N_36913,N_34263,N_35989);
nand U36914 (N_36914,N_35509,N_34977);
nand U36915 (N_36915,N_34776,N_34918);
nor U36916 (N_36916,N_35081,N_34758);
or U36917 (N_36917,N_34182,N_34639);
or U36918 (N_36918,N_35742,N_34835);
or U36919 (N_36919,N_34019,N_34492);
nor U36920 (N_36920,N_35203,N_35664);
and U36921 (N_36921,N_34871,N_34271);
nand U36922 (N_36922,N_34198,N_34368);
or U36923 (N_36923,N_35187,N_35730);
xor U36924 (N_36924,N_34869,N_34070);
or U36925 (N_36925,N_35911,N_35223);
nand U36926 (N_36926,N_34295,N_35892);
or U36927 (N_36927,N_34691,N_35504);
xor U36928 (N_36928,N_34726,N_34211);
xnor U36929 (N_36929,N_34355,N_34606);
and U36930 (N_36930,N_35997,N_35264);
and U36931 (N_36931,N_34818,N_34964);
nand U36932 (N_36932,N_34699,N_34555);
nand U36933 (N_36933,N_35750,N_35088);
nor U36934 (N_36934,N_34589,N_35622);
nand U36935 (N_36935,N_34022,N_34742);
xnor U36936 (N_36936,N_35139,N_35990);
and U36937 (N_36937,N_35072,N_34344);
and U36938 (N_36938,N_35456,N_34786);
nor U36939 (N_36939,N_34516,N_35674);
or U36940 (N_36940,N_35286,N_34434);
nor U36941 (N_36941,N_35808,N_35283);
xnor U36942 (N_36942,N_34864,N_34247);
or U36943 (N_36943,N_34593,N_35347);
or U36944 (N_36944,N_34802,N_34436);
nand U36945 (N_36945,N_34280,N_34266);
and U36946 (N_36946,N_34361,N_35693);
xnor U36947 (N_36947,N_34545,N_35625);
or U36948 (N_36948,N_35806,N_34769);
xor U36949 (N_36949,N_35067,N_35837);
xor U36950 (N_36950,N_34547,N_35909);
and U36951 (N_36951,N_34921,N_35940);
or U36952 (N_36952,N_34290,N_35222);
nand U36953 (N_36953,N_35174,N_34193);
nor U36954 (N_36954,N_34695,N_35883);
xor U36955 (N_36955,N_34734,N_34905);
nand U36956 (N_36956,N_35318,N_34163);
or U36957 (N_36957,N_35018,N_35148);
or U36958 (N_36958,N_34240,N_35435);
xor U36959 (N_36959,N_35575,N_35184);
nand U36960 (N_36960,N_34546,N_34842);
nand U36961 (N_36961,N_34707,N_35638);
and U36962 (N_36962,N_34686,N_34447);
or U36963 (N_36963,N_34120,N_35333);
or U36964 (N_36964,N_34652,N_34558);
nand U36965 (N_36965,N_34795,N_34774);
nand U36966 (N_36966,N_34762,N_35376);
nor U36967 (N_36967,N_35572,N_34649);
xor U36968 (N_36968,N_35408,N_35046);
xor U36969 (N_36969,N_35986,N_34282);
xnor U36970 (N_36970,N_35491,N_34928);
nor U36971 (N_36971,N_34568,N_35927);
nand U36972 (N_36972,N_34642,N_35065);
xnor U36973 (N_36973,N_34820,N_35201);
nand U36974 (N_36974,N_34430,N_35208);
and U36975 (N_36975,N_35130,N_34058);
xor U36976 (N_36976,N_34137,N_34276);
nor U36977 (N_36977,N_34023,N_34513);
and U36978 (N_36978,N_35751,N_34823);
and U36979 (N_36979,N_34849,N_35448);
or U36980 (N_36980,N_34272,N_35517);
nand U36981 (N_36981,N_34343,N_35968);
nor U36982 (N_36982,N_35217,N_35066);
or U36983 (N_36983,N_34765,N_35634);
xor U36984 (N_36984,N_34521,N_35984);
xnor U36985 (N_36985,N_35399,N_35460);
xnor U36986 (N_36986,N_34635,N_34724);
nor U36987 (N_36987,N_34341,N_35706);
nor U36988 (N_36988,N_34889,N_34146);
or U36989 (N_36989,N_34131,N_34506);
xnor U36990 (N_36990,N_35044,N_34462);
xnor U36991 (N_36991,N_35948,N_34005);
xnor U36992 (N_36992,N_35149,N_35891);
nor U36993 (N_36993,N_34906,N_35119);
nand U36994 (N_36994,N_35665,N_35125);
and U36995 (N_36995,N_34571,N_35269);
xnor U36996 (N_36996,N_34986,N_34072);
or U36997 (N_36997,N_34024,N_35757);
nand U36998 (N_36998,N_35221,N_34701);
nor U36999 (N_36999,N_34962,N_34085);
xnor U37000 (N_37000,N_35856,N_34750);
nor U37001 (N_37001,N_34514,N_35309);
or U37002 (N_37002,N_34408,N_34503);
nor U37003 (N_37003,N_35494,N_35864);
nand U37004 (N_37004,N_35841,N_35759);
and U37005 (N_37005,N_34035,N_35403);
xnor U37006 (N_37006,N_34993,N_35339);
nand U37007 (N_37007,N_34208,N_35884);
and U37008 (N_37008,N_35477,N_35917);
nor U37009 (N_37009,N_35809,N_35876);
and U37010 (N_37010,N_34082,N_34691);
nand U37011 (N_37011,N_35935,N_35148);
xor U37012 (N_37012,N_34339,N_34072);
nor U37013 (N_37013,N_34204,N_34108);
and U37014 (N_37014,N_35405,N_35681);
or U37015 (N_37015,N_34982,N_35944);
or U37016 (N_37016,N_34939,N_35720);
nand U37017 (N_37017,N_34865,N_35744);
nand U37018 (N_37018,N_34852,N_35263);
nand U37019 (N_37019,N_34854,N_34365);
nor U37020 (N_37020,N_35501,N_34490);
nor U37021 (N_37021,N_35701,N_34877);
nor U37022 (N_37022,N_35895,N_34068);
nand U37023 (N_37023,N_35309,N_35676);
nor U37024 (N_37024,N_35236,N_35274);
xor U37025 (N_37025,N_34645,N_34564);
and U37026 (N_37026,N_35961,N_34192);
nor U37027 (N_37027,N_34963,N_34575);
nand U37028 (N_37028,N_34048,N_35463);
xor U37029 (N_37029,N_34770,N_35629);
nand U37030 (N_37030,N_35802,N_34378);
xnor U37031 (N_37031,N_35574,N_35234);
nor U37032 (N_37032,N_34230,N_34889);
or U37033 (N_37033,N_35721,N_35348);
or U37034 (N_37034,N_35514,N_34082);
or U37035 (N_37035,N_35174,N_34028);
and U37036 (N_37036,N_35497,N_34864);
nand U37037 (N_37037,N_35752,N_35530);
or U37038 (N_37038,N_34744,N_35998);
xnor U37039 (N_37039,N_35802,N_34913);
and U37040 (N_37040,N_35907,N_35054);
nand U37041 (N_37041,N_35221,N_34070);
or U37042 (N_37042,N_35528,N_35455);
nand U37043 (N_37043,N_34703,N_34439);
nand U37044 (N_37044,N_34207,N_35884);
or U37045 (N_37045,N_35846,N_34088);
and U37046 (N_37046,N_35904,N_35243);
nor U37047 (N_37047,N_34646,N_35797);
and U37048 (N_37048,N_35926,N_34766);
xor U37049 (N_37049,N_35997,N_35713);
xor U37050 (N_37050,N_34718,N_34127);
nand U37051 (N_37051,N_34661,N_35708);
xnor U37052 (N_37052,N_35155,N_35630);
and U37053 (N_37053,N_35067,N_35491);
and U37054 (N_37054,N_34789,N_34799);
xor U37055 (N_37055,N_34942,N_35809);
xnor U37056 (N_37056,N_35843,N_34792);
and U37057 (N_37057,N_35475,N_35705);
nor U37058 (N_37058,N_34319,N_34282);
or U37059 (N_37059,N_35292,N_34245);
or U37060 (N_37060,N_34069,N_35212);
nor U37061 (N_37061,N_34831,N_34577);
nand U37062 (N_37062,N_34396,N_34102);
xnor U37063 (N_37063,N_34937,N_34169);
nand U37064 (N_37064,N_35976,N_35817);
nor U37065 (N_37065,N_34770,N_35281);
xor U37066 (N_37066,N_35738,N_34289);
and U37067 (N_37067,N_34719,N_35666);
nand U37068 (N_37068,N_34336,N_34785);
nor U37069 (N_37069,N_35346,N_34251);
nand U37070 (N_37070,N_34579,N_35931);
or U37071 (N_37071,N_34928,N_34125);
nor U37072 (N_37072,N_35809,N_34298);
or U37073 (N_37073,N_34319,N_34234);
xor U37074 (N_37074,N_35710,N_34595);
xor U37075 (N_37075,N_34463,N_35764);
nand U37076 (N_37076,N_34033,N_34452);
xnor U37077 (N_37077,N_34831,N_35648);
nand U37078 (N_37078,N_35800,N_34672);
xnor U37079 (N_37079,N_34530,N_35335);
nor U37080 (N_37080,N_34698,N_35810);
or U37081 (N_37081,N_35636,N_34733);
nand U37082 (N_37082,N_35479,N_35134);
nor U37083 (N_37083,N_35372,N_34778);
nand U37084 (N_37084,N_34784,N_35785);
or U37085 (N_37085,N_35081,N_34527);
and U37086 (N_37086,N_35836,N_35185);
xor U37087 (N_37087,N_35098,N_35722);
xor U37088 (N_37088,N_35428,N_34873);
nor U37089 (N_37089,N_34186,N_34454);
or U37090 (N_37090,N_34041,N_35689);
or U37091 (N_37091,N_35628,N_35648);
or U37092 (N_37092,N_35208,N_35387);
nand U37093 (N_37093,N_35890,N_34799);
or U37094 (N_37094,N_34446,N_35913);
nand U37095 (N_37095,N_35664,N_35765);
nand U37096 (N_37096,N_35838,N_35121);
xnor U37097 (N_37097,N_35613,N_34794);
nor U37098 (N_37098,N_34081,N_35972);
xor U37099 (N_37099,N_34585,N_35479);
and U37100 (N_37100,N_34218,N_35705);
nand U37101 (N_37101,N_35940,N_34838);
xnor U37102 (N_37102,N_34068,N_35749);
or U37103 (N_37103,N_34463,N_35234);
and U37104 (N_37104,N_35452,N_34851);
and U37105 (N_37105,N_34821,N_35030);
nand U37106 (N_37106,N_35924,N_35634);
nand U37107 (N_37107,N_35517,N_34700);
nand U37108 (N_37108,N_35050,N_34981);
nand U37109 (N_37109,N_34816,N_35207);
xor U37110 (N_37110,N_34247,N_34197);
and U37111 (N_37111,N_35837,N_35493);
nor U37112 (N_37112,N_35816,N_34001);
and U37113 (N_37113,N_35711,N_35351);
and U37114 (N_37114,N_34634,N_35237);
or U37115 (N_37115,N_35159,N_35646);
or U37116 (N_37116,N_34160,N_35406);
nand U37117 (N_37117,N_34241,N_34032);
nand U37118 (N_37118,N_34410,N_35800);
nor U37119 (N_37119,N_35407,N_35034);
or U37120 (N_37120,N_34872,N_34735);
nor U37121 (N_37121,N_35754,N_35532);
nand U37122 (N_37122,N_34855,N_35534);
or U37123 (N_37123,N_35002,N_35488);
and U37124 (N_37124,N_34020,N_34338);
nand U37125 (N_37125,N_34919,N_35608);
or U37126 (N_37126,N_35756,N_34091);
nand U37127 (N_37127,N_35418,N_34214);
nor U37128 (N_37128,N_35305,N_34387);
nor U37129 (N_37129,N_35932,N_34044);
and U37130 (N_37130,N_35130,N_34467);
xnor U37131 (N_37131,N_35261,N_35902);
xnor U37132 (N_37132,N_35246,N_34230);
nand U37133 (N_37133,N_35923,N_35702);
nand U37134 (N_37134,N_34745,N_34626);
xor U37135 (N_37135,N_35922,N_34939);
nor U37136 (N_37136,N_34710,N_35610);
or U37137 (N_37137,N_34937,N_34186);
and U37138 (N_37138,N_34528,N_35441);
nand U37139 (N_37139,N_34459,N_35982);
nand U37140 (N_37140,N_35528,N_34509);
xor U37141 (N_37141,N_34501,N_35744);
and U37142 (N_37142,N_35571,N_34081);
xnor U37143 (N_37143,N_34055,N_35717);
xor U37144 (N_37144,N_35982,N_35691);
or U37145 (N_37145,N_34083,N_34765);
xor U37146 (N_37146,N_35565,N_34145);
nand U37147 (N_37147,N_35766,N_34246);
or U37148 (N_37148,N_35986,N_34754);
and U37149 (N_37149,N_35182,N_34903);
xnor U37150 (N_37150,N_35617,N_34770);
and U37151 (N_37151,N_34051,N_34229);
nor U37152 (N_37152,N_35008,N_35237);
and U37153 (N_37153,N_35232,N_34856);
xnor U37154 (N_37154,N_35116,N_35942);
or U37155 (N_37155,N_35955,N_35349);
nand U37156 (N_37156,N_35269,N_34447);
or U37157 (N_37157,N_34009,N_35146);
nor U37158 (N_37158,N_35003,N_35254);
and U37159 (N_37159,N_34020,N_34872);
or U37160 (N_37160,N_35665,N_34501);
or U37161 (N_37161,N_34122,N_35407);
nand U37162 (N_37162,N_35131,N_35876);
xnor U37163 (N_37163,N_35312,N_34425);
nor U37164 (N_37164,N_35441,N_34007);
xnor U37165 (N_37165,N_34201,N_34455);
or U37166 (N_37166,N_34813,N_34132);
xnor U37167 (N_37167,N_35516,N_35294);
and U37168 (N_37168,N_35672,N_35294);
or U37169 (N_37169,N_35764,N_34789);
xor U37170 (N_37170,N_34497,N_35403);
nor U37171 (N_37171,N_34052,N_35407);
and U37172 (N_37172,N_35851,N_35728);
nor U37173 (N_37173,N_35505,N_35555);
nor U37174 (N_37174,N_35560,N_35861);
or U37175 (N_37175,N_35711,N_34974);
xor U37176 (N_37176,N_35561,N_34964);
or U37177 (N_37177,N_34498,N_34527);
xnor U37178 (N_37178,N_34190,N_34061);
or U37179 (N_37179,N_34893,N_35508);
nand U37180 (N_37180,N_35253,N_35838);
or U37181 (N_37181,N_34128,N_35949);
nor U37182 (N_37182,N_34950,N_35967);
and U37183 (N_37183,N_34826,N_35462);
and U37184 (N_37184,N_35635,N_35118);
nand U37185 (N_37185,N_34576,N_34196);
or U37186 (N_37186,N_35387,N_34729);
xnor U37187 (N_37187,N_35011,N_34732);
nor U37188 (N_37188,N_35492,N_34601);
nor U37189 (N_37189,N_34057,N_34182);
xor U37190 (N_37190,N_35772,N_34954);
and U37191 (N_37191,N_35679,N_35452);
and U37192 (N_37192,N_34768,N_35316);
nand U37193 (N_37193,N_34752,N_34149);
nand U37194 (N_37194,N_34246,N_35500);
or U37195 (N_37195,N_34370,N_34941);
nor U37196 (N_37196,N_35914,N_35124);
xnor U37197 (N_37197,N_35060,N_34895);
and U37198 (N_37198,N_35764,N_35163);
or U37199 (N_37199,N_35525,N_34320);
nor U37200 (N_37200,N_35122,N_34228);
xnor U37201 (N_37201,N_34096,N_34777);
nor U37202 (N_37202,N_35411,N_35905);
and U37203 (N_37203,N_35713,N_35319);
nand U37204 (N_37204,N_34007,N_34651);
nor U37205 (N_37205,N_35089,N_35160);
and U37206 (N_37206,N_34254,N_34379);
nand U37207 (N_37207,N_35426,N_35364);
or U37208 (N_37208,N_34591,N_34999);
and U37209 (N_37209,N_35512,N_35797);
nor U37210 (N_37210,N_35144,N_35097);
and U37211 (N_37211,N_34162,N_35478);
and U37212 (N_37212,N_35862,N_35071);
nor U37213 (N_37213,N_35274,N_34677);
or U37214 (N_37214,N_34693,N_35200);
nand U37215 (N_37215,N_35216,N_35610);
and U37216 (N_37216,N_35143,N_35930);
nor U37217 (N_37217,N_35563,N_35588);
and U37218 (N_37218,N_34559,N_35527);
nand U37219 (N_37219,N_34796,N_34418);
or U37220 (N_37220,N_35868,N_34256);
and U37221 (N_37221,N_34290,N_35011);
nor U37222 (N_37222,N_34604,N_35251);
nor U37223 (N_37223,N_35463,N_35210);
and U37224 (N_37224,N_34145,N_35410);
nor U37225 (N_37225,N_34361,N_35078);
xnor U37226 (N_37226,N_34350,N_35502);
nand U37227 (N_37227,N_34529,N_34260);
or U37228 (N_37228,N_35642,N_35055);
nand U37229 (N_37229,N_34444,N_35879);
nand U37230 (N_37230,N_35771,N_34204);
and U37231 (N_37231,N_34786,N_34265);
nand U37232 (N_37232,N_34391,N_34816);
nand U37233 (N_37233,N_34602,N_34228);
nor U37234 (N_37234,N_35582,N_34011);
xnor U37235 (N_37235,N_34735,N_34458);
nor U37236 (N_37236,N_35172,N_35611);
and U37237 (N_37237,N_35927,N_35749);
and U37238 (N_37238,N_34253,N_35982);
and U37239 (N_37239,N_35842,N_35521);
xor U37240 (N_37240,N_35938,N_34333);
nor U37241 (N_37241,N_34190,N_35013);
nand U37242 (N_37242,N_34407,N_34949);
nor U37243 (N_37243,N_35650,N_34621);
nand U37244 (N_37244,N_34127,N_34751);
nand U37245 (N_37245,N_35834,N_35154);
or U37246 (N_37246,N_34113,N_34923);
or U37247 (N_37247,N_35649,N_35258);
or U37248 (N_37248,N_35567,N_35135);
nand U37249 (N_37249,N_34441,N_34572);
nor U37250 (N_37250,N_34638,N_35073);
and U37251 (N_37251,N_34978,N_35003);
or U37252 (N_37252,N_34193,N_35080);
or U37253 (N_37253,N_35138,N_35317);
or U37254 (N_37254,N_34386,N_35168);
nor U37255 (N_37255,N_34781,N_34003);
and U37256 (N_37256,N_34066,N_35762);
xnor U37257 (N_37257,N_35015,N_35755);
xnor U37258 (N_37258,N_34091,N_35436);
or U37259 (N_37259,N_35005,N_35884);
nor U37260 (N_37260,N_34775,N_35542);
nand U37261 (N_37261,N_34954,N_35398);
or U37262 (N_37262,N_35794,N_35730);
or U37263 (N_37263,N_34678,N_35690);
and U37264 (N_37264,N_34471,N_34777);
xor U37265 (N_37265,N_34660,N_34174);
and U37266 (N_37266,N_35243,N_34303);
and U37267 (N_37267,N_34246,N_34382);
nor U37268 (N_37268,N_34573,N_35938);
nand U37269 (N_37269,N_34538,N_35485);
and U37270 (N_37270,N_34580,N_34846);
nor U37271 (N_37271,N_35746,N_34102);
and U37272 (N_37272,N_35426,N_35766);
or U37273 (N_37273,N_34154,N_34836);
xnor U37274 (N_37274,N_34040,N_34407);
or U37275 (N_37275,N_35435,N_34443);
xnor U37276 (N_37276,N_34149,N_35029);
and U37277 (N_37277,N_34478,N_34450);
nor U37278 (N_37278,N_34997,N_35270);
or U37279 (N_37279,N_34918,N_34778);
nor U37280 (N_37280,N_35697,N_35341);
and U37281 (N_37281,N_34480,N_35479);
and U37282 (N_37282,N_35228,N_34669);
or U37283 (N_37283,N_34732,N_34302);
nand U37284 (N_37284,N_34880,N_35868);
and U37285 (N_37285,N_34638,N_35256);
nand U37286 (N_37286,N_34934,N_35329);
and U37287 (N_37287,N_35543,N_35772);
nand U37288 (N_37288,N_35663,N_34572);
xnor U37289 (N_37289,N_35844,N_34016);
nand U37290 (N_37290,N_34126,N_35988);
and U37291 (N_37291,N_35696,N_35968);
or U37292 (N_37292,N_34061,N_35984);
nand U37293 (N_37293,N_35485,N_35385);
or U37294 (N_37294,N_35887,N_35756);
nor U37295 (N_37295,N_35663,N_35701);
and U37296 (N_37296,N_35218,N_34022);
and U37297 (N_37297,N_35495,N_35635);
or U37298 (N_37298,N_35307,N_34464);
nor U37299 (N_37299,N_34699,N_34505);
xor U37300 (N_37300,N_34172,N_35532);
xor U37301 (N_37301,N_35709,N_34251);
nor U37302 (N_37302,N_35007,N_35164);
nand U37303 (N_37303,N_35293,N_35361);
or U37304 (N_37304,N_34139,N_34303);
nor U37305 (N_37305,N_35415,N_35188);
xnor U37306 (N_37306,N_35958,N_34648);
or U37307 (N_37307,N_34649,N_35321);
nand U37308 (N_37308,N_35659,N_34910);
and U37309 (N_37309,N_34669,N_35524);
nor U37310 (N_37310,N_34956,N_34350);
nor U37311 (N_37311,N_35665,N_34472);
or U37312 (N_37312,N_35367,N_34115);
nand U37313 (N_37313,N_34507,N_34606);
nor U37314 (N_37314,N_34191,N_34202);
and U37315 (N_37315,N_35617,N_34201);
and U37316 (N_37316,N_35597,N_35536);
xor U37317 (N_37317,N_35387,N_34320);
xor U37318 (N_37318,N_35558,N_34770);
nor U37319 (N_37319,N_35265,N_35585);
or U37320 (N_37320,N_34293,N_35906);
nor U37321 (N_37321,N_35088,N_34098);
xnor U37322 (N_37322,N_34471,N_35886);
xor U37323 (N_37323,N_35907,N_34326);
and U37324 (N_37324,N_34645,N_34225);
xnor U37325 (N_37325,N_34385,N_34959);
or U37326 (N_37326,N_35591,N_34275);
or U37327 (N_37327,N_34126,N_34617);
xor U37328 (N_37328,N_34393,N_34697);
nor U37329 (N_37329,N_35559,N_35472);
nor U37330 (N_37330,N_34824,N_35173);
nor U37331 (N_37331,N_34486,N_35940);
or U37332 (N_37332,N_34070,N_35194);
or U37333 (N_37333,N_34443,N_34570);
and U37334 (N_37334,N_34632,N_34024);
xor U37335 (N_37335,N_35316,N_35468);
nand U37336 (N_37336,N_34879,N_35400);
or U37337 (N_37337,N_34178,N_35575);
or U37338 (N_37338,N_34742,N_35604);
and U37339 (N_37339,N_35761,N_35577);
nand U37340 (N_37340,N_35202,N_34924);
nand U37341 (N_37341,N_35224,N_34932);
and U37342 (N_37342,N_34093,N_34330);
and U37343 (N_37343,N_34950,N_35147);
nor U37344 (N_37344,N_35964,N_34141);
nand U37345 (N_37345,N_34371,N_35225);
nand U37346 (N_37346,N_34905,N_34521);
or U37347 (N_37347,N_35501,N_35932);
nand U37348 (N_37348,N_35521,N_35009);
nor U37349 (N_37349,N_34947,N_35428);
xor U37350 (N_37350,N_34121,N_34496);
nand U37351 (N_37351,N_34788,N_34068);
nand U37352 (N_37352,N_35620,N_34074);
or U37353 (N_37353,N_35249,N_35264);
or U37354 (N_37354,N_35316,N_34699);
or U37355 (N_37355,N_35669,N_35182);
and U37356 (N_37356,N_34504,N_34777);
xor U37357 (N_37357,N_34423,N_35061);
nand U37358 (N_37358,N_34547,N_34697);
nand U37359 (N_37359,N_35691,N_35767);
nor U37360 (N_37360,N_34594,N_35762);
nor U37361 (N_37361,N_34313,N_34372);
xnor U37362 (N_37362,N_34554,N_34608);
and U37363 (N_37363,N_35805,N_34247);
and U37364 (N_37364,N_35356,N_34058);
or U37365 (N_37365,N_35145,N_34226);
nand U37366 (N_37366,N_35256,N_34941);
and U37367 (N_37367,N_34769,N_34139);
xor U37368 (N_37368,N_34543,N_34782);
nand U37369 (N_37369,N_35142,N_35347);
nand U37370 (N_37370,N_34977,N_34474);
nand U37371 (N_37371,N_34662,N_34204);
nor U37372 (N_37372,N_35926,N_35762);
nor U37373 (N_37373,N_35229,N_35751);
nor U37374 (N_37374,N_34917,N_35888);
xor U37375 (N_37375,N_35494,N_34697);
nand U37376 (N_37376,N_34225,N_35249);
nor U37377 (N_37377,N_34639,N_35789);
nand U37378 (N_37378,N_34542,N_35450);
nand U37379 (N_37379,N_35364,N_35010);
xnor U37380 (N_37380,N_34950,N_35299);
xnor U37381 (N_37381,N_35238,N_35148);
and U37382 (N_37382,N_35502,N_35874);
nand U37383 (N_37383,N_34284,N_35380);
nor U37384 (N_37384,N_34645,N_35151);
nor U37385 (N_37385,N_34081,N_35959);
nand U37386 (N_37386,N_35636,N_34370);
nor U37387 (N_37387,N_35010,N_34869);
or U37388 (N_37388,N_34467,N_34299);
or U37389 (N_37389,N_35986,N_34796);
or U37390 (N_37390,N_35286,N_34476);
or U37391 (N_37391,N_34850,N_35309);
or U37392 (N_37392,N_34427,N_34044);
and U37393 (N_37393,N_35451,N_34170);
or U37394 (N_37394,N_35269,N_35225);
xnor U37395 (N_37395,N_34262,N_35793);
or U37396 (N_37396,N_35552,N_35332);
nand U37397 (N_37397,N_35511,N_34809);
or U37398 (N_37398,N_35204,N_35540);
xnor U37399 (N_37399,N_34648,N_34343);
nand U37400 (N_37400,N_34832,N_34122);
and U37401 (N_37401,N_35728,N_35253);
nand U37402 (N_37402,N_35382,N_35131);
nor U37403 (N_37403,N_34238,N_34159);
nor U37404 (N_37404,N_34595,N_34122);
or U37405 (N_37405,N_35511,N_34857);
and U37406 (N_37406,N_34360,N_35498);
or U37407 (N_37407,N_34365,N_35719);
or U37408 (N_37408,N_34475,N_34009);
and U37409 (N_37409,N_34652,N_34785);
nand U37410 (N_37410,N_35341,N_35899);
nor U37411 (N_37411,N_35218,N_34842);
nand U37412 (N_37412,N_35006,N_35691);
and U37413 (N_37413,N_35487,N_34895);
nor U37414 (N_37414,N_34238,N_34198);
and U37415 (N_37415,N_35688,N_35840);
nand U37416 (N_37416,N_34847,N_34789);
nand U37417 (N_37417,N_35905,N_35111);
xor U37418 (N_37418,N_34617,N_35080);
nand U37419 (N_37419,N_35232,N_34948);
xor U37420 (N_37420,N_35234,N_34648);
or U37421 (N_37421,N_35012,N_34474);
nor U37422 (N_37422,N_35226,N_35457);
nor U37423 (N_37423,N_34088,N_35806);
or U37424 (N_37424,N_35929,N_35057);
nor U37425 (N_37425,N_35552,N_35132);
nand U37426 (N_37426,N_35200,N_34717);
nand U37427 (N_37427,N_35307,N_35493);
nor U37428 (N_37428,N_35388,N_34657);
nand U37429 (N_37429,N_34817,N_34307);
xnor U37430 (N_37430,N_34828,N_35388);
or U37431 (N_37431,N_35825,N_35141);
and U37432 (N_37432,N_34000,N_35220);
nor U37433 (N_37433,N_34702,N_34160);
nand U37434 (N_37434,N_35268,N_34504);
nor U37435 (N_37435,N_34733,N_34160);
xor U37436 (N_37436,N_34817,N_35745);
xnor U37437 (N_37437,N_34250,N_34416);
nor U37438 (N_37438,N_34808,N_35393);
and U37439 (N_37439,N_35707,N_35082);
nand U37440 (N_37440,N_34754,N_34908);
or U37441 (N_37441,N_35842,N_34185);
and U37442 (N_37442,N_34836,N_34899);
xor U37443 (N_37443,N_35090,N_34220);
nand U37444 (N_37444,N_34388,N_34650);
or U37445 (N_37445,N_35683,N_34284);
xnor U37446 (N_37446,N_34618,N_35590);
and U37447 (N_37447,N_34513,N_35528);
xnor U37448 (N_37448,N_35116,N_34312);
or U37449 (N_37449,N_34599,N_35906);
nand U37450 (N_37450,N_35358,N_34907);
nand U37451 (N_37451,N_34372,N_35727);
nand U37452 (N_37452,N_34598,N_34465);
or U37453 (N_37453,N_34072,N_35039);
nand U37454 (N_37454,N_34878,N_35066);
nand U37455 (N_37455,N_34815,N_34043);
nor U37456 (N_37456,N_34267,N_34198);
and U37457 (N_37457,N_34711,N_34094);
nand U37458 (N_37458,N_35638,N_34701);
xnor U37459 (N_37459,N_34150,N_34392);
nand U37460 (N_37460,N_34602,N_34903);
and U37461 (N_37461,N_35357,N_34115);
or U37462 (N_37462,N_34174,N_35755);
and U37463 (N_37463,N_34419,N_35787);
or U37464 (N_37464,N_35094,N_34164);
or U37465 (N_37465,N_35582,N_35108);
and U37466 (N_37466,N_35778,N_35908);
nor U37467 (N_37467,N_34538,N_35099);
xnor U37468 (N_37468,N_34755,N_34550);
nand U37469 (N_37469,N_35503,N_35095);
or U37470 (N_37470,N_35928,N_34475);
or U37471 (N_37471,N_35879,N_35781);
nand U37472 (N_37472,N_34221,N_34918);
nor U37473 (N_37473,N_34842,N_35529);
nor U37474 (N_37474,N_35936,N_35891);
and U37475 (N_37475,N_34589,N_35387);
xor U37476 (N_37476,N_34637,N_34989);
nor U37477 (N_37477,N_35886,N_35725);
and U37478 (N_37478,N_34851,N_35956);
nor U37479 (N_37479,N_34897,N_35360);
nor U37480 (N_37480,N_35222,N_35162);
xor U37481 (N_37481,N_34436,N_34906);
xor U37482 (N_37482,N_35958,N_34236);
and U37483 (N_37483,N_35193,N_35602);
xor U37484 (N_37484,N_34138,N_35015);
or U37485 (N_37485,N_34846,N_34129);
or U37486 (N_37486,N_34208,N_34833);
or U37487 (N_37487,N_34442,N_34063);
xor U37488 (N_37488,N_34406,N_35346);
or U37489 (N_37489,N_35887,N_35730);
xnor U37490 (N_37490,N_35088,N_35897);
or U37491 (N_37491,N_34945,N_34188);
and U37492 (N_37492,N_35246,N_34179);
xnor U37493 (N_37493,N_34450,N_34775);
nand U37494 (N_37494,N_35411,N_35477);
or U37495 (N_37495,N_35206,N_34083);
or U37496 (N_37496,N_34452,N_34515);
or U37497 (N_37497,N_34598,N_34922);
and U37498 (N_37498,N_35340,N_35490);
or U37499 (N_37499,N_35293,N_35714);
nand U37500 (N_37500,N_34021,N_34351);
xnor U37501 (N_37501,N_34251,N_34824);
nor U37502 (N_37502,N_35406,N_34502);
nor U37503 (N_37503,N_34748,N_35527);
nor U37504 (N_37504,N_35406,N_34738);
xnor U37505 (N_37505,N_35729,N_35929);
nand U37506 (N_37506,N_34060,N_34673);
nand U37507 (N_37507,N_34735,N_35032);
and U37508 (N_37508,N_34718,N_35081);
nor U37509 (N_37509,N_35514,N_34921);
or U37510 (N_37510,N_34516,N_35454);
nand U37511 (N_37511,N_35195,N_34302);
nand U37512 (N_37512,N_35438,N_35021);
xnor U37513 (N_37513,N_34883,N_35645);
xnor U37514 (N_37514,N_34993,N_35859);
xnor U37515 (N_37515,N_34767,N_34812);
nor U37516 (N_37516,N_34634,N_34137);
nor U37517 (N_37517,N_34239,N_35916);
nor U37518 (N_37518,N_34962,N_34944);
nand U37519 (N_37519,N_35601,N_35971);
and U37520 (N_37520,N_35225,N_35709);
and U37521 (N_37521,N_35689,N_35428);
or U37522 (N_37522,N_35435,N_34436);
nor U37523 (N_37523,N_34918,N_34123);
nor U37524 (N_37524,N_34494,N_35608);
nand U37525 (N_37525,N_35399,N_34711);
and U37526 (N_37526,N_35191,N_35543);
nand U37527 (N_37527,N_35337,N_35622);
xnor U37528 (N_37528,N_34938,N_35117);
nand U37529 (N_37529,N_34607,N_35605);
nor U37530 (N_37530,N_34275,N_34845);
or U37531 (N_37531,N_35063,N_35720);
or U37532 (N_37532,N_34636,N_35348);
nand U37533 (N_37533,N_35446,N_35351);
nand U37534 (N_37534,N_34182,N_34204);
or U37535 (N_37535,N_35902,N_35864);
nand U37536 (N_37536,N_34621,N_35307);
and U37537 (N_37537,N_35383,N_34064);
xor U37538 (N_37538,N_35532,N_35973);
and U37539 (N_37539,N_34028,N_35572);
nor U37540 (N_37540,N_35785,N_34956);
xor U37541 (N_37541,N_35987,N_34164);
xor U37542 (N_37542,N_35706,N_35681);
or U37543 (N_37543,N_34826,N_34594);
and U37544 (N_37544,N_35272,N_34952);
or U37545 (N_37545,N_34173,N_35792);
nand U37546 (N_37546,N_34012,N_34757);
nor U37547 (N_37547,N_35321,N_35633);
nand U37548 (N_37548,N_34944,N_35327);
or U37549 (N_37549,N_35302,N_35630);
or U37550 (N_37550,N_35732,N_35749);
and U37551 (N_37551,N_34908,N_35037);
or U37552 (N_37552,N_35327,N_35800);
nand U37553 (N_37553,N_34280,N_35703);
nand U37554 (N_37554,N_34488,N_34415);
nor U37555 (N_37555,N_35352,N_34304);
nor U37556 (N_37556,N_35360,N_35289);
nand U37557 (N_37557,N_34876,N_35007);
and U37558 (N_37558,N_34715,N_35818);
or U37559 (N_37559,N_35371,N_35144);
xor U37560 (N_37560,N_35961,N_34369);
nand U37561 (N_37561,N_34383,N_34907);
nand U37562 (N_37562,N_34098,N_35508);
nand U37563 (N_37563,N_35625,N_35445);
xnor U37564 (N_37564,N_35697,N_34177);
or U37565 (N_37565,N_34782,N_35661);
and U37566 (N_37566,N_34124,N_34277);
or U37567 (N_37567,N_35697,N_35534);
or U37568 (N_37568,N_34230,N_35856);
nand U37569 (N_37569,N_34719,N_35941);
nand U37570 (N_37570,N_34126,N_35300);
xor U37571 (N_37571,N_35802,N_35284);
nor U37572 (N_37572,N_34137,N_35749);
and U37573 (N_37573,N_34837,N_35615);
and U37574 (N_37574,N_35569,N_35425);
and U37575 (N_37575,N_34526,N_35886);
nand U37576 (N_37576,N_34983,N_34495);
or U37577 (N_37577,N_35956,N_34569);
nand U37578 (N_37578,N_35065,N_35693);
xor U37579 (N_37579,N_35887,N_35556);
nor U37580 (N_37580,N_34913,N_34002);
nand U37581 (N_37581,N_34141,N_35327);
and U37582 (N_37582,N_35251,N_34548);
xor U37583 (N_37583,N_35502,N_34706);
and U37584 (N_37584,N_34371,N_35406);
or U37585 (N_37585,N_34895,N_34391);
or U37586 (N_37586,N_35945,N_34588);
xor U37587 (N_37587,N_34612,N_35215);
nand U37588 (N_37588,N_34142,N_34725);
or U37589 (N_37589,N_35401,N_35317);
and U37590 (N_37590,N_35868,N_35585);
nor U37591 (N_37591,N_34745,N_34825);
nand U37592 (N_37592,N_35394,N_35813);
nor U37593 (N_37593,N_35672,N_35040);
or U37594 (N_37594,N_34728,N_35036);
nand U37595 (N_37595,N_35063,N_35745);
and U37596 (N_37596,N_34459,N_34789);
nor U37597 (N_37597,N_34913,N_35757);
and U37598 (N_37598,N_34436,N_34559);
or U37599 (N_37599,N_35669,N_35549);
xor U37600 (N_37600,N_34566,N_35193);
and U37601 (N_37601,N_35342,N_35444);
nor U37602 (N_37602,N_35111,N_35323);
or U37603 (N_37603,N_34107,N_34509);
or U37604 (N_37604,N_34791,N_34381);
nand U37605 (N_37605,N_35649,N_35244);
and U37606 (N_37606,N_35092,N_35536);
or U37607 (N_37607,N_34845,N_35065);
or U37608 (N_37608,N_35799,N_35311);
nor U37609 (N_37609,N_34406,N_35500);
and U37610 (N_37610,N_35141,N_35268);
and U37611 (N_37611,N_34091,N_35149);
or U37612 (N_37612,N_34792,N_34821);
nor U37613 (N_37613,N_35507,N_35876);
nor U37614 (N_37614,N_35054,N_35391);
xor U37615 (N_37615,N_34398,N_35270);
xor U37616 (N_37616,N_35510,N_35116);
or U37617 (N_37617,N_34878,N_35026);
nor U37618 (N_37618,N_35087,N_35245);
and U37619 (N_37619,N_35121,N_35248);
nand U37620 (N_37620,N_35714,N_34332);
nand U37621 (N_37621,N_34223,N_35336);
nor U37622 (N_37622,N_35858,N_35826);
xnor U37623 (N_37623,N_35911,N_34579);
nand U37624 (N_37624,N_35830,N_34855);
and U37625 (N_37625,N_34987,N_35494);
nor U37626 (N_37626,N_34762,N_34740);
or U37627 (N_37627,N_34230,N_35870);
xnor U37628 (N_37628,N_35137,N_35492);
nand U37629 (N_37629,N_35062,N_35003);
xnor U37630 (N_37630,N_34862,N_35431);
xnor U37631 (N_37631,N_34195,N_34498);
or U37632 (N_37632,N_34669,N_34297);
and U37633 (N_37633,N_35183,N_35022);
and U37634 (N_37634,N_34278,N_35600);
nor U37635 (N_37635,N_35478,N_35769);
nand U37636 (N_37636,N_35436,N_34579);
nand U37637 (N_37637,N_35294,N_35903);
nand U37638 (N_37638,N_34554,N_35663);
or U37639 (N_37639,N_35544,N_35923);
nand U37640 (N_37640,N_35019,N_35397);
nand U37641 (N_37641,N_34254,N_35431);
nor U37642 (N_37642,N_34039,N_35585);
nor U37643 (N_37643,N_35232,N_35419);
or U37644 (N_37644,N_34753,N_34966);
or U37645 (N_37645,N_34965,N_35654);
or U37646 (N_37646,N_34296,N_34164);
xor U37647 (N_37647,N_34702,N_35456);
and U37648 (N_37648,N_35352,N_35750);
nand U37649 (N_37649,N_34844,N_35557);
nand U37650 (N_37650,N_34257,N_34504);
and U37651 (N_37651,N_35075,N_35582);
nor U37652 (N_37652,N_34784,N_35519);
or U37653 (N_37653,N_34013,N_34465);
nand U37654 (N_37654,N_34304,N_35501);
and U37655 (N_37655,N_35377,N_35700);
nor U37656 (N_37656,N_35765,N_34824);
nand U37657 (N_37657,N_34815,N_35584);
or U37658 (N_37658,N_35379,N_34502);
and U37659 (N_37659,N_35279,N_34205);
nand U37660 (N_37660,N_35548,N_35046);
and U37661 (N_37661,N_34013,N_34826);
and U37662 (N_37662,N_35263,N_34043);
xor U37663 (N_37663,N_34316,N_35243);
and U37664 (N_37664,N_35154,N_35502);
or U37665 (N_37665,N_34662,N_35933);
and U37666 (N_37666,N_34724,N_35763);
nor U37667 (N_37667,N_35223,N_34091);
or U37668 (N_37668,N_35226,N_34018);
nand U37669 (N_37669,N_35009,N_35480);
or U37670 (N_37670,N_35034,N_35661);
xnor U37671 (N_37671,N_34572,N_34077);
xnor U37672 (N_37672,N_34036,N_35648);
xor U37673 (N_37673,N_34007,N_35343);
xnor U37674 (N_37674,N_35553,N_35617);
xor U37675 (N_37675,N_35815,N_34290);
nor U37676 (N_37676,N_34117,N_35395);
nor U37677 (N_37677,N_35708,N_34918);
xor U37678 (N_37678,N_35942,N_35266);
nand U37679 (N_37679,N_34736,N_34028);
xor U37680 (N_37680,N_35438,N_35630);
and U37681 (N_37681,N_35771,N_35055);
and U37682 (N_37682,N_35096,N_35203);
xnor U37683 (N_37683,N_35789,N_34174);
nor U37684 (N_37684,N_34198,N_34350);
nor U37685 (N_37685,N_35972,N_34358);
and U37686 (N_37686,N_35952,N_35776);
nand U37687 (N_37687,N_34483,N_35611);
nand U37688 (N_37688,N_35488,N_34544);
nor U37689 (N_37689,N_35139,N_35163);
or U37690 (N_37690,N_35655,N_34277);
xor U37691 (N_37691,N_34276,N_34906);
nor U37692 (N_37692,N_35551,N_35802);
xnor U37693 (N_37693,N_35085,N_34381);
nand U37694 (N_37694,N_35690,N_35815);
and U37695 (N_37695,N_34382,N_34150);
xor U37696 (N_37696,N_34901,N_34110);
and U37697 (N_37697,N_35693,N_34765);
nand U37698 (N_37698,N_35444,N_35956);
xor U37699 (N_37699,N_34639,N_35868);
and U37700 (N_37700,N_34481,N_34842);
xnor U37701 (N_37701,N_35575,N_34190);
xnor U37702 (N_37702,N_34265,N_34920);
nor U37703 (N_37703,N_34662,N_34925);
and U37704 (N_37704,N_34457,N_35523);
or U37705 (N_37705,N_35632,N_35355);
xor U37706 (N_37706,N_34139,N_35293);
nor U37707 (N_37707,N_34664,N_35343);
xor U37708 (N_37708,N_34777,N_35363);
or U37709 (N_37709,N_34499,N_34335);
xor U37710 (N_37710,N_35635,N_34758);
nor U37711 (N_37711,N_34191,N_35694);
nand U37712 (N_37712,N_35018,N_34427);
nand U37713 (N_37713,N_35700,N_35055);
nor U37714 (N_37714,N_34740,N_35001);
or U37715 (N_37715,N_34740,N_35656);
and U37716 (N_37716,N_34389,N_35388);
or U37717 (N_37717,N_34093,N_34274);
xor U37718 (N_37718,N_34924,N_35058);
and U37719 (N_37719,N_35229,N_34053);
nor U37720 (N_37720,N_34259,N_34552);
nor U37721 (N_37721,N_35779,N_34671);
nor U37722 (N_37722,N_34732,N_35443);
nor U37723 (N_37723,N_35170,N_34662);
xnor U37724 (N_37724,N_34188,N_34302);
or U37725 (N_37725,N_34594,N_35842);
or U37726 (N_37726,N_35800,N_35948);
xor U37727 (N_37727,N_35600,N_34202);
xnor U37728 (N_37728,N_34887,N_34390);
xor U37729 (N_37729,N_34868,N_35507);
or U37730 (N_37730,N_35043,N_35478);
nor U37731 (N_37731,N_34355,N_34545);
or U37732 (N_37732,N_34955,N_34306);
nand U37733 (N_37733,N_34460,N_35732);
and U37734 (N_37734,N_35337,N_34525);
xnor U37735 (N_37735,N_35304,N_35233);
or U37736 (N_37736,N_34690,N_35234);
nand U37737 (N_37737,N_35401,N_34360);
or U37738 (N_37738,N_34926,N_35367);
nand U37739 (N_37739,N_34713,N_35723);
and U37740 (N_37740,N_35517,N_35611);
nor U37741 (N_37741,N_34928,N_35197);
nor U37742 (N_37742,N_35370,N_34941);
nor U37743 (N_37743,N_35168,N_35180);
or U37744 (N_37744,N_34016,N_34464);
xor U37745 (N_37745,N_35753,N_34541);
xor U37746 (N_37746,N_35519,N_34790);
or U37747 (N_37747,N_34056,N_34175);
or U37748 (N_37748,N_34191,N_34851);
xnor U37749 (N_37749,N_35696,N_35258);
nand U37750 (N_37750,N_34039,N_35954);
nor U37751 (N_37751,N_34087,N_34109);
nor U37752 (N_37752,N_34745,N_35729);
xor U37753 (N_37753,N_34630,N_35150);
xor U37754 (N_37754,N_35049,N_35533);
or U37755 (N_37755,N_34951,N_35923);
xor U37756 (N_37756,N_35577,N_34556);
nand U37757 (N_37757,N_34589,N_34489);
nand U37758 (N_37758,N_34180,N_35376);
nor U37759 (N_37759,N_35058,N_35100);
nor U37760 (N_37760,N_35557,N_35085);
or U37761 (N_37761,N_34769,N_35783);
nand U37762 (N_37762,N_34160,N_35934);
nand U37763 (N_37763,N_34692,N_35454);
nand U37764 (N_37764,N_34133,N_34547);
xor U37765 (N_37765,N_34118,N_34730);
xnor U37766 (N_37766,N_34033,N_34820);
and U37767 (N_37767,N_35812,N_35717);
and U37768 (N_37768,N_35047,N_34209);
or U37769 (N_37769,N_35608,N_35988);
nor U37770 (N_37770,N_34225,N_35693);
or U37771 (N_37771,N_34068,N_35191);
or U37772 (N_37772,N_35336,N_35988);
and U37773 (N_37773,N_34164,N_35312);
or U37774 (N_37774,N_35698,N_34970);
nand U37775 (N_37775,N_34188,N_34102);
nor U37776 (N_37776,N_34746,N_35496);
nor U37777 (N_37777,N_35837,N_35745);
and U37778 (N_37778,N_34439,N_34233);
or U37779 (N_37779,N_35706,N_35333);
nor U37780 (N_37780,N_35004,N_34709);
or U37781 (N_37781,N_34125,N_34002);
nand U37782 (N_37782,N_35675,N_34963);
xor U37783 (N_37783,N_35022,N_35995);
or U37784 (N_37784,N_35398,N_35711);
and U37785 (N_37785,N_35210,N_35439);
nor U37786 (N_37786,N_35101,N_34567);
and U37787 (N_37787,N_34151,N_34174);
nor U37788 (N_37788,N_35532,N_34690);
xor U37789 (N_37789,N_34431,N_35027);
and U37790 (N_37790,N_34472,N_35767);
or U37791 (N_37791,N_35177,N_34248);
xnor U37792 (N_37792,N_34801,N_34025);
nand U37793 (N_37793,N_35560,N_35443);
or U37794 (N_37794,N_34497,N_34081);
xor U37795 (N_37795,N_35167,N_34008);
xnor U37796 (N_37796,N_34016,N_35087);
nand U37797 (N_37797,N_35018,N_35935);
xor U37798 (N_37798,N_34124,N_34994);
or U37799 (N_37799,N_35672,N_35659);
and U37800 (N_37800,N_35581,N_34250);
or U37801 (N_37801,N_34395,N_34175);
nand U37802 (N_37802,N_35200,N_34886);
and U37803 (N_37803,N_35432,N_35335);
xor U37804 (N_37804,N_34915,N_35533);
or U37805 (N_37805,N_34346,N_35357);
xnor U37806 (N_37806,N_35097,N_34242);
and U37807 (N_37807,N_34643,N_35282);
nor U37808 (N_37808,N_35262,N_34656);
nand U37809 (N_37809,N_34029,N_35510);
or U37810 (N_37810,N_35943,N_34278);
nand U37811 (N_37811,N_34206,N_35947);
nor U37812 (N_37812,N_35008,N_35224);
and U37813 (N_37813,N_34504,N_35597);
nor U37814 (N_37814,N_35128,N_35728);
nor U37815 (N_37815,N_34630,N_35126);
nand U37816 (N_37816,N_34803,N_35169);
xnor U37817 (N_37817,N_35674,N_35355);
nor U37818 (N_37818,N_35328,N_34099);
and U37819 (N_37819,N_34707,N_35071);
nor U37820 (N_37820,N_34153,N_35135);
and U37821 (N_37821,N_35693,N_34226);
or U37822 (N_37822,N_34496,N_34708);
nand U37823 (N_37823,N_35734,N_35471);
and U37824 (N_37824,N_34293,N_34497);
or U37825 (N_37825,N_35099,N_35765);
nand U37826 (N_37826,N_34184,N_35519);
or U37827 (N_37827,N_34350,N_34587);
nor U37828 (N_37828,N_34402,N_34806);
xor U37829 (N_37829,N_34105,N_34549);
nor U37830 (N_37830,N_35746,N_34155);
and U37831 (N_37831,N_34601,N_34939);
or U37832 (N_37832,N_34716,N_35970);
nand U37833 (N_37833,N_35479,N_35220);
and U37834 (N_37834,N_34366,N_35324);
nor U37835 (N_37835,N_35005,N_35467);
nor U37836 (N_37836,N_35328,N_35380);
nor U37837 (N_37837,N_35894,N_35252);
or U37838 (N_37838,N_34041,N_34226);
xor U37839 (N_37839,N_35717,N_34227);
or U37840 (N_37840,N_35969,N_34047);
xnor U37841 (N_37841,N_34747,N_35681);
xor U37842 (N_37842,N_35569,N_35472);
or U37843 (N_37843,N_34280,N_34412);
nor U37844 (N_37844,N_35399,N_34535);
nand U37845 (N_37845,N_35832,N_35451);
xor U37846 (N_37846,N_34358,N_35451);
and U37847 (N_37847,N_35834,N_34608);
nor U37848 (N_37848,N_35427,N_34622);
xor U37849 (N_37849,N_35925,N_35218);
nand U37850 (N_37850,N_35180,N_34269);
and U37851 (N_37851,N_35750,N_34739);
nor U37852 (N_37852,N_34827,N_35311);
xnor U37853 (N_37853,N_35250,N_34828);
nor U37854 (N_37854,N_34065,N_34132);
xor U37855 (N_37855,N_35608,N_34127);
and U37856 (N_37856,N_34177,N_34524);
or U37857 (N_37857,N_34522,N_34814);
or U37858 (N_37858,N_35611,N_35598);
and U37859 (N_37859,N_35186,N_34433);
nand U37860 (N_37860,N_34661,N_34682);
or U37861 (N_37861,N_35102,N_34243);
or U37862 (N_37862,N_34753,N_34324);
and U37863 (N_37863,N_35619,N_34747);
and U37864 (N_37864,N_35928,N_34103);
xnor U37865 (N_37865,N_35576,N_34681);
and U37866 (N_37866,N_35523,N_35561);
xor U37867 (N_37867,N_34201,N_35195);
nand U37868 (N_37868,N_35053,N_34697);
nor U37869 (N_37869,N_35342,N_34144);
and U37870 (N_37870,N_34114,N_34178);
xor U37871 (N_37871,N_35299,N_34744);
xnor U37872 (N_37872,N_34359,N_34281);
xor U37873 (N_37873,N_35096,N_34181);
nor U37874 (N_37874,N_35956,N_35811);
and U37875 (N_37875,N_34354,N_34920);
or U37876 (N_37876,N_34336,N_35806);
or U37877 (N_37877,N_34689,N_34891);
xor U37878 (N_37878,N_35303,N_35775);
xnor U37879 (N_37879,N_35514,N_35401);
xnor U37880 (N_37880,N_34488,N_34535);
or U37881 (N_37881,N_34119,N_34206);
nor U37882 (N_37882,N_34153,N_35619);
or U37883 (N_37883,N_34079,N_35892);
or U37884 (N_37884,N_35044,N_35870);
or U37885 (N_37885,N_34723,N_34427);
nand U37886 (N_37886,N_34292,N_35001);
or U37887 (N_37887,N_34093,N_35883);
nand U37888 (N_37888,N_35086,N_35619);
nor U37889 (N_37889,N_35191,N_34338);
nor U37890 (N_37890,N_34958,N_35257);
nor U37891 (N_37891,N_34731,N_34404);
xnor U37892 (N_37892,N_35986,N_35564);
and U37893 (N_37893,N_34651,N_35111);
nor U37894 (N_37894,N_34166,N_35684);
or U37895 (N_37895,N_34089,N_35044);
and U37896 (N_37896,N_34303,N_35839);
or U37897 (N_37897,N_35113,N_35808);
and U37898 (N_37898,N_34013,N_34244);
and U37899 (N_37899,N_34048,N_35061);
nor U37900 (N_37900,N_35354,N_34219);
and U37901 (N_37901,N_34359,N_34207);
and U37902 (N_37902,N_34973,N_34956);
xor U37903 (N_37903,N_34935,N_34526);
xnor U37904 (N_37904,N_35248,N_35697);
nand U37905 (N_37905,N_35682,N_35598);
nand U37906 (N_37906,N_34880,N_34543);
nand U37907 (N_37907,N_34268,N_35931);
xor U37908 (N_37908,N_34492,N_34826);
nor U37909 (N_37909,N_35283,N_35953);
nand U37910 (N_37910,N_35878,N_34769);
nor U37911 (N_37911,N_34824,N_35261);
xnor U37912 (N_37912,N_35039,N_35930);
nor U37913 (N_37913,N_35513,N_35203);
and U37914 (N_37914,N_34635,N_34677);
nand U37915 (N_37915,N_35373,N_35314);
nor U37916 (N_37916,N_34925,N_34690);
or U37917 (N_37917,N_34436,N_35682);
nor U37918 (N_37918,N_35297,N_34662);
nand U37919 (N_37919,N_34109,N_34236);
xor U37920 (N_37920,N_34889,N_35019);
nor U37921 (N_37921,N_35440,N_35615);
or U37922 (N_37922,N_34648,N_34131);
or U37923 (N_37923,N_34134,N_34688);
xor U37924 (N_37924,N_34835,N_34910);
xor U37925 (N_37925,N_35643,N_35698);
or U37926 (N_37926,N_35923,N_35036);
nor U37927 (N_37927,N_35685,N_35313);
xor U37928 (N_37928,N_35405,N_35421);
nor U37929 (N_37929,N_34634,N_35811);
nand U37930 (N_37930,N_34901,N_35143);
nand U37931 (N_37931,N_35732,N_34312);
nand U37932 (N_37932,N_34531,N_35723);
and U37933 (N_37933,N_34028,N_35633);
or U37934 (N_37934,N_34445,N_35266);
or U37935 (N_37935,N_34836,N_34822);
nor U37936 (N_37936,N_35852,N_34794);
nand U37937 (N_37937,N_34869,N_34356);
and U37938 (N_37938,N_35363,N_35913);
xor U37939 (N_37939,N_35951,N_34472);
nand U37940 (N_37940,N_35884,N_35875);
nor U37941 (N_37941,N_35872,N_35285);
or U37942 (N_37942,N_35865,N_34966);
and U37943 (N_37943,N_35359,N_35232);
nand U37944 (N_37944,N_35296,N_35483);
xnor U37945 (N_37945,N_34453,N_35186);
nand U37946 (N_37946,N_35645,N_34891);
nor U37947 (N_37947,N_35131,N_34883);
and U37948 (N_37948,N_34478,N_34120);
nand U37949 (N_37949,N_35025,N_35247);
or U37950 (N_37950,N_35951,N_34718);
and U37951 (N_37951,N_34342,N_34068);
nand U37952 (N_37952,N_35857,N_34563);
and U37953 (N_37953,N_34063,N_35071);
and U37954 (N_37954,N_34821,N_35231);
xor U37955 (N_37955,N_35554,N_34473);
and U37956 (N_37956,N_34143,N_35631);
nor U37957 (N_37957,N_34534,N_35696);
nor U37958 (N_37958,N_35894,N_35942);
or U37959 (N_37959,N_34453,N_34444);
or U37960 (N_37960,N_35830,N_35323);
or U37961 (N_37961,N_34014,N_34970);
xnor U37962 (N_37962,N_35823,N_34523);
nor U37963 (N_37963,N_34993,N_34947);
and U37964 (N_37964,N_34212,N_35418);
nand U37965 (N_37965,N_35815,N_34428);
nand U37966 (N_37966,N_35191,N_34993);
nor U37967 (N_37967,N_34430,N_34306);
nand U37968 (N_37968,N_34775,N_35194);
or U37969 (N_37969,N_34585,N_34354);
nand U37970 (N_37970,N_34979,N_34801);
and U37971 (N_37971,N_34179,N_34593);
or U37972 (N_37972,N_35914,N_35852);
nor U37973 (N_37973,N_35370,N_34903);
or U37974 (N_37974,N_35591,N_34762);
and U37975 (N_37975,N_35497,N_34470);
and U37976 (N_37976,N_35769,N_35067);
nand U37977 (N_37977,N_34915,N_35116);
xor U37978 (N_37978,N_35957,N_34687);
xnor U37979 (N_37979,N_35180,N_35847);
and U37980 (N_37980,N_34565,N_34629);
and U37981 (N_37981,N_35591,N_34829);
nand U37982 (N_37982,N_35182,N_34937);
xor U37983 (N_37983,N_34158,N_35697);
xnor U37984 (N_37984,N_34338,N_34090);
or U37985 (N_37985,N_34602,N_34368);
nor U37986 (N_37986,N_35374,N_35024);
or U37987 (N_37987,N_35360,N_34121);
nand U37988 (N_37988,N_35706,N_35777);
or U37989 (N_37989,N_34259,N_34636);
and U37990 (N_37990,N_35004,N_34423);
nand U37991 (N_37991,N_34202,N_34435);
or U37992 (N_37992,N_34965,N_35730);
nand U37993 (N_37993,N_35709,N_34137);
or U37994 (N_37994,N_34770,N_34414);
nand U37995 (N_37995,N_35302,N_35689);
xnor U37996 (N_37996,N_35803,N_35302);
and U37997 (N_37997,N_35413,N_35677);
xor U37998 (N_37998,N_34521,N_34655);
or U37999 (N_37999,N_35789,N_35600);
xor U38000 (N_38000,N_37785,N_37691);
or U38001 (N_38001,N_36149,N_36876);
nand U38002 (N_38002,N_37492,N_37346);
and U38003 (N_38003,N_36628,N_36317);
nor U38004 (N_38004,N_36698,N_37729);
xnor U38005 (N_38005,N_36042,N_37875);
nand U38006 (N_38006,N_37893,N_36569);
and U38007 (N_38007,N_36140,N_37982);
nand U38008 (N_38008,N_37139,N_36986);
xnor U38009 (N_38009,N_37291,N_36534);
and U38010 (N_38010,N_36286,N_37929);
nand U38011 (N_38011,N_36898,N_37626);
nor U38012 (N_38012,N_37207,N_37718);
or U38013 (N_38013,N_36475,N_36394);
or U38014 (N_38014,N_36764,N_37411);
nand U38015 (N_38015,N_36830,N_36875);
nand U38016 (N_38016,N_37822,N_36298);
xor U38017 (N_38017,N_36603,N_37027);
nand U38018 (N_38018,N_36491,N_36770);
nand U38019 (N_38019,N_37337,N_36520);
and U38020 (N_38020,N_37656,N_37274);
nor U38021 (N_38021,N_37111,N_37939);
or U38022 (N_38022,N_36863,N_36581);
and U38023 (N_38023,N_36307,N_36154);
nor U38024 (N_38024,N_36881,N_37428);
nand U38025 (N_38025,N_36445,N_37062);
nand U38026 (N_38026,N_36841,N_36405);
nand U38027 (N_38027,N_36783,N_36952);
nand U38028 (N_38028,N_37572,N_37366);
nor U38029 (N_38029,N_36991,N_37717);
or U38030 (N_38030,N_36277,N_37142);
nor U38031 (N_38031,N_36145,N_36413);
or U38032 (N_38032,N_36153,N_36275);
and U38033 (N_38033,N_36195,N_36867);
xor U38034 (N_38034,N_36811,N_37906);
or U38035 (N_38035,N_37059,N_37852);
and U38036 (N_38036,N_37349,N_36339);
or U38037 (N_38037,N_37077,N_37424);
or U38038 (N_38038,N_36172,N_37132);
xor U38039 (N_38039,N_37553,N_36329);
and U38040 (N_38040,N_36296,N_37797);
nor U38041 (N_38041,N_36548,N_36449);
nand U38042 (N_38042,N_37234,N_36415);
nand U38043 (N_38043,N_36654,N_36079);
and U38044 (N_38044,N_37280,N_37767);
nand U38045 (N_38045,N_36142,N_37360);
and U38046 (N_38046,N_36926,N_37598);
or U38047 (N_38047,N_36285,N_36860);
nor U38048 (N_38048,N_37526,N_37092);
xor U38049 (N_38049,N_37934,N_37272);
and U38050 (N_38050,N_37375,N_37335);
and U38051 (N_38051,N_37815,N_36980);
and U38052 (N_38052,N_37447,N_36459);
nor U38053 (N_38053,N_37556,N_37429);
xnor U38054 (N_38054,N_37477,N_36139);
xnor U38055 (N_38055,N_36141,N_36385);
nand U38056 (N_38056,N_37339,N_37867);
xnor U38057 (N_38057,N_37571,N_36144);
xnor U38058 (N_38058,N_36780,N_36564);
nor U38059 (N_38059,N_36211,N_36524);
and U38060 (N_38060,N_37136,N_36801);
and U38061 (N_38061,N_36466,N_36041);
xor U38062 (N_38062,N_36454,N_36559);
or U38063 (N_38063,N_37780,N_36955);
nor U38064 (N_38064,N_37392,N_36210);
or U38065 (N_38065,N_36773,N_36412);
nor U38066 (N_38066,N_36127,N_36810);
nor U38067 (N_38067,N_36176,N_37200);
xnor U38068 (N_38068,N_37277,N_36993);
and U38069 (N_38069,N_36276,N_36212);
nand U38070 (N_38070,N_36798,N_37282);
or U38071 (N_38071,N_36664,N_36113);
or U38072 (N_38072,N_37009,N_36486);
nor U38073 (N_38073,N_37568,N_36814);
nand U38074 (N_38074,N_37472,N_37849);
xor U38075 (N_38075,N_37733,N_36477);
nor U38076 (N_38076,N_37823,N_36974);
and U38077 (N_38077,N_37805,N_37298);
nand U38078 (N_38078,N_36049,N_36168);
or U38079 (N_38079,N_36938,N_36723);
xnor U38080 (N_38080,N_36761,N_37180);
and U38081 (N_38081,N_36273,N_37205);
xnor U38082 (N_38082,N_36341,N_37373);
nor U38083 (N_38083,N_36021,N_37258);
nor U38084 (N_38084,N_37854,N_36853);
and U38085 (N_38085,N_37026,N_36418);
xnor U38086 (N_38086,N_36743,N_36312);
nor U38087 (N_38087,N_36242,N_36512);
nor U38088 (N_38088,N_36604,N_36782);
or U38089 (N_38089,N_36992,N_36779);
nor U38090 (N_38090,N_37203,N_37348);
nor U38091 (N_38091,N_37932,N_36998);
xor U38092 (N_38092,N_36589,N_37061);
nand U38093 (N_38093,N_36771,N_37157);
or U38094 (N_38094,N_36766,N_37618);
and U38095 (N_38095,N_37523,N_37511);
xnor U38096 (N_38096,N_37228,N_36774);
xor U38097 (N_38097,N_36636,N_37028);
xnor U38098 (N_38098,N_36557,N_37218);
or U38099 (N_38099,N_36487,N_36895);
and U38100 (N_38100,N_37992,N_36631);
nand U38101 (N_38101,N_36692,N_37172);
nor U38102 (N_38102,N_37538,N_37145);
and U38103 (N_38103,N_36816,N_37701);
xnor U38104 (N_38104,N_36778,N_36015);
xor U38105 (N_38105,N_36889,N_36755);
nand U38106 (N_38106,N_36874,N_36805);
and U38107 (N_38107,N_37605,N_37476);
nor U38108 (N_38108,N_37094,N_36130);
nor U38109 (N_38109,N_37898,N_36157);
nand U38110 (N_38110,N_37403,N_37487);
nor U38111 (N_38111,N_37400,N_36790);
or U38112 (N_38112,N_36505,N_37922);
and U38113 (N_38113,N_37301,N_37935);
nand U38114 (N_38114,N_37819,N_37249);
or U38115 (N_38115,N_36960,N_36202);
nand U38116 (N_38116,N_37226,N_36733);
and U38117 (N_38117,N_36851,N_36036);
and U38118 (N_38118,N_37548,N_36767);
and U38119 (N_38119,N_37612,N_36138);
nor U38120 (N_38120,N_36359,N_36367);
or U38121 (N_38121,N_36084,N_36769);
or U38122 (N_38122,N_37999,N_37760);
or U38123 (N_38123,N_37319,N_36326);
and U38124 (N_38124,N_36468,N_36802);
nor U38125 (N_38125,N_36201,N_36833);
nor U38126 (N_38126,N_37372,N_37166);
or U38127 (N_38127,N_37897,N_36279);
and U38128 (N_38128,N_36575,N_36229);
and U38129 (N_38129,N_37918,N_36431);
nor U38130 (N_38130,N_36797,N_37243);
nor U38131 (N_38131,N_37821,N_36885);
or U38132 (N_38132,N_37161,N_36701);
nand U38133 (N_38133,N_37536,N_36726);
nor U38134 (N_38134,N_36350,N_36082);
or U38135 (N_38135,N_36132,N_37387);
nand U38136 (N_38136,N_36111,N_36072);
xor U38137 (N_38137,N_36147,N_37021);
or U38138 (N_38138,N_36563,N_36725);
xor U38139 (N_38139,N_37160,N_37017);
nor U38140 (N_38140,N_36002,N_37834);
nand U38141 (N_38141,N_37457,N_36682);
xor U38142 (N_38142,N_37962,N_36781);
nor U38143 (N_38143,N_36092,N_37383);
and U38144 (N_38144,N_36194,N_37738);
and U38145 (N_38145,N_36513,N_36035);
or U38146 (N_38146,N_37037,N_36788);
or U38147 (N_38147,N_37762,N_36492);
nor U38148 (N_38148,N_36862,N_37546);
or U38149 (N_38149,N_37911,N_37155);
and U38150 (N_38150,N_37613,N_36186);
or U38151 (N_38151,N_37238,N_37471);
xor U38152 (N_38152,N_37550,N_36443);
nand U38153 (N_38153,N_37545,N_37997);
xnor U38154 (N_38154,N_36947,N_37789);
nor U38155 (N_38155,N_36489,N_36568);
and U38156 (N_38156,N_37745,N_37475);
nand U38157 (N_38157,N_36228,N_36984);
nand U38158 (N_38158,N_36458,N_36966);
nor U38159 (N_38159,N_36989,N_37557);
xnor U38160 (N_38160,N_37287,N_36572);
and U38161 (N_38161,N_37670,N_36836);
nor U38162 (N_38162,N_36691,N_37576);
nand U38163 (N_38163,N_36261,N_37253);
or U38164 (N_38164,N_36735,N_37667);
nor U38165 (N_38165,N_37498,N_36705);
and U38166 (N_38166,N_36732,N_36452);
nand U38167 (N_38167,N_36839,N_37371);
or U38168 (N_38168,N_36233,N_37955);
xor U38169 (N_38169,N_37352,N_37215);
nand U38170 (N_38170,N_37254,N_36806);
nand U38171 (N_38171,N_36180,N_37079);
nor U38172 (N_38172,N_36406,N_36050);
nor U38173 (N_38173,N_37835,N_36820);
or U38174 (N_38174,N_36346,N_37883);
xnor U38175 (N_38175,N_36511,N_37659);
nor U38176 (N_38176,N_36174,N_36185);
or U38177 (N_38177,N_37799,N_37887);
nor U38178 (N_38178,N_36029,N_37844);
xor U38179 (N_38179,N_36845,N_36920);
xor U38180 (N_38180,N_37378,N_36944);
and U38181 (N_38181,N_36122,N_36541);
xnor U38182 (N_38182,N_36358,N_36422);
nand U38183 (N_38183,N_36754,N_36638);
nand U38184 (N_38184,N_37022,N_37574);
and U38185 (N_38185,N_36582,N_36982);
or U38186 (N_38186,N_36686,N_37578);
xor U38187 (N_38187,N_36794,N_36590);
and U38188 (N_38188,N_36197,N_36073);
xor U38189 (N_38189,N_36223,N_37833);
and U38190 (N_38190,N_36646,N_37053);
nor U38191 (N_38191,N_37169,N_37953);
xnor U38192 (N_38192,N_37096,N_37227);
xnor U38193 (N_38193,N_36995,N_36643);
xnor U38194 (N_38194,N_37908,N_36509);
and U38195 (N_38195,N_37904,N_36265);
xnor U38196 (N_38196,N_36598,N_37007);
nand U38197 (N_38197,N_36518,N_36450);
xor U38198 (N_38198,N_36252,N_37485);
nor U38199 (N_38199,N_36403,N_37871);
nor U38200 (N_38200,N_37812,N_36561);
and U38201 (N_38201,N_36759,N_36745);
xnor U38202 (N_38202,N_37882,N_36245);
nor U38203 (N_38203,N_36463,N_37879);
and U38204 (N_38204,N_37054,N_37630);
and U38205 (N_38205,N_37134,N_37240);
nand U38206 (N_38206,N_37531,N_36493);
xnor U38207 (N_38207,N_36043,N_37845);
or U38208 (N_38208,N_36374,N_37664);
nor U38209 (N_38209,N_36118,N_36900);
and U38210 (N_38210,N_37299,N_37281);
nor U38211 (N_38211,N_36813,N_36356);
xor U38212 (N_38212,N_37537,N_37303);
or U38213 (N_38213,N_37996,N_37310);
and U38214 (N_38214,N_36430,N_36940);
nand U38215 (N_38215,N_37231,N_36232);
xor U38216 (N_38216,N_37003,N_37005);
nor U38217 (N_38217,N_37636,N_37316);
or U38218 (N_38218,N_36973,N_37338);
xnor U38219 (N_38219,N_36488,N_36361);
nor U38220 (N_38220,N_37236,N_36439);
and U38221 (N_38221,N_37391,N_37314);
xnor U38222 (N_38222,N_37412,N_36784);
and U38223 (N_38223,N_36155,N_36856);
nor U38224 (N_38224,N_37580,N_37486);
and U38225 (N_38225,N_37792,N_36469);
nor U38226 (N_38226,N_36181,N_36190);
nand U38227 (N_38227,N_36251,N_36303);
xnor U38228 (N_38228,N_37355,N_37719);
nand U38229 (N_38229,N_36268,N_36409);
nor U38230 (N_38230,N_36227,N_37500);
or U38231 (N_38231,N_37210,N_36007);
or U38232 (N_38232,N_37095,N_37270);
nor U38233 (N_38233,N_37924,N_37067);
or U38234 (N_38234,N_36510,N_37680);
xor U38235 (N_38235,N_37588,N_36667);
or U38236 (N_38236,N_36347,N_37004);
nor U38237 (N_38237,N_37824,N_36397);
nand U38238 (N_38238,N_37133,N_36230);
nand U38239 (N_38239,N_36234,N_36956);
xor U38240 (N_38240,N_36474,N_36380);
and U38241 (N_38241,N_36437,N_36967);
nand U38242 (N_38242,N_36205,N_37229);
nand U38243 (N_38243,N_36479,N_36095);
nor U38244 (N_38244,N_36017,N_36320);
or U38245 (N_38245,N_36090,N_37857);
and U38246 (N_38246,N_36131,N_36057);
nor U38247 (N_38247,N_36150,N_37149);
nor U38248 (N_38248,N_37599,N_36419);
or U38249 (N_38249,N_37765,N_36535);
or U38250 (N_38250,N_37436,N_36997);
nor U38251 (N_38251,N_36004,N_37611);
xor U38252 (N_38252,N_36121,N_37730);
xnor U38253 (N_38253,N_36522,N_36602);
xnor U38254 (N_38254,N_37945,N_36679);
nand U38255 (N_38255,N_36546,N_36968);
or U38256 (N_38256,N_37665,N_37855);
and U38257 (N_38257,N_37195,N_36096);
xor U38258 (N_38258,N_36390,N_36316);
nand U38259 (N_38259,N_36278,N_36653);
and U38260 (N_38260,N_36872,N_36508);
nand U38261 (N_38261,N_37582,N_37441);
or U38262 (N_38262,N_37478,N_37164);
nor U38263 (N_38263,N_37581,N_37863);
or U38264 (N_38264,N_36829,N_36503);
nand U38265 (N_38265,N_36013,N_36565);
and U38266 (N_38266,N_36681,N_36873);
and U38267 (N_38267,N_36584,N_36869);
nand U38268 (N_38268,N_36442,N_37980);
nand U38269 (N_38269,N_36687,N_36832);
nand U38270 (N_38270,N_37802,N_37137);
nand U38271 (N_38271,N_37330,N_36941);
or U38272 (N_38272,N_36948,N_36399);
and U38273 (N_38273,N_37858,N_37127);
and U38274 (N_38274,N_37451,N_36351);
nor U38275 (N_38275,N_36617,N_37547);
and U38276 (N_38276,N_36507,N_36531);
nor U38277 (N_38277,N_36169,N_36578);
nand U38278 (N_38278,N_36901,N_37023);
nor U38279 (N_38279,N_37551,N_37591);
nand U38280 (N_38280,N_36614,N_36124);
xnor U38281 (N_38281,N_37920,N_37047);
and U38282 (N_38282,N_37178,N_36388);
or U38283 (N_38283,N_36777,N_37596);
or U38284 (N_38284,N_36987,N_36461);
and U38285 (N_38285,N_37088,N_36842);
nor U38286 (N_38286,N_37484,N_36537);
xor U38287 (N_38287,N_36824,N_37367);
nand U38288 (N_38288,N_36718,N_37758);
or U38289 (N_38289,N_36069,N_37524);
xnor U38290 (N_38290,N_36971,N_37933);
and U38291 (N_38291,N_36758,N_36396);
and U38292 (N_38292,N_37099,N_36818);
xnor U38293 (N_38293,N_36495,N_37621);
nand U38294 (N_38294,N_37552,N_37187);
nor U38295 (N_38295,N_36676,N_37831);
xor U38296 (N_38296,N_37135,N_37756);
or U38297 (N_38297,N_37516,N_37507);
xor U38298 (N_38298,N_36498,N_36056);
nor U38299 (N_38299,N_36914,N_37827);
xor U38300 (N_38300,N_37791,N_37422);
and U38301 (N_38301,N_36293,N_37057);
or U38302 (N_38302,N_37888,N_36429);
nand U38303 (N_38303,N_37752,N_37525);
or U38304 (N_38304,N_36360,N_37936);
nor U38305 (N_38305,N_37016,N_36099);
nand U38306 (N_38306,N_36594,N_37640);
nand U38307 (N_38307,N_37940,N_37695);
or U38308 (N_38308,N_36378,N_36663);
nor U38309 (N_38309,N_36158,N_37259);
and U38310 (N_38310,N_36903,N_36203);
or U38311 (N_38311,N_36465,N_37952);
or U38312 (N_38312,N_36135,N_36864);
or U38313 (N_38313,N_36707,N_37419);
and U38314 (N_38314,N_36193,N_36595);
or U38315 (N_38315,N_36068,N_36440);
or U38316 (N_38316,N_36206,N_37326);
or U38317 (N_38317,N_37862,N_36384);
nor U38318 (N_38318,N_36609,N_37423);
nand U38319 (N_38319,N_37570,N_36476);
xnor U38320 (N_38320,N_36250,N_37396);
nand U38321 (N_38321,N_36803,N_37151);
or U38322 (N_38322,N_37600,N_36456);
or U38323 (N_38323,N_37344,N_37084);
nor U38324 (N_38324,N_36807,N_36527);
xnor U38325 (N_38325,N_37150,N_36763);
or U38326 (N_38326,N_36151,N_37290);
nor U38327 (N_38327,N_36648,N_36426);
or U38328 (N_38328,N_36455,N_36100);
or U38329 (N_38329,N_37465,N_36792);
nand U38330 (N_38330,N_37579,N_36672);
and U38331 (N_38331,N_36933,N_36787);
or U38332 (N_38332,N_37090,N_36846);
and U38333 (N_38333,N_36173,N_37710);
nand U38334 (N_38334,N_36752,N_37499);
nand U38335 (N_38335,N_36539,N_36785);
nand U38336 (N_38336,N_36552,N_37774);
and U38337 (N_38337,N_37121,N_36645);
nor U38338 (N_38338,N_37928,N_37244);
xnor U38339 (N_38339,N_36460,N_37113);
xnor U38340 (N_38340,N_37171,N_37881);
nor U38341 (N_38341,N_37702,N_37850);
xor U38342 (N_38342,N_36331,N_37644);
or U38343 (N_38343,N_37284,N_37811);
or U38344 (N_38344,N_36936,N_37608);
nor U38345 (N_38345,N_37035,N_37211);
and U38346 (N_38346,N_36289,N_36930);
and U38347 (N_38347,N_37394,N_36854);
xnor U38348 (N_38348,N_36272,N_36420);
nand U38349 (N_38349,N_37329,N_37575);
nand U38350 (N_38350,N_37619,N_37075);
or U38351 (N_38351,N_36655,N_36529);
and U38352 (N_38352,N_36625,N_37777);
nor U38353 (N_38353,N_36526,N_36402);
nand U38354 (N_38354,N_37223,N_37304);
xnor U38355 (N_38355,N_36046,N_37617);
nor U38356 (N_38356,N_37770,N_37241);
nor U38357 (N_38357,N_36961,N_37709);
and U38358 (N_38358,N_37776,N_37165);
or U38359 (N_38359,N_36975,N_36204);
xnor U38360 (N_38360,N_37444,N_36152);
nor U38361 (N_38361,N_37216,N_37179);
xor U38362 (N_38362,N_37185,N_37721);
and U38363 (N_38363,N_37430,N_36184);
nand U38364 (N_38364,N_36170,N_37753);
xnor U38365 (N_38365,N_36985,N_37638);
or U38366 (N_38366,N_37377,N_37724);
xnor U38367 (N_38367,N_37828,N_36040);
nor U38368 (N_38368,N_37464,N_37981);
nor U38369 (N_38369,N_36677,N_37884);
nand U38370 (N_38370,N_37779,N_36086);
xnor U38371 (N_38371,N_36462,N_36299);
or U38372 (N_38372,N_37832,N_37554);
xnor U38373 (N_38373,N_37331,N_37439);
nor U38374 (N_38374,N_37184,N_37517);
nand U38375 (N_38375,N_37450,N_37983);
or U38376 (N_38376,N_37808,N_37105);
nor U38377 (N_38377,N_36922,N_37109);
and U38378 (N_38378,N_36586,N_36244);
or U38379 (N_38379,N_37255,N_37217);
nor U38380 (N_38380,N_36239,N_36321);
nor U38381 (N_38381,N_36349,N_36747);
nor U38382 (N_38382,N_36262,N_36642);
and U38383 (N_38383,N_36847,N_37182);
and U38384 (N_38384,N_37707,N_36815);
and U38385 (N_38385,N_37183,N_37083);
nand U38386 (N_38386,N_36030,N_36545);
or U38387 (N_38387,N_36247,N_37562);
and U38388 (N_38388,N_36963,N_37878);
and U38389 (N_38389,N_36633,N_36480);
nor U38390 (N_38390,N_36470,N_36407);
xnor U38391 (N_38391,N_37409,N_36125);
nand U38392 (N_38392,N_36668,N_37325);
xor U38393 (N_38393,N_37196,N_37972);
or U38394 (N_38394,N_37452,N_37842);
nand U38395 (N_38395,N_36037,N_36685);
nand U38396 (N_38396,N_37503,N_37045);
nand U38397 (N_38397,N_36704,N_36435);
or U38398 (N_38398,N_37690,N_37804);
nand U38399 (N_38399,N_36292,N_36490);
nor U38400 (N_38400,N_37896,N_36156);
nor U38401 (N_38401,N_36608,N_37408);
or U38402 (N_38402,N_36301,N_37984);
nor U38403 (N_38403,N_36722,N_36644);
nor U38404 (N_38404,N_36696,N_36106);
nand U38405 (N_38405,N_36219,N_36884);
or U38406 (N_38406,N_37432,N_36924);
nor U38407 (N_38407,N_36300,N_37964);
nand U38408 (N_38408,N_37629,N_37610);
and U38409 (N_38409,N_36280,N_36721);
nor U38410 (N_38410,N_37720,N_36626);
xnor U38411 (N_38411,N_37589,N_36207);
xnor U38412 (N_38412,N_36621,N_37220);
nand U38413 (N_38413,N_36762,N_36238);
or U38414 (N_38414,N_36728,N_36994);
xnor U38415 (N_38415,N_37773,N_37642);
nor U38416 (N_38416,N_36379,N_36432);
nor U38417 (N_38417,N_37489,N_36371);
or U38418 (N_38418,N_36757,N_36905);
xor U38419 (N_38419,N_36965,N_36632);
and U38420 (N_38420,N_36327,N_37769);
and U38421 (N_38421,N_36249,N_36870);
xnor U38422 (N_38422,N_37052,N_37836);
nand U38423 (N_38423,N_37081,N_37469);
and U38424 (N_38424,N_37410,N_36817);
or U38425 (N_38425,N_37624,N_36161);
or U38426 (N_38426,N_37970,N_36673);
xnor U38427 (N_38427,N_36949,N_37232);
and U38428 (N_38428,N_36266,N_37388);
or U38429 (N_38429,N_37941,N_36005);
nor U38430 (N_38430,N_36964,N_37625);
and U38431 (N_38431,N_37675,N_36906);
and U38432 (N_38432,N_36362,N_37189);
xor U38433 (N_38433,N_36908,N_36925);
or U38434 (N_38434,N_37341,N_36216);
xnor U38435 (N_38435,N_37307,N_37239);
nand U38436 (N_38436,N_37968,N_36683);
or U38437 (N_38437,N_36983,N_37063);
nor U38438 (N_38438,N_36850,N_37816);
nor U38439 (N_38439,N_36753,N_37010);
and U38440 (N_38440,N_36026,N_36220);
or U38441 (N_38441,N_37191,N_37129);
nand U38442 (N_38442,N_36795,N_36182);
or U38443 (N_38443,N_37944,N_37861);
and U38444 (N_38444,N_36235,N_36164);
nor U38445 (N_38445,N_36979,N_36143);
and U38446 (N_38446,N_37990,N_37639);
and U38447 (N_38447,N_36613,N_36697);
nor U38448 (N_38448,N_37114,N_37930);
and U38449 (N_38449,N_36381,N_36583);
and U38450 (N_38450,N_37379,N_36776);
nand U38451 (N_38451,N_36283,N_36434);
xor U38452 (N_38452,N_36011,N_36256);
or U38453 (N_38453,N_36953,N_36464);
and U38454 (N_38454,N_37085,N_36404);
nor U38455 (N_38455,N_36916,N_36751);
nor U38456 (N_38456,N_36800,N_36352);
or U38457 (N_38457,N_37544,N_37755);
nor U38458 (N_38458,N_37851,N_37885);
nand U38459 (N_38459,N_36684,N_37480);
and U38460 (N_38460,N_37015,N_37839);
and U38461 (N_38461,N_36714,N_37697);
nand U38462 (N_38462,N_36091,N_37495);
nor U38463 (N_38463,N_36886,N_36446);
xor U38464 (N_38464,N_37199,N_37462);
or U38465 (N_38465,N_36083,N_37097);
and U38466 (N_38466,N_36198,N_36647);
nor U38467 (N_38467,N_36045,N_36738);
nor U38468 (N_38468,N_37632,N_37306);
and U38469 (N_38469,N_37006,N_37497);
xor U38470 (N_38470,N_37402,N_37604);
and U38471 (N_38471,N_37772,N_36260);
and U38472 (N_38472,N_37332,N_37261);
nor U38473 (N_38473,N_36313,N_36809);
nand U38474 (N_38474,N_37748,N_37198);
nand U38475 (N_38475,N_36291,N_36427);
and U38476 (N_38476,N_36731,N_37741);
xnor U38477 (N_38477,N_36009,N_36627);
nor U38478 (N_38478,N_36544,N_37567);
nand U38479 (N_38479,N_37156,N_37682);
nand U38480 (N_38480,N_36003,N_36183);
nand U38481 (N_38481,N_36727,N_37584);
nor U38482 (N_38482,N_36592,N_37159);
nor U38483 (N_38483,N_37643,N_37583);
xor U38484 (N_38484,N_37627,N_37740);
nand U38485 (N_38485,N_36913,N_36719);
nand U38486 (N_38486,N_37672,N_36369);
or U38487 (N_38487,N_36191,N_36530);
or U38488 (N_38488,N_36689,N_36890);
nor U38489 (N_38489,N_36616,N_37807);
and U38490 (N_38490,N_37494,N_36093);
xor U38491 (N_38491,N_36052,N_37687);
xnor U38492 (N_38492,N_36615,N_37201);
nor U38493 (N_38493,N_36451,N_37739);
nand U38494 (N_38494,N_36772,N_36547);
or U38495 (N_38495,N_37312,N_36218);
xor U38496 (N_38496,N_37263,N_37957);
and U38497 (N_38497,N_36253,N_36319);
nor U38498 (N_38498,N_37946,N_37998);
nor U38499 (N_38499,N_37676,N_37974);
nor U38500 (N_38500,N_36146,N_37175);
nor U38501 (N_38501,N_36416,N_36958);
and U38502 (N_38502,N_36942,N_36659);
and U38503 (N_38503,N_37374,N_36240);
xor U38504 (N_38504,N_37786,N_36760);
or U38505 (N_38505,N_37705,N_37445);
xnor U38506 (N_38506,N_36775,N_36827);
nor U38507 (N_38507,N_37837,N_37043);
nand U38508 (N_38508,N_37224,N_36536);
xor U38509 (N_38509,N_36306,N_36333);
xor U38510 (N_38510,N_37810,N_37768);
and U38511 (N_38511,N_37206,N_36107);
nor U38512 (N_38512,N_36226,N_36678);
nand U38513 (N_38513,N_36573,N_37628);
nor U38514 (N_38514,N_36259,N_36571);
xnor U38515 (N_38515,N_37986,N_37110);
xnor U38516 (N_38516,N_36109,N_37712);
nor U38517 (N_38517,N_37395,N_37747);
nor U38518 (N_38518,N_37937,N_37385);
nor U38519 (N_38519,N_37141,N_36022);
or U38520 (N_38520,N_36270,N_37317);
or U38521 (N_38521,N_37685,N_36500);
and U38522 (N_38522,N_36389,N_36902);
nor U38523 (N_38523,N_37509,N_36533);
and U38524 (N_38524,N_36742,N_36893);
or U38525 (N_38525,N_37123,N_37293);
and U38526 (N_38526,N_36910,N_36789);
nand U38527 (N_38527,N_36858,N_36282);
nor U38528 (N_38528,N_36935,N_36504);
nor U38529 (N_38529,N_37907,N_37460);
or U38530 (N_38530,N_36484,N_36657);
nand U38531 (N_38531,N_36756,N_36264);
and U38532 (N_38532,N_36823,N_36467);
or U38533 (N_38533,N_37654,N_36551);
xnor U38534 (N_38534,N_36322,N_37308);
and U38535 (N_38535,N_36651,N_37848);
and U38536 (N_38536,N_36661,N_36115);
nand U38537 (N_38537,N_37176,N_37784);
and U38538 (N_38538,N_36000,N_36295);
xor U38539 (N_38539,N_37264,N_36162);
or U38540 (N_38540,N_36243,N_36088);
nand U38541 (N_38541,N_37260,N_37000);
or U38542 (N_38542,N_36137,N_37056);
nand U38543 (N_38543,N_36310,N_37222);
nand U38544 (N_38544,N_37091,N_37534);
nand U38545 (N_38545,N_37154,N_36969);
or U38546 (N_38546,N_36410,N_37434);
nor U38547 (N_38547,N_36062,N_37798);
nor U38548 (N_38548,N_36354,N_37530);
nor U38549 (N_38549,N_37448,N_37369);
and U38550 (N_38550,N_36528,N_36365);
nor U38551 (N_38551,N_36712,N_36217);
nand U38552 (N_38552,N_37637,N_36209);
xor U38553 (N_38553,N_36515,N_37662);
nand U38554 (N_38554,N_37783,N_36167);
and U38555 (N_38555,N_36812,N_37148);
nand U38556 (N_38556,N_37873,N_37728);
nor U38557 (N_38557,N_37603,N_36222);
xor U38558 (N_38558,N_36257,N_36724);
nor U38559 (N_38559,N_37267,N_37734);
and U38560 (N_38560,N_36302,N_37488);
xnor U38561 (N_38561,N_36748,N_37988);
or U38562 (N_38562,N_36671,N_36032);
and U38563 (N_38563,N_36213,N_36166);
and U38564 (N_38564,N_36117,N_37197);
or U38565 (N_38565,N_37788,N_37917);
nor U38566 (N_38566,N_37324,N_36258);
xor U38567 (N_38567,N_37221,N_36129);
and U38568 (N_38568,N_36104,N_36972);
nor U38569 (N_38569,N_36255,N_36236);
xnor U38570 (N_38570,N_37311,N_37292);
nor U38571 (N_38571,N_36324,N_36074);
nand U38572 (N_38572,N_36880,N_37120);
nor U38573 (N_38573,N_37297,N_36383);
nor U38574 (N_38574,N_37468,N_37066);
nand U38575 (N_38575,N_36148,N_37302);
nand U38576 (N_38576,N_37796,N_36819);
or U38577 (N_38577,N_37188,N_37969);
and U38578 (N_38578,N_36835,N_36134);
nand U38579 (N_38579,N_36108,N_37322);
and U38580 (N_38580,N_36408,N_37749);
and U38581 (N_38581,N_37723,N_36308);
xnor U38582 (N_38582,N_37426,N_37731);
xor U38583 (N_38583,N_36221,N_36611);
nand U38584 (N_38584,N_37595,N_37615);
nor U38585 (N_38585,N_37458,N_37529);
xor U38586 (N_38586,N_36502,N_37233);
or U38587 (N_38587,N_37496,N_36826);
nor U38588 (N_38588,N_37295,N_36919);
nand U38589 (N_38589,N_36523,N_37563);
or U38590 (N_38590,N_37735,N_37473);
nor U38591 (N_38591,N_36060,N_36281);
or U38592 (N_38592,N_36020,N_36336);
or U38593 (N_38593,N_37493,N_37902);
and U38594 (N_38594,N_37153,N_37813);
xnor U38595 (N_38595,N_37686,N_37128);
or U38596 (N_38596,N_37616,N_37961);
or U38597 (N_38597,N_37989,N_36746);
nand U38598 (N_38598,N_36305,N_36345);
nand U38599 (N_38599,N_37407,N_36662);
xor U38600 (N_38600,N_36428,N_36943);
xor U38601 (N_38601,N_36178,N_36976);
xnor U38602 (N_38602,N_37118,N_36635);
nor U38603 (N_38603,N_36694,N_37041);
nand U38604 (N_38604,N_37903,N_37116);
or U38605 (N_38605,N_37177,N_37696);
nand U38606 (N_38606,N_37520,N_36838);
xor U38607 (N_38607,N_37271,N_36897);
nand U38608 (N_38608,N_37087,N_36912);
and U38609 (N_38609,N_36921,N_36840);
nand U38610 (N_38610,N_36640,N_37869);
nand U38611 (N_38611,N_37384,N_36622);
or U38612 (N_38612,N_37895,N_36453);
nand U38613 (N_38613,N_36039,N_36363);
or U38614 (N_38614,N_37703,N_37050);
nand U38615 (N_38615,N_37014,N_37300);
and U38616 (N_38616,N_37759,N_37449);
and U38617 (N_38617,N_37590,N_37751);
xnor U38618 (N_38618,N_37518,N_37973);
xnor U38619 (N_38619,N_37162,N_36749);
nand U38620 (N_38620,N_37560,N_36928);
xnor U38621 (N_38621,N_36868,N_36457);
and U38622 (N_38622,N_36999,N_37040);
nor U38623 (N_38623,N_37512,N_36549);
and U38624 (N_38624,N_36496,N_37782);
or U38625 (N_38625,N_37726,N_37649);
and U38626 (N_38626,N_36087,N_37029);
or U38627 (N_38627,N_36641,N_37289);
and U38628 (N_38628,N_36699,N_37305);
nand U38629 (N_38629,N_37381,N_37020);
nand U38630 (N_38630,N_36931,N_36423);
nand U38631 (N_38631,N_37661,N_36330);
and U38632 (N_38632,N_37513,N_36016);
nor U38633 (N_38633,N_36497,N_37283);
nor U38634 (N_38634,N_37757,N_36377);
or U38635 (N_38635,N_37651,N_36481);
and U38636 (N_38636,N_36825,N_37931);
xnor U38637 (N_38637,N_36702,N_37692);
nand U38638 (N_38638,N_36297,N_37514);
or U38639 (N_38639,N_36828,N_37795);
nor U38640 (N_38640,N_36950,N_36438);
nor U38641 (N_38641,N_37089,N_36652);
nor U38642 (N_38642,N_36294,N_36105);
xnor U38643 (N_38643,N_37947,N_36514);
or U38644 (N_38644,N_37925,N_36978);
xor U38645 (N_38645,N_37086,N_36175);
nand U38646 (N_38646,N_36580,N_37713);
nand U38647 (N_38647,N_37323,N_37192);
nand U38648 (N_38648,N_36623,N_37362);
xnor U38649 (N_38649,N_37204,N_37737);
and U38650 (N_38650,N_36945,N_37678);
and U38651 (N_38651,N_37257,N_36558);
and U38652 (N_38652,N_37108,N_37645);
nor U38653 (N_38653,N_36048,N_37586);
or U38654 (N_38654,N_37031,N_37490);
nor U38655 (N_38655,N_37328,N_36012);
xor U38656 (N_38656,N_37569,N_37318);
or U38657 (N_38657,N_37076,N_37843);
xor U38658 (N_38658,N_37971,N_37361);
nand U38659 (N_38659,N_36038,N_36525);
nor U38660 (N_38660,N_37506,N_37242);
or U38661 (N_38661,N_37481,N_37034);
xnor U38662 (N_38662,N_37985,N_37838);
and U38663 (N_38663,N_37761,N_36287);
xnor U38664 (N_38664,N_36822,N_36542);
xor U38665 (N_38665,N_36934,N_37158);
or U38666 (N_38666,N_37533,N_36601);
nor U38667 (N_38667,N_37414,N_36123);
nand U38668 (N_38668,N_37886,N_37454);
xor U38669 (N_38669,N_37251,N_36075);
nor U38670 (N_38670,N_37711,N_37543);
nand U38671 (N_38671,N_37112,N_37461);
xnor U38672 (N_38672,N_37995,N_36494);
or U38673 (N_38673,N_37978,N_36160);
xnor U38674 (N_38674,N_36391,N_37979);
and U38675 (N_38675,N_37146,N_37510);
or U38676 (N_38676,N_36857,N_37073);
nor U38677 (N_38677,N_36911,N_36077);
nor U38678 (N_38678,N_36887,N_37943);
nor U38679 (N_38679,N_36344,N_37340);
and U38680 (N_38680,N_37987,N_36215);
xor U38681 (N_38681,N_36114,N_36448);
xnor U38682 (N_38682,N_37437,N_36044);
or U38683 (N_38683,N_37446,N_37008);
and U38684 (N_38684,N_36499,N_36703);
nand U38685 (N_38685,N_37397,N_36649);
nand U38686 (N_38686,N_37601,N_37956);
nand U38687 (N_38687,N_36550,N_37549);
nand U38688 (N_38688,N_37652,N_36120);
nand U38689 (N_38689,N_36006,N_37082);
nor U38690 (N_38690,N_36852,N_37746);
and U38691 (N_38691,N_37074,N_36744);
nand U38692 (N_38692,N_37942,N_37435);
and U38693 (N_38693,N_37100,N_37459);
xnor U38694 (N_38694,N_37890,N_36866);
nor U38695 (N_38695,N_36101,N_36717);
or U38696 (N_38696,N_37647,N_36577);
or U38697 (N_38697,N_36959,N_36192);
nand U38698 (N_38698,N_37285,N_37343);
xnor U38699 (N_38699,N_37708,N_36517);
nand U38700 (N_38700,N_37275,N_37781);
and U38701 (N_38701,N_37794,N_36768);
and U38702 (N_38702,N_36666,N_36325);
and U38703 (N_38703,N_37669,N_36907);
and U38704 (N_38704,N_36553,N_37927);
or U38705 (N_38705,N_37248,N_36214);
and U38706 (N_38706,N_37900,N_36353);
and U38707 (N_38707,N_36165,N_36690);
or U38708 (N_38708,N_37829,N_36877);
and U38709 (N_38709,N_36849,N_36425);
or U38710 (N_38710,N_36368,N_37803);
or U38711 (N_38711,N_36051,N_36962);
or U38712 (N_38712,N_37225,N_37899);
nor U38713 (N_38713,N_36656,N_36386);
nand U38714 (N_38714,N_36695,N_37463);
xnor U38715 (N_38715,N_37826,N_37213);
nand U38716 (N_38716,N_36567,N_37870);
nand U38717 (N_38717,N_36163,N_37064);
nand U38718 (N_38718,N_37566,N_36471);
and U38719 (N_38719,N_37541,N_36177);
and U38720 (N_38720,N_37269,N_37181);
xor U38721 (N_38721,N_37609,N_37778);
xnor U38722 (N_38722,N_37186,N_37049);
nand U38723 (N_38723,N_37440,N_36065);
nor U38724 (N_38724,N_37048,N_37237);
nand U38725 (N_38725,N_37889,N_37115);
nor U38726 (N_38726,N_37102,N_36740);
and U38727 (N_38727,N_36606,N_37359);
nor U38728 (N_38728,N_36364,N_37024);
nand U38729 (N_38729,N_37001,N_37764);
nor U38730 (N_38730,N_37347,N_37646);
or U38731 (N_38731,N_37358,N_36630);
xor U38732 (N_38732,N_36597,N_37700);
or U38733 (N_38733,N_36008,N_36562);
nor U38734 (N_38734,N_37688,N_36472);
xnor U38735 (N_38735,N_36711,N_37483);
and U38736 (N_38736,N_36896,N_36025);
nor U38737 (N_38737,N_37704,N_36225);
and U38738 (N_38738,N_37012,N_36579);
nand U38739 (N_38739,N_36923,N_36808);
and U38740 (N_38740,N_37648,N_36882);
and U38741 (N_38741,N_37294,N_37501);
and U38742 (N_38742,N_36179,N_36883);
xnor U38743 (N_38743,N_37190,N_36071);
nor U38744 (N_38744,N_36990,N_37607);
nand U38745 (N_38745,N_37744,N_36387);
and U38746 (N_38746,N_36338,N_36085);
xnor U38747 (N_38747,N_37390,N_37975);
or U38748 (N_38748,N_36027,N_36791);
or U38749 (N_38749,N_36076,N_36658);
xnor U38750 (N_38750,N_37321,N_36599);
and U38751 (N_38751,N_36574,N_37673);
nand U38752 (N_38752,N_37800,N_36878);
or U38753 (N_38753,N_37715,N_37587);
nand U38754 (N_38754,N_37698,N_37106);
or U38755 (N_38755,N_37716,N_37252);
nand U38756 (N_38756,N_36376,N_36392);
nor U38757 (N_38757,N_36014,N_36447);
and U38758 (N_38758,N_37393,N_37539);
nor U38759 (N_38759,N_37872,N_37679);
nand U38760 (N_38760,N_37958,N_36254);
nor U38761 (N_38761,N_37069,N_36957);
or U38762 (N_38762,N_37143,N_36532);
and U38763 (N_38763,N_37399,N_37011);
nand U38764 (N_38764,N_37954,N_36996);
xnor U38765 (N_38765,N_36034,N_36892);
xor U38766 (N_38766,N_37320,N_36538);
or U38767 (N_38767,N_37370,N_36588);
xnor U38768 (N_38768,N_36591,N_36634);
or U38769 (N_38769,N_37809,N_37431);
and U38770 (N_38770,N_37965,N_37002);
xnor U38771 (N_38771,N_36501,N_36939);
nor U38772 (N_38772,N_37212,N_36373);
nand U38773 (N_38773,N_37820,N_36821);
xor U38774 (N_38774,N_36248,N_36607);
nor U38775 (N_38775,N_37265,N_37658);
nor U38776 (N_38776,N_37013,N_37193);
and U38777 (N_38777,N_36398,N_36954);
nand U38778 (N_38778,N_37138,N_37505);
and U38779 (N_38779,N_37174,N_37532);
nand U38780 (N_38780,N_36554,N_37683);
nor U38781 (N_38781,N_37597,N_37401);
xnor U38782 (N_38782,N_37479,N_36375);
nand U38783 (N_38783,N_36917,N_37754);
nor U38784 (N_38784,N_36669,N_36786);
and U38785 (N_38785,N_37877,N_37606);
nand U38786 (N_38786,N_37959,N_36929);
xnor U38787 (N_38787,N_36382,N_36102);
nand U38788 (N_38788,N_36555,N_37684);
and U38789 (N_38789,N_36482,N_36485);
nand U38790 (N_38790,N_36843,N_36516);
nor U38791 (N_38791,N_36332,N_37219);
xor U38792 (N_38792,N_37351,N_37039);
xnor U38793 (N_38793,N_37327,N_37235);
or U38794 (N_38794,N_37433,N_36660);
xnor U38795 (N_38795,N_37279,N_36620);
nor U38796 (N_38796,N_36937,N_37963);
or U38797 (N_38797,N_36417,N_37967);
nand U38798 (N_38798,N_36436,N_36054);
nand U38799 (N_38799,N_36372,N_37790);
xor U38800 (N_38800,N_36328,N_36519);
nand U38801 (N_38801,N_36737,N_37418);
xor U38802 (N_38802,N_36837,N_36348);
and U38803 (N_38803,N_36224,N_36366);
and U38804 (N_38804,N_36909,N_36444);
or U38805 (N_38805,N_36309,N_37742);
or U38806 (N_38806,N_36675,N_36033);
xor U38807 (N_38807,N_37515,N_36946);
and U38808 (N_38808,N_36116,N_37060);
nand U38809 (N_38809,N_37421,N_36750);
xnor U38810 (N_38810,N_37699,N_37055);
nand U38811 (N_38811,N_37140,N_36018);
nand U38812 (N_38812,N_37353,N_37333);
nand U38813 (N_38813,N_37763,N_36424);
nor U38814 (N_38814,N_37345,N_37288);
nor U38815 (N_38815,N_37976,N_37266);
and U38816 (N_38816,N_37966,N_37044);
and U38817 (N_38817,N_36395,N_37689);
nor U38818 (N_38818,N_37030,N_37107);
and U38819 (N_38819,N_37919,N_37038);
xnor U38820 (N_38820,N_37376,N_37951);
nand U38821 (N_38821,N_37504,N_37960);
nor U38822 (N_38822,N_37309,N_36688);
nand U38823 (N_38823,N_37923,N_37948);
or U38824 (N_38824,N_37025,N_37268);
xnor U38825 (N_38825,N_37577,N_37910);
nor U38826 (N_38826,N_37144,N_36891);
and U38827 (N_38827,N_37818,N_37602);
and U38828 (N_38828,N_37666,N_37380);
or U38829 (N_38829,N_37866,N_36556);
nor U38830 (N_38830,N_36337,N_36831);
or U38831 (N_38831,N_36064,N_37214);
xor U38832 (N_38832,N_36483,N_37650);
or U38833 (N_38833,N_37455,N_36894);
and U38834 (N_38834,N_37714,N_36237);
or U38835 (N_38835,N_37771,N_37722);
and U38836 (N_38836,N_37262,N_36094);
or U38837 (N_38837,N_36540,N_36058);
nand U38838 (N_38838,N_37901,N_37286);
nor U38839 (N_38839,N_37938,N_37442);
or U38840 (N_38840,N_36411,N_36393);
and U38841 (N_38841,N_37585,N_37564);
and U38842 (N_38842,N_37732,N_37736);
and U38843 (N_38843,N_37817,N_37273);
nand U38844 (N_38844,N_36081,N_36600);
nand U38845 (N_38845,N_37467,N_36576);
nand U38846 (N_38846,N_36693,N_37846);
and U38847 (N_38847,N_37101,N_37806);
nor U38848 (N_38848,N_37250,N_36290);
nand U38849 (N_38849,N_37926,N_36729);
nand U38850 (N_38850,N_36355,N_37993);
xnor U38851 (N_38851,N_36357,N_36665);
xnor U38852 (N_38852,N_37663,N_36799);
and U38853 (N_38853,N_37787,N_37830);
xor U38854 (N_38854,N_36031,N_37046);
nand U38855 (N_38855,N_36433,N_37559);
and U38856 (N_38856,N_37657,N_37865);
nand U38857 (N_38857,N_36706,N_37905);
xor U38858 (N_38858,N_37389,N_36716);
xnor U38859 (N_38859,N_36401,N_37914);
and U38860 (N_38860,N_36263,N_37404);
and U38861 (N_38861,N_37296,N_37415);
and U38862 (N_38862,N_37635,N_37634);
xor U38863 (N_38863,N_37766,N_36055);
and U38864 (N_38864,N_37173,N_37167);
xor U38865 (N_38865,N_37246,N_36865);
and U38866 (N_38866,N_36674,N_36899);
or U38867 (N_38867,N_36323,N_36066);
xnor U38868 (N_38868,N_36340,N_36624);
nor U38869 (N_38869,N_37417,N_37368);
nand U38870 (N_38870,N_37491,N_37051);
and U38871 (N_38871,N_36189,N_37949);
or U38872 (N_38872,N_36473,N_37864);
or U38873 (N_38873,N_37018,N_36342);
or U38874 (N_38874,N_37727,N_37042);
nand U38875 (N_38875,N_36560,N_37070);
xnor U38876 (N_38876,N_37443,N_36311);
xnor U38877 (N_38877,N_37398,N_36932);
xnor U38878 (N_38878,N_37122,N_36241);
nand U38879 (N_38879,N_37124,N_36521);
nor U38880 (N_38880,N_37356,N_36915);
and U38881 (N_38881,N_37693,N_36848);
xnor U38882 (N_38882,N_37152,N_36053);
nor U38883 (N_38883,N_37202,N_36023);
nand U38884 (N_38884,N_37036,N_37098);
nor U38885 (N_38885,N_37542,N_37168);
nand U38886 (N_38886,N_37033,N_36610);
nor U38887 (N_38887,N_37977,N_36136);
nor U38888 (N_38888,N_37750,N_36187);
xnor U38889 (N_38889,N_36128,N_36133);
nor U38890 (N_38890,N_36269,N_36981);
xnor U38891 (N_38891,N_36713,N_37365);
nor U38892 (N_38892,N_37880,N_36639);
nor U38893 (N_38893,N_37453,N_37793);
xor U38894 (N_38894,N_36315,N_36304);
and U38895 (N_38895,N_37438,N_37655);
or U38896 (N_38896,N_37382,N_36708);
xnor U38897 (N_38897,N_37425,N_36441);
nand U38898 (N_38898,N_37482,N_37119);
xnor U38899 (N_38899,N_36080,N_37386);
nor U38900 (N_38900,N_36741,N_37117);
xor U38901 (N_38901,N_37668,N_37334);
or U38902 (N_38902,N_37653,N_37405);
or U38903 (N_38903,N_37406,N_36119);
nor U38904 (N_38904,N_36288,N_36231);
nor U38905 (N_38905,N_36804,N_36047);
or U38906 (N_38906,N_37775,N_36970);
xor U38907 (N_38907,N_36200,N_37071);
xor U38908 (N_38908,N_37104,N_36629);
nor U38909 (N_38909,N_36859,N_37573);
xnor U38910 (N_38910,N_36793,N_37694);
and U38911 (N_38911,N_36566,N_37522);
nand U38912 (N_38912,N_36059,N_36736);
xnor U38913 (N_38913,N_37555,N_36343);
nor U38914 (N_38914,N_37991,N_37994);
or U38915 (N_38915,N_36274,N_37413);
nand U38916 (N_38916,N_37093,N_37671);
nand U38917 (N_38917,N_37677,N_37230);
xor U38918 (N_38918,N_37660,N_36271);
xnor U38919 (N_38919,N_36506,N_36927);
nand U38920 (N_38920,N_37276,N_37508);
nand U38921 (N_38921,N_36715,N_37527);
xor U38922 (N_38922,N_37065,N_36605);
nand U38923 (N_38923,N_37950,N_36977);
or U38924 (N_38924,N_37072,N_36596);
nand U38925 (N_38925,N_36024,N_37058);
and U38926 (N_38926,N_37194,N_37594);
xor U38927 (N_38927,N_36834,N_37470);
nand U38928 (N_38928,N_36888,N_36196);
or U38929 (N_38929,N_37558,N_37078);
nand U38930 (N_38930,N_37354,N_36861);
nand U38931 (N_38931,N_37892,N_37725);
nand U38932 (N_38932,N_36739,N_36112);
xnor U38933 (N_38933,N_37350,N_37247);
nor U38934 (N_38934,N_36585,N_37633);
and U38935 (N_38935,N_36335,N_37620);
nor U38936 (N_38936,N_37521,N_37915);
and U38937 (N_38937,N_37623,N_37131);
nand U38938 (N_38938,N_37921,N_36570);
and U38939 (N_38939,N_37313,N_37519);
nor U38940 (N_38940,N_36680,N_36951);
nor U38941 (N_38941,N_36734,N_37641);
nand U38942 (N_38942,N_37080,N_37364);
and U38943 (N_38943,N_36612,N_36414);
nor U38944 (N_38944,N_37681,N_36318);
nand U38945 (N_38945,N_37336,N_36171);
nor U38946 (N_38946,N_36267,N_36670);
nor U38947 (N_38947,N_36019,N_36097);
and U38948 (N_38948,N_36063,N_37163);
and U38949 (N_38949,N_36543,N_36314);
and U38950 (N_38950,N_36126,N_36844);
and U38951 (N_38951,N_37622,N_37840);
nand U38952 (N_38952,N_36796,N_36110);
nand U38953 (N_38953,N_37456,N_37209);
nor U38954 (N_38954,N_36370,N_36010);
or U38955 (N_38955,N_37125,N_36618);
or U38956 (N_38956,N_37474,N_37357);
nand U38957 (N_38957,N_37416,N_36089);
xnor U38958 (N_38958,N_36918,N_36067);
nand U38959 (N_38959,N_37706,N_36208);
xor U38960 (N_38960,N_37466,N_37593);
nor U38961 (N_38961,N_36855,N_36078);
xor U38962 (N_38962,N_37502,N_37891);
nor U38963 (N_38963,N_36400,N_37860);
xnor U38964 (N_38964,N_36001,N_36904);
and U38965 (N_38965,N_36988,N_36710);
or U38966 (N_38966,N_37874,N_36061);
xor U38967 (N_38967,N_37894,N_37853);
nor U38968 (N_38968,N_37535,N_37814);
xnor U38969 (N_38969,N_37801,N_36593);
or U38970 (N_38970,N_36637,N_36284);
nand U38971 (N_38971,N_36098,N_37825);
or U38972 (N_38972,N_36478,N_37561);
xnor U38973 (N_38973,N_37859,N_37130);
nand U38974 (N_38974,N_37614,N_36619);
nand U38975 (N_38975,N_36199,N_37565);
or U38976 (N_38976,N_36720,N_37847);
nor U38977 (N_38977,N_36070,N_37278);
and U38978 (N_38978,N_37876,N_36730);
nand U38979 (N_38979,N_36421,N_37841);
nor U38980 (N_38980,N_37743,N_37909);
xor U38981 (N_38981,N_37528,N_36871);
nand U38982 (N_38982,N_37170,N_37068);
xnor U38983 (N_38983,N_37631,N_36334);
xnor U38984 (N_38984,N_37147,N_37315);
nor U38985 (N_38985,N_37245,N_36765);
or U38986 (N_38986,N_37032,N_37674);
and U38987 (N_38987,N_37868,N_37126);
or U38988 (N_38988,N_36650,N_36159);
nand U38989 (N_38989,N_37592,N_37540);
or U38990 (N_38990,N_36028,N_36700);
xnor U38991 (N_38991,N_37420,N_37916);
xor U38992 (N_38992,N_37363,N_37019);
nand U38993 (N_38993,N_36188,N_36879);
nor U38994 (N_38994,N_37856,N_36246);
and U38995 (N_38995,N_37256,N_37427);
nand U38996 (N_38996,N_37342,N_37103);
xnor U38997 (N_38997,N_37913,N_36103);
nor U38998 (N_38998,N_37208,N_37912);
nand U38999 (N_38999,N_36587,N_36709);
and U39000 (N_39000,N_36936,N_37571);
xnor U39001 (N_39001,N_36747,N_37890);
xor U39002 (N_39002,N_36871,N_37849);
or U39003 (N_39003,N_36474,N_36635);
and U39004 (N_39004,N_37691,N_37429);
and U39005 (N_39005,N_37895,N_36201);
or U39006 (N_39006,N_36534,N_36022);
nor U39007 (N_39007,N_37541,N_36720);
xnor U39008 (N_39008,N_36617,N_37525);
and U39009 (N_39009,N_36897,N_36492);
nand U39010 (N_39010,N_36958,N_37239);
nor U39011 (N_39011,N_36024,N_36015);
or U39012 (N_39012,N_37976,N_37555);
and U39013 (N_39013,N_36231,N_36273);
nand U39014 (N_39014,N_36468,N_36499);
or U39015 (N_39015,N_36193,N_37461);
nand U39016 (N_39016,N_36970,N_37818);
and U39017 (N_39017,N_37469,N_36419);
xnor U39018 (N_39018,N_37002,N_36848);
xor U39019 (N_39019,N_37934,N_37444);
xor U39020 (N_39020,N_36566,N_37921);
nand U39021 (N_39021,N_37382,N_36395);
and U39022 (N_39022,N_36068,N_37680);
and U39023 (N_39023,N_37713,N_36239);
xnor U39024 (N_39024,N_36112,N_37004);
and U39025 (N_39025,N_37603,N_36560);
xnor U39026 (N_39026,N_37318,N_36814);
or U39027 (N_39027,N_36946,N_36934);
nor U39028 (N_39028,N_37425,N_37399);
xnor U39029 (N_39029,N_37066,N_36892);
xnor U39030 (N_39030,N_37465,N_37606);
nand U39031 (N_39031,N_36843,N_37567);
nand U39032 (N_39032,N_37161,N_36533);
nor U39033 (N_39033,N_37642,N_37981);
or U39034 (N_39034,N_36241,N_36531);
and U39035 (N_39035,N_37285,N_37355);
and U39036 (N_39036,N_37216,N_36805);
nand U39037 (N_39037,N_37335,N_37614);
xnor U39038 (N_39038,N_37145,N_36107);
xnor U39039 (N_39039,N_37226,N_37410);
nor U39040 (N_39040,N_37991,N_36823);
and U39041 (N_39041,N_36237,N_36780);
and U39042 (N_39042,N_37442,N_36992);
nand U39043 (N_39043,N_37486,N_36665);
nor U39044 (N_39044,N_36214,N_36750);
nand U39045 (N_39045,N_37862,N_37342);
nand U39046 (N_39046,N_37557,N_37330);
nand U39047 (N_39047,N_37923,N_37576);
and U39048 (N_39048,N_36969,N_37479);
nor U39049 (N_39049,N_37561,N_37464);
nor U39050 (N_39050,N_37129,N_36102);
xnor U39051 (N_39051,N_36829,N_37427);
or U39052 (N_39052,N_37138,N_37187);
or U39053 (N_39053,N_37618,N_37387);
or U39054 (N_39054,N_36215,N_37866);
nand U39055 (N_39055,N_37517,N_36271);
xnor U39056 (N_39056,N_36241,N_36867);
nand U39057 (N_39057,N_36385,N_36665);
xor U39058 (N_39058,N_37345,N_37782);
nand U39059 (N_39059,N_36759,N_36996);
nand U39060 (N_39060,N_37316,N_36857);
nor U39061 (N_39061,N_36826,N_36079);
nor U39062 (N_39062,N_37572,N_37054);
and U39063 (N_39063,N_36501,N_37631);
nor U39064 (N_39064,N_37903,N_36041);
nand U39065 (N_39065,N_37147,N_36519);
or U39066 (N_39066,N_37001,N_36624);
or U39067 (N_39067,N_37709,N_37948);
and U39068 (N_39068,N_37936,N_37208);
xor U39069 (N_39069,N_37244,N_37558);
xor U39070 (N_39070,N_36614,N_36054);
xnor U39071 (N_39071,N_36478,N_36993);
or U39072 (N_39072,N_36692,N_36945);
nor U39073 (N_39073,N_37746,N_36954);
nand U39074 (N_39074,N_36735,N_36203);
xor U39075 (N_39075,N_37050,N_36922);
and U39076 (N_39076,N_37979,N_36247);
nor U39077 (N_39077,N_37585,N_37138);
and U39078 (N_39078,N_37024,N_36038);
nor U39079 (N_39079,N_36675,N_36413);
and U39080 (N_39080,N_36066,N_36571);
nand U39081 (N_39081,N_37937,N_37225);
and U39082 (N_39082,N_36459,N_36713);
and U39083 (N_39083,N_37471,N_36995);
or U39084 (N_39084,N_36879,N_36888);
nor U39085 (N_39085,N_37927,N_37502);
and U39086 (N_39086,N_37482,N_37659);
or U39087 (N_39087,N_37962,N_37981);
xnor U39088 (N_39088,N_37973,N_37093);
nand U39089 (N_39089,N_36093,N_36561);
xor U39090 (N_39090,N_37302,N_36238);
xnor U39091 (N_39091,N_37000,N_36491);
nor U39092 (N_39092,N_37008,N_37063);
or U39093 (N_39093,N_36428,N_37907);
and U39094 (N_39094,N_37394,N_37849);
or U39095 (N_39095,N_37795,N_36954);
nand U39096 (N_39096,N_37043,N_37970);
xnor U39097 (N_39097,N_36116,N_37316);
xnor U39098 (N_39098,N_36126,N_37573);
or U39099 (N_39099,N_37121,N_36248);
or U39100 (N_39100,N_36925,N_37054);
nand U39101 (N_39101,N_36828,N_37128);
nand U39102 (N_39102,N_36669,N_36232);
nand U39103 (N_39103,N_36503,N_37828);
and U39104 (N_39104,N_36338,N_36404);
nor U39105 (N_39105,N_37312,N_37573);
and U39106 (N_39106,N_36747,N_36499);
xor U39107 (N_39107,N_37293,N_37143);
nand U39108 (N_39108,N_36114,N_36000);
and U39109 (N_39109,N_37985,N_37372);
xor U39110 (N_39110,N_36549,N_37096);
or U39111 (N_39111,N_36529,N_37244);
nor U39112 (N_39112,N_37654,N_36523);
nor U39113 (N_39113,N_36888,N_37208);
or U39114 (N_39114,N_37730,N_37660);
xnor U39115 (N_39115,N_37167,N_36814);
nand U39116 (N_39116,N_36096,N_36007);
or U39117 (N_39117,N_37664,N_36780);
xnor U39118 (N_39118,N_37735,N_37121);
nor U39119 (N_39119,N_37175,N_36099);
xnor U39120 (N_39120,N_36642,N_37918);
nor U39121 (N_39121,N_36172,N_37061);
and U39122 (N_39122,N_36618,N_37235);
nor U39123 (N_39123,N_36305,N_37394);
or U39124 (N_39124,N_36139,N_36121);
and U39125 (N_39125,N_36528,N_36758);
and U39126 (N_39126,N_37304,N_37551);
nand U39127 (N_39127,N_37022,N_36599);
or U39128 (N_39128,N_36892,N_37377);
xor U39129 (N_39129,N_37056,N_36185);
xnor U39130 (N_39130,N_37566,N_37366);
nand U39131 (N_39131,N_36973,N_37662);
xnor U39132 (N_39132,N_37429,N_36548);
nor U39133 (N_39133,N_36323,N_37668);
and U39134 (N_39134,N_37419,N_36812);
and U39135 (N_39135,N_36389,N_36073);
nor U39136 (N_39136,N_37518,N_37712);
nand U39137 (N_39137,N_37908,N_36135);
or U39138 (N_39138,N_36974,N_36454);
and U39139 (N_39139,N_36980,N_37004);
xor U39140 (N_39140,N_36750,N_37390);
nand U39141 (N_39141,N_37555,N_37301);
xnor U39142 (N_39142,N_36230,N_37131);
or U39143 (N_39143,N_37002,N_37338);
xnor U39144 (N_39144,N_37993,N_36165);
or U39145 (N_39145,N_36924,N_36284);
or U39146 (N_39146,N_37563,N_37197);
nor U39147 (N_39147,N_37943,N_37952);
nand U39148 (N_39148,N_36315,N_36132);
or U39149 (N_39149,N_37765,N_37953);
xnor U39150 (N_39150,N_37560,N_36268);
and U39151 (N_39151,N_36005,N_36135);
nand U39152 (N_39152,N_37192,N_36474);
and U39153 (N_39153,N_36476,N_37240);
nor U39154 (N_39154,N_36885,N_36173);
xor U39155 (N_39155,N_37588,N_36030);
and U39156 (N_39156,N_36347,N_36640);
or U39157 (N_39157,N_36225,N_36887);
xor U39158 (N_39158,N_37047,N_37041);
nor U39159 (N_39159,N_37743,N_37842);
nand U39160 (N_39160,N_36871,N_37541);
nor U39161 (N_39161,N_36531,N_37116);
nor U39162 (N_39162,N_37929,N_36193);
xor U39163 (N_39163,N_36988,N_36769);
nor U39164 (N_39164,N_37469,N_37562);
xor U39165 (N_39165,N_36688,N_37556);
nand U39166 (N_39166,N_36710,N_37177);
nand U39167 (N_39167,N_37824,N_36685);
nor U39168 (N_39168,N_37869,N_36209);
nand U39169 (N_39169,N_36060,N_36150);
and U39170 (N_39170,N_36141,N_37171);
xnor U39171 (N_39171,N_37182,N_36276);
and U39172 (N_39172,N_37421,N_37728);
nor U39173 (N_39173,N_37927,N_36264);
xnor U39174 (N_39174,N_37416,N_36252);
xor U39175 (N_39175,N_36246,N_36247);
nand U39176 (N_39176,N_37242,N_37864);
and U39177 (N_39177,N_36259,N_37930);
and U39178 (N_39178,N_36131,N_37086);
and U39179 (N_39179,N_36509,N_36484);
nor U39180 (N_39180,N_37082,N_37075);
or U39181 (N_39181,N_36113,N_37875);
xor U39182 (N_39182,N_37860,N_37272);
nand U39183 (N_39183,N_37825,N_37457);
and U39184 (N_39184,N_36623,N_37293);
nor U39185 (N_39185,N_37898,N_37232);
xor U39186 (N_39186,N_36075,N_36003);
xor U39187 (N_39187,N_36743,N_36172);
nand U39188 (N_39188,N_37444,N_36198);
xor U39189 (N_39189,N_37210,N_37086);
nand U39190 (N_39190,N_36285,N_36378);
and U39191 (N_39191,N_36802,N_36893);
and U39192 (N_39192,N_36090,N_36055);
or U39193 (N_39193,N_37681,N_37804);
xnor U39194 (N_39194,N_37652,N_36159);
nand U39195 (N_39195,N_37666,N_37932);
and U39196 (N_39196,N_37116,N_37443);
xor U39197 (N_39197,N_36577,N_36244);
xor U39198 (N_39198,N_36311,N_36064);
and U39199 (N_39199,N_36144,N_37677);
nand U39200 (N_39200,N_36158,N_37154);
or U39201 (N_39201,N_37286,N_36678);
and U39202 (N_39202,N_36723,N_36714);
or U39203 (N_39203,N_37932,N_36717);
or U39204 (N_39204,N_36407,N_37562);
xnor U39205 (N_39205,N_36812,N_36491);
and U39206 (N_39206,N_36301,N_36169);
nor U39207 (N_39207,N_37755,N_36306);
nor U39208 (N_39208,N_37585,N_36596);
and U39209 (N_39209,N_37440,N_36414);
and U39210 (N_39210,N_36023,N_36053);
or U39211 (N_39211,N_36539,N_37152);
or U39212 (N_39212,N_36036,N_36577);
xor U39213 (N_39213,N_36859,N_37275);
nand U39214 (N_39214,N_36057,N_36227);
and U39215 (N_39215,N_37504,N_36261);
and U39216 (N_39216,N_36800,N_36428);
nor U39217 (N_39217,N_37652,N_37083);
and U39218 (N_39218,N_37273,N_37982);
or U39219 (N_39219,N_36228,N_36234);
nand U39220 (N_39220,N_36998,N_36037);
or U39221 (N_39221,N_37085,N_37354);
nand U39222 (N_39222,N_36979,N_37253);
xor U39223 (N_39223,N_36265,N_36899);
xnor U39224 (N_39224,N_36688,N_37318);
and U39225 (N_39225,N_37000,N_36837);
and U39226 (N_39226,N_37823,N_36237);
or U39227 (N_39227,N_37243,N_37656);
xor U39228 (N_39228,N_36251,N_37471);
nor U39229 (N_39229,N_37172,N_37254);
xnor U39230 (N_39230,N_37009,N_36527);
nor U39231 (N_39231,N_36934,N_37489);
or U39232 (N_39232,N_36415,N_36372);
or U39233 (N_39233,N_36671,N_37009);
nor U39234 (N_39234,N_36703,N_36890);
xor U39235 (N_39235,N_37930,N_37699);
nand U39236 (N_39236,N_37176,N_36537);
and U39237 (N_39237,N_37118,N_37829);
and U39238 (N_39238,N_37667,N_36655);
nand U39239 (N_39239,N_37387,N_37990);
and U39240 (N_39240,N_36462,N_37638);
nand U39241 (N_39241,N_36119,N_36647);
and U39242 (N_39242,N_37566,N_36902);
or U39243 (N_39243,N_37539,N_36407);
nor U39244 (N_39244,N_36003,N_36484);
and U39245 (N_39245,N_37221,N_36581);
and U39246 (N_39246,N_37537,N_36054);
and U39247 (N_39247,N_37636,N_36356);
and U39248 (N_39248,N_36917,N_37233);
xor U39249 (N_39249,N_37822,N_36380);
or U39250 (N_39250,N_36708,N_36143);
or U39251 (N_39251,N_36731,N_37229);
xor U39252 (N_39252,N_36274,N_37908);
nor U39253 (N_39253,N_37546,N_37387);
xor U39254 (N_39254,N_37309,N_37699);
or U39255 (N_39255,N_37156,N_36358);
xnor U39256 (N_39256,N_36613,N_36967);
nand U39257 (N_39257,N_36945,N_37364);
xor U39258 (N_39258,N_36352,N_36817);
xnor U39259 (N_39259,N_36315,N_37829);
or U39260 (N_39260,N_36107,N_36486);
nor U39261 (N_39261,N_36486,N_37966);
xor U39262 (N_39262,N_36257,N_36045);
xnor U39263 (N_39263,N_37874,N_37608);
or U39264 (N_39264,N_37591,N_37897);
and U39265 (N_39265,N_36432,N_36562);
xnor U39266 (N_39266,N_36582,N_37628);
nand U39267 (N_39267,N_37098,N_37731);
xor U39268 (N_39268,N_37940,N_37407);
xnor U39269 (N_39269,N_37925,N_36419);
or U39270 (N_39270,N_37952,N_36410);
nor U39271 (N_39271,N_37088,N_36594);
or U39272 (N_39272,N_36618,N_36672);
nand U39273 (N_39273,N_36141,N_37029);
nor U39274 (N_39274,N_36486,N_36254);
xor U39275 (N_39275,N_36923,N_37589);
or U39276 (N_39276,N_37105,N_37872);
or U39277 (N_39277,N_36889,N_37867);
nor U39278 (N_39278,N_36571,N_36070);
nor U39279 (N_39279,N_36754,N_37246);
and U39280 (N_39280,N_36882,N_37824);
nand U39281 (N_39281,N_37563,N_36697);
xnor U39282 (N_39282,N_36878,N_36365);
or U39283 (N_39283,N_36907,N_36215);
nand U39284 (N_39284,N_36694,N_36483);
nor U39285 (N_39285,N_36777,N_37499);
nand U39286 (N_39286,N_36036,N_36070);
nor U39287 (N_39287,N_36175,N_37048);
xor U39288 (N_39288,N_36566,N_36490);
or U39289 (N_39289,N_36370,N_37142);
nor U39290 (N_39290,N_36054,N_37885);
xor U39291 (N_39291,N_37152,N_36655);
nand U39292 (N_39292,N_36498,N_36444);
nor U39293 (N_39293,N_37699,N_36581);
nor U39294 (N_39294,N_37200,N_36193);
or U39295 (N_39295,N_37078,N_36353);
xor U39296 (N_39296,N_37462,N_36935);
or U39297 (N_39297,N_37139,N_37942);
nor U39298 (N_39298,N_37799,N_37281);
nor U39299 (N_39299,N_37263,N_37162);
xor U39300 (N_39300,N_37748,N_36494);
xnor U39301 (N_39301,N_36404,N_36671);
xnor U39302 (N_39302,N_37167,N_36272);
and U39303 (N_39303,N_37234,N_36133);
nor U39304 (N_39304,N_37496,N_36142);
nand U39305 (N_39305,N_37455,N_37496);
xnor U39306 (N_39306,N_36089,N_36710);
nor U39307 (N_39307,N_36676,N_37227);
nor U39308 (N_39308,N_36255,N_36343);
and U39309 (N_39309,N_37251,N_36317);
xnor U39310 (N_39310,N_36686,N_37797);
nand U39311 (N_39311,N_36577,N_37789);
nand U39312 (N_39312,N_36165,N_36198);
xnor U39313 (N_39313,N_37633,N_36063);
or U39314 (N_39314,N_37476,N_36319);
nand U39315 (N_39315,N_36122,N_37167);
nor U39316 (N_39316,N_36458,N_36275);
and U39317 (N_39317,N_37734,N_37439);
xor U39318 (N_39318,N_37616,N_36212);
nand U39319 (N_39319,N_37687,N_37747);
nor U39320 (N_39320,N_37230,N_36493);
or U39321 (N_39321,N_36770,N_37312);
or U39322 (N_39322,N_37498,N_36443);
and U39323 (N_39323,N_37703,N_36760);
nand U39324 (N_39324,N_37954,N_36156);
and U39325 (N_39325,N_37609,N_37535);
xnor U39326 (N_39326,N_37358,N_37413);
nand U39327 (N_39327,N_37190,N_36215);
nor U39328 (N_39328,N_36825,N_36750);
and U39329 (N_39329,N_36506,N_36122);
nand U39330 (N_39330,N_37858,N_36781);
or U39331 (N_39331,N_37292,N_37655);
nor U39332 (N_39332,N_36214,N_36037);
nor U39333 (N_39333,N_36318,N_36337);
nand U39334 (N_39334,N_36873,N_36828);
or U39335 (N_39335,N_37989,N_36933);
nand U39336 (N_39336,N_37351,N_37825);
nand U39337 (N_39337,N_36246,N_36224);
or U39338 (N_39338,N_37053,N_36393);
xnor U39339 (N_39339,N_36700,N_36262);
and U39340 (N_39340,N_36688,N_36114);
nor U39341 (N_39341,N_37048,N_37514);
xor U39342 (N_39342,N_36730,N_36298);
or U39343 (N_39343,N_36612,N_37135);
and U39344 (N_39344,N_36328,N_37194);
and U39345 (N_39345,N_36238,N_37886);
xnor U39346 (N_39346,N_36761,N_37279);
nand U39347 (N_39347,N_37002,N_37047);
and U39348 (N_39348,N_37054,N_37287);
xor U39349 (N_39349,N_36586,N_37871);
or U39350 (N_39350,N_36036,N_37539);
or U39351 (N_39351,N_37701,N_36700);
and U39352 (N_39352,N_37827,N_36629);
and U39353 (N_39353,N_36127,N_36454);
and U39354 (N_39354,N_37176,N_37834);
and U39355 (N_39355,N_37524,N_37925);
and U39356 (N_39356,N_37492,N_37291);
nand U39357 (N_39357,N_37222,N_36276);
or U39358 (N_39358,N_37254,N_37866);
and U39359 (N_39359,N_36564,N_37985);
or U39360 (N_39360,N_36715,N_37914);
nor U39361 (N_39361,N_37314,N_36227);
nand U39362 (N_39362,N_36591,N_36156);
nand U39363 (N_39363,N_37107,N_37773);
nor U39364 (N_39364,N_36960,N_36608);
xor U39365 (N_39365,N_36518,N_36907);
and U39366 (N_39366,N_36420,N_37384);
or U39367 (N_39367,N_37219,N_36622);
and U39368 (N_39368,N_36223,N_37237);
xor U39369 (N_39369,N_37716,N_36577);
and U39370 (N_39370,N_37361,N_36969);
or U39371 (N_39371,N_37990,N_36952);
nor U39372 (N_39372,N_36136,N_37722);
xnor U39373 (N_39373,N_36898,N_36847);
nand U39374 (N_39374,N_36668,N_36814);
nor U39375 (N_39375,N_37366,N_37879);
xor U39376 (N_39376,N_36098,N_36352);
nand U39377 (N_39377,N_37481,N_37645);
and U39378 (N_39378,N_36559,N_36900);
and U39379 (N_39379,N_36034,N_36440);
nor U39380 (N_39380,N_36477,N_36425);
and U39381 (N_39381,N_36733,N_36992);
xnor U39382 (N_39382,N_36109,N_36060);
xnor U39383 (N_39383,N_37457,N_36088);
nand U39384 (N_39384,N_36783,N_36234);
xor U39385 (N_39385,N_37016,N_37458);
xnor U39386 (N_39386,N_36001,N_36774);
nor U39387 (N_39387,N_36845,N_36531);
xnor U39388 (N_39388,N_36057,N_36426);
nor U39389 (N_39389,N_36684,N_36491);
nor U39390 (N_39390,N_37713,N_36867);
nand U39391 (N_39391,N_36901,N_36999);
or U39392 (N_39392,N_36666,N_36883);
nor U39393 (N_39393,N_36700,N_36458);
or U39394 (N_39394,N_36005,N_36351);
nand U39395 (N_39395,N_37674,N_37083);
nor U39396 (N_39396,N_36341,N_37876);
xor U39397 (N_39397,N_36139,N_37682);
and U39398 (N_39398,N_37293,N_36076);
nor U39399 (N_39399,N_36011,N_36710);
nand U39400 (N_39400,N_36607,N_37477);
nor U39401 (N_39401,N_36316,N_37830);
or U39402 (N_39402,N_36342,N_37268);
nand U39403 (N_39403,N_36129,N_36589);
nand U39404 (N_39404,N_37185,N_37466);
nand U39405 (N_39405,N_36988,N_37442);
and U39406 (N_39406,N_37904,N_37617);
xnor U39407 (N_39407,N_37022,N_36423);
nand U39408 (N_39408,N_37598,N_37793);
nor U39409 (N_39409,N_36420,N_37577);
nand U39410 (N_39410,N_36401,N_36733);
or U39411 (N_39411,N_37654,N_36314);
xor U39412 (N_39412,N_37549,N_36148);
or U39413 (N_39413,N_37356,N_37239);
nor U39414 (N_39414,N_37814,N_36199);
or U39415 (N_39415,N_37521,N_36416);
xor U39416 (N_39416,N_36640,N_37360);
or U39417 (N_39417,N_37846,N_37113);
or U39418 (N_39418,N_37795,N_36406);
and U39419 (N_39419,N_37042,N_37883);
xor U39420 (N_39420,N_36378,N_36592);
nand U39421 (N_39421,N_37853,N_37008);
xor U39422 (N_39422,N_37742,N_37687);
xnor U39423 (N_39423,N_36881,N_37259);
nor U39424 (N_39424,N_36004,N_36495);
nand U39425 (N_39425,N_37746,N_36030);
xor U39426 (N_39426,N_37847,N_36335);
and U39427 (N_39427,N_37071,N_37677);
nand U39428 (N_39428,N_36759,N_37449);
nor U39429 (N_39429,N_37731,N_37083);
nor U39430 (N_39430,N_36387,N_37332);
nand U39431 (N_39431,N_37054,N_37721);
nor U39432 (N_39432,N_36641,N_37281);
and U39433 (N_39433,N_37645,N_37701);
nor U39434 (N_39434,N_37107,N_37558);
or U39435 (N_39435,N_37768,N_36768);
or U39436 (N_39436,N_36113,N_36512);
or U39437 (N_39437,N_36018,N_36100);
nand U39438 (N_39438,N_36758,N_36710);
nand U39439 (N_39439,N_36536,N_37605);
and U39440 (N_39440,N_36787,N_36105);
nand U39441 (N_39441,N_37827,N_37154);
xor U39442 (N_39442,N_37094,N_37849);
or U39443 (N_39443,N_36116,N_37784);
xnor U39444 (N_39444,N_36261,N_37782);
xor U39445 (N_39445,N_36490,N_36540);
xor U39446 (N_39446,N_37479,N_36803);
xor U39447 (N_39447,N_36296,N_36321);
and U39448 (N_39448,N_37584,N_36833);
and U39449 (N_39449,N_36012,N_37521);
and U39450 (N_39450,N_36220,N_36201);
xor U39451 (N_39451,N_37875,N_36841);
and U39452 (N_39452,N_36351,N_36170);
or U39453 (N_39453,N_37458,N_36197);
xnor U39454 (N_39454,N_36094,N_36386);
or U39455 (N_39455,N_37410,N_36994);
nor U39456 (N_39456,N_37268,N_37020);
nor U39457 (N_39457,N_36606,N_36830);
and U39458 (N_39458,N_37950,N_37139);
or U39459 (N_39459,N_36439,N_36168);
xnor U39460 (N_39460,N_37487,N_36926);
nor U39461 (N_39461,N_36645,N_36624);
xor U39462 (N_39462,N_37608,N_37947);
nor U39463 (N_39463,N_37531,N_36616);
and U39464 (N_39464,N_36310,N_36082);
or U39465 (N_39465,N_37191,N_36032);
xnor U39466 (N_39466,N_36714,N_37810);
nor U39467 (N_39467,N_36617,N_36067);
or U39468 (N_39468,N_36491,N_36135);
nor U39469 (N_39469,N_37712,N_36961);
or U39470 (N_39470,N_36682,N_37192);
or U39471 (N_39471,N_37698,N_37786);
or U39472 (N_39472,N_36932,N_37687);
nor U39473 (N_39473,N_37880,N_37700);
nor U39474 (N_39474,N_36757,N_36776);
nand U39475 (N_39475,N_36506,N_36778);
nand U39476 (N_39476,N_37872,N_36421);
or U39477 (N_39477,N_37889,N_36906);
nor U39478 (N_39478,N_37309,N_37861);
xor U39479 (N_39479,N_37371,N_36239);
nand U39480 (N_39480,N_36003,N_36483);
nor U39481 (N_39481,N_36859,N_36645);
or U39482 (N_39482,N_36079,N_37359);
or U39483 (N_39483,N_36501,N_37861);
or U39484 (N_39484,N_36803,N_37813);
xnor U39485 (N_39485,N_36987,N_36906);
nor U39486 (N_39486,N_36363,N_36157);
or U39487 (N_39487,N_36367,N_37016);
and U39488 (N_39488,N_36462,N_37199);
and U39489 (N_39489,N_37428,N_36270);
and U39490 (N_39490,N_36242,N_37780);
or U39491 (N_39491,N_36495,N_36196);
xnor U39492 (N_39492,N_37116,N_36989);
nand U39493 (N_39493,N_36155,N_37138);
and U39494 (N_39494,N_36608,N_37294);
nor U39495 (N_39495,N_36070,N_36396);
nor U39496 (N_39496,N_36222,N_37922);
or U39497 (N_39497,N_36702,N_37202);
nand U39498 (N_39498,N_37179,N_37293);
or U39499 (N_39499,N_36639,N_37336);
nor U39500 (N_39500,N_36983,N_36054);
or U39501 (N_39501,N_36778,N_37179);
and U39502 (N_39502,N_36710,N_36026);
or U39503 (N_39503,N_36226,N_37635);
and U39504 (N_39504,N_37895,N_37741);
and U39505 (N_39505,N_36265,N_36313);
xor U39506 (N_39506,N_36392,N_37720);
and U39507 (N_39507,N_36510,N_36700);
nand U39508 (N_39508,N_36858,N_36009);
nand U39509 (N_39509,N_37382,N_37701);
xor U39510 (N_39510,N_36548,N_36990);
nor U39511 (N_39511,N_36032,N_37341);
nor U39512 (N_39512,N_36257,N_36832);
nor U39513 (N_39513,N_36654,N_37737);
xor U39514 (N_39514,N_37280,N_37847);
nor U39515 (N_39515,N_36740,N_37248);
and U39516 (N_39516,N_37101,N_37536);
xnor U39517 (N_39517,N_37311,N_36996);
nor U39518 (N_39518,N_36077,N_37312);
xnor U39519 (N_39519,N_37044,N_37294);
or U39520 (N_39520,N_36834,N_36972);
or U39521 (N_39521,N_37821,N_36199);
nand U39522 (N_39522,N_36361,N_36254);
or U39523 (N_39523,N_37830,N_37473);
and U39524 (N_39524,N_36383,N_36117);
and U39525 (N_39525,N_36258,N_36118);
and U39526 (N_39526,N_36858,N_36341);
xor U39527 (N_39527,N_36813,N_37243);
xor U39528 (N_39528,N_36066,N_37263);
nor U39529 (N_39529,N_36263,N_36465);
nor U39530 (N_39530,N_37880,N_37004);
nor U39531 (N_39531,N_37781,N_37084);
and U39532 (N_39532,N_36324,N_37439);
or U39533 (N_39533,N_36982,N_37153);
xor U39534 (N_39534,N_37356,N_37923);
and U39535 (N_39535,N_37001,N_37970);
xor U39536 (N_39536,N_36567,N_36918);
xnor U39537 (N_39537,N_37659,N_37069);
and U39538 (N_39538,N_37132,N_36256);
or U39539 (N_39539,N_36390,N_36324);
and U39540 (N_39540,N_36661,N_36644);
or U39541 (N_39541,N_36936,N_37627);
nor U39542 (N_39542,N_36901,N_37916);
or U39543 (N_39543,N_36474,N_36828);
or U39544 (N_39544,N_36366,N_37226);
xnor U39545 (N_39545,N_36382,N_36510);
and U39546 (N_39546,N_36503,N_37071);
and U39547 (N_39547,N_36000,N_37153);
and U39548 (N_39548,N_36362,N_37343);
and U39549 (N_39549,N_37071,N_37860);
nor U39550 (N_39550,N_37267,N_37555);
and U39551 (N_39551,N_36936,N_37132);
and U39552 (N_39552,N_36604,N_36396);
and U39553 (N_39553,N_37675,N_36330);
or U39554 (N_39554,N_37844,N_37863);
nand U39555 (N_39555,N_37091,N_37252);
nand U39556 (N_39556,N_37317,N_37901);
xor U39557 (N_39557,N_37472,N_37580);
xnor U39558 (N_39558,N_37984,N_37017);
and U39559 (N_39559,N_36018,N_37955);
xnor U39560 (N_39560,N_37265,N_36731);
and U39561 (N_39561,N_36618,N_37593);
or U39562 (N_39562,N_37531,N_37046);
xor U39563 (N_39563,N_36101,N_37435);
nor U39564 (N_39564,N_36836,N_37726);
or U39565 (N_39565,N_37562,N_37318);
or U39566 (N_39566,N_36746,N_36653);
xnor U39567 (N_39567,N_36967,N_36383);
nand U39568 (N_39568,N_36169,N_37057);
or U39569 (N_39569,N_36233,N_36370);
and U39570 (N_39570,N_37136,N_36994);
xor U39571 (N_39571,N_37729,N_37706);
nor U39572 (N_39572,N_36680,N_37970);
or U39573 (N_39573,N_37689,N_36941);
or U39574 (N_39574,N_36096,N_36562);
xnor U39575 (N_39575,N_36018,N_37651);
xor U39576 (N_39576,N_36754,N_36663);
and U39577 (N_39577,N_37043,N_36143);
or U39578 (N_39578,N_36084,N_37696);
nor U39579 (N_39579,N_36317,N_36719);
xnor U39580 (N_39580,N_36246,N_36211);
or U39581 (N_39581,N_37695,N_37213);
nand U39582 (N_39582,N_37905,N_37339);
xor U39583 (N_39583,N_36955,N_36754);
and U39584 (N_39584,N_36655,N_36151);
or U39585 (N_39585,N_37902,N_36442);
nand U39586 (N_39586,N_37646,N_36275);
xnor U39587 (N_39587,N_37555,N_37846);
and U39588 (N_39588,N_36370,N_37266);
xor U39589 (N_39589,N_37235,N_37176);
xor U39590 (N_39590,N_37024,N_37265);
and U39591 (N_39591,N_36410,N_37683);
xnor U39592 (N_39592,N_36671,N_37505);
nand U39593 (N_39593,N_36690,N_37882);
xor U39594 (N_39594,N_36885,N_36322);
nor U39595 (N_39595,N_36631,N_36213);
nand U39596 (N_39596,N_37669,N_37181);
or U39597 (N_39597,N_36878,N_37870);
or U39598 (N_39598,N_37082,N_36254);
nor U39599 (N_39599,N_36423,N_37398);
xnor U39600 (N_39600,N_37552,N_37632);
and U39601 (N_39601,N_37125,N_36514);
or U39602 (N_39602,N_37006,N_37053);
nor U39603 (N_39603,N_37543,N_37565);
and U39604 (N_39604,N_36252,N_37064);
nor U39605 (N_39605,N_36994,N_36778);
and U39606 (N_39606,N_37311,N_36162);
and U39607 (N_39607,N_36147,N_36752);
xor U39608 (N_39608,N_36011,N_36483);
nand U39609 (N_39609,N_36165,N_36272);
xnor U39610 (N_39610,N_36530,N_37551);
xor U39611 (N_39611,N_36906,N_37335);
nor U39612 (N_39612,N_36767,N_36747);
nor U39613 (N_39613,N_36074,N_36137);
nand U39614 (N_39614,N_37167,N_37030);
xnor U39615 (N_39615,N_36149,N_37158);
or U39616 (N_39616,N_36521,N_36183);
and U39617 (N_39617,N_37723,N_37631);
and U39618 (N_39618,N_37830,N_37346);
or U39619 (N_39619,N_37233,N_36925);
and U39620 (N_39620,N_36501,N_36853);
nand U39621 (N_39621,N_37761,N_37074);
or U39622 (N_39622,N_36668,N_36360);
xnor U39623 (N_39623,N_37092,N_36884);
or U39624 (N_39624,N_37720,N_36229);
or U39625 (N_39625,N_37037,N_37540);
and U39626 (N_39626,N_36040,N_37955);
nand U39627 (N_39627,N_37249,N_36211);
nand U39628 (N_39628,N_37347,N_37494);
or U39629 (N_39629,N_37941,N_36570);
nor U39630 (N_39630,N_37908,N_37250);
nor U39631 (N_39631,N_36409,N_37127);
nor U39632 (N_39632,N_37448,N_36000);
or U39633 (N_39633,N_37739,N_36157);
nand U39634 (N_39634,N_37800,N_36769);
and U39635 (N_39635,N_36415,N_37663);
nor U39636 (N_39636,N_37517,N_37283);
nor U39637 (N_39637,N_37253,N_36908);
xor U39638 (N_39638,N_36392,N_36629);
nor U39639 (N_39639,N_37751,N_37465);
xnor U39640 (N_39640,N_36070,N_36579);
or U39641 (N_39641,N_36444,N_36957);
xnor U39642 (N_39642,N_36167,N_37127);
nand U39643 (N_39643,N_36997,N_36312);
xor U39644 (N_39644,N_37176,N_37389);
nand U39645 (N_39645,N_36439,N_36848);
nand U39646 (N_39646,N_36845,N_37729);
nand U39647 (N_39647,N_37567,N_37531);
xor U39648 (N_39648,N_36151,N_36510);
and U39649 (N_39649,N_37130,N_37619);
nor U39650 (N_39650,N_37320,N_36833);
and U39651 (N_39651,N_37799,N_36354);
and U39652 (N_39652,N_36864,N_37659);
or U39653 (N_39653,N_37797,N_36904);
nor U39654 (N_39654,N_36459,N_37225);
xor U39655 (N_39655,N_37274,N_36946);
and U39656 (N_39656,N_36205,N_36406);
xor U39657 (N_39657,N_37758,N_37847);
nor U39658 (N_39658,N_36107,N_37442);
nor U39659 (N_39659,N_37009,N_36348);
nor U39660 (N_39660,N_37017,N_36685);
or U39661 (N_39661,N_36550,N_37421);
and U39662 (N_39662,N_36096,N_36366);
or U39663 (N_39663,N_36182,N_37436);
or U39664 (N_39664,N_37292,N_37318);
nor U39665 (N_39665,N_36148,N_37705);
and U39666 (N_39666,N_37922,N_36597);
nor U39667 (N_39667,N_37208,N_37053);
or U39668 (N_39668,N_36756,N_36621);
or U39669 (N_39669,N_36697,N_36123);
and U39670 (N_39670,N_37843,N_37488);
xnor U39671 (N_39671,N_37521,N_36838);
and U39672 (N_39672,N_36983,N_36403);
xnor U39673 (N_39673,N_37654,N_36044);
xor U39674 (N_39674,N_37909,N_36179);
xnor U39675 (N_39675,N_37305,N_36204);
xnor U39676 (N_39676,N_36408,N_37339);
xnor U39677 (N_39677,N_36911,N_37068);
nor U39678 (N_39678,N_36446,N_36308);
nand U39679 (N_39679,N_37376,N_36595);
nor U39680 (N_39680,N_36734,N_36663);
or U39681 (N_39681,N_36559,N_37896);
nand U39682 (N_39682,N_37312,N_36051);
nor U39683 (N_39683,N_36533,N_37763);
nor U39684 (N_39684,N_37572,N_37190);
nand U39685 (N_39685,N_36662,N_36203);
and U39686 (N_39686,N_36969,N_36319);
or U39687 (N_39687,N_37259,N_36501);
nand U39688 (N_39688,N_37511,N_36177);
nor U39689 (N_39689,N_36246,N_36188);
or U39690 (N_39690,N_36063,N_36724);
xor U39691 (N_39691,N_36954,N_37680);
nand U39692 (N_39692,N_36314,N_36950);
or U39693 (N_39693,N_37097,N_37497);
or U39694 (N_39694,N_37811,N_36706);
nand U39695 (N_39695,N_37341,N_37038);
nand U39696 (N_39696,N_37846,N_36767);
xor U39697 (N_39697,N_37638,N_37360);
nor U39698 (N_39698,N_36533,N_36987);
or U39699 (N_39699,N_37032,N_37093);
nor U39700 (N_39700,N_37172,N_36740);
or U39701 (N_39701,N_36609,N_36199);
xnor U39702 (N_39702,N_36955,N_36829);
and U39703 (N_39703,N_36600,N_36908);
nor U39704 (N_39704,N_36811,N_37292);
nor U39705 (N_39705,N_37461,N_37786);
nor U39706 (N_39706,N_36160,N_37786);
nand U39707 (N_39707,N_37569,N_37793);
and U39708 (N_39708,N_36797,N_37621);
and U39709 (N_39709,N_36267,N_37076);
or U39710 (N_39710,N_37922,N_37480);
or U39711 (N_39711,N_36981,N_36544);
xnor U39712 (N_39712,N_37763,N_37260);
or U39713 (N_39713,N_36179,N_36435);
or U39714 (N_39714,N_36931,N_37887);
nor U39715 (N_39715,N_37771,N_36522);
nand U39716 (N_39716,N_37040,N_37889);
and U39717 (N_39717,N_36938,N_36339);
xnor U39718 (N_39718,N_37642,N_37248);
and U39719 (N_39719,N_37053,N_37260);
xnor U39720 (N_39720,N_36294,N_36076);
nor U39721 (N_39721,N_36102,N_37699);
or U39722 (N_39722,N_37009,N_36124);
xnor U39723 (N_39723,N_36612,N_36805);
or U39724 (N_39724,N_37317,N_37611);
nor U39725 (N_39725,N_37802,N_36154);
xnor U39726 (N_39726,N_36887,N_36411);
or U39727 (N_39727,N_37220,N_37123);
nand U39728 (N_39728,N_37275,N_36642);
nor U39729 (N_39729,N_36814,N_36325);
nand U39730 (N_39730,N_36238,N_37743);
xor U39731 (N_39731,N_36999,N_36695);
xnor U39732 (N_39732,N_36616,N_37437);
and U39733 (N_39733,N_37316,N_37783);
and U39734 (N_39734,N_36227,N_36044);
xor U39735 (N_39735,N_36467,N_36056);
nand U39736 (N_39736,N_36240,N_37230);
nor U39737 (N_39737,N_37217,N_37702);
nor U39738 (N_39738,N_36719,N_36098);
nor U39739 (N_39739,N_36022,N_36341);
and U39740 (N_39740,N_36308,N_37501);
xnor U39741 (N_39741,N_37422,N_37178);
or U39742 (N_39742,N_37399,N_37800);
nor U39743 (N_39743,N_36770,N_36586);
nor U39744 (N_39744,N_37545,N_36081);
xor U39745 (N_39745,N_36084,N_37261);
and U39746 (N_39746,N_36402,N_37582);
nand U39747 (N_39747,N_37725,N_36791);
nor U39748 (N_39748,N_37107,N_36378);
nand U39749 (N_39749,N_37381,N_36634);
xnor U39750 (N_39750,N_37672,N_37075);
nand U39751 (N_39751,N_37934,N_37917);
nor U39752 (N_39752,N_36565,N_36856);
xor U39753 (N_39753,N_36112,N_37967);
or U39754 (N_39754,N_36153,N_36963);
or U39755 (N_39755,N_36034,N_37040);
nand U39756 (N_39756,N_36745,N_36699);
nand U39757 (N_39757,N_37890,N_36737);
nor U39758 (N_39758,N_36281,N_36146);
xor U39759 (N_39759,N_36637,N_37813);
xor U39760 (N_39760,N_37803,N_37191);
nor U39761 (N_39761,N_36997,N_37254);
nand U39762 (N_39762,N_36976,N_37688);
nor U39763 (N_39763,N_36912,N_37126);
nor U39764 (N_39764,N_37556,N_36736);
xor U39765 (N_39765,N_37431,N_37524);
or U39766 (N_39766,N_37979,N_37623);
and U39767 (N_39767,N_37318,N_36411);
or U39768 (N_39768,N_36879,N_37631);
and U39769 (N_39769,N_36719,N_36728);
xnor U39770 (N_39770,N_37387,N_37620);
nor U39771 (N_39771,N_36934,N_36923);
nand U39772 (N_39772,N_37563,N_36348);
and U39773 (N_39773,N_37111,N_37990);
and U39774 (N_39774,N_37665,N_36351);
and U39775 (N_39775,N_36452,N_36645);
and U39776 (N_39776,N_36811,N_36538);
nor U39777 (N_39777,N_36231,N_36194);
xnor U39778 (N_39778,N_37142,N_36272);
or U39779 (N_39779,N_36890,N_36335);
nand U39780 (N_39780,N_37213,N_37659);
or U39781 (N_39781,N_37942,N_37525);
nand U39782 (N_39782,N_37327,N_37970);
nor U39783 (N_39783,N_37543,N_37862);
and U39784 (N_39784,N_36336,N_37970);
and U39785 (N_39785,N_36475,N_37639);
nor U39786 (N_39786,N_36790,N_37997);
nor U39787 (N_39787,N_37176,N_37447);
nand U39788 (N_39788,N_36424,N_36886);
and U39789 (N_39789,N_36231,N_36105);
xnor U39790 (N_39790,N_36432,N_36656);
xor U39791 (N_39791,N_36402,N_37140);
nor U39792 (N_39792,N_37478,N_37137);
nor U39793 (N_39793,N_36843,N_36410);
nor U39794 (N_39794,N_36016,N_36249);
and U39795 (N_39795,N_37838,N_37396);
nor U39796 (N_39796,N_36787,N_37049);
or U39797 (N_39797,N_36635,N_36726);
nand U39798 (N_39798,N_36402,N_37119);
or U39799 (N_39799,N_37475,N_37346);
or U39800 (N_39800,N_36535,N_36788);
nor U39801 (N_39801,N_36968,N_37833);
nand U39802 (N_39802,N_37716,N_37713);
xor U39803 (N_39803,N_37689,N_37301);
xnor U39804 (N_39804,N_36048,N_36998);
nor U39805 (N_39805,N_37938,N_37483);
nor U39806 (N_39806,N_36129,N_37303);
nand U39807 (N_39807,N_37682,N_37601);
nor U39808 (N_39808,N_37376,N_37954);
xnor U39809 (N_39809,N_37284,N_37955);
nor U39810 (N_39810,N_37409,N_37847);
and U39811 (N_39811,N_37636,N_36219);
xor U39812 (N_39812,N_37447,N_36413);
or U39813 (N_39813,N_37561,N_36368);
or U39814 (N_39814,N_36123,N_36837);
nor U39815 (N_39815,N_37728,N_36021);
nor U39816 (N_39816,N_36534,N_36662);
nand U39817 (N_39817,N_36042,N_36792);
nand U39818 (N_39818,N_36276,N_37388);
xnor U39819 (N_39819,N_36648,N_37964);
xnor U39820 (N_39820,N_37997,N_37218);
and U39821 (N_39821,N_37969,N_37696);
nor U39822 (N_39822,N_36808,N_37698);
xor U39823 (N_39823,N_37237,N_36230);
xnor U39824 (N_39824,N_36899,N_36730);
nor U39825 (N_39825,N_37728,N_36142);
or U39826 (N_39826,N_37938,N_37940);
xor U39827 (N_39827,N_37445,N_37605);
nor U39828 (N_39828,N_36960,N_36125);
nor U39829 (N_39829,N_36445,N_37956);
nand U39830 (N_39830,N_37608,N_37353);
and U39831 (N_39831,N_36207,N_37365);
or U39832 (N_39832,N_36826,N_37610);
nor U39833 (N_39833,N_36743,N_36860);
or U39834 (N_39834,N_36613,N_36050);
or U39835 (N_39835,N_36305,N_36632);
nor U39836 (N_39836,N_36973,N_36173);
and U39837 (N_39837,N_37376,N_36219);
and U39838 (N_39838,N_37993,N_37923);
nand U39839 (N_39839,N_36850,N_36350);
nand U39840 (N_39840,N_37087,N_36455);
xnor U39841 (N_39841,N_36327,N_36418);
or U39842 (N_39842,N_36415,N_37885);
nor U39843 (N_39843,N_36200,N_36065);
or U39844 (N_39844,N_36589,N_37797);
nor U39845 (N_39845,N_36857,N_36735);
xnor U39846 (N_39846,N_36456,N_37424);
nor U39847 (N_39847,N_37584,N_37012);
or U39848 (N_39848,N_36825,N_36466);
and U39849 (N_39849,N_36556,N_36042);
or U39850 (N_39850,N_37829,N_36142);
xor U39851 (N_39851,N_36838,N_37150);
or U39852 (N_39852,N_37148,N_37564);
or U39853 (N_39853,N_37253,N_37199);
or U39854 (N_39854,N_37497,N_37222);
nand U39855 (N_39855,N_36768,N_36267);
and U39856 (N_39856,N_37879,N_37804);
nor U39857 (N_39857,N_37387,N_37550);
xor U39858 (N_39858,N_37649,N_36880);
or U39859 (N_39859,N_37275,N_37484);
or U39860 (N_39860,N_36252,N_37110);
nor U39861 (N_39861,N_37080,N_37474);
nor U39862 (N_39862,N_37975,N_37775);
nor U39863 (N_39863,N_36853,N_37896);
or U39864 (N_39864,N_37077,N_37073);
nand U39865 (N_39865,N_37169,N_36269);
nor U39866 (N_39866,N_36654,N_36727);
nor U39867 (N_39867,N_37801,N_37329);
xor U39868 (N_39868,N_37649,N_37764);
and U39869 (N_39869,N_36701,N_37953);
and U39870 (N_39870,N_37983,N_37932);
xnor U39871 (N_39871,N_37454,N_36406);
nand U39872 (N_39872,N_36930,N_36426);
and U39873 (N_39873,N_37404,N_36760);
and U39874 (N_39874,N_37030,N_36191);
and U39875 (N_39875,N_37963,N_36941);
or U39876 (N_39876,N_36272,N_36296);
nand U39877 (N_39877,N_37002,N_37873);
nand U39878 (N_39878,N_37629,N_36656);
nand U39879 (N_39879,N_37407,N_37647);
nor U39880 (N_39880,N_36210,N_37270);
or U39881 (N_39881,N_37836,N_37214);
or U39882 (N_39882,N_37805,N_37563);
nor U39883 (N_39883,N_36686,N_36930);
and U39884 (N_39884,N_37367,N_36434);
and U39885 (N_39885,N_36188,N_36596);
xor U39886 (N_39886,N_36213,N_37937);
xnor U39887 (N_39887,N_36552,N_37969);
or U39888 (N_39888,N_37057,N_36756);
and U39889 (N_39889,N_37023,N_36851);
nand U39890 (N_39890,N_36008,N_36586);
xor U39891 (N_39891,N_36808,N_36395);
nor U39892 (N_39892,N_36213,N_36683);
nor U39893 (N_39893,N_37226,N_37431);
xnor U39894 (N_39894,N_37192,N_36788);
nor U39895 (N_39895,N_37345,N_36299);
xnor U39896 (N_39896,N_37106,N_37326);
nor U39897 (N_39897,N_37313,N_36214);
xnor U39898 (N_39898,N_37612,N_37671);
or U39899 (N_39899,N_37369,N_37744);
or U39900 (N_39900,N_36356,N_37124);
nand U39901 (N_39901,N_36929,N_36129);
xor U39902 (N_39902,N_37197,N_36797);
or U39903 (N_39903,N_36840,N_36001);
or U39904 (N_39904,N_37995,N_36363);
and U39905 (N_39905,N_36316,N_36306);
xor U39906 (N_39906,N_37291,N_37771);
nor U39907 (N_39907,N_37021,N_36170);
xor U39908 (N_39908,N_36919,N_36393);
xnor U39909 (N_39909,N_36393,N_36077);
xnor U39910 (N_39910,N_37933,N_36890);
nor U39911 (N_39911,N_37827,N_36616);
xor U39912 (N_39912,N_37317,N_37995);
xor U39913 (N_39913,N_36038,N_36599);
and U39914 (N_39914,N_37166,N_37990);
nand U39915 (N_39915,N_36797,N_37945);
or U39916 (N_39916,N_37884,N_36424);
nor U39917 (N_39917,N_36350,N_36667);
nor U39918 (N_39918,N_37187,N_36191);
xnor U39919 (N_39919,N_36542,N_37852);
xor U39920 (N_39920,N_36908,N_37995);
nor U39921 (N_39921,N_36802,N_36895);
or U39922 (N_39922,N_36441,N_37496);
nor U39923 (N_39923,N_36858,N_37562);
xor U39924 (N_39924,N_36952,N_37241);
xor U39925 (N_39925,N_36979,N_36790);
and U39926 (N_39926,N_37479,N_37279);
nand U39927 (N_39927,N_36897,N_37901);
and U39928 (N_39928,N_36473,N_36010);
nand U39929 (N_39929,N_37455,N_36122);
xor U39930 (N_39930,N_36627,N_37359);
xnor U39931 (N_39931,N_36177,N_36891);
xnor U39932 (N_39932,N_36966,N_37159);
or U39933 (N_39933,N_37377,N_36495);
nor U39934 (N_39934,N_36486,N_36677);
nand U39935 (N_39935,N_36253,N_36798);
xnor U39936 (N_39936,N_36881,N_37613);
nor U39937 (N_39937,N_36960,N_37251);
or U39938 (N_39938,N_37044,N_37800);
nand U39939 (N_39939,N_36081,N_36423);
nand U39940 (N_39940,N_36102,N_37187);
nand U39941 (N_39941,N_37402,N_36599);
and U39942 (N_39942,N_36065,N_37914);
nand U39943 (N_39943,N_36046,N_36198);
xor U39944 (N_39944,N_37586,N_37908);
or U39945 (N_39945,N_36945,N_37847);
nand U39946 (N_39946,N_36681,N_37271);
nand U39947 (N_39947,N_36923,N_37539);
and U39948 (N_39948,N_36057,N_36387);
or U39949 (N_39949,N_37609,N_37150);
xnor U39950 (N_39950,N_36534,N_37717);
and U39951 (N_39951,N_37445,N_37259);
or U39952 (N_39952,N_37956,N_36624);
xnor U39953 (N_39953,N_36200,N_36296);
nand U39954 (N_39954,N_36794,N_37454);
nor U39955 (N_39955,N_36490,N_37844);
nor U39956 (N_39956,N_37500,N_36978);
xnor U39957 (N_39957,N_37669,N_36838);
and U39958 (N_39958,N_37684,N_36880);
nor U39959 (N_39959,N_36271,N_36667);
or U39960 (N_39960,N_36177,N_36704);
and U39961 (N_39961,N_36358,N_36356);
nand U39962 (N_39962,N_37201,N_36892);
nor U39963 (N_39963,N_36583,N_37665);
xnor U39964 (N_39964,N_37940,N_37344);
nand U39965 (N_39965,N_36050,N_37819);
or U39966 (N_39966,N_36575,N_36827);
and U39967 (N_39967,N_37467,N_37770);
xor U39968 (N_39968,N_36519,N_37052);
xnor U39969 (N_39969,N_36639,N_37804);
nand U39970 (N_39970,N_36029,N_37580);
nand U39971 (N_39971,N_37817,N_37222);
or U39972 (N_39972,N_36721,N_37001);
xnor U39973 (N_39973,N_37509,N_37250);
nand U39974 (N_39974,N_37732,N_36505);
xor U39975 (N_39975,N_37271,N_36207);
or U39976 (N_39976,N_37140,N_37436);
nand U39977 (N_39977,N_37611,N_37086);
and U39978 (N_39978,N_37632,N_37600);
nor U39979 (N_39979,N_36701,N_37664);
and U39980 (N_39980,N_36888,N_36230);
nand U39981 (N_39981,N_37718,N_36421);
nor U39982 (N_39982,N_36989,N_37276);
or U39983 (N_39983,N_37998,N_37987);
xnor U39984 (N_39984,N_37323,N_37304);
nor U39985 (N_39985,N_36301,N_37964);
or U39986 (N_39986,N_37955,N_36015);
xnor U39987 (N_39987,N_37695,N_37407);
or U39988 (N_39988,N_37579,N_36547);
or U39989 (N_39989,N_36475,N_37366);
and U39990 (N_39990,N_36291,N_37716);
nand U39991 (N_39991,N_37272,N_36092);
and U39992 (N_39992,N_37798,N_36895);
xnor U39993 (N_39993,N_36768,N_37607);
xnor U39994 (N_39994,N_37981,N_36449);
nor U39995 (N_39995,N_37669,N_36961);
xor U39996 (N_39996,N_37491,N_37766);
and U39997 (N_39997,N_37261,N_36651);
xor U39998 (N_39998,N_37114,N_36247);
or U39999 (N_39999,N_37774,N_36103);
and U40000 (N_40000,N_38121,N_38469);
xnor U40001 (N_40001,N_38857,N_39384);
xor U40002 (N_40002,N_38774,N_39005);
nor U40003 (N_40003,N_38297,N_38790);
xnor U40004 (N_40004,N_39655,N_38265);
and U40005 (N_40005,N_38796,N_39348);
xor U40006 (N_40006,N_39635,N_39863);
nor U40007 (N_40007,N_38600,N_38041);
or U40008 (N_40008,N_38997,N_38667);
or U40009 (N_40009,N_38665,N_39639);
or U40010 (N_40010,N_38888,N_38019);
or U40011 (N_40011,N_39389,N_39745);
nor U40012 (N_40012,N_39299,N_38974);
or U40013 (N_40013,N_39754,N_38229);
or U40014 (N_40014,N_39315,N_38275);
nor U40015 (N_40015,N_38151,N_39708);
nor U40016 (N_40016,N_38718,N_38850);
and U40017 (N_40017,N_38598,N_38399);
and U40018 (N_40018,N_39910,N_38379);
or U40019 (N_40019,N_38903,N_38002);
nor U40020 (N_40020,N_38914,N_39105);
nor U40021 (N_40021,N_38506,N_38881);
and U40022 (N_40022,N_38291,N_39727);
and U40023 (N_40023,N_39515,N_38818);
and U40024 (N_40024,N_38022,N_38423);
and U40025 (N_40025,N_38919,N_38473);
and U40026 (N_40026,N_38089,N_39711);
and U40027 (N_40027,N_38754,N_38846);
xnor U40028 (N_40028,N_39466,N_38367);
xnor U40029 (N_40029,N_39646,N_39660);
xor U40030 (N_40030,N_39004,N_39517);
xnor U40031 (N_40031,N_38226,N_38648);
nor U40032 (N_40032,N_38276,N_38452);
and U40033 (N_40033,N_38928,N_38514);
and U40034 (N_40034,N_39246,N_38905);
xnor U40035 (N_40035,N_38823,N_38621);
and U40036 (N_40036,N_38738,N_39632);
nor U40037 (N_40037,N_39447,N_38509);
xor U40038 (N_40038,N_38875,N_39191);
nor U40039 (N_40039,N_38432,N_39484);
and U40040 (N_40040,N_39792,N_38688);
nand U40041 (N_40041,N_38462,N_38781);
xor U40042 (N_40042,N_39379,N_38840);
nand U40043 (N_40043,N_38540,N_39850);
and U40044 (N_40044,N_39149,N_38983);
nor U40045 (N_40045,N_39464,N_39420);
xor U40046 (N_40046,N_39067,N_39394);
or U40047 (N_40047,N_38256,N_39796);
and U40048 (N_40048,N_38885,N_38434);
and U40049 (N_40049,N_38938,N_38567);
nor U40050 (N_40050,N_38264,N_39081);
or U40051 (N_40051,N_38477,N_38483);
or U40052 (N_40052,N_39425,N_38366);
xnor U40053 (N_40053,N_39500,N_39165);
nand U40054 (N_40054,N_39586,N_38731);
nand U40055 (N_40055,N_39018,N_39166);
and U40056 (N_40056,N_38664,N_38582);
nor U40057 (N_40057,N_38179,N_38181);
xnor U40058 (N_40058,N_39038,N_38126);
or U40059 (N_40059,N_39088,N_38383);
xor U40060 (N_40060,N_39352,N_38119);
or U40061 (N_40061,N_38628,N_39519);
nand U40062 (N_40062,N_38597,N_38729);
xnor U40063 (N_40063,N_38095,N_38713);
xor U40064 (N_40064,N_39504,N_38958);
or U40065 (N_40065,N_39961,N_39229);
nand U40066 (N_40066,N_38936,N_39121);
xor U40067 (N_40067,N_38015,N_38541);
xor U40068 (N_40068,N_39082,N_39257);
or U40069 (N_40069,N_39617,N_38314);
nand U40070 (N_40070,N_38703,N_39022);
nor U40071 (N_40071,N_38955,N_39955);
or U40072 (N_40072,N_38058,N_39087);
xnor U40073 (N_40073,N_39865,N_38085);
xnor U40074 (N_40074,N_39702,N_38609);
nand U40075 (N_40075,N_39558,N_38829);
and U40076 (N_40076,N_39232,N_38944);
and U40077 (N_40077,N_38956,N_38136);
nand U40078 (N_40078,N_38158,N_39901);
or U40079 (N_40079,N_39092,N_38373);
xor U40080 (N_40080,N_38555,N_39684);
xor U40081 (N_40081,N_38087,N_38173);
and U40082 (N_40082,N_39450,N_38508);
nor U40083 (N_40083,N_38494,N_38932);
nand U40084 (N_40084,N_39279,N_39306);
xnor U40085 (N_40085,N_38464,N_38312);
nor U40086 (N_40086,N_39426,N_39124);
xnor U40087 (N_40087,N_38460,N_39759);
nand U40088 (N_40088,N_39360,N_38951);
and U40089 (N_40089,N_39951,N_38671);
xnor U40090 (N_40090,N_39520,N_38822);
nor U40091 (N_40091,N_39679,N_39095);
nand U40092 (N_40092,N_39355,N_38835);
nand U40093 (N_40093,N_39612,N_39904);
or U40094 (N_40094,N_39002,N_39623);
nand U40095 (N_40095,N_38893,N_39024);
or U40096 (N_40096,N_39561,N_38934);
nor U40097 (N_40097,N_39267,N_39753);
or U40098 (N_40098,N_38242,N_39099);
nor U40099 (N_40099,N_38200,N_38468);
xnor U40100 (N_40100,N_39505,N_39581);
and U40101 (N_40101,N_38415,N_39643);
nor U40102 (N_40102,N_38605,N_39486);
nor U40103 (N_40103,N_39887,N_39738);
nand U40104 (N_40104,N_39443,N_39377);
nand U40105 (N_40105,N_38153,N_38140);
xor U40106 (N_40106,N_38505,N_39465);
nor U40107 (N_40107,N_38907,N_38225);
and U40108 (N_40108,N_38203,N_38182);
xnor U40109 (N_40109,N_38478,N_38204);
xor U40110 (N_40110,N_39532,N_38524);
or U40111 (N_40111,N_39181,N_39113);
or U40112 (N_40112,N_39335,N_38248);
nor U40113 (N_40113,N_38219,N_39178);
nor U40114 (N_40114,N_38685,N_39490);
nand U40115 (N_40115,N_38396,N_38877);
nand U40116 (N_40116,N_38224,N_38359);
nor U40117 (N_40117,N_38583,N_39122);
or U40118 (N_40118,N_38694,N_39179);
or U40119 (N_40119,N_38674,N_39950);
xor U40120 (N_40120,N_39999,N_39816);
xor U40121 (N_40121,N_38213,N_38602);
nand U40122 (N_40122,N_39260,N_38608);
or U40123 (N_40123,N_38116,N_38520);
or U40124 (N_40124,N_38209,N_39441);
xor U40125 (N_40125,N_38240,N_39336);
or U40126 (N_40126,N_38308,N_39563);
nand U40127 (N_40127,N_39198,N_39776);
or U40128 (N_40128,N_38254,N_38145);
nor U40129 (N_40129,N_39442,N_39980);
nand U40130 (N_40130,N_39968,N_38438);
nand U40131 (N_40131,N_39469,N_39603);
and U40132 (N_40132,N_38719,N_39296);
nand U40133 (N_40133,N_39316,N_38198);
xor U40134 (N_40134,N_39750,N_38660);
nand U40135 (N_40135,N_38963,N_39765);
nand U40136 (N_40136,N_39930,N_39010);
nor U40137 (N_40137,N_38640,N_38737);
or U40138 (N_40138,N_38160,N_38528);
or U40139 (N_40139,N_39368,N_38645);
nor U40140 (N_40140,N_39917,N_38734);
nand U40141 (N_40141,N_39035,N_39799);
nor U40142 (N_40142,N_38354,N_38606);
or U40143 (N_40143,N_39280,N_39042);
xor U40144 (N_40144,N_39763,N_39046);
nor U40145 (N_40145,N_38206,N_39359);
or U40146 (N_40146,N_38966,N_38770);
or U40147 (N_40147,N_39560,N_38953);
xnor U40148 (N_40148,N_39777,N_38487);
or U40149 (N_40149,N_39044,N_38252);
and U40150 (N_40150,N_39848,N_38066);
nor U40151 (N_40151,N_39626,N_39023);
or U40152 (N_40152,N_39268,N_38266);
nor U40153 (N_40153,N_38316,N_38842);
and U40154 (N_40154,N_39458,N_39089);
nand U40155 (N_40155,N_39784,N_39262);
and U40156 (N_40156,N_39180,N_38696);
or U40157 (N_40157,N_38457,N_39456);
or U40158 (N_40158,N_38595,N_38050);
nand U40159 (N_40159,N_38003,N_38642);
and U40160 (N_40160,N_38725,N_38326);
nand U40161 (N_40161,N_38954,N_39544);
nand U40162 (N_40162,N_39036,N_38115);
and U40163 (N_40163,N_39924,N_39404);
or U40164 (N_40164,N_38976,N_38243);
xnor U40165 (N_40165,N_39548,N_38616);
and U40166 (N_40166,N_38573,N_39245);
nand U40167 (N_40167,N_39638,N_39615);
nor U40168 (N_40168,N_39125,N_38247);
xor U40169 (N_40169,N_38750,N_39290);
and U40170 (N_40170,N_39721,N_39749);
or U40171 (N_40171,N_39291,N_39964);
and U40172 (N_40172,N_39707,N_38388);
nor U40173 (N_40173,N_39851,N_39199);
xnor U40174 (N_40174,N_39417,N_39475);
or U40175 (N_40175,N_38552,N_39827);
nor U40176 (N_40176,N_38658,N_38189);
or U40177 (N_40177,N_38287,N_39704);
nor U40178 (N_40178,N_38049,N_38537);
nand U40179 (N_40179,N_38566,N_38199);
xor U40180 (N_40180,N_39568,N_39528);
nand U40181 (N_40181,N_38480,N_38786);
or U40182 (N_40182,N_38693,N_38346);
and U40183 (N_40183,N_38307,N_39885);
nor U40184 (N_40184,N_38286,N_39907);
xnor U40185 (N_40185,N_38249,N_39886);
nand U40186 (N_40186,N_38281,N_39772);
nand U40187 (N_40187,N_38724,N_39369);
or U40188 (N_40188,N_39782,N_38129);
xor U40189 (N_40189,N_38607,N_39758);
nand U40190 (N_40190,N_39650,N_39473);
and U40191 (N_40191,N_39193,N_39706);
nor U40192 (N_40192,N_39593,N_39733);
and U40193 (N_40193,N_39200,N_39699);
and U40194 (N_40194,N_39616,N_39818);
nand U40195 (N_40195,N_39476,N_38594);
and U40196 (N_40196,N_38649,N_39401);
nor U40197 (N_40197,N_38887,N_39471);
nor U40198 (N_40198,N_39567,N_38960);
and U40199 (N_40199,N_38639,N_39011);
nand U40200 (N_40200,N_39026,N_38064);
and U40201 (N_40201,N_39808,N_39506);
nand U40202 (N_40202,N_39152,N_39841);
or U40203 (N_40203,N_39562,N_39957);
or U40204 (N_40204,N_38666,N_38358);
nor U40205 (N_40205,N_38092,N_39353);
and U40206 (N_40206,N_38815,N_39694);
or U40207 (N_40207,N_38939,N_39527);
nor U40208 (N_40208,N_39977,N_39640);
or U40209 (N_40209,N_38838,N_39284);
nand U40210 (N_40210,N_38557,N_39872);
or U40211 (N_40211,N_38011,N_39631);
or U40212 (N_40212,N_39888,N_39894);
nor U40213 (N_40213,N_39761,N_39947);
or U40214 (N_40214,N_38183,N_39371);
and U40215 (N_40215,N_39480,N_39677);
xnor U40216 (N_40216,N_39669,N_39256);
nor U40217 (N_40217,N_38981,N_38854);
and U40218 (N_40218,N_39895,N_38561);
nor U40219 (N_40219,N_39676,N_38894);
and U40220 (N_40220,N_39331,N_39015);
and U40221 (N_40221,N_38086,N_39112);
nor U40222 (N_40222,N_39196,N_39009);
nand U40223 (N_40223,N_38037,N_39342);
xor U40224 (N_40224,N_39222,N_39387);
nand U40225 (N_40225,N_38704,N_39667);
xor U40226 (N_40226,N_38698,N_39236);
nand U40227 (N_40227,N_38592,N_38617);
nand U40228 (N_40228,N_38337,N_39569);
nor U40229 (N_40229,N_39062,N_39255);
nand U40230 (N_40230,N_39963,N_38395);
nor U40231 (N_40231,N_39867,N_39053);
xnor U40232 (N_40232,N_39974,N_39604);
and U40233 (N_40233,N_38467,N_39893);
xnor U40234 (N_40234,N_39918,N_39844);
nor U40235 (N_40235,N_39083,N_38496);
or U40236 (N_40236,N_39177,N_38924);
nand U40237 (N_40237,N_38122,N_39582);
and U40238 (N_40238,N_39071,N_38884);
and U40239 (N_40239,N_38341,N_39167);
or U40240 (N_40240,N_39878,N_38917);
nor U40241 (N_40241,N_39195,N_39800);
nor U40242 (N_40242,N_38593,N_38930);
nor U40243 (N_40243,N_38044,N_38262);
nor U40244 (N_40244,N_38634,N_38339);
or U40245 (N_40245,N_39109,N_38589);
or U40246 (N_40246,N_38431,N_38440);
or U40247 (N_40247,N_38652,N_38739);
nand U40248 (N_40248,N_38948,N_39382);
xor U40249 (N_40249,N_38865,N_39295);
xor U40250 (N_40250,N_39739,N_38171);
or U40251 (N_40251,N_39407,N_39148);
or U40252 (N_40252,N_38004,N_39409);
or U40253 (N_40253,N_39147,N_39680);
and U40254 (N_40254,N_38522,N_39857);
or U40255 (N_40255,N_39760,N_38051);
nand U40256 (N_40256,N_39543,N_39127);
nor U40257 (N_40257,N_38028,N_38220);
nand U40258 (N_40258,N_39644,N_38079);
xnor U40259 (N_40259,N_38527,N_38836);
and U40260 (N_40260,N_38891,N_39224);
nand U40261 (N_40261,N_39607,N_39115);
nor U40262 (N_40262,N_39111,N_39883);
or U40263 (N_40263,N_39959,N_38073);
xnor U40264 (N_40264,N_38449,N_38825);
nor U40265 (N_40265,N_38682,N_39186);
nand U40266 (N_40266,N_39956,N_38993);
or U40267 (N_40267,N_38251,N_39662);
xor U40268 (N_40268,N_38510,N_39118);
or U40269 (N_40269,N_39933,N_39884);
xnor U40270 (N_40270,N_39430,N_38344);
or U40271 (N_40271,N_39602,N_38328);
nor U40272 (N_40272,N_38563,N_39498);
nor U40273 (N_40273,N_39503,N_39275);
nand U40274 (N_40274,N_39228,N_39597);
nand U40275 (N_40275,N_39381,N_38493);
or U40276 (N_40276,N_38302,N_39438);
xnor U40277 (N_40277,N_39319,N_38858);
or U40278 (N_40278,N_39648,N_39986);
nand U40279 (N_40279,N_38728,N_38751);
xor U40280 (N_40280,N_38172,N_38402);
or U40281 (N_40281,N_38157,N_38808);
xor U40282 (N_40282,N_38238,N_38217);
xor U40283 (N_40283,N_38047,N_38138);
nand U40284 (N_40284,N_39789,N_39451);
nor U40285 (N_40285,N_39090,N_39059);
xor U40286 (N_40286,N_39274,N_39055);
and U40287 (N_40287,N_38068,N_38657);
nand U40288 (N_40288,N_39743,N_38856);
xor U40289 (N_40289,N_39129,N_38706);
or U40290 (N_40290,N_39052,N_39462);
nor U40291 (N_40291,N_39821,N_39217);
xnor U40292 (N_40292,N_39672,N_38042);
xor U40293 (N_40293,N_39658,N_38873);
nor U40294 (N_40294,N_38872,N_38123);
or U40295 (N_40295,N_39367,N_38654);
or U40296 (N_40296,N_38813,N_39590);
nand U40297 (N_40297,N_39823,N_38659);
and U40298 (N_40298,N_38986,N_39169);
nand U40299 (N_40299,N_39031,N_39244);
and U40300 (N_40300,N_39960,N_39880);
nor U40301 (N_40301,N_39334,N_38629);
nand U40302 (N_40302,N_38627,N_39550);
nor U40303 (N_40303,N_39097,N_39117);
xnor U40304 (N_40304,N_38847,N_38717);
or U40305 (N_40305,N_39405,N_39058);
nand U40306 (N_40306,N_38029,N_38531);
or U40307 (N_40307,N_38715,N_38851);
xnor U40308 (N_40308,N_39728,N_38832);
and U40309 (N_40309,N_39920,N_38476);
nand U40310 (N_40310,N_39170,N_39131);
or U40311 (N_40311,N_39211,N_39233);
nor U40312 (N_40312,N_38231,N_39254);
xor U40313 (N_40313,N_39554,N_38347);
xnor U40314 (N_40314,N_38127,N_38779);
or U40315 (N_40315,N_39637,N_38979);
or U40316 (N_40316,N_39459,N_38756);
or U40317 (N_40317,N_39340,N_39390);
xnor U40318 (N_40318,N_38331,N_39019);
xnor U40319 (N_40319,N_38961,N_39984);
xnor U40320 (N_40320,N_38964,N_39049);
nand U40321 (N_40321,N_38996,N_38711);
nand U40322 (N_40322,N_38599,N_39987);
or U40323 (N_40323,N_38973,N_38484);
and U40324 (N_40324,N_38879,N_38013);
nand U40325 (N_40325,N_39029,N_39156);
and U40326 (N_40326,N_38982,N_38864);
nand U40327 (N_40327,N_39145,N_38439);
and U40328 (N_40328,N_38309,N_39689);
xnor U40329 (N_40329,N_39123,N_39080);
or U40330 (N_40330,N_38192,N_38290);
xor U40331 (N_40331,N_39197,N_39483);
nand U40332 (N_40332,N_38775,N_39110);
nand U40333 (N_40333,N_38804,N_38435);
xnor U40334 (N_40334,N_38169,N_39512);
or U40335 (N_40335,N_39847,N_39300);
nand U40336 (N_40336,N_39742,N_39396);
nand U40337 (N_40337,N_39424,N_38662);
nor U40338 (N_40338,N_38397,N_38548);
or U40339 (N_40339,N_39478,N_38700);
xnor U40340 (N_40340,N_38603,N_38017);
xor U40341 (N_40341,N_38369,N_39997);
nor U40342 (N_40342,N_39696,N_38099);
or U40343 (N_40343,N_39511,N_39715);
or U40344 (N_40344,N_38980,N_38195);
and U40345 (N_40345,N_38735,N_39909);
xor U40346 (N_40346,N_39712,N_39549);
nand U40347 (N_40347,N_39205,N_38445);
and U40348 (N_40348,N_38147,N_38523);
nand U40349 (N_40349,N_38760,N_39374);
nor U40350 (N_40350,N_38472,N_38056);
xor U40351 (N_40351,N_39130,N_39678);
nand U40352 (N_40352,N_38677,N_38260);
xnor U40353 (N_40353,N_38353,N_39846);
and U40354 (N_40354,N_38826,N_39204);
nand U40355 (N_40355,N_38408,N_39454);
and U40356 (N_40356,N_39891,N_39429);
nor U40357 (N_40357,N_38912,N_39618);
nand U40358 (N_40358,N_39120,N_38504);
xnor U40359 (N_40359,N_38726,N_38797);
xnor U40360 (N_40360,N_38673,N_39819);
and U40361 (N_40361,N_39435,N_38257);
nor U40362 (N_40362,N_38533,N_39444);
nor U40363 (N_40363,N_39399,N_39713);
and U40364 (N_40364,N_39251,N_38994);
nand U40365 (N_40365,N_39014,N_39903);
nor U40366 (N_40366,N_39864,N_39155);
nand U40367 (N_40367,N_38536,N_39460);
nand U40368 (N_40368,N_39954,N_39051);
and U40369 (N_40369,N_39237,N_39173);
and U40370 (N_40370,N_39326,N_38581);
nor U40371 (N_40371,N_38987,N_38419);
or U40372 (N_40372,N_38190,N_39656);
and U40373 (N_40373,N_38057,N_38232);
and U40374 (N_40374,N_38390,N_39214);
nor U40375 (N_40375,N_38783,N_38280);
or U40376 (N_40376,N_38277,N_38901);
xor U40377 (N_40377,N_38456,N_39665);
nor U40378 (N_40378,N_39989,N_38810);
xor U40379 (N_40379,N_38448,N_38176);
nand U40380 (N_40380,N_39832,N_38896);
xnor U40381 (N_40381,N_38097,N_39411);
and U40382 (N_40382,N_39273,N_38132);
or U40383 (N_40383,N_38799,N_38356);
xnor U40384 (N_40384,N_39731,N_39578);
and U40385 (N_40385,N_39277,N_38422);
and U40386 (N_40386,N_39645,N_39240);
or U40387 (N_40387,N_38384,N_38026);
or U40388 (N_40388,N_38038,N_38902);
and U40389 (N_40389,N_39363,N_38428);
and U40390 (N_40390,N_39730,N_38625);
and U40391 (N_40391,N_39470,N_39943);
nor U40392 (N_40392,N_39627,N_38519);
or U40393 (N_40393,N_38210,N_38845);
or U40394 (N_40394,N_38992,N_39323);
xnor U40395 (N_40395,N_38759,N_39613);
or U40396 (N_40396,N_39128,N_39585);
xnor U40397 (N_40397,N_38773,N_38168);
and U40398 (N_40398,N_39289,N_39724);
or U40399 (N_40399,N_38672,N_38118);
and U40400 (N_40400,N_38162,N_39595);
or U40401 (N_40401,N_38320,N_38348);
nor U40402 (N_40402,N_39154,N_38580);
and U40403 (N_40403,N_39915,N_38733);
and U40404 (N_40404,N_38646,N_38860);
nand U40405 (N_40405,N_39033,N_38977);
xor U40406 (N_40406,N_39219,N_39346);
or U40407 (N_40407,N_38793,N_38134);
or U40408 (N_40408,N_39188,N_38370);
xor U40409 (N_40409,N_38084,N_38638);
or U40410 (N_40410,N_39116,N_39041);
nand U40411 (N_40411,N_39716,N_39175);
and U40412 (N_40412,N_39858,N_39096);
nor U40413 (N_40413,N_38572,N_39762);
nand U40414 (N_40414,N_38539,N_38117);
nand U40415 (N_40415,N_38710,N_39061);
xnor U40416 (N_40416,N_38604,N_39820);
nand U40417 (N_40417,N_39270,N_39370);
nor U40418 (N_40418,N_38062,N_39767);
xor U40419 (N_40419,N_39845,N_39171);
or U40420 (N_40420,N_39892,N_38636);
nand U40421 (N_40421,N_39013,N_38904);
nand U40422 (N_40422,N_39812,N_39467);
nand U40423 (N_40423,N_39533,N_38125);
xor U40424 (N_40424,N_38485,N_39376);
nor U40425 (N_40425,N_38362,N_39970);
nand U40426 (N_40426,N_38430,N_39412);
and U40427 (N_40427,N_38152,N_39868);
or U40428 (N_40428,N_39440,N_38322);
nand U40429 (N_40429,N_39911,N_38036);
nor U40430 (N_40430,N_39771,N_39834);
or U40431 (N_40431,N_39735,N_39069);
xor U40432 (N_40432,N_39630,N_38795);
nand U40433 (N_40433,N_39075,N_39591);
or U40434 (N_40434,N_39570,N_39555);
or U40435 (N_40435,N_39263,N_38765);
and U40436 (N_40436,N_38149,N_39988);
nand U40437 (N_40437,N_38789,N_38416);
xnor U40438 (N_40438,N_38538,N_38244);
nand U40439 (N_40439,N_39770,N_39189);
nand U40440 (N_40440,N_39744,N_38495);
or U40441 (N_40441,N_38687,N_38867);
and U40442 (N_40442,N_39373,N_38197);
and U40443 (N_40443,N_39012,N_38692);
and U40444 (N_40444,N_38223,N_39305);
or U40445 (N_40445,N_39962,N_38767);
and U40446 (N_40446,N_38663,N_39837);
nor U40447 (N_40447,N_38909,N_39830);
xnor U40448 (N_40448,N_38294,N_39135);
xor U40449 (N_40449,N_39203,N_38361);
and U40450 (N_40450,N_39380,N_38043);
and U40451 (N_40451,N_39521,N_39815);
or U40452 (N_40452,N_38270,N_38543);
xnor U40453 (N_40453,N_39971,N_38551);
or U40454 (N_40454,N_38880,N_39755);
xnor U40455 (N_40455,N_39328,N_38820);
and U40456 (N_40456,N_38046,N_38550);
xnor U40457 (N_40457,N_39151,N_39047);
nor U40458 (N_40458,N_38910,N_38070);
or U40459 (N_40459,N_38278,N_38908);
xor U40460 (N_40460,N_39213,N_39144);
nand U40461 (N_40461,N_38807,N_38191);
or U40462 (N_40462,N_39421,N_39862);
xnor U40463 (N_40463,N_39861,N_39372);
and U40464 (N_40464,N_38377,N_38131);
nor U40465 (N_40465,N_39361,N_39701);
nand U40466 (N_40466,N_38641,N_38313);
and U40467 (N_40467,N_38686,N_39098);
or U40468 (N_40468,N_38516,N_39139);
nand U40469 (N_40469,N_38985,N_39094);
or U40470 (N_40470,N_39803,N_38385);
xor U40471 (N_40471,N_39877,N_38106);
nand U40472 (N_40472,N_38827,N_38007);
and U40473 (N_40473,N_38651,N_39671);
xor U40474 (N_40474,N_38915,N_39001);
xnor U40475 (N_40475,N_39788,N_38586);
xnor U40476 (N_40476,N_39542,N_39241);
nand U40477 (N_40477,N_39302,N_39060);
or U40478 (N_40478,N_39007,N_39327);
and U40479 (N_40479,N_39086,N_39106);
and U40480 (N_40480,N_39525,N_39248);
or U40481 (N_40481,N_39101,N_39691);
or U40482 (N_40482,N_38926,N_39798);
and U40483 (N_40483,N_38632,N_38707);
and U40484 (N_40484,N_39449,N_39551);
nor U40485 (N_40485,N_38762,N_38025);
or U40486 (N_40486,N_39419,N_38072);
nand U40487 (N_40487,N_38098,N_39108);
xnor U40488 (N_40488,N_38819,N_38761);
xnor U40489 (N_40489,N_38777,N_38420);
or U40490 (N_40490,N_38021,N_38833);
or U40491 (N_40491,N_39806,N_39566);
or U40492 (N_40492,N_39313,N_39889);
or U40493 (N_40493,N_39916,N_38295);
xnor U40494 (N_40494,N_39364,N_39393);
nand U40495 (N_40495,N_39032,N_38215);
or U40496 (N_40496,N_39298,N_39698);
xnor U40497 (N_40497,N_38890,N_39596);
nor U40498 (N_40498,N_39497,N_39526);
xnor U40499 (N_40499,N_38030,N_39184);
nand U40500 (N_40500,N_39985,N_38869);
and U40501 (N_40501,N_38998,N_38655);
and U40502 (N_40502,N_38900,N_38529);
xnor U40503 (N_40503,N_38090,N_39338);
nor U40504 (N_40504,N_39201,N_38755);
xnor U40505 (N_40505,N_38500,N_38273);
and U40506 (N_40506,N_38006,N_39783);
xor U40507 (N_40507,N_38336,N_39822);
nor U40508 (N_40508,N_39378,N_39687);
and U40509 (N_40509,N_38637,N_39693);
nand U40510 (N_40510,N_39428,N_38568);
and U40511 (N_40511,N_39463,N_39995);
and U40512 (N_40512,N_38113,N_38412);
or U40513 (N_40513,N_39981,N_39766);
nor U40514 (N_40514,N_38757,N_39785);
nand U40515 (N_40515,N_38497,N_39247);
nand U40516 (N_40516,N_39900,N_39668);
nand U40517 (N_40517,N_38338,N_38352);
and U40518 (N_40518,N_38413,N_38764);
and U40519 (N_40519,N_39472,N_38296);
and U40520 (N_40520,N_38906,N_39934);
or U40521 (N_40521,N_38031,N_38027);
nor U40522 (N_40522,N_39842,N_38556);
nor U40523 (N_40523,N_39453,N_39423);
xnor U40524 (N_40524,N_39079,N_38241);
nand U40525 (N_40525,N_38405,N_38436);
nor U40526 (N_40526,N_39375,N_39119);
nand U40527 (N_40527,N_38268,N_39932);
xnor U40528 (N_40528,N_38768,N_38988);
xnor U40529 (N_40529,N_38427,N_39418);
or U40530 (N_40530,N_39043,N_38475);
and U40531 (N_40531,N_39831,N_38156);
and U40532 (N_40532,N_39529,N_39606);
nor U40533 (N_40533,N_39242,N_38619);
nor U40534 (N_40534,N_38702,N_39153);
or U40535 (N_40535,N_39252,N_39935);
nor U40536 (N_40536,N_38758,N_38853);
nor U40537 (N_40537,N_39301,N_39666);
and U40538 (N_40538,N_38878,N_39620);
nand U40539 (N_40539,N_38554,N_39446);
or U40540 (N_40540,N_38800,N_39925);
nand U40541 (N_40541,N_38562,N_39317);
and U40542 (N_40542,N_38736,N_38357);
nand U40543 (N_40543,N_39264,N_39619);
xnor U40544 (N_40544,N_38005,N_38585);
nand U40545 (N_40545,N_39580,N_38942);
or U40546 (N_40546,N_38305,N_39634);
and U40547 (N_40547,N_38670,N_38798);
xnor U40548 (N_40548,N_39577,N_38871);
nor U40549 (N_40549,N_38424,N_39881);
xor U40550 (N_40550,N_38916,N_39781);
and U40551 (N_40551,N_38716,N_39879);
or U40552 (N_40552,N_38576,N_39732);
xnor U40553 (N_40553,N_38180,N_39415);
nor U40554 (N_40554,N_38623,N_39875);
and U40555 (N_40555,N_39685,N_38389);
or U40556 (N_40556,N_39439,N_38184);
xnor U40557 (N_40557,N_38380,N_38697);
and U40558 (N_40558,N_39905,N_39809);
and U40559 (N_40559,N_39161,N_38989);
xnor U40560 (N_40560,N_39157,N_38343);
and U40561 (N_40561,N_38364,N_38839);
nand U40562 (N_40562,N_38048,N_38055);
or U40563 (N_40563,N_38237,N_38018);
nand U40564 (N_40564,N_38253,N_38558);
or U40565 (N_40565,N_39065,N_38681);
nor U40566 (N_40566,N_39350,N_38000);
nand U40567 (N_40567,N_38633,N_39286);
or U40568 (N_40568,N_38656,N_38749);
or U40569 (N_40569,N_39039,N_38111);
or U40570 (N_40570,N_39652,N_38560);
xor U40571 (N_40571,N_38675,N_38078);
nor U40572 (N_40572,N_38526,N_39945);
nor U40573 (N_40573,N_39940,N_38263);
nor U40574 (N_40574,N_39902,N_39736);
xnor U40575 (N_40575,N_39223,N_38946);
nor U40576 (N_40576,N_38684,N_39941);
nand U40577 (N_40577,N_39654,N_38311);
or U40578 (N_40578,N_38455,N_38208);
nand U40579 (N_40579,N_39912,N_39780);
xnor U40580 (N_40580,N_39982,N_39998);
nor U40581 (N_40581,N_39791,N_38318);
xnor U40582 (N_40582,N_39748,N_38014);
xor U40583 (N_40583,N_38785,N_38001);
and U40584 (N_40584,N_38848,N_39825);
xor U40585 (N_40585,N_38110,N_39574);
xnor U40586 (N_40586,N_38292,N_38577);
or U40587 (N_40587,N_39673,N_39400);
nand U40588 (N_40588,N_39801,N_38876);
nand U40589 (N_40589,N_38144,N_39534);
and U40590 (N_40590,N_39057,N_38150);
nor U40591 (N_40591,N_38109,N_38852);
or U40592 (N_40592,N_39091,N_38447);
nand U40593 (N_40593,N_38474,N_38425);
xnor U40594 (N_40594,N_38283,N_38112);
or U40595 (N_40595,N_38747,N_38288);
and U40596 (N_40596,N_38742,N_39692);
and U40597 (N_40597,N_38368,N_39564);
or U40598 (N_40598,N_38763,N_38991);
nor U40599 (N_40599,N_38778,N_39448);
xnor U40600 (N_40600,N_38730,N_39134);
nand U40601 (N_40601,N_39628,N_39729);
nor U40602 (N_40602,N_38542,N_38471);
nand U40603 (N_40603,N_39045,N_39690);
xor U40604 (N_40604,N_39869,N_38574);
and U40605 (N_40605,N_38479,N_38020);
nor U40606 (N_40606,N_39584,N_38401);
and U40607 (N_40607,N_38952,N_38794);
nand U40608 (N_40608,N_38193,N_39949);
nor U40609 (N_40609,N_39269,N_38709);
nand U40610 (N_40610,N_38969,N_39967);
or U40611 (N_40611,N_39572,N_39538);
or U40612 (N_40612,N_39502,N_39852);
xor U40613 (N_40613,N_38745,N_38486);
or U40614 (N_40614,N_39972,N_39757);
and U40615 (N_40615,N_38083,N_39162);
and U40616 (N_40616,N_39598,N_39826);
and U40617 (N_40617,N_39675,N_38805);
nand U40618 (N_40618,N_38889,N_39397);
nor U40619 (N_40619,N_38788,N_38535);
and U40620 (N_40620,N_38727,N_38016);
or U40621 (N_40621,N_38441,N_38792);
or U40622 (N_40622,N_39674,N_39908);
and U40623 (N_40623,N_39536,N_38481);
or U40624 (N_40624,N_38925,N_39764);
and U40625 (N_40625,N_38584,N_39332);
nand U40626 (N_40626,N_39705,N_38146);
nand U40627 (N_40627,N_39541,N_39365);
and U40628 (N_40628,N_39416,N_39003);
nor U40629 (N_40629,N_38301,N_39385);
nor U40630 (N_40630,N_38837,N_39890);
and U40631 (N_40631,N_38207,N_39769);
nand U40632 (N_40632,N_38211,N_39293);
and U40633 (N_40633,N_39016,N_39114);
nand U40634 (N_40634,N_39017,N_39592);
or U40635 (N_40635,N_39461,N_38033);
nand U40636 (N_40636,N_38780,N_38414);
and U40637 (N_40637,N_39913,N_38534);
and U40638 (N_40638,N_38678,N_38451);
or U40639 (N_40639,N_39164,N_38114);
or U40640 (N_40640,N_38345,N_39714);
and U40641 (N_40641,N_39659,N_38299);
nand U40642 (N_40642,N_39817,N_38130);
or U40643 (N_40643,N_38679,N_39922);
nor U40644 (N_40644,N_38886,N_38899);
or U40645 (N_40645,N_38221,N_38590);
nand U40646 (N_40646,N_38272,N_38032);
and U40647 (N_40647,N_39259,N_39492);
and U40648 (N_40648,N_38446,N_39507);
and U40649 (N_40649,N_38463,N_39482);
or U40650 (N_40650,N_38972,N_38714);
nor U40651 (N_40651,N_39192,N_39395);
nor U40652 (N_40652,N_38075,N_39100);
and U40653 (N_40653,N_39383,N_38784);
and U40654 (N_40654,N_39174,N_39583);
nand U40655 (N_40655,N_38250,N_38545);
nand U40656 (N_40656,N_38498,N_38061);
or U40657 (N_40657,N_39457,N_39339);
nand U40658 (N_40658,N_39265,N_39034);
nor U40659 (N_40659,N_38334,N_39859);
xor U40660 (N_40660,N_39787,N_39261);
nand U40661 (N_40661,N_38721,N_39138);
or U40662 (N_40662,N_39354,N_39006);
and U40663 (N_40663,N_39828,N_38315);
and U40664 (N_40664,N_38613,N_39746);
nand U40665 (N_40665,N_38404,N_38323);
nor U40666 (N_40666,N_39663,N_39605);
or U40667 (N_40667,N_39392,N_39856);
xnor U40668 (N_40668,N_39571,N_39073);
nor U40669 (N_40669,N_38063,N_39386);
or U40670 (N_40670,N_38874,N_38300);
xor U40671 (N_40671,N_38398,N_38748);
xnor U40672 (N_40672,N_38482,N_39076);
nor U40673 (N_40673,N_39432,N_39427);
and U40674 (N_40674,N_39351,N_38258);
or U40675 (N_40675,N_39522,N_39294);
nand U40676 (N_40676,N_39176,N_39066);
nand U40677 (N_40677,N_39107,N_39768);
xor U40678 (N_40678,N_39594,N_38587);
nor U40679 (N_40679,N_38630,N_39140);
and U40680 (N_40680,N_38959,N_38082);
or U40681 (N_40681,N_39547,N_39720);
nand U40682 (N_40682,N_38166,N_39838);
or U40683 (N_40683,N_39206,N_39751);
and U40684 (N_40684,N_38546,N_39683);
xor U40685 (N_40685,N_38935,N_38165);
nor U40686 (N_40686,N_39068,N_38647);
and U40687 (N_40687,N_38547,N_39102);
or U40688 (N_40688,N_39487,N_38045);
and U40689 (N_40689,N_38330,N_39281);
xor U40690 (N_40690,N_38394,N_38965);
or U40691 (N_40691,N_39309,N_39182);
nor U40692 (N_40692,N_39194,N_38863);
and U40693 (N_40693,N_39695,N_38950);
and U40694 (N_40694,N_38614,N_38120);
or U40695 (N_40695,N_39717,N_38205);
and U40696 (N_40696,N_39686,N_39579);
and U40697 (N_40697,N_38806,N_39215);
xnor U40698 (N_40698,N_38228,N_39501);
nand U40699 (N_40699,N_38411,N_39413);
nand U40700 (N_40700,N_39843,N_38553);
nor U40701 (N_40701,N_38393,N_39855);
nand U40702 (N_40702,N_38569,N_39790);
or U40703 (N_40703,N_39477,N_39833);
nor U40704 (N_40704,N_39938,N_39347);
xor U40705 (N_40705,N_39994,N_38712);
and U40706 (N_40706,N_38861,N_38544);
or U40707 (N_40707,N_38306,N_39285);
or U40708 (N_40708,N_39697,N_38107);
and U40709 (N_40709,N_38053,N_39990);
nand U40710 (N_40710,N_38752,N_39468);
nand U40711 (N_40711,N_39485,N_38859);
and U40712 (N_40712,N_39871,N_38382);
or U40713 (N_40713,N_38444,N_39709);
nand U40714 (N_40714,N_39357,N_38769);
xor U40715 (N_40715,N_38175,N_39545);
nor U40716 (N_40716,N_38511,N_39249);
xnor U40717 (N_40717,N_38105,N_39649);
nand U40718 (N_40718,N_39642,N_38060);
xor U40719 (N_40719,N_39559,N_38327);
xnor U40720 (N_40720,N_38378,N_39137);
or U40721 (N_40721,N_39288,N_39797);
or U40722 (N_40722,N_38501,N_39936);
and U40723 (N_40723,N_39927,N_38920);
nor U40724 (N_40724,N_39235,N_38317);
nor U40725 (N_40725,N_39163,N_39054);
or U40726 (N_40726,N_38024,N_38142);
and U40727 (N_40727,N_39048,N_38532);
xor U40728 (N_40728,N_38695,N_39314);
or U40729 (N_40729,N_38088,N_39814);
xnor U40730 (N_40730,N_38077,N_39366);
xor U40731 (N_40731,N_38776,N_39734);
xnor U40732 (N_40732,N_38069,N_39499);
xor U40733 (N_40733,N_39939,N_39190);
and U40734 (N_40734,N_38094,N_38100);
or U40735 (N_40735,N_39513,N_38236);
xor U40736 (N_40736,N_39756,N_39272);
or U40737 (N_40737,N_39150,N_38104);
nand U40738 (N_40738,N_38990,N_39775);
and U40739 (N_40739,N_39608,N_39625);
and U40740 (N_40740,N_38284,N_38618);
and U40741 (N_40741,N_39992,N_38012);
or U40742 (N_40742,N_38631,N_39216);
and U40743 (N_40743,N_38403,N_38421);
nand U40744 (N_40744,N_38040,N_39811);
or U40745 (N_40745,N_38669,N_38321);
and U40746 (N_40746,N_38304,N_39085);
nand U40747 (N_40747,N_38610,N_38913);
nor U40748 (N_40748,N_38791,N_39965);
nor U40749 (N_40749,N_39243,N_39330);
nand U40750 (N_40750,N_38978,N_38081);
or U40751 (N_40751,N_38143,N_38185);
and U40752 (N_40752,N_38588,N_39208);
nand U40753 (N_40753,N_39388,N_39839);
or U40754 (N_40754,N_39810,N_38644);
xnor U40755 (N_40755,N_39303,N_39614);
nand U40756 (N_40756,N_39737,N_39931);
nand U40757 (N_40757,N_38676,N_38340);
nor U40758 (N_40758,N_39942,N_38035);
or U40759 (N_40759,N_39588,N_39641);
and U40760 (N_40760,N_39282,N_38933);
nor U40761 (N_40761,N_38271,N_38201);
xnor U40762 (N_40762,N_38999,N_39896);
nand U40763 (N_40763,N_39882,N_39836);
or U40764 (N_40764,N_39345,N_39168);
or U40765 (N_40765,N_39937,N_38261);
or U40766 (N_40766,N_38870,N_38521);
or U40767 (N_40767,N_39874,N_38626);
or U40768 (N_40768,N_38816,N_39278);
xor U40769 (N_40769,N_39258,N_38940);
or U40770 (N_40770,N_38124,N_38701);
and U40771 (N_40771,N_38376,N_38255);
nand U40772 (N_40772,N_38689,N_39723);
and U40773 (N_40773,N_38705,N_38289);
or U40774 (N_40774,N_38372,N_39509);
or U40775 (N_40775,N_39725,N_39431);
nand U40776 (N_40776,N_38844,N_39813);
xor U40777 (N_40777,N_38849,N_38407);
or U40778 (N_40778,N_39653,N_39921);
nand U40779 (N_40779,N_39070,N_39966);
xor U40780 (N_40780,N_38923,N_38831);
and U40781 (N_40781,N_39324,N_39718);
or U40782 (N_40782,N_38054,N_38429);
or U40783 (N_40783,N_38387,N_38234);
nand U40784 (N_40784,N_39050,N_38202);
or U40785 (N_40785,N_39218,N_39741);
nand U40786 (N_40786,N_38096,N_38488);
xor U40787 (N_40787,N_39946,N_38661);
and U40788 (N_40788,N_39853,N_39078);
nor U40789 (N_40789,N_39975,N_38635);
or U40790 (N_40790,N_39494,N_39752);
or U40791 (N_40791,N_38067,N_38194);
xor U40792 (N_40792,N_38285,N_39320);
nor U40793 (N_40793,N_38921,N_38620);
or U40794 (N_40794,N_39926,N_39344);
or U40795 (N_40795,N_39919,N_39530);
and U40796 (N_40796,N_38892,N_38571);
nor U40797 (N_40797,N_39958,N_39661);
and U40798 (N_40798,N_39953,N_39866);
xnor U40799 (N_40799,N_39207,N_38039);
or U40800 (N_40800,N_38525,N_38499);
and U40801 (N_40801,N_38188,N_39403);
xnor U40802 (N_40802,N_38732,N_39433);
xnor U40803 (N_40803,N_39493,N_38967);
nand U40804 (N_40804,N_39297,N_38458);
and U40805 (N_40805,N_39056,N_39325);
nand U40806 (N_40806,N_38489,N_38450);
or U40807 (N_40807,N_38466,N_39231);
and U40808 (N_40808,N_39629,N_39020);
xor U40809 (N_40809,N_38154,N_39906);
nand U40810 (N_40810,N_39209,N_38491);
nor U40811 (N_40811,N_38332,N_38319);
or U40812 (N_40812,N_38492,N_39146);
nor U40813 (N_40813,N_39710,N_39944);
nand U40814 (N_40814,N_39074,N_39037);
and U40815 (N_40815,N_39793,N_39508);
nand U40816 (N_40816,N_39681,N_38259);
and U40817 (N_40817,N_38417,N_38298);
nor U40818 (N_40818,N_38828,N_39126);
nor U40819 (N_40819,N_38239,N_39021);
and U40820 (N_40820,N_39807,N_39774);
nor U40821 (N_40821,N_39553,N_38882);
or U40822 (N_40822,N_39805,N_39829);
nand U40823 (N_40823,N_38374,N_39158);
and U40824 (N_40824,N_39133,N_39539);
nor U40825 (N_40825,N_39778,N_39495);
nand U40826 (N_40826,N_39804,N_39979);
and U40827 (N_40827,N_39983,N_39136);
or U40828 (N_40828,N_38787,N_39000);
nor U40829 (N_40829,N_39027,N_38668);
and U40830 (N_40830,N_39341,N_38490);
or U40831 (N_40831,N_39311,N_39310);
and U40832 (N_40832,N_39524,N_38155);
xor U40833 (N_40833,N_39343,N_39063);
xor U40834 (N_40834,N_39266,N_38650);
nor U40835 (N_40835,N_39740,N_39546);
or U40836 (N_40836,N_38643,N_38911);
nand U40837 (N_40837,N_39250,N_38400);
xnor U40838 (N_40838,N_39565,N_38148);
and U40839 (N_40839,N_38222,N_38164);
and U40840 (N_40840,N_39406,N_39491);
nor U40841 (N_40841,N_38371,N_39601);
nand U40842 (N_40842,N_38690,N_38578);
xnor U40843 (N_40843,N_38392,N_38918);
or U40844 (N_40844,N_39141,N_39437);
xnor U40845 (N_40845,N_38766,N_38931);
nand U40846 (N_40846,N_39028,N_38834);
nor U40847 (N_40847,N_38459,N_38929);
xnor U40848 (N_40848,N_38862,N_39422);
xor U40849 (N_40849,N_38802,N_39225);
nor U40850 (N_40850,N_38365,N_39622);
nor U40851 (N_40851,N_39025,N_38461);
and U40852 (N_40852,N_38059,N_39898);
nand U40853 (N_40853,N_38897,N_38269);
nand U40854 (N_40854,N_38615,N_39899);
nor U40855 (N_40855,N_38381,N_38186);
or U40856 (N_40856,N_39040,N_38611);
or U40857 (N_40857,N_38009,N_38821);
and U40858 (N_40858,N_38159,N_38233);
and U40859 (N_40859,N_38128,N_39227);
or U40860 (N_40860,N_39271,N_39488);
or U40861 (N_40861,N_39160,N_38406);
nor U40862 (N_40862,N_39030,N_39587);
and U40863 (N_40863,N_38937,N_38741);
or U40864 (N_40864,N_39329,N_39321);
xnor U40865 (N_40865,N_39292,N_38282);
and U40866 (N_40866,N_39103,N_39952);
and U40867 (N_40867,N_38133,N_39307);
nand U40868 (N_40868,N_38071,N_39337);
nand U40869 (N_40869,N_38898,N_38811);
or U40870 (N_40870,N_39747,N_39794);
nand U40871 (N_40871,N_39172,N_38245);
and U40872 (N_40872,N_38325,N_38895);
nor U40873 (N_40873,N_39308,N_38949);
nand U40874 (N_40874,N_39455,N_39234);
and U40875 (N_40875,N_38418,N_39479);
nor U40876 (N_40876,N_38782,N_39786);
nor U40877 (N_40877,N_39978,N_38442);
nand U40878 (N_40878,N_39287,N_38470);
and U40879 (N_40879,N_39221,N_38279);
and U40880 (N_40880,N_39973,N_38995);
nand U40881 (N_40881,N_39514,N_38801);
or U40882 (N_40882,N_38680,N_38622);
nand U40883 (N_40883,N_38093,N_39860);
nor U40884 (N_40884,N_38947,N_38517);
or U40885 (N_40885,N_38386,N_38922);
or U40886 (N_40886,N_38962,N_39651);
and U40887 (N_40887,N_39333,N_39996);
and U40888 (N_40888,N_39398,N_38355);
nor U40889 (N_40889,N_38363,N_38034);
nand U40890 (N_40890,N_39540,N_38803);
nand U40891 (N_40891,N_38214,N_39226);
xnor U40892 (N_40892,N_38722,N_39434);
xnor U40893 (N_40893,N_38503,N_38216);
and U40894 (N_40894,N_38855,N_38699);
or U40895 (N_40895,N_38753,N_38968);
nand U40896 (N_40896,N_38246,N_39084);
nor U40897 (N_40897,N_39312,N_38927);
and U40898 (N_40898,N_39187,N_38426);
xnor U40899 (N_40899,N_39633,N_38601);
nor U40900 (N_40900,N_38518,N_39557);
and U40901 (N_40901,N_38163,N_38218);
or U40902 (N_40902,N_39220,N_39349);
and U40903 (N_40903,N_39185,N_39993);
nor U40904 (N_40904,N_39779,N_38437);
xnor U40905 (N_40905,N_38108,N_39132);
and U40906 (N_40906,N_39238,N_38744);
nor U40907 (N_40907,N_39230,N_38513);
xnor U40908 (N_40908,N_39854,N_38102);
xnor U40909 (N_40909,N_38809,N_39703);
nor U40910 (N_40910,N_38570,N_39445);
xnor U40911 (N_40911,N_38772,N_38212);
nand U40912 (N_40912,N_38101,N_38196);
xnor U40913 (N_40913,N_39824,N_38943);
xor U40914 (N_40914,N_38230,N_39795);
and U40915 (N_40915,N_39948,N_38008);
nand U40916 (N_40916,N_39304,N_38023);
xor U40917 (N_40917,N_38167,N_38624);
or U40918 (N_40918,N_39391,N_38074);
xnor U40919 (N_40919,N_39402,N_39664);
nand U40920 (N_40920,N_39210,N_38342);
nor U40921 (N_40921,N_39876,N_39212);
or U40922 (N_40922,N_39682,N_39408);
nor U40923 (N_40923,N_38824,N_38814);
or U40924 (N_40924,N_39077,N_39436);
nand U40925 (N_40925,N_38324,N_38335);
nor U40926 (N_40926,N_38137,N_38723);
or U40927 (N_40927,N_39610,N_38135);
xor U40928 (N_40928,N_38443,N_39523);
nor U40929 (N_40929,N_39928,N_39414);
nor U40930 (N_40930,N_38720,N_38830);
nor U40931 (N_40931,N_39589,N_38596);
and U40932 (N_40932,N_38274,N_38351);
and U40933 (N_40933,N_39474,N_39802);
or U40934 (N_40934,N_38515,N_39611);
or U40935 (N_40935,N_39670,N_38743);
or U40936 (N_40936,N_38984,N_39362);
and U40937 (N_40937,N_39142,N_38052);
or U40938 (N_40938,N_38957,N_39923);
xnor U40939 (N_40939,N_39835,N_38375);
or U40940 (N_40940,N_39276,N_38350);
xnor U40941 (N_40941,N_39991,N_39576);
or U40942 (N_40942,N_38293,N_39093);
and U40943 (N_40943,N_39700,N_39283);
and U40944 (N_40944,N_38310,N_38971);
xnor U40945 (N_40945,N_39573,N_38174);
or U40946 (N_40946,N_39537,N_39647);
and U40947 (N_40947,N_39599,N_38883);
nor U40948 (N_40948,N_39356,N_38575);
or U40949 (N_40949,N_39318,N_39722);
and U40950 (N_40950,N_39489,N_39600);
and U40951 (N_40951,N_39969,N_39008);
or U40952 (N_40952,N_39873,N_38683);
and U40953 (N_40953,N_39556,N_38653);
nor U40954 (N_40954,N_38391,N_38303);
nand U40955 (N_40955,N_38360,N_39253);
nand U40956 (N_40956,N_38841,N_39183);
nor U40957 (N_40957,N_39531,N_38235);
or U40958 (N_40958,N_39636,N_38454);
and U40959 (N_40959,N_39064,N_39239);
and U40960 (N_40960,N_38433,N_38349);
and U40961 (N_40961,N_39358,N_38076);
xnor U40962 (N_40962,N_38817,N_38746);
or U40963 (N_40963,N_38945,N_38080);
xor U40964 (N_40964,N_39072,N_38065);
or U40965 (N_40965,N_38559,N_38227);
and U40966 (N_40966,N_39535,N_38843);
nor U40967 (N_40967,N_39516,N_38267);
nor U40968 (N_40968,N_38161,N_38691);
xnor U40969 (N_40969,N_38564,N_39719);
or U40970 (N_40970,N_38465,N_38141);
nand U40971 (N_40971,N_38502,N_38579);
xor U40972 (N_40972,N_39929,N_38612);
or U40973 (N_40973,N_38975,N_39657);
nor U40974 (N_40974,N_39688,N_38091);
nor U40975 (N_40975,N_39726,N_39976);
nand U40976 (N_40976,N_38866,N_38178);
and U40977 (N_40977,N_39510,N_39624);
nand U40978 (N_40978,N_39609,N_39496);
and U40979 (N_40979,N_38530,N_38549);
nor U40980 (N_40980,N_39143,N_38941);
xor U40981 (N_40981,N_39552,N_39322);
xor U40982 (N_40982,N_38812,N_38771);
and U40983 (N_40983,N_39840,N_38740);
and U40984 (N_40984,N_38177,N_38565);
nor U40985 (N_40985,N_38970,N_38453);
nor U40986 (N_40986,N_38170,N_38333);
xnor U40987 (N_40987,N_39575,N_38512);
nor U40988 (N_40988,N_38187,N_38329);
nand U40989 (N_40989,N_38409,N_39104);
xor U40990 (N_40990,N_38591,N_39621);
or U40991 (N_40991,N_38103,N_39202);
xnor U40992 (N_40992,N_39897,N_38010);
xnor U40993 (N_40993,N_38410,N_39410);
nor U40994 (N_40994,N_38507,N_39159);
or U40995 (N_40995,N_39452,N_38708);
nand U40996 (N_40996,N_39849,N_39773);
nand U40997 (N_40997,N_39518,N_39870);
or U40998 (N_40998,N_39914,N_38139);
and U40999 (N_40999,N_39481,N_38868);
nand U41000 (N_41000,N_38555,N_38809);
nand U41001 (N_41001,N_39567,N_39192);
nor U41002 (N_41002,N_38622,N_39650);
nand U41003 (N_41003,N_38212,N_39065);
and U41004 (N_41004,N_38075,N_38383);
and U41005 (N_41005,N_38970,N_39919);
xor U41006 (N_41006,N_39331,N_39414);
and U41007 (N_41007,N_38768,N_38495);
and U41008 (N_41008,N_38209,N_39289);
or U41009 (N_41009,N_39083,N_39717);
and U41010 (N_41010,N_38476,N_39869);
xor U41011 (N_41011,N_38193,N_38986);
nand U41012 (N_41012,N_39283,N_39911);
nand U41013 (N_41013,N_39754,N_39200);
nand U41014 (N_41014,N_39755,N_39931);
nor U41015 (N_41015,N_38497,N_39968);
nor U41016 (N_41016,N_38605,N_39731);
or U41017 (N_41017,N_38264,N_39498);
nand U41018 (N_41018,N_39947,N_39345);
xnor U41019 (N_41019,N_38887,N_38807);
and U41020 (N_41020,N_38675,N_38880);
and U41021 (N_41021,N_38317,N_38772);
or U41022 (N_41022,N_38245,N_39409);
nand U41023 (N_41023,N_38401,N_38974);
or U41024 (N_41024,N_39976,N_38729);
nor U41025 (N_41025,N_39012,N_39193);
and U41026 (N_41026,N_39837,N_38513);
nor U41027 (N_41027,N_38791,N_39744);
nand U41028 (N_41028,N_39486,N_39995);
xor U41029 (N_41029,N_38112,N_39854);
or U41030 (N_41030,N_39320,N_39268);
and U41031 (N_41031,N_38443,N_38646);
nor U41032 (N_41032,N_38101,N_38167);
nand U41033 (N_41033,N_38941,N_38484);
and U41034 (N_41034,N_39165,N_39130);
nand U41035 (N_41035,N_38460,N_39080);
nor U41036 (N_41036,N_39008,N_38258);
nor U41037 (N_41037,N_38097,N_38624);
xnor U41038 (N_41038,N_38750,N_39241);
xnor U41039 (N_41039,N_38665,N_38164);
or U41040 (N_41040,N_38638,N_38650);
xnor U41041 (N_41041,N_39649,N_38539);
nand U41042 (N_41042,N_39541,N_39785);
xnor U41043 (N_41043,N_39879,N_39288);
xnor U41044 (N_41044,N_38697,N_38816);
or U41045 (N_41045,N_39975,N_39152);
and U41046 (N_41046,N_39239,N_38487);
nor U41047 (N_41047,N_38785,N_38964);
and U41048 (N_41048,N_38091,N_38182);
and U41049 (N_41049,N_39567,N_38282);
xnor U41050 (N_41050,N_39459,N_38283);
nand U41051 (N_41051,N_38296,N_39079);
or U41052 (N_41052,N_38732,N_38147);
and U41053 (N_41053,N_38518,N_39134);
and U41054 (N_41054,N_39138,N_39896);
nand U41055 (N_41055,N_39912,N_38386);
nand U41056 (N_41056,N_39403,N_39601);
nor U41057 (N_41057,N_39112,N_39534);
and U41058 (N_41058,N_38471,N_38140);
and U41059 (N_41059,N_39396,N_39456);
or U41060 (N_41060,N_38172,N_39858);
xor U41061 (N_41061,N_38224,N_38094);
or U41062 (N_41062,N_38339,N_38330);
xor U41063 (N_41063,N_39700,N_38660);
xnor U41064 (N_41064,N_39181,N_39858);
and U41065 (N_41065,N_38508,N_38082);
xor U41066 (N_41066,N_38979,N_38213);
xor U41067 (N_41067,N_39967,N_39440);
and U41068 (N_41068,N_38327,N_39880);
xnor U41069 (N_41069,N_38001,N_38526);
xor U41070 (N_41070,N_38706,N_38066);
nand U41071 (N_41071,N_39860,N_39414);
nand U41072 (N_41072,N_38633,N_39583);
nor U41073 (N_41073,N_38236,N_38488);
or U41074 (N_41074,N_38991,N_38662);
nand U41075 (N_41075,N_38483,N_39257);
nand U41076 (N_41076,N_38817,N_38365);
nor U41077 (N_41077,N_39811,N_39587);
xor U41078 (N_41078,N_39916,N_38274);
xnor U41079 (N_41079,N_38467,N_39094);
xor U41080 (N_41080,N_38346,N_39356);
and U41081 (N_41081,N_39636,N_39835);
xnor U41082 (N_41082,N_38130,N_39244);
and U41083 (N_41083,N_38447,N_39032);
nor U41084 (N_41084,N_38896,N_39995);
and U41085 (N_41085,N_39162,N_38699);
and U41086 (N_41086,N_39139,N_39378);
nand U41087 (N_41087,N_39725,N_38782);
nor U41088 (N_41088,N_38843,N_38116);
nand U41089 (N_41089,N_39445,N_39045);
or U41090 (N_41090,N_38799,N_39494);
nand U41091 (N_41091,N_38054,N_39657);
xnor U41092 (N_41092,N_38531,N_39381);
or U41093 (N_41093,N_39493,N_38013);
nor U41094 (N_41094,N_38036,N_39286);
or U41095 (N_41095,N_38810,N_38115);
nand U41096 (N_41096,N_38465,N_38941);
nor U41097 (N_41097,N_38080,N_38835);
and U41098 (N_41098,N_39583,N_39276);
xor U41099 (N_41099,N_38032,N_39522);
or U41100 (N_41100,N_38107,N_38784);
nand U41101 (N_41101,N_38667,N_39843);
xnor U41102 (N_41102,N_39313,N_39634);
and U41103 (N_41103,N_39518,N_39379);
xnor U41104 (N_41104,N_39814,N_38503);
xnor U41105 (N_41105,N_38552,N_38370);
nand U41106 (N_41106,N_39835,N_38168);
nor U41107 (N_41107,N_38243,N_39197);
nand U41108 (N_41108,N_39053,N_38286);
or U41109 (N_41109,N_38185,N_39003);
nand U41110 (N_41110,N_39921,N_38830);
nand U41111 (N_41111,N_38521,N_39133);
xnor U41112 (N_41112,N_39986,N_38354);
and U41113 (N_41113,N_39992,N_39084);
and U41114 (N_41114,N_39473,N_38785);
or U41115 (N_41115,N_38669,N_38196);
and U41116 (N_41116,N_38230,N_38072);
or U41117 (N_41117,N_38391,N_38215);
nand U41118 (N_41118,N_39723,N_39499);
nand U41119 (N_41119,N_38015,N_39721);
or U41120 (N_41120,N_39620,N_39418);
nor U41121 (N_41121,N_39619,N_39533);
or U41122 (N_41122,N_38258,N_39589);
and U41123 (N_41123,N_39854,N_38416);
xor U41124 (N_41124,N_39706,N_39328);
and U41125 (N_41125,N_39793,N_38080);
nand U41126 (N_41126,N_38331,N_39171);
xor U41127 (N_41127,N_38356,N_38513);
nor U41128 (N_41128,N_39742,N_39031);
nand U41129 (N_41129,N_38590,N_39733);
and U41130 (N_41130,N_38554,N_38121);
and U41131 (N_41131,N_38414,N_39599);
xor U41132 (N_41132,N_38267,N_39935);
nand U41133 (N_41133,N_39746,N_38856);
nor U41134 (N_41134,N_38568,N_38985);
xnor U41135 (N_41135,N_38424,N_38307);
nor U41136 (N_41136,N_38154,N_39825);
nor U41137 (N_41137,N_38074,N_38259);
xnor U41138 (N_41138,N_39614,N_38428);
xor U41139 (N_41139,N_39250,N_38431);
nor U41140 (N_41140,N_38083,N_38848);
or U41141 (N_41141,N_38016,N_39012);
nor U41142 (N_41142,N_38792,N_38130);
or U41143 (N_41143,N_38088,N_38523);
and U41144 (N_41144,N_38855,N_38445);
nor U41145 (N_41145,N_38910,N_38677);
xor U41146 (N_41146,N_39702,N_38051);
nand U41147 (N_41147,N_38752,N_38822);
nor U41148 (N_41148,N_38640,N_39537);
nand U41149 (N_41149,N_39864,N_39048);
nor U41150 (N_41150,N_39303,N_39825);
or U41151 (N_41151,N_39545,N_38299);
or U41152 (N_41152,N_38370,N_38473);
nand U41153 (N_41153,N_39870,N_39735);
and U41154 (N_41154,N_39075,N_38524);
or U41155 (N_41155,N_39422,N_39768);
or U41156 (N_41156,N_38882,N_38429);
and U41157 (N_41157,N_38698,N_39193);
or U41158 (N_41158,N_38712,N_38631);
or U41159 (N_41159,N_38395,N_39771);
nor U41160 (N_41160,N_38029,N_39582);
nand U41161 (N_41161,N_38943,N_38494);
or U41162 (N_41162,N_38381,N_38493);
or U41163 (N_41163,N_39074,N_38938);
nor U41164 (N_41164,N_39295,N_38523);
nor U41165 (N_41165,N_39342,N_38854);
xor U41166 (N_41166,N_39696,N_38975);
or U41167 (N_41167,N_38239,N_38387);
and U41168 (N_41168,N_38668,N_38448);
nand U41169 (N_41169,N_38601,N_39855);
nor U41170 (N_41170,N_38419,N_39941);
or U41171 (N_41171,N_38217,N_39160);
nor U41172 (N_41172,N_38903,N_38545);
and U41173 (N_41173,N_39441,N_38539);
nand U41174 (N_41174,N_39213,N_39230);
xnor U41175 (N_41175,N_39815,N_39193);
or U41176 (N_41176,N_39303,N_39292);
nor U41177 (N_41177,N_38334,N_38897);
xnor U41178 (N_41178,N_38777,N_39848);
nand U41179 (N_41179,N_38731,N_39419);
nand U41180 (N_41180,N_38795,N_38558);
and U41181 (N_41181,N_38782,N_38521);
or U41182 (N_41182,N_38134,N_38549);
nand U41183 (N_41183,N_39292,N_38509);
and U41184 (N_41184,N_39729,N_39610);
nor U41185 (N_41185,N_39741,N_39590);
and U41186 (N_41186,N_39018,N_39072);
xnor U41187 (N_41187,N_39149,N_39035);
xnor U41188 (N_41188,N_38779,N_39328);
and U41189 (N_41189,N_38236,N_38535);
or U41190 (N_41190,N_38540,N_39748);
nand U41191 (N_41191,N_38555,N_38162);
nor U41192 (N_41192,N_39792,N_39762);
and U41193 (N_41193,N_38960,N_38588);
and U41194 (N_41194,N_39271,N_38674);
nand U41195 (N_41195,N_38169,N_38085);
or U41196 (N_41196,N_38207,N_39295);
and U41197 (N_41197,N_38298,N_39226);
nand U41198 (N_41198,N_39422,N_39711);
or U41199 (N_41199,N_39447,N_38445);
xnor U41200 (N_41200,N_39511,N_38808);
and U41201 (N_41201,N_38950,N_38340);
or U41202 (N_41202,N_38981,N_38208);
xor U41203 (N_41203,N_38226,N_39707);
or U41204 (N_41204,N_39949,N_38132);
nor U41205 (N_41205,N_39186,N_38886);
nor U41206 (N_41206,N_39946,N_39084);
and U41207 (N_41207,N_38099,N_39217);
xor U41208 (N_41208,N_38735,N_39797);
or U41209 (N_41209,N_38223,N_39765);
xnor U41210 (N_41210,N_39668,N_38378);
and U41211 (N_41211,N_38975,N_38852);
nand U41212 (N_41212,N_39901,N_38717);
nor U41213 (N_41213,N_39369,N_39503);
and U41214 (N_41214,N_38255,N_38322);
or U41215 (N_41215,N_39532,N_38941);
nor U41216 (N_41216,N_38505,N_38821);
or U41217 (N_41217,N_38446,N_39917);
xnor U41218 (N_41218,N_38318,N_38287);
and U41219 (N_41219,N_39353,N_38955);
or U41220 (N_41220,N_38357,N_39991);
and U41221 (N_41221,N_39014,N_39557);
nand U41222 (N_41222,N_39774,N_39679);
nand U41223 (N_41223,N_38169,N_38608);
nand U41224 (N_41224,N_38879,N_38091);
nor U41225 (N_41225,N_39439,N_38764);
xor U41226 (N_41226,N_38875,N_39972);
or U41227 (N_41227,N_39767,N_38215);
nand U41228 (N_41228,N_38185,N_39476);
and U41229 (N_41229,N_39603,N_39033);
xnor U41230 (N_41230,N_39919,N_39905);
nor U41231 (N_41231,N_38655,N_39315);
xnor U41232 (N_41232,N_38885,N_38100);
and U41233 (N_41233,N_39601,N_38633);
nor U41234 (N_41234,N_39032,N_39994);
nor U41235 (N_41235,N_38274,N_38166);
and U41236 (N_41236,N_38957,N_38409);
nand U41237 (N_41237,N_38308,N_38439);
nand U41238 (N_41238,N_38088,N_38020);
nor U41239 (N_41239,N_39330,N_39927);
nor U41240 (N_41240,N_38356,N_38343);
or U41241 (N_41241,N_39238,N_38573);
nand U41242 (N_41242,N_39736,N_39501);
xnor U41243 (N_41243,N_39355,N_38121);
and U41244 (N_41244,N_38438,N_39622);
xnor U41245 (N_41245,N_39794,N_38548);
or U41246 (N_41246,N_39166,N_38236);
nand U41247 (N_41247,N_39930,N_39608);
xor U41248 (N_41248,N_39440,N_38459);
or U41249 (N_41249,N_38867,N_38831);
or U41250 (N_41250,N_38867,N_38035);
nor U41251 (N_41251,N_39106,N_39783);
nor U41252 (N_41252,N_39738,N_39280);
nor U41253 (N_41253,N_39843,N_38425);
and U41254 (N_41254,N_38639,N_38527);
and U41255 (N_41255,N_39174,N_39756);
nand U41256 (N_41256,N_38868,N_38821);
and U41257 (N_41257,N_38769,N_38124);
nand U41258 (N_41258,N_39462,N_38081);
xnor U41259 (N_41259,N_39613,N_38560);
nor U41260 (N_41260,N_39893,N_39512);
xor U41261 (N_41261,N_38386,N_39895);
or U41262 (N_41262,N_38671,N_39399);
or U41263 (N_41263,N_38242,N_39721);
nand U41264 (N_41264,N_38299,N_39913);
and U41265 (N_41265,N_38780,N_39558);
or U41266 (N_41266,N_39422,N_39287);
nand U41267 (N_41267,N_38302,N_39910);
nor U41268 (N_41268,N_38257,N_39598);
or U41269 (N_41269,N_38381,N_39968);
nand U41270 (N_41270,N_39716,N_38507);
or U41271 (N_41271,N_38777,N_38764);
xnor U41272 (N_41272,N_38701,N_39503);
xor U41273 (N_41273,N_39407,N_39431);
nand U41274 (N_41274,N_38785,N_39357);
nand U41275 (N_41275,N_39731,N_38925);
nand U41276 (N_41276,N_39203,N_39639);
xnor U41277 (N_41277,N_38227,N_39910);
xnor U41278 (N_41278,N_39192,N_38529);
and U41279 (N_41279,N_38139,N_38971);
and U41280 (N_41280,N_38512,N_38191);
nor U41281 (N_41281,N_38703,N_39664);
xor U41282 (N_41282,N_38612,N_38905);
xor U41283 (N_41283,N_38351,N_38835);
nand U41284 (N_41284,N_38379,N_38593);
or U41285 (N_41285,N_38617,N_39088);
xnor U41286 (N_41286,N_39172,N_39005);
and U41287 (N_41287,N_38157,N_39502);
or U41288 (N_41288,N_38649,N_39546);
or U41289 (N_41289,N_38510,N_39560);
or U41290 (N_41290,N_39835,N_38986);
or U41291 (N_41291,N_39385,N_39971);
nor U41292 (N_41292,N_38778,N_38922);
nor U41293 (N_41293,N_39892,N_39572);
or U41294 (N_41294,N_38311,N_39336);
xor U41295 (N_41295,N_38157,N_39090);
xor U41296 (N_41296,N_39555,N_39984);
and U41297 (N_41297,N_38378,N_39169);
nand U41298 (N_41298,N_39583,N_39423);
xor U41299 (N_41299,N_38408,N_39797);
and U41300 (N_41300,N_39549,N_38510);
or U41301 (N_41301,N_39796,N_38258);
nand U41302 (N_41302,N_39970,N_39319);
and U41303 (N_41303,N_38727,N_38222);
nand U41304 (N_41304,N_39320,N_39373);
nand U41305 (N_41305,N_39286,N_38042);
and U41306 (N_41306,N_39533,N_38114);
nand U41307 (N_41307,N_38854,N_38623);
nand U41308 (N_41308,N_39793,N_39370);
or U41309 (N_41309,N_38634,N_38654);
and U41310 (N_41310,N_39989,N_39415);
or U41311 (N_41311,N_38644,N_38169);
nand U41312 (N_41312,N_38354,N_39139);
nand U41313 (N_41313,N_38910,N_38938);
or U41314 (N_41314,N_38806,N_39135);
xor U41315 (N_41315,N_39633,N_39281);
xor U41316 (N_41316,N_38266,N_39178);
xor U41317 (N_41317,N_38527,N_39717);
xnor U41318 (N_41318,N_38759,N_39672);
nor U41319 (N_41319,N_38130,N_38289);
nand U41320 (N_41320,N_39344,N_38633);
xor U41321 (N_41321,N_38215,N_38277);
and U41322 (N_41322,N_39355,N_39213);
and U41323 (N_41323,N_39306,N_39601);
nand U41324 (N_41324,N_38156,N_38723);
nor U41325 (N_41325,N_39307,N_39752);
and U41326 (N_41326,N_39624,N_38724);
xor U41327 (N_41327,N_38483,N_39295);
nand U41328 (N_41328,N_39587,N_38648);
and U41329 (N_41329,N_38030,N_38620);
nor U41330 (N_41330,N_38903,N_38384);
nor U41331 (N_41331,N_39823,N_39453);
or U41332 (N_41332,N_38994,N_39883);
and U41333 (N_41333,N_38298,N_38740);
nor U41334 (N_41334,N_39224,N_39543);
nor U41335 (N_41335,N_39469,N_39297);
xnor U41336 (N_41336,N_38381,N_39720);
nor U41337 (N_41337,N_39403,N_39533);
nor U41338 (N_41338,N_38728,N_38863);
nand U41339 (N_41339,N_39240,N_38570);
and U41340 (N_41340,N_38281,N_39257);
xnor U41341 (N_41341,N_38235,N_38576);
and U41342 (N_41342,N_39547,N_39779);
or U41343 (N_41343,N_39754,N_38982);
xor U41344 (N_41344,N_39524,N_38245);
or U41345 (N_41345,N_38842,N_39867);
nor U41346 (N_41346,N_38484,N_38313);
nand U41347 (N_41347,N_39454,N_39133);
nor U41348 (N_41348,N_38463,N_38170);
xor U41349 (N_41349,N_39173,N_38882);
nor U41350 (N_41350,N_39681,N_38862);
and U41351 (N_41351,N_38361,N_39942);
xor U41352 (N_41352,N_38541,N_39789);
nand U41353 (N_41353,N_39145,N_38303);
nor U41354 (N_41354,N_38905,N_39503);
nand U41355 (N_41355,N_38434,N_39962);
xnor U41356 (N_41356,N_39995,N_38827);
xor U41357 (N_41357,N_38742,N_39790);
xnor U41358 (N_41358,N_38686,N_39586);
or U41359 (N_41359,N_38327,N_39963);
xor U41360 (N_41360,N_39809,N_39943);
xor U41361 (N_41361,N_38240,N_38943);
nor U41362 (N_41362,N_39286,N_39830);
and U41363 (N_41363,N_39361,N_38470);
nor U41364 (N_41364,N_39350,N_38959);
xnor U41365 (N_41365,N_38864,N_39805);
or U41366 (N_41366,N_38841,N_39727);
or U41367 (N_41367,N_39465,N_39193);
or U41368 (N_41368,N_39810,N_38158);
nand U41369 (N_41369,N_39424,N_38408);
xor U41370 (N_41370,N_38701,N_38909);
or U41371 (N_41371,N_38189,N_38347);
xnor U41372 (N_41372,N_39297,N_39753);
or U41373 (N_41373,N_38810,N_38019);
and U41374 (N_41374,N_38717,N_39113);
and U41375 (N_41375,N_38494,N_39889);
or U41376 (N_41376,N_38615,N_39695);
xnor U41377 (N_41377,N_38797,N_38088);
xnor U41378 (N_41378,N_38142,N_39639);
nor U41379 (N_41379,N_39697,N_38643);
xor U41380 (N_41380,N_38493,N_39353);
and U41381 (N_41381,N_39302,N_38840);
or U41382 (N_41382,N_38497,N_38845);
or U41383 (N_41383,N_38672,N_38880);
or U41384 (N_41384,N_38642,N_39652);
and U41385 (N_41385,N_39511,N_38547);
xnor U41386 (N_41386,N_38088,N_38739);
nand U41387 (N_41387,N_38075,N_38277);
xnor U41388 (N_41388,N_38327,N_38608);
or U41389 (N_41389,N_39277,N_39036);
or U41390 (N_41390,N_38382,N_39162);
xor U41391 (N_41391,N_39290,N_38723);
or U41392 (N_41392,N_39629,N_38909);
and U41393 (N_41393,N_39817,N_39693);
and U41394 (N_41394,N_39890,N_39840);
nor U41395 (N_41395,N_39052,N_39045);
nand U41396 (N_41396,N_38652,N_39105);
or U41397 (N_41397,N_39582,N_39625);
xnor U41398 (N_41398,N_38960,N_39527);
and U41399 (N_41399,N_39665,N_39813);
or U41400 (N_41400,N_38128,N_38327);
xor U41401 (N_41401,N_38148,N_39034);
and U41402 (N_41402,N_39169,N_38790);
xor U41403 (N_41403,N_39554,N_38375);
and U41404 (N_41404,N_38214,N_38501);
xnor U41405 (N_41405,N_39374,N_38917);
xnor U41406 (N_41406,N_39115,N_38766);
xnor U41407 (N_41407,N_38455,N_38165);
nand U41408 (N_41408,N_39683,N_38011);
or U41409 (N_41409,N_39878,N_39644);
and U41410 (N_41410,N_39026,N_39041);
nand U41411 (N_41411,N_38289,N_38463);
nand U41412 (N_41412,N_38144,N_38954);
and U41413 (N_41413,N_38078,N_38926);
or U41414 (N_41414,N_39199,N_39347);
nand U41415 (N_41415,N_39593,N_38701);
nor U41416 (N_41416,N_39094,N_39896);
or U41417 (N_41417,N_39051,N_38087);
and U41418 (N_41418,N_39678,N_39464);
and U41419 (N_41419,N_38377,N_39402);
nor U41420 (N_41420,N_39164,N_39124);
nor U41421 (N_41421,N_38559,N_38238);
or U41422 (N_41422,N_38424,N_38345);
or U41423 (N_41423,N_39264,N_38798);
nand U41424 (N_41424,N_39868,N_39283);
or U41425 (N_41425,N_39138,N_38353);
or U41426 (N_41426,N_39334,N_38473);
nor U41427 (N_41427,N_39321,N_38566);
xnor U41428 (N_41428,N_38940,N_38565);
or U41429 (N_41429,N_39860,N_38027);
and U41430 (N_41430,N_38212,N_38892);
nor U41431 (N_41431,N_39093,N_38239);
and U41432 (N_41432,N_39058,N_38499);
and U41433 (N_41433,N_39635,N_38610);
or U41434 (N_41434,N_39396,N_38049);
nor U41435 (N_41435,N_38742,N_38052);
nand U41436 (N_41436,N_39662,N_39064);
xor U41437 (N_41437,N_39481,N_39005);
and U41438 (N_41438,N_38336,N_39128);
or U41439 (N_41439,N_39181,N_39055);
or U41440 (N_41440,N_39158,N_39457);
or U41441 (N_41441,N_39254,N_39027);
or U41442 (N_41442,N_39864,N_38904);
or U41443 (N_41443,N_38053,N_39662);
nor U41444 (N_41444,N_39370,N_39143);
nor U41445 (N_41445,N_38223,N_39052);
xor U41446 (N_41446,N_39172,N_38024);
xnor U41447 (N_41447,N_38073,N_39801);
nor U41448 (N_41448,N_39512,N_38817);
nor U41449 (N_41449,N_39368,N_39728);
nor U41450 (N_41450,N_38588,N_38514);
nor U41451 (N_41451,N_38601,N_39942);
nor U41452 (N_41452,N_39433,N_39251);
and U41453 (N_41453,N_38540,N_38650);
nor U41454 (N_41454,N_38964,N_38447);
or U41455 (N_41455,N_39320,N_38460);
xnor U41456 (N_41456,N_39899,N_39000);
nor U41457 (N_41457,N_38811,N_39611);
nor U41458 (N_41458,N_38850,N_38612);
nand U41459 (N_41459,N_38177,N_38861);
and U41460 (N_41460,N_38120,N_39712);
and U41461 (N_41461,N_39288,N_38282);
nand U41462 (N_41462,N_38445,N_39297);
xor U41463 (N_41463,N_38593,N_38793);
xnor U41464 (N_41464,N_39885,N_38364);
and U41465 (N_41465,N_38361,N_38260);
or U41466 (N_41466,N_38960,N_39715);
and U41467 (N_41467,N_38233,N_39186);
and U41468 (N_41468,N_39872,N_39966);
and U41469 (N_41469,N_38071,N_39269);
nor U41470 (N_41470,N_38694,N_39321);
and U41471 (N_41471,N_38574,N_38803);
xnor U41472 (N_41472,N_39238,N_38663);
nor U41473 (N_41473,N_38352,N_38924);
xnor U41474 (N_41474,N_38112,N_38294);
xnor U41475 (N_41475,N_38246,N_38057);
nor U41476 (N_41476,N_38379,N_39951);
or U41477 (N_41477,N_38094,N_39956);
nor U41478 (N_41478,N_38743,N_38256);
or U41479 (N_41479,N_38456,N_38064);
nor U41480 (N_41480,N_38788,N_39297);
nand U41481 (N_41481,N_39462,N_39348);
or U41482 (N_41482,N_39283,N_38143);
xnor U41483 (N_41483,N_39121,N_39167);
xor U41484 (N_41484,N_38252,N_38082);
nor U41485 (N_41485,N_38265,N_39371);
and U41486 (N_41486,N_38665,N_39048);
nand U41487 (N_41487,N_39070,N_39772);
and U41488 (N_41488,N_39800,N_39789);
and U41489 (N_41489,N_39970,N_39218);
and U41490 (N_41490,N_38040,N_39966);
nor U41491 (N_41491,N_39602,N_38489);
and U41492 (N_41492,N_38281,N_39718);
or U41493 (N_41493,N_38456,N_39885);
or U41494 (N_41494,N_38402,N_39591);
nor U41495 (N_41495,N_38940,N_39291);
nand U41496 (N_41496,N_39128,N_38728);
nand U41497 (N_41497,N_38810,N_38108);
xor U41498 (N_41498,N_39439,N_39070);
and U41499 (N_41499,N_39191,N_39485);
xor U41500 (N_41500,N_38360,N_39084);
xnor U41501 (N_41501,N_39626,N_38385);
xor U41502 (N_41502,N_39242,N_39518);
nand U41503 (N_41503,N_38253,N_38039);
xor U41504 (N_41504,N_38757,N_38931);
and U41505 (N_41505,N_38146,N_39606);
xnor U41506 (N_41506,N_38035,N_38905);
and U41507 (N_41507,N_39462,N_39854);
xnor U41508 (N_41508,N_39456,N_39874);
and U41509 (N_41509,N_38978,N_39839);
nor U41510 (N_41510,N_38618,N_38827);
and U41511 (N_41511,N_39549,N_39051);
nor U41512 (N_41512,N_39075,N_39910);
nand U41513 (N_41513,N_38219,N_39243);
nor U41514 (N_41514,N_39026,N_38088);
nand U41515 (N_41515,N_38343,N_39864);
and U41516 (N_41516,N_39632,N_39920);
nand U41517 (N_41517,N_39135,N_39922);
nand U41518 (N_41518,N_38953,N_38594);
xor U41519 (N_41519,N_38268,N_39362);
or U41520 (N_41520,N_38920,N_38938);
xnor U41521 (N_41521,N_39320,N_38798);
and U41522 (N_41522,N_39476,N_39647);
and U41523 (N_41523,N_38307,N_39953);
nand U41524 (N_41524,N_39201,N_38451);
xnor U41525 (N_41525,N_38845,N_39112);
and U41526 (N_41526,N_38078,N_38986);
nor U41527 (N_41527,N_39022,N_39981);
nor U41528 (N_41528,N_39363,N_38738);
nand U41529 (N_41529,N_38835,N_38370);
nor U41530 (N_41530,N_38790,N_39960);
or U41531 (N_41531,N_39319,N_38995);
or U41532 (N_41532,N_39348,N_39430);
nand U41533 (N_41533,N_38844,N_38392);
or U41534 (N_41534,N_39864,N_39630);
nor U41535 (N_41535,N_38866,N_39239);
or U41536 (N_41536,N_38511,N_39855);
or U41537 (N_41537,N_39433,N_38727);
xor U41538 (N_41538,N_39349,N_38244);
nand U41539 (N_41539,N_39260,N_39402);
and U41540 (N_41540,N_39725,N_39648);
nand U41541 (N_41541,N_38878,N_39804);
or U41542 (N_41542,N_39392,N_38909);
nand U41543 (N_41543,N_38477,N_39165);
and U41544 (N_41544,N_38749,N_39943);
nor U41545 (N_41545,N_38671,N_39577);
and U41546 (N_41546,N_38193,N_39188);
nor U41547 (N_41547,N_38239,N_39679);
or U41548 (N_41548,N_39808,N_39505);
and U41549 (N_41549,N_38708,N_38966);
nor U41550 (N_41550,N_38671,N_38709);
nor U41551 (N_41551,N_38464,N_38474);
nor U41552 (N_41552,N_39846,N_39305);
xor U41553 (N_41553,N_39529,N_39306);
nor U41554 (N_41554,N_38156,N_39682);
nand U41555 (N_41555,N_38598,N_38619);
nor U41556 (N_41556,N_38281,N_39695);
xor U41557 (N_41557,N_38004,N_39481);
xor U41558 (N_41558,N_38595,N_38045);
or U41559 (N_41559,N_39953,N_39889);
or U41560 (N_41560,N_39333,N_39271);
nand U41561 (N_41561,N_38222,N_38509);
nand U41562 (N_41562,N_39505,N_39221);
nor U41563 (N_41563,N_39925,N_39969);
nand U41564 (N_41564,N_39553,N_39911);
xnor U41565 (N_41565,N_39167,N_38413);
and U41566 (N_41566,N_38026,N_38557);
nor U41567 (N_41567,N_38460,N_39093);
and U41568 (N_41568,N_39264,N_38203);
and U41569 (N_41569,N_38510,N_39652);
nand U41570 (N_41570,N_39617,N_38179);
and U41571 (N_41571,N_39288,N_39386);
or U41572 (N_41572,N_39206,N_39441);
and U41573 (N_41573,N_38003,N_39316);
or U41574 (N_41574,N_39602,N_39502);
xnor U41575 (N_41575,N_39916,N_38284);
nand U41576 (N_41576,N_38608,N_39134);
and U41577 (N_41577,N_38981,N_38194);
nand U41578 (N_41578,N_39419,N_38651);
nand U41579 (N_41579,N_39912,N_38466);
nor U41580 (N_41580,N_39488,N_39906);
nor U41581 (N_41581,N_38578,N_39486);
nor U41582 (N_41582,N_39939,N_39492);
or U41583 (N_41583,N_39421,N_38603);
nand U41584 (N_41584,N_38634,N_38597);
and U41585 (N_41585,N_39268,N_39436);
and U41586 (N_41586,N_39536,N_39841);
or U41587 (N_41587,N_39982,N_39143);
or U41588 (N_41588,N_39156,N_38283);
or U41589 (N_41589,N_38245,N_39701);
or U41590 (N_41590,N_39348,N_39094);
and U41591 (N_41591,N_39737,N_38251);
xor U41592 (N_41592,N_38936,N_38241);
nor U41593 (N_41593,N_39097,N_38354);
nand U41594 (N_41594,N_38731,N_39172);
nor U41595 (N_41595,N_39913,N_39514);
nor U41596 (N_41596,N_38781,N_39508);
nor U41597 (N_41597,N_38961,N_38784);
nor U41598 (N_41598,N_39838,N_39769);
nand U41599 (N_41599,N_38023,N_39603);
nand U41600 (N_41600,N_39333,N_39569);
and U41601 (N_41601,N_38894,N_38875);
or U41602 (N_41602,N_38811,N_39473);
nand U41603 (N_41603,N_39562,N_38177);
or U41604 (N_41604,N_39919,N_38110);
or U41605 (N_41605,N_38285,N_38127);
xor U41606 (N_41606,N_38796,N_39456);
xnor U41607 (N_41607,N_38360,N_39876);
xnor U41608 (N_41608,N_38053,N_39217);
nand U41609 (N_41609,N_38943,N_39578);
nor U41610 (N_41610,N_39341,N_38600);
and U41611 (N_41611,N_39687,N_38110);
or U41612 (N_41612,N_38188,N_38861);
nor U41613 (N_41613,N_39346,N_38856);
and U41614 (N_41614,N_38292,N_38475);
nand U41615 (N_41615,N_38426,N_39468);
nand U41616 (N_41616,N_39359,N_38832);
and U41617 (N_41617,N_38134,N_39693);
and U41618 (N_41618,N_38314,N_38522);
nand U41619 (N_41619,N_38416,N_38775);
nor U41620 (N_41620,N_39155,N_38327);
nor U41621 (N_41621,N_38444,N_39159);
and U41622 (N_41622,N_39764,N_38068);
nand U41623 (N_41623,N_39560,N_38912);
xor U41624 (N_41624,N_39421,N_38827);
nor U41625 (N_41625,N_38960,N_38346);
or U41626 (N_41626,N_38781,N_39284);
and U41627 (N_41627,N_39997,N_38276);
nand U41628 (N_41628,N_38374,N_39964);
nand U41629 (N_41629,N_39039,N_38166);
and U41630 (N_41630,N_38092,N_38087);
nor U41631 (N_41631,N_38162,N_39930);
or U41632 (N_41632,N_39143,N_38637);
nor U41633 (N_41633,N_39190,N_39368);
xnor U41634 (N_41634,N_39505,N_38662);
nor U41635 (N_41635,N_38607,N_39711);
xor U41636 (N_41636,N_39835,N_39185);
nor U41637 (N_41637,N_38371,N_38721);
or U41638 (N_41638,N_38050,N_38656);
nand U41639 (N_41639,N_38300,N_38196);
nand U41640 (N_41640,N_38681,N_38511);
xnor U41641 (N_41641,N_39573,N_38711);
nor U41642 (N_41642,N_39347,N_38759);
or U41643 (N_41643,N_38031,N_39420);
nand U41644 (N_41644,N_38733,N_39480);
nor U41645 (N_41645,N_38994,N_38135);
nor U41646 (N_41646,N_39439,N_39978);
or U41647 (N_41647,N_38306,N_38105);
nor U41648 (N_41648,N_38202,N_39156);
nand U41649 (N_41649,N_38694,N_38903);
xnor U41650 (N_41650,N_38503,N_38777);
nand U41651 (N_41651,N_38617,N_39502);
nand U41652 (N_41652,N_38750,N_39578);
nand U41653 (N_41653,N_39010,N_38707);
and U41654 (N_41654,N_39846,N_39385);
xor U41655 (N_41655,N_39419,N_38668);
or U41656 (N_41656,N_39516,N_38484);
nor U41657 (N_41657,N_38001,N_38818);
nand U41658 (N_41658,N_38104,N_39277);
xnor U41659 (N_41659,N_38947,N_38861);
xnor U41660 (N_41660,N_39143,N_39694);
nor U41661 (N_41661,N_39548,N_39004);
nand U41662 (N_41662,N_39227,N_38548);
xnor U41663 (N_41663,N_39604,N_39333);
or U41664 (N_41664,N_39123,N_38050);
nand U41665 (N_41665,N_39407,N_39294);
xnor U41666 (N_41666,N_38084,N_39221);
nor U41667 (N_41667,N_39763,N_39793);
or U41668 (N_41668,N_39964,N_39305);
nor U41669 (N_41669,N_39398,N_38396);
and U41670 (N_41670,N_39596,N_38637);
and U41671 (N_41671,N_38658,N_38431);
and U41672 (N_41672,N_39424,N_39352);
nor U41673 (N_41673,N_38208,N_39925);
nand U41674 (N_41674,N_38907,N_39078);
nor U41675 (N_41675,N_39469,N_38290);
nand U41676 (N_41676,N_38766,N_39313);
or U41677 (N_41677,N_38359,N_39015);
xor U41678 (N_41678,N_38243,N_38250);
nand U41679 (N_41679,N_38535,N_39751);
nand U41680 (N_41680,N_38259,N_39395);
nand U41681 (N_41681,N_38613,N_38961);
and U41682 (N_41682,N_39919,N_39385);
nand U41683 (N_41683,N_39573,N_39870);
and U41684 (N_41684,N_38206,N_38981);
or U41685 (N_41685,N_39496,N_38041);
and U41686 (N_41686,N_38177,N_39135);
and U41687 (N_41687,N_39912,N_38600);
nor U41688 (N_41688,N_38204,N_38160);
nand U41689 (N_41689,N_39052,N_39545);
xnor U41690 (N_41690,N_39231,N_38332);
and U41691 (N_41691,N_39338,N_39298);
and U41692 (N_41692,N_39070,N_38233);
or U41693 (N_41693,N_38604,N_38631);
or U41694 (N_41694,N_38658,N_38683);
or U41695 (N_41695,N_39679,N_38982);
or U41696 (N_41696,N_38893,N_39992);
nand U41697 (N_41697,N_38815,N_39332);
nand U41698 (N_41698,N_39240,N_39900);
nor U41699 (N_41699,N_39271,N_39936);
or U41700 (N_41700,N_39037,N_38511);
and U41701 (N_41701,N_38515,N_39755);
and U41702 (N_41702,N_38982,N_39346);
nand U41703 (N_41703,N_39408,N_39374);
xor U41704 (N_41704,N_38179,N_39562);
nand U41705 (N_41705,N_39496,N_38202);
nand U41706 (N_41706,N_39966,N_38400);
nor U41707 (N_41707,N_39507,N_39731);
nand U41708 (N_41708,N_39703,N_39074);
or U41709 (N_41709,N_38576,N_38919);
nand U41710 (N_41710,N_39388,N_39575);
nor U41711 (N_41711,N_38466,N_39662);
nor U41712 (N_41712,N_38294,N_39224);
nor U41713 (N_41713,N_39066,N_38556);
nand U41714 (N_41714,N_38148,N_39906);
nor U41715 (N_41715,N_38000,N_38911);
nand U41716 (N_41716,N_39517,N_38955);
nor U41717 (N_41717,N_38067,N_39902);
xnor U41718 (N_41718,N_39665,N_39150);
nand U41719 (N_41719,N_39405,N_38649);
and U41720 (N_41720,N_38979,N_39907);
nor U41721 (N_41721,N_38886,N_38802);
xor U41722 (N_41722,N_39632,N_38876);
nand U41723 (N_41723,N_38378,N_38332);
xor U41724 (N_41724,N_38494,N_38322);
nand U41725 (N_41725,N_38073,N_38405);
or U41726 (N_41726,N_39297,N_39793);
nor U41727 (N_41727,N_39973,N_39956);
xnor U41728 (N_41728,N_38794,N_39967);
nor U41729 (N_41729,N_39852,N_39606);
and U41730 (N_41730,N_38138,N_38876);
and U41731 (N_41731,N_39085,N_39049);
nand U41732 (N_41732,N_39741,N_39908);
nand U41733 (N_41733,N_39054,N_39176);
or U41734 (N_41734,N_38988,N_39027);
or U41735 (N_41735,N_39812,N_39172);
nor U41736 (N_41736,N_39310,N_38593);
and U41737 (N_41737,N_38377,N_38283);
nor U41738 (N_41738,N_38535,N_38388);
nor U41739 (N_41739,N_39445,N_38682);
nor U41740 (N_41740,N_39841,N_38138);
xor U41741 (N_41741,N_38902,N_38814);
xnor U41742 (N_41742,N_38495,N_38207);
nand U41743 (N_41743,N_39073,N_39564);
nand U41744 (N_41744,N_38980,N_38681);
nor U41745 (N_41745,N_38998,N_39959);
or U41746 (N_41746,N_39516,N_38142);
or U41747 (N_41747,N_38901,N_39365);
nor U41748 (N_41748,N_38001,N_38248);
and U41749 (N_41749,N_39172,N_38667);
and U41750 (N_41750,N_38423,N_39757);
nand U41751 (N_41751,N_39767,N_38113);
xor U41752 (N_41752,N_39516,N_39565);
xnor U41753 (N_41753,N_39828,N_39084);
xnor U41754 (N_41754,N_38744,N_38388);
xor U41755 (N_41755,N_39641,N_38170);
or U41756 (N_41756,N_39080,N_38395);
and U41757 (N_41757,N_39267,N_38419);
or U41758 (N_41758,N_39618,N_39038);
nor U41759 (N_41759,N_38053,N_39718);
xnor U41760 (N_41760,N_39195,N_39235);
and U41761 (N_41761,N_39983,N_39474);
nor U41762 (N_41762,N_38330,N_38181);
nand U41763 (N_41763,N_39373,N_39509);
nand U41764 (N_41764,N_38907,N_39967);
nor U41765 (N_41765,N_38218,N_39089);
or U41766 (N_41766,N_38959,N_38019);
nor U41767 (N_41767,N_39773,N_38968);
nor U41768 (N_41768,N_39145,N_39844);
xor U41769 (N_41769,N_38266,N_38591);
and U41770 (N_41770,N_38747,N_39725);
or U41771 (N_41771,N_39385,N_38264);
nor U41772 (N_41772,N_38738,N_38065);
nand U41773 (N_41773,N_39220,N_38116);
xor U41774 (N_41774,N_39808,N_39730);
nand U41775 (N_41775,N_39738,N_38128);
or U41776 (N_41776,N_39005,N_38805);
nor U41777 (N_41777,N_38759,N_39568);
xor U41778 (N_41778,N_39002,N_38168);
and U41779 (N_41779,N_39804,N_38501);
and U41780 (N_41780,N_39305,N_38676);
or U41781 (N_41781,N_38858,N_38294);
nor U41782 (N_41782,N_38892,N_38097);
or U41783 (N_41783,N_39946,N_38107);
nand U41784 (N_41784,N_39022,N_39827);
xor U41785 (N_41785,N_38494,N_38090);
nor U41786 (N_41786,N_39018,N_38972);
nor U41787 (N_41787,N_38525,N_39886);
xor U41788 (N_41788,N_38168,N_38564);
nand U41789 (N_41789,N_39713,N_39774);
nand U41790 (N_41790,N_38935,N_39671);
xor U41791 (N_41791,N_39725,N_38663);
nor U41792 (N_41792,N_38949,N_38756);
nor U41793 (N_41793,N_39491,N_39991);
nor U41794 (N_41794,N_39007,N_38212);
xor U41795 (N_41795,N_38482,N_39194);
or U41796 (N_41796,N_38908,N_38887);
xor U41797 (N_41797,N_39611,N_38808);
nor U41798 (N_41798,N_39546,N_38625);
nor U41799 (N_41799,N_38620,N_39453);
or U41800 (N_41800,N_39001,N_39203);
or U41801 (N_41801,N_38020,N_38226);
nor U41802 (N_41802,N_38172,N_39694);
or U41803 (N_41803,N_38736,N_38319);
nand U41804 (N_41804,N_39906,N_39390);
or U41805 (N_41805,N_38028,N_39448);
nand U41806 (N_41806,N_39698,N_38565);
nor U41807 (N_41807,N_39670,N_38805);
nor U41808 (N_41808,N_38696,N_38755);
or U41809 (N_41809,N_38830,N_39007);
nand U41810 (N_41810,N_39825,N_39172);
nor U41811 (N_41811,N_39359,N_39102);
or U41812 (N_41812,N_39580,N_38392);
nor U41813 (N_41813,N_39613,N_39412);
nand U41814 (N_41814,N_39011,N_38942);
nand U41815 (N_41815,N_39013,N_39463);
or U41816 (N_41816,N_38137,N_39612);
or U41817 (N_41817,N_38424,N_38769);
nand U41818 (N_41818,N_38164,N_38446);
nor U41819 (N_41819,N_39797,N_38971);
and U41820 (N_41820,N_39234,N_39187);
and U41821 (N_41821,N_39336,N_39488);
nand U41822 (N_41822,N_39450,N_39388);
xor U41823 (N_41823,N_39232,N_39503);
nand U41824 (N_41824,N_39778,N_39178);
or U41825 (N_41825,N_38382,N_38218);
or U41826 (N_41826,N_38548,N_38482);
or U41827 (N_41827,N_39878,N_39307);
nor U41828 (N_41828,N_39585,N_38309);
and U41829 (N_41829,N_38595,N_39772);
xnor U41830 (N_41830,N_39898,N_38108);
or U41831 (N_41831,N_38756,N_39336);
and U41832 (N_41832,N_39859,N_39056);
nand U41833 (N_41833,N_38079,N_38962);
or U41834 (N_41834,N_39427,N_38031);
nand U41835 (N_41835,N_39474,N_38932);
nand U41836 (N_41836,N_38297,N_39353);
xnor U41837 (N_41837,N_39662,N_38228);
and U41838 (N_41838,N_38617,N_38005);
and U41839 (N_41839,N_38235,N_38660);
xnor U41840 (N_41840,N_38834,N_39508);
xor U41841 (N_41841,N_38789,N_38725);
nor U41842 (N_41842,N_39501,N_38653);
nand U41843 (N_41843,N_38260,N_38299);
xnor U41844 (N_41844,N_38925,N_39621);
and U41845 (N_41845,N_38940,N_39623);
xnor U41846 (N_41846,N_39423,N_39016);
or U41847 (N_41847,N_39407,N_38118);
nor U41848 (N_41848,N_39340,N_39765);
nand U41849 (N_41849,N_38211,N_39245);
nand U41850 (N_41850,N_38051,N_38265);
or U41851 (N_41851,N_38724,N_38155);
nor U41852 (N_41852,N_39935,N_38299);
and U41853 (N_41853,N_38876,N_38462);
xor U41854 (N_41854,N_38648,N_39838);
nor U41855 (N_41855,N_39939,N_39245);
nand U41856 (N_41856,N_38429,N_38994);
nand U41857 (N_41857,N_38947,N_38949);
and U41858 (N_41858,N_38197,N_38386);
nor U41859 (N_41859,N_38901,N_39140);
nand U41860 (N_41860,N_38086,N_39702);
and U41861 (N_41861,N_39532,N_38360);
or U41862 (N_41862,N_38580,N_38881);
and U41863 (N_41863,N_39847,N_39639);
nand U41864 (N_41864,N_39311,N_39608);
nand U41865 (N_41865,N_39713,N_38240);
nor U41866 (N_41866,N_39320,N_38880);
xor U41867 (N_41867,N_39899,N_39946);
or U41868 (N_41868,N_38018,N_39706);
nand U41869 (N_41869,N_39011,N_38827);
xor U41870 (N_41870,N_38453,N_38449);
nand U41871 (N_41871,N_39697,N_38611);
nor U41872 (N_41872,N_38582,N_39130);
and U41873 (N_41873,N_38019,N_38378);
nand U41874 (N_41874,N_39087,N_39042);
and U41875 (N_41875,N_38570,N_39745);
xor U41876 (N_41876,N_39425,N_38193);
and U41877 (N_41877,N_38946,N_39818);
or U41878 (N_41878,N_38859,N_38616);
nand U41879 (N_41879,N_38029,N_38696);
and U41880 (N_41880,N_39337,N_39253);
or U41881 (N_41881,N_39883,N_38807);
or U41882 (N_41882,N_38193,N_39985);
nor U41883 (N_41883,N_39745,N_38199);
and U41884 (N_41884,N_38470,N_38118);
or U41885 (N_41885,N_38146,N_38325);
nand U41886 (N_41886,N_39989,N_38337);
nor U41887 (N_41887,N_39991,N_38377);
nor U41888 (N_41888,N_38537,N_39496);
nand U41889 (N_41889,N_38531,N_39251);
nand U41890 (N_41890,N_38561,N_39291);
xor U41891 (N_41891,N_38361,N_38224);
nand U41892 (N_41892,N_38717,N_39422);
nand U41893 (N_41893,N_38957,N_39967);
nand U41894 (N_41894,N_39234,N_38115);
xnor U41895 (N_41895,N_39522,N_39328);
nor U41896 (N_41896,N_38794,N_38622);
nor U41897 (N_41897,N_39524,N_39045);
or U41898 (N_41898,N_39218,N_39935);
xnor U41899 (N_41899,N_38799,N_38827);
nand U41900 (N_41900,N_38775,N_39439);
or U41901 (N_41901,N_38683,N_38721);
xnor U41902 (N_41902,N_38087,N_38327);
and U41903 (N_41903,N_39941,N_39676);
or U41904 (N_41904,N_39766,N_38905);
nand U41905 (N_41905,N_39997,N_39498);
xor U41906 (N_41906,N_38174,N_39077);
nor U41907 (N_41907,N_38669,N_39729);
nand U41908 (N_41908,N_39725,N_39236);
nand U41909 (N_41909,N_39859,N_39364);
nand U41910 (N_41910,N_38449,N_38811);
xor U41911 (N_41911,N_39085,N_39638);
and U41912 (N_41912,N_38426,N_39105);
xor U41913 (N_41913,N_38778,N_38479);
nor U41914 (N_41914,N_39145,N_38348);
and U41915 (N_41915,N_39707,N_38405);
nor U41916 (N_41916,N_38023,N_39926);
and U41917 (N_41917,N_39106,N_38438);
nor U41918 (N_41918,N_38605,N_39861);
and U41919 (N_41919,N_39835,N_39032);
nor U41920 (N_41920,N_38498,N_39211);
xnor U41921 (N_41921,N_39933,N_39331);
nor U41922 (N_41922,N_38379,N_39393);
nand U41923 (N_41923,N_38149,N_39153);
or U41924 (N_41924,N_39426,N_39887);
nand U41925 (N_41925,N_38800,N_39491);
nand U41926 (N_41926,N_38984,N_39903);
nand U41927 (N_41927,N_39118,N_38901);
xnor U41928 (N_41928,N_38822,N_39557);
nand U41929 (N_41929,N_38435,N_38811);
xnor U41930 (N_41930,N_38784,N_39907);
and U41931 (N_41931,N_39536,N_39359);
and U41932 (N_41932,N_38640,N_38713);
and U41933 (N_41933,N_38204,N_39783);
nand U41934 (N_41934,N_39960,N_39168);
xnor U41935 (N_41935,N_38008,N_38983);
and U41936 (N_41936,N_39043,N_38608);
xnor U41937 (N_41937,N_38479,N_39159);
nand U41938 (N_41938,N_38670,N_39389);
or U41939 (N_41939,N_38440,N_38029);
and U41940 (N_41940,N_39354,N_38420);
and U41941 (N_41941,N_38946,N_39064);
and U41942 (N_41942,N_38695,N_39400);
and U41943 (N_41943,N_39202,N_38128);
or U41944 (N_41944,N_38352,N_39980);
xnor U41945 (N_41945,N_38775,N_38874);
nor U41946 (N_41946,N_39361,N_39920);
nor U41947 (N_41947,N_38842,N_39602);
xnor U41948 (N_41948,N_39608,N_38267);
or U41949 (N_41949,N_39110,N_39940);
or U41950 (N_41950,N_38086,N_39793);
xnor U41951 (N_41951,N_38394,N_39042);
or U41952 (N_41952,N_38064,N_39988);
nor U41953 (N_41953,N_39271,N_39572);
or U41954 (N_41954,N_39258,N_38011);
and U41955 (N_41955,N_39740,N_38366);
nand U41956 (N_41956,N_38633,N_38681);
xnor U41957 (N_41957,N_39895,N_38589);
or U41958 (N_41958,N_39782,N_39138);
and U41959 (N_41959,N_39643,N_39791);
and U41960 (N_41960,N_39299,N_39932);
and U41961 (N_41961,N_38779,N_38848);
or U41962 (N_41962,N_38334,N_38019);
and U41963 (N_41963,N_39917,N_39012);
nand U41964 (N_41964,N_38753,N_38174);
and U41965 (N_41965,N_39895,N_38286);
and U41966 (N_41966,N_39829,N_39391);
xor U41967 (N_41967,N_39847,N_38183);
and U41968 (N_41968,N_38236,N_38423);
and U41969 (N_41969,N_39605,N_39553);
nand U41970 (N_41970,N_38498,N_38319);
nand U41971 (N_41971,N_38873,N_38720);
and U41972 (N_41972,N_39147,N_39787);
and U41973 (N_41973,N_38909,N_39499);
or U41974 (N_41974,N_39446,N_39250);
xor U41975 (N_41975,N_39947,N_38462);
xnor U41976 (N_41976,N_38757,N_38279);
and U41977 (N_41977,N_38709,N_39270);
or U41978 (N_41978,N_39922,N_38269);
xnor U41979 (N_41979,N_38947,N_39644);
and U41980 (N_41980,N_39169,N_39137);
and U41981 (N_41981,N_38605,N_38451);
and U41982 (N_41982,N_38228,N_38262);
xnor U41983 (N_41983,N_38152,N_39108);
nor U41984 (N_41984,N_39093,N_39693);
nor U41985 (N_41985,N_39717,N_38800);
nor U41986 (N_41986,N_38265,N_39217);
nor U41987 (N_41987,N_38058,N_39913);
and U41988 (N_41988,N_38423,N_38555);
and U41989 (N_41989,N_38198,N_38245);
and U41990 (N_41990,N_39834,N_38964);
nand U41991 (N_41991,N_39626,N_38810);
xnor U41992 (N_41992,N_39412,N_38096);
nor U41993 (N_41993,N_38010,N_38019);
or U41994 (N_41994,N_39906,N_38764);
and U41995 (N_41995,N_39120,N_39567);
nand U41996 (N_41996,N_38320,N_39105);
or U41997 (N_41997,N_38309,N_38761);
and U41998 (N_41998,N_38210,N_39956);
xor U41999 (N_41999,N_38802,N_39199);
nor U42000 (N_42000,N_41987,N_40793);
nor U42001 (N_42001,N_40179,N_41455);
and U42002 (N_42002,N_41434,N_40153);
or U42003 (N_42003,N_40876,N_40394);
and U42004 (N_42004,N_41275,N_41057);
nand U42005 (N_42005,N_40148,N_40655);
nand U42006 (N_42006,N_41509,N_40170);
nor U42007 (N_42007,N_40889,N_40919);
and U42008 (N_42008,N_41986,N_40715);
and U42009 (N_42009,N_41380,N_40670);
nor U42010 (N_42010,N_40171,N_40528);
xor U42011 (N_42011,N_41179,N_40074);
and U42012 (N_42012,N_41655,N_41675);
or U42013 (N_42013,N_40961,N_41387);
nand U42014 (N_42014,N_40452,N_41828);
and U42015 (N_42015,N_41044,N_40802);
nor U42016 (N_42016,N_40969,N_41627);
or U42017 (N_42017,N_41467,N_41264);
or U42018 (N_42018,N_41652,N_40262);
or U42019 (N_42019,N_41431,N_40861);
nor U42020 (N_42020,N_40230,N_41874);
nor U42021 (N_42021,N_41092,N_41790);
nand U42022 (N_42022,N_40258,N_40450);
xnor U42023 (N_42023,N_41802,N_40075);
xor U42024 (N_42024,N_41424,N_40747);
nand U42025 (N_42025,N_41925,N_41500);
and U42026 (N_42026,N_40281,N_40009);
and U42027 (N_42027,N_40509,N_41938);
xnor U42028 (N_42028,N_41018,N_40098);
and U42029 (N_42029,N_40240,N_41633);
or U42030 (N_42030,N_41451,N_41969);
or U42031 (N_42031,N_41714,N_40077);
nor U42032 (N_42032,N_40701,N_41889);
xor U42033 (N_42033,N_40959,N_41862);
xor U42034 (N_42034,N_40843,N_41609);
or U42035 (N_42035,N_41965,N_40614);
xnor U42036 (N_42036,N_40297,N_40242);
or U42037 (N_42037,N_40921,N_41197);
or U42038 (N_42038,N_41845,N_40834);
xor U42039 (N_42039,N_40584,N_40072);
or U42040 (N_42040,N_41447,N_40836);
xor U42041 (N_42041,N_40298,N_41180);
and U42042 (N_42042,N_40723,N_40273);
or U42043 (N_42043,N_40488,N_41383);
nand U42044 (N_42044,N_40480,N_41558);
nand U42045 (N_42045,N_41647,N_40182);
or U42046 (N_42046,N_41854,N_40388);
and U42047 (N_42047,N_41242,N_41477);
nand U42048 (N_42048,N_41167,N_40566);
or U42049 (N_42049,N_41523,N_41660);
nand U42050 (N_42050,N_41379,N_41397);
nor U42051 (N_42051,N_41728,N_41530);
and U42052 (N_42052,N_41235,N_41677);
and U42053 (N_42053,N_40574,N_41581);
nand U42054 (N_42054,N_40223,N_41086);
xnor U42055 (N_42055,N_41634,N_40222);
nor U42056 (N_42056,N_41462,N_41396);
nor U42057 (N_42057,N_41875,N_41545);
xor U42058 (N_42058,N_41706,N_41183);
or U42059 (N_42059,N_41270,N_41782);
or U42060 (N_42060,N_40947,N_40735);
xnor U42061 (N_42061,N_41446,N_40904);
xnor U42062 (N_42062,N_41592,N_41411);
and U42063 (N_42063,N_41959,N_41740);
and U42064 (N_42064,N_40219,N_41074);
and U42065 (N_42065,N_40526,N_41843);
nand U42066 (N_42066,N_41886,N_41911);
or U42067 (N_42067,N_41869,N_41865);
and U42068 (N_42068,N_41697,N_40397);
nand U42069 (N_42069,N_41166,N_41830);
or U42070 (N_42070,N_40940,N_40638);
or U42071 (N_42071,N_41529,N_41405);
and U42072 (N_42072,N_40031,N_40410);
or U42073 (N_42073,N_41499,N_40785);
nand U42074 (N_42074,N_41328,N_41468);
nand U42075 (N_42075,N_40546,N_40726);
or U42076 (N_42076,N_40825,N_41810);
xnor U42077 (N_42077,N_41531,N_41619);
nor U42078 (N_42078,N_40381,N_40286);
or U42079 (N_42079,N_41739,N_40781);
nor U42080 (N_42080,N_40897,N_40491);
or U42081 (N_42081,N_41217,N_41471);
nand U42082 (N_42082,N_41248,N_40453);
nand U42083 (N_42083,N_41518,N_41227);
nor U42084 (N_42084,N_40444,N_40702);
nand U42085 (N_42085,N_40913,N_41491);
and U42086 (N_42086,N_40169,N_41335);
and U42087 (N_42087,N_41290,N_40740);
or U42088 (N_42088,N_40982,N_41804);
nor U42089 (N_42089,N_41011,N_41209);
xor U42090 (N_42090,N_40656,N_41564);
and U42091 (N_42091,N_41409,N_41600);
nand U42092 (N_42092,N_41768,N_40300);
nor U42093 (N_42093,N_41878,N_40192);
nor U42094 (N_42094,N_41587,N_41686);
nor U42095 (N_42095,N_40172,N_41648);
nand U42096 (N_42096,N_41436,N_41576);
nor U42097 (N_42097,N_41897,N_40421);
nand U42098 (N_42098,N_41694,N_40336);
nand U42099 (N_42099,N_41220,N_41761);
and U42100 (N_42100,N_40120,N_40900);
nor U42101 (N_42101,N_40161,N_40254);
and U42102 (N_42102,N_41617,N_41165);
xor U42103 (N_42103,N_41414,N_41422);
and U42104 (N_42104,N_40607,N_41813);
nor U42105 (N_42105,N_40977,N_41992);
or U42106 (N_42106,N_41962,N_41563);
nor U42107 (N_42107,N_40379,N_41051);
xnor U42108 (N_42108,N_40313,N_40440);
nor U42109 (N_42109,N_41452,N_40877);
xor U42110 (N_42110,N_41734,N_41249);
and U42111 (N_42111,N_40885,N_40253);
nand U42112 (N_42112,N_40360,N_40511);
and U42113 (N_42113,N_40034,N_40618);
and U42114 (N_42114,N_40902,N_41006);
and U42115 (N_42115,N_40090,N_41549);
nand U42116 (N_42116,N_41901,N_41138);
and U42117 (N_42117,N_40689,N_41053);
and U42118 (N_42118,N_41341,N_40048);
and U42119 (N_42119,N_40291,N_40774);
xnor U42120 (N_42120,N_40532,N_41352);
nand U42121 (N_42121,N_41187,N_40003);
or U42122 (N_42122,N_41147,N_40576);
xnor U42123 (N_42123,N_40682,N_40502);
and U42124 (N_42124,N_41474,N_40026);
xnor U42125 (N_42125,N_41780,N_41663);
or U42126 (N_42126,N_41015,N_40251);
or U42127 (N_42127,N_41759,N_40610);
nor U42128 (N_42128,N_41542,N_41635);
or U42129 (N_42129,N_41861,N_41124);
xnor U42130 (N_42130,N_41887,N_40632);
xor U42131 (N_42131,N_41963,N_41200);
nand U42132 (N_42132,N_41292,N_40542);
xnor U42133 (N_42133,N_41514,N_41787);
xor U42134 (N_42134,N_40901,N_41099);
xnor U42135 (N_42135,N_41507,N_41184);
nor U42136 (N_42136,N_40772,N_41713);
or U42137 (N_42137,N_40773,N_40830);
and U42138 (N_42138,N_41244,N_40318);
nand U42139 (N_42139,N_40974,N_41920);
nor U42140 (N_42140,N_40661,N_40863);
and U42141 (N_42141,N_41737,N_40184);
xor U42142 (N_42142,N_40046,N_41076);
nor U42143 (N_42143,N_41082,N_40493);
nor U42144 (N_42144,N_40150,N_40699);
nor U42145 (N_42145,N_41113,N_40916);
nor U42146 (N_42146,N_40272,N_41503);
nor U42147 (N_42147,N_41762,N_41090);
xor U42148 (N_42148,N_41385,N_41261);
nand U42149 (N_42149,N_40296,N_40369);
nand U42150 (N_42150,N_40418,N_41597);
xor U42151 (N_42151,N_40282,N_41373);
nor U42152 (N_42152,N_40758,N_40938);
and U42153 (N_42153,N_40976,N_41116);
nand U42154 (N_42154,N_40335,N_41610);
nor U42155 (N_42155,N_40896,N_41173);
and U42156 (N_42156,N_40260,N_41551);
xnor U42157 (N_42157,N_41644,N_41691);
xor U42158 (N_42158,N_41747,N_41561);
or U42159 (N_42159,N_40965,N_41594);
and U42160 (N_42160,N_41584,N_40978);
xnor U42161 (N_42161,N_40108,N_41339);
and U42162 (N_42162,N_41094,N_41289);
and U42163 (N_42163,N_41151,N_40842);
and U42164 (N_42164,N_41818,N_41135);
xor U42165 (N_42165,N_41316,N_40685);
or U42166 (N_42166,N_41286,N_41501);
and U42167 (N_42167,N_41596,N_41950);
nor U42168 (N_42168,N_40988,N_40555);
or U42169 (N_42169,N_41738,N_41505);
nand U42170 (N_42170,N_40665,N_40713);
xor U42171 (N_42171,N_40430,N_41528);
or U42172 (N_42172,N_41727,N_40693);
or U42173 (N_42173,N_41871,N_40152);
and U42174 (N_42174,N_40243,N_40137);
nand U42175 (N_42175,N_41265,N_40441);
and U42176 (N_42176,N_40552,N_40166);
or U42177 (N_42177,N_41976,N_41517);
nor U42178 (N_42178,N_40415,N_40798);
or U42179 (N_42179,N_40795,N_40276);
nand U42180 (N_42180,N_40845,N_40070);
nor U42181 (N_42181,N_40017,N_41899);
nor U42182 (N_42182,N_41671,N_41924);
nor U42183 (N_42183,N_41918,N_40789);
nor U42184 (N_42184,N_41495,N_40920);
and U42185 (N_42185,N_41836,N_41771);
nor U42186 (N_42186,N_41742,N_40043);
xnor U42187 (N_42187,N_40141,N_41510);
or U42188 (N_42188,N_41071,N_40371);
nor U42189 (N_42189,N_41073,N_41022);
and U42190 (N_42190,N_41281,N_41196);
nor U42191 (N_42191,N_41990,N_40256);
nor U42192 (N_42192,N_41702,N_41985);
or U42193 (N_42193,N_40392,N_41372);
or U42194 (N_42194,N_40571,N_40745);
and U42195 (N_42195,N_40719,N_41351);
or U42196 (N_42196,N_41294,N_40563);
nor U42197 (N_42197,N_41114,N_41668);
or U42198 (N_42198,N_41287,N_41858);
or U42199 (N_42199,N_41107,N_41700);
and U42200 (N_42200,N_41161,N_40886);
nand U42201 (N_42201,N_40824,N_41588);
nor U42202 (N_42202,N_40892,N_41623);
nor U42203 (N_42203,N_40157,N_40229);
nand U42204 (N_42204,N_41715,N_40432);
and U42205 (N_42205,N_40577,N_40218);
or U42206 (N_42206,N_41021,N_40206);
and U42207 (N_42207,N_41932,N_41350);
or U42208 (N_42208,N_41391,N_40249);
or U42209 (N_42209,N_40014,N_41176);
or U42210 (N_42210,N_40210,N_41636);
or U42211 (N_42211,N_41615,N_41954);
xor U42212 (N_42212,N_40626,N_40342);
xnor U42213 (N_42213,N_40694,N_41357);
or U42214 (N_42214,N_41376,N_40633);
nor U42215 (N_42215,N_41801,N_40942);
or U42216 (N_42216,N_40927,N_41544);
xor U42217 (N_42217,N_41958,N_41100);
nor U42218 (N_42218,N_40568,N_41488);
or U42219 (N_42219,N_40439,N_40115);
nand U42220 (N_42220,N_41896,N_41829);
xor U42221 (N_42221,N_40466,N_41565);
xnor U42222 (N_42222,N_41237,N_41809);
xor U42223 (N_42223,N_40391,N_41935);
and U42224 (N_42224,N_40826,N_41148);
nor U42225 (N_42225,N_41185,N_41522);
xnor U42226 (N_42226,N_40064,N_40967);
and U42227 (N_42227,N_41582,N_40448);
nand U42228 (N_42228,N_40998,N_41075);
nand U42229 (N_42229,N_41273,N_41979);
nor U42230 (N_42230,N_41560,N_40245);
nand U42231 (N_42231,N_40145,N_40905);
or U42232 (N_42232,N_41322,N_41382);
nor U42233 (N_42233,N_41957,N_41624);
nor U42234 (N_42234,N_40645,N_40779);
or U42235 (N_42235,N_40419,N_41749);
nor U42236 (N_42236,N_40517,N_41068);
or U42237 (N_42237,N_41877,N_41163);
or U42238 (N_42238,N_41916,N_41601);
or U42239 (N_42239,N_41122,N_41253);
nor U42240 (N_42240,N_41628,N_40068);
nand U42241 (N_42241,N_40302,N_40540);
or U42242 (N_42242,N_40549,N_41310);
or U42243 (N_42243,N_41750,N_41562);
nand U42244 (N_42244,N_41527,N_41554);
and U42245 (N_42245,N_41543,N_40541);
or U42246 (N_42246,N_40736,N_40197);
and U42247 (N_42247,N_40878,N_40939);
nand U42248 (N_42248,N_40992,N_40387);
nand U42249 (N_42249,N_41442,N_40044);
and U42250 (N_42250,N_41162,N_41219);
and U42251 (N_42251,N_40525,N_40033);
or U42252 (N_42252,N_40029,N_40690);
or U42253 (N_42253,N_40429,N_40246);
or U42254 (N_42254,N_41947,N_40784);
and U42255 (N_42255,N_40981,N_41506);
or U42256 (N_42256,N_41586,N_40013);
nand U42257 (N_42257,N_41437,N_41520);
nor U42258 (N_42258,N_40483,N_40874);
xnor U42259 (N_42259,N_41908,N_40748);
nor U42260 (N_42260,N_40007,N_40567);
nand U42261 (N_42261,N_40482,N_40579);
nor U42262 (N_42262,N_40237,N_41394);
nor U42263 (N_42263,N_40551,N_41998);
xor U42264 (N_42264,N_41643,N_41078);
or U42265 (N_42265,N_40314,N_41997);
and U42266 (N_42266,N_40193,N_41995);
xor U42267 (N_42267,N_41944,N_41898);
xnor U42268 (N_42268,N_40550,N_41744);
xnor U42269 (N_42269,N_40850,N_40175);
and U42270 (N_42270,N_40716,N_41428);
and U42271 (N_42271,N_41566,N_40573);
and U42272 (N_42272,N_41064,N_41573);
or U42273 (N_42273,N_41095,N_40635);
xor U42274 (N_42274,N_41892,N_40316);
nand U42275 (N_42275,N_40703,N_40040);
xnor U42276 (N_42276,N_41680,N_40548);
and U42277 (N_42277,N_40340,N_41052);
or U42278 (N_42278,N_41880,N_41188);
or U42279 (N_42279,N_40099,N_40136);
nand U42280 (N_42280,N_40964,N_40127);
xor U42281 (N_42281,N_40416,N_40220);
and U42282 (N_42282,N_41296,N_40803);
and U42283 (N_42283,N_41313,N_41288);
xor U42284 (N_42284,N_41241,N_41484);
nor U42285 (N_42285,N_40820,N_40377);
and U42286 (N_42286,N_40692,N_40671);
or U42287 (N_42287,N_41685,N_40285);
and U42288 (N_42288,N_41541,N_40505);
xnor U42289 (N_42289,N_40492,N_41764);
nor U42290 (N_42290,N_40792,N_41651);
or U42291 (N_42291,N_41333,N_41433);
nor U42292 (N_42292,N_40188,N_40923);
xor U42293 (N_42293,N_41479,N_40816);
or U42294 (N_42294,N_40815,N_40451);
or U42295 (N_42295,N_41795,N_41699);
xor U42296 (N_42296,N_40644,N_41045);
and U42297 (N_42297,N_40497,N_40827);
xnor U42298 (N_42298,N_40212,N_40250);
xnor U42299 (N_42299,N_41608,N_41207);
nand U42300 (N_42300,N_40104,N_40899);
xor U42301 (N_42301,N_41841,N_40761);
nand U42302 (N_42302,N_40751,N_41621);
nor U42303 (N_42303,N_40983,N_41360);
nand U42304 (N_42304,N_41630,N_41260);
nor U42305 (N_42305,N_41577,N_40585);
xor U42306 (N_42306,N_41005,N_41323);
and U42307 (N_42307,N_40378,N_40456);
or U42308 (N_42308,N_41967,N_40651);
xnor U42309 (N_42309,N_40531,N_41141);
or U42310 (N_42310,N_40217,N_41758);
nor U42311 (N_42311,N_41791,N_40760);
xnor U42312 (N_42312,N_41010,N_40831);
nand U42313 (N_42313,N_40997,N_40195);
nand U42314 (N_42314,N_41991,N_41524);
nand U42315 (N_42315,N_40722,N_40156);
nand U42316 (N_42316,N_41711,N_40201);
and U42317 (N_42317,N_41109,N_40753);
nand U42318 (N_42318,N_41720,N_41888);
nand U42319 (N_42319,N_41312,N_41614);
and U42320 (N_42320,N_40770,N_41401);
nor U42321 (N_42321,N_40461,N_41656);
and U42322 (N_42322,N_40045,N_40849);
xnor U42323 (N_42323,N_41695,N_41306);
and U42324 (N_42324,N_40624,N_41756);
and U42325 (N_42325,N_40399,N_40473);
and U42326 (N_42326,N_40319,N_40829);
xnor U42327 (N_42327,N_41681,N_40084);
and U42328 (N_42328,N_41283,N_41295);
xor U42329 (N_42329,N_40343,N_41133);
nand U42330 (N_42330,N_40085,N_41805);
xnor U42331 (N_42331,N_40489,N_41640);
and U42332 (N_42332,N_40706,N_41012);
or U42333 (N_42333,N_41489,N_40729);
nand U42334 (N_42334,N_40686,N_41672);
nor U42335 (N_42335,N_40389,N_41732);
or U42336 (N_42336,N_41980,N_40600);
and U42337 (N_42337,N_40928,N_40603);
nand U42338 (N_42338,N_40123,N_41872);
xnor U42339 (N_42339,N_40320,N_41314);
or U42340 (N_42340,N_41039,N_40231);
xnor U42341 (N_42341,N_40535,N_40167);
xnor U42342 (N_42342,N_40518,N_41381);
nand U42343 (N_42343,N_40543,N_40420);
nand U42344 (N_42344,N_40255,N_40067);
nor U42345 (N_42345,N_41578,N_41811);
xor U42346 (N_42346,N_41123,N_41859);
xnor U42347 (N_42347,N_40675,N_40930);
nor U42348 (N_42348,N_40209,N_41481);
and U42349 (N_42349,N_40022,N_40971);
and U42350 (N_42350,N_40353,N_41449);
xnor U42351 (N_42351,N_40890,N_41426);
nand U42352 (N_42352,N_41278,N_40883);
xnor U42353 (N_42353,N_40700,N_41160);
nor U42354 (N_42354,N_41302,N_41081);
nor U42355 (N_42355,N_41902,N_40943);
xnor U42356 (N_42356,N_40951,N_41384);
or U42357 (N_42357,N_41538,N_41735);
and U42358 (N_42358,N_41326,N_40813);
or U42359 (N_42359,N_41091,N_40768);
nand U42360 (N_42360,N_41718,N_41701);
nor U42361 (N_42361,N_41108,N_40687);
and U42362 (N_42362,N_41632,N_41069);
xor U42363 (N_42363,N_40879,N_41687);
nand U42364 (N_42364,N_40130,N_41689);
or U42365 (N_42365,N_40739,N_41355);
or U42366 (N_42366,N_41398,N_41927);
and U42367 (N_42367,N_40559,N_40608);
xnor U42368 (N_42368,N_41425,N_41407);
xor U42369 (N_42369,N_40800,N_40054);
and U42370 (N_42370,N_41978,N_41906);
nor U42371 (N_42371,N_41246,N_41026);
nor U42372 (N_42372,N_41438,N_41450);
and U42373 (N_42373,N_41848,N_41238);
or U42374 (N_42374,N_40484,N_40235);
or U42375 (N_42375,N_41585,N_40357);
and U42376 (N_42376,N_40105,N_40398);
xnor U42377 (N_42377,N_41463,N_40125);
or U42378 (N_42378,N_41937,N_41548);
nand U42379 (N_42379,N_41493,N_41393);
xnor U42380 (N_42380,N_40786,N_41882);
or U42381 (N_42381,N_40208,N_40909);
xnor U42382 (N_42382,N_40593,N_41798);
or U42383 (N_42383,N_40037,N_41868);
nor U42384 (N_42384,N_40578,N_40906);
nor U42385 (N_42385,N_41793,N_40322);
nor U42386 (N_42386,N_41303,N_41480);
and U42387 (N_42387,N_41338,N_41783);
xor U42388 (N_42388,N_40944,N_40323);
nor U42389 (N_42389,N_41956,N_41612);
and U42390 (N_42390,N_40674,N_40288);
or U42391 (N_42391,N_41773,N_40957);
nand U42392 (N_42392,N_40583,N_41905);
and U42393 (N_42393,N_40490,N_41126);
nor U42394 (N_42394,N_41894,N_41827);
xnor U42395 (N_42395,N_40647,N_41110);
xor U42396 (N_42396,N_40814,N_41002);
xnor U42397 (N_42397,N_41860,N_40936);
and U42398 (N_42398,N_40190,N_41840);
or U42399 (N_42399,N_41191,N_41629);
xnor U42400 (N_42400,N_41301,N_41465);
nand U42401 (N_42401,N_41717,N_41456);
and U42402 (N_42402,N_40838,N_41061);
xnor U42403 (N_42403,N_40080,N_40459);
xnor U42404 (N_42404,N_41308,N_40177);
nor U42405 (N_42405,N_41800,N_40612);
and U42406 (N_42406,N_41754,N_40326);
nor U42407 (N_42407,N_41525,N_40362);
nand U42408 (N_42408,N_40376,N_40908);
or U42409 (N_42409,N_41366,N_40116);
xor U42410 (N_42410,N_41280,N_40390);
and U42411 (N_42411,N_41626,N_40854);
and U42412 (N_42412,N_40766,N_40018);
and U42413 (N_42413,N_41821,N_40447);
nor U42414 (N_42414,N_41098,N_41508);
xnor U42415 (N_42415,N_41175,N_40063);
nand U42416 (N_42416,N_41359,N_41224);
or U42417 (N_42417,N_40061,N_40306);
and U42418 (N_42418,N_40228,N_41400);
nand U42419 (N_42419,N_41569,N_41096);
nand U42420 (N_42420,N_41483,N_40259);
or U42421 (N_42421,N_40062,N_40324);
nor U42422 (N_42422,N_40287,N_41067);
xor U42423 (N_42423,N_41353,N_41922);
or U42424 (N_42424,N_41311,N_40910);
xnor U42425 (N_42425,N_41150,N_40859);
nor U42426 (N_42426,N_41218,N_41816);
xnor U42427 (N_42427,N_41103,N_41658);
or U42428 (N_42428,N_40370,N_41469);
or U42429 (N_42429,N_40503,N_41111);
and U42430 (N_42430,N_41690,N_41072);
and U42431 (N_42431,N_41516,N_41129);
or U42432 (N_42432,N_41172,N_40539);
xor U42433 (N_42433,N_40350,N_40096);
or U42434 (N_42434,N_40666,N_41943);
and U42435 (N_42435,N_41374,N_40409);
and U42436 (N_42436,N_40966,N_41034);
and U42437 (N_42437,N_40134,N_40069);
xnor U42438 (N_42438,N_40621,N_41667);
and U42439 (N_42439,N_40189,N_40294);
xor U42440 (N_42440,N_40934,N_40864);
or U42441 (N_42441,N_41033,N_41984);
nor U42442 (N_42442,N_41535,N_41533);
or U42443 (N_42443,N_41050,N_41420);
nor U42444 (N_42444,N_41662,N_41060);
or U42445 (N_42445,N_41657,N_41419);
or U42446 (N_42446,N_41825,N_40737);
nor U42447 (N_42447,N_41960,N_40979);
xnor U42448 (N_42448,N_41190,N_40299);
and U42449 (N_42449,N_40019,N_40968);
or U42450 (N_42450,N_40331,N_40688);
nor U42451 (N_42451,N_40224,N_41631);
nor U42452 (N_42452,N_41709,N_41364);
or U42453 (N_42453,N_41181,N_40305);
and U42454 (N_42454,N_40637,N_40140);
nor U42455 (N_42455,N_40349,N_41362);
nand U42456 (N_42456,N_40263,N_41251);
or U42457 (N_42457,N_40464,N_41772);
and U42458 (N_42458,N_40393,N_41591);
nor U42459 (N_42459,N_41233,N_41460);
and U42460 (N_42460,N_40727,N_41305);
nand U42461 (N_42461,N_41826,N_41404);
nand U42462 (N_42462,N_40196,N_40292);
xnor U42463 (N_42463,N_41752,N_40762);
and U42464 (N_42464,N_40799,N_40643);
nand U42465 (N_42465,N_40780,N_41966);
or U42466 (N_42466,N_41014,N_41247);
and U42467 (N_42467,N_40428,N_40524);
nand U42468 (N_42468,N_40274,N_41440);
nor U42469 (N_42469,N_40512,N_40283);
nand U42470 (N_42470,N_41169,N_40499);
and U42471 (N_42471,N_41349,N_40352);
or U42472 (N_42472,N_40659,N_41620);
nand U42473 (N_42473,N_40384,N_41413);
nand U42474 (N_42474,N_41453,N_40562);
nor U42475 (N_42475,N_40307,N_40131);
nand U42476 (N_42476,N_41120,N_41445);
nor U42477 (N_42477,N_40993,N_40832);
xor U42478 (N_42478,N_40422,N_41174);
xnor U42479 (N_42479,N_40118,N_40405);
nor U42480 (N_42480,N_41839,N_40623);
and U42481 (N_42481,N_41893,N_40893);
or U42482 (N_42482,N_40520,N_40213);
or U42483 (N_42483,N_41746,N_41649);
and U42484 (N_42484,N_40903,N_41595);
and U42485 (N_42485,N_41639,N_41299);
nor U42486 (N_42486,N_41598,N_41796);
xnor U42487 (N_42487,N_40641,N_40955);
xor U42488 (N_42488,N_41575,N_40289);
nor U42489 (N_42489,N_41767,N_40382);
and U42490 (N_42490,N_40308,N_40049);
or U42491 (N_42491,N_41354,N_40066);
nand U42492 (N_42492,N_41139,N_41766);
nand U42493 (N_42493,N_41638,N_40165);
and U42494 (N_42494,N_41583,N_40657);
xnor U42495 (N_42495,N_41037,N_41776);
and U42496 (N_42496,N_41923,N_41537);
and U42497 (N_42497,N_40144,N_40962);
and U42498 (N_42498,N_40588,N_40315);
xnor U42499 (N_42499,N_41134,N_40460);
nand U42500 (N_42500,N_41526,N_40199);
nor U42501 (N_42501,N_40478,N_40865);
nor U42502 (N_42502,N_40759,N_40536);
nand U42503 (N_42503,N_40327,N_40364);
or U42504 (N_42504,N_40203,N_41786);
nor U42505 (N_42505,N_40782,N_41547);
and U42506 (N_42506,N_40207,N_41891);
or U42507 (N_42507,N_40006,N_40275);
or U42508 (N_42508,N_40039,N_41863);
and U42509 (N_42509,N_40672,N_40047);
or U42510 (N_42510,N_41031,N_41476);
xnor U42511 (N_42511,N_40403,N_40216);
nor U42512 (N_42512,N_41723,N_41808);
and U42513 (N_42513,N_41763,N_40496);
nor U42514 (N_42514,N_40128,N_40367);
xor U42515 (N_42515,N_40021,N_41721);
nor U42516 (N_42516,N_40173,N_41850);
nand U42517 (N_42517,N_41613,N_40366);
nand U42518 (N_42518,N_41410,N_41267);
nand U42519 (N_42519,N_40474,N_40114);
xnor U42520 (N_42520,N_41198,N_40119);
xor U42521 (N_42521,N_41605,N_41676);
nor U42522 (N_42522,N_40677,N_40572);
nand U42523 (N_42523,N_41940,N_41047);
or U42524 (N_42524,N_40720,N_40504);
or U42525 (N_42525,N_41781,N_40261);
or U42526 (N_42526,N_41490,N_40586);
and U42527 (N_42527,N_40857,N_40710);
nor U42528 (N_42528,N_41994,N_41929);
nand U42529 (N_42529,N_40581,N_40221);
nor U42530 (N_42530,N_40818,N_40875);
or U42531 (N_42531,N_41567,N_41291);
xor U42532 (N_42532,N_40835,N_41222);
nand U42533 (N_42533,N_41832,N_41939);
xor U42534 (N_42534,N_40400,N_41370);
nand U42535 (N_42535,N_40673,N_41102);
or U42536 (N_42536,N_40527,N_40778);
nor U42537 (N_42537,N_40427,N_41152);
or U42538 (N_42538,N_41448,N_41604);
nand U42539 (N_42539,N_41926,N_40925);
and U42540 (N_42540,N_41189,N_41903);
or U42541 (N_42541,N_41087,N_41089);
xnor U42542 (N_42542,N_40368,N_41703);
nand U42543 (N_42543,N_40035,N_41945);
nor U42544 (N_42544,N_41856,N_41088);
xnor U42545 (N_42545,N_40508,N_41325);
nor U42546 (N_42546,N_41029,N_41368);
or U42547 (N_42547,N_40598,N_40545);
and U42548 (N_42548,N_41221,N_40538);
and U42549 (N_42549,N_41334,N_41665);
and U42550 (N_42550,N_41606,N_40252);
and U42551 (N_42551,N_41127,N_41741);
xor U42552 (N_42552,N_40653,N_40247);
xnor U42553 (N_42553,N_41032,N_40958);
xor U42554 (N_42554,N_41777,N_41981);
nor U42555 (N_42555,N_40414,N_41914);
and U42556 (N_42556,N_41427,N_40946);
xor U42557 (N_42557,N_41023,N_41177);
or U42558 (N_42558,N_41659,N_41343);
xnor U42559 (N_42559,N_40051,N_41847);
or U42560 (N_42560,N_41852,N_40788);
or U42561 (N_42561,N_41482,N_40174);
xor U42562 (N_42562,N_40953,N_40180);
nor U42563 (N_42563,N_40107,N_40479);
and U42564 (N_42564,N_40027,N_40147);
nor U42565 (N_42565,N_41853,N_40941);
xor U42566 (N_42566,N_40164,N_40858);
nand U42567 (N_42567,N_40055,N_41277);
nand U42568 (N_42568,N_41432,N_40821);
and U42569 (N_42569,N_41038,N_40746);
nor U42570 (N_42570,N_40985,N_41955);
nand U42571 (N_42571,N_40372,N_40351);
nor U42572 (N_42572,N_41968,N_40590);
and U42573 (N_42573,N_41155,N_41153);
xor U42574 (N_42574,N_40500,N_41900);
or U42575 (N_42575,N_40363,N_40423);
xnor U42576 (N_42576,N_41835,N_40926);
nand U42577 (N_42577,N_40616,N_40731);
nor U42578 (N_42578,N_40856,N_41678);
nand U42579 (N_42579,N_40560,N_41866);
nand U42580 (N_42580,N_41274,N_40000);
or U42581 (N_42581,N_40091,N_41498);
and U42582 (N_42582,N_40065,N_40094);
nand U42583 (N_42583,N_40956,N_40712);
nor U42584 (N_42584,N_40485,N_40554);
nor U42585 (N_42585,N_40058,N_40667);
or U42586 (N_42586,N_41030,N_41930);
nor U42587 (N_42587,N_40733,N_40817);
xnor U42588 (N_42588,N_41194,N_41329);
xor U42589 (N_42589,N_40662,N_40695);
xor U42590 (N_42590,N_40468,N_41371);
nand U42591 (N_42591,N_40436,N_41646);
nor U42592 (N_42592,N_41730,N_41951);
nor U42593 (N_42593,N_41970,N_40794);
nand U42594 (N_42594,N_40604,N_40787);
nor U42595 (N_42595,N_40698,N_40912);
and U42596 (N_42596,N_40862,N_40634);
and U42597 (N_42597,N_40767,N_41806);
or U42598 (N_42598,N_41430,N_41912);
and U42599 (N_42599,N_40954,N_40852);
xnor U42600 (N_42600,N_41386,N_40135);
xnor U42601 (N_42601,N_40443,N_40487);
xor U42602 (N_42602,N_40728,N_40776);
and U42603 (N_42603,N_40741,N_41679);
and U42604 (N_42604,N_40683,N_41403);
and U42605 (N_42605,N_40442,N_41000);
nand U42606 (N_42606,N_41170,N_40984);
or U42607 (N_42607,N_40109,N_40122);
nand U42608 (N_42608,N_41315,N_40005);
xnor U42609 (N_42609,N_40486,N_40293);
and U42610 (N_42610,N_40149,N_41225);
and U42611 (N_42611,N_41988,N_40556);
or U42612 (N_42612,N_41178,N_41550);
xor U42613 (N_42613,N_40176,N_40155);
or U42614 (N_42614,N_41855,N_40001);
nor U42615 (N_42615,N_41004,N_41654);
or U42616 (N_42616,N_41348,N_40454);
and U42617 (N_42617,N_40396,N_40073);
xnor U42618 (N_42618,N_40211,N_41146);
nand U42619 (N_42619,N_41814,N_41070);
and U42620 (N_42620,N_40679,N_41625);
nor U42621 (N_42621,N_41049,N_40570);
and U42622 (N_42622,N_41820,N_40154);
xor U42623 (N_42623,N_40663,N_41933);
nor U42624 (N_42624,N_41212,N_41269);
nor U42625 (N_42625,N_40402,N_41603);
nand U42626 (N_42626,N_41895,N_40241);
xnor U42627 (N_42627,N_41683,N_40991);
nor U42628 (N_42628,N_41693,N_41485);
xnor U42629 (N_42629,N_41534,N_40952);
or U42630 (N_42630,N_41757,N_40648);
nand U42631 (N_42631,N_40016,N_40848);
and U42632 (N_42632,N_40880,N_40117);
and U42633 (N_42633,N_40752,N_40110);
nor U42634 (N_42634,N_40804,N_40232);
nor U42635 (N_42635,N_41692,N_40872);
nand U42636 (N_42636,N_40204,N_40406);
or U42637 (N_42637,N_40911,N_40718);
and U42638 (N_42638,N_41571,N_40994);
and U42639 (N_42639,N_40714,N_41948);
or U42640 (N_42640,N_41321,N_40625);
nand U42641 (N_42641,N_40380,N_40704);
nor U42642 (N_42642,N_41252,N_40279);
xor U42643 (N_42643,N_40810,N_40086);
xor U42644 (N_42644,N_41815,N_40519);
nand U42645 (N_42645,N_40295,N_40092);
and U42646 (N_42646,N_40317,N_40649);
or U42647 (N_42647,N_40095,N_40544);
and U42648 (N_42648,N_41186,N_40042);
nand U42649 (N_42649,N_41504,N_40076);
and U42650 (N_42650,N_40569,N_40438);
and U42651 (N_42651,N_41536,N_40162);
nand U42652 (N_42652,N_41344,N_40321);
or U42653 (N_42653,N_40434,N_40895);
or U42654 (N_42654,N_41331,N_40613);
and U42655 (N_42655,N_41140,N_41682);
nand U42656 (N_42656,N_41797,N_40960);
and U42657 (N_42657,N_40888,N_41036);
nor U42658 (N_42658,N_41572,N_40158);
xnor U42659 (N_42659,N_41412,N_40929);
xnor U42660 (N_42660,N_41769,N_40972);
xor U42661 (N_42661,N_41399,N_40304);
nand U42662 (N_42662,N_40412,N_41199);
or U42663 (N_42663,N_41936,N_41794);
or U42664 (N_42664,N_40765,N_40589);
xnor U42665 (N_42665,N_40124,N_40278);
and U42666 (N_42666,N_41356,N_40530);
xor U42667 (N_42667,N_41673,N_41705);
nand U42668 (N_42668,N_40594,N_40894);
nand U42669 (N_42669,N_40617,N_40113);
or U42670 (N_42670,N_41416,N_40404);
nor U42671 (N_42671,N_41719,N_41066);
nand U42672 (N_42672,N_41054,N_41833);
nand U42673 (N_42673,N_40853,N_41842);
nor U42674 (N_42674,N_40884,N_40796);
nand U42675 (N_42675,N_40111,N_41736);
or U42676 (N_42676,N_40631,N_40822);
nor U42677 (N_42677,N_41009,N_40931);
nor U42678 (N_42678,N_41046,N_41213);
nand U42679 (N_42679,N_41519,N_40112);
and U42680 (N_42680,N_40494,N_41059);
nor U42681 (N_42681,N_41496,N_41760);
xor U42682 (N_42682,N_41570,N_40980);
xnor U42683 (N_42683,N_41993,N_41048);
or U42684 (N_42684,N_40652,N_41559);
xnor U42685 (N_42685,N_41712,N_41317);
and U42686 (N_42686,N_40756,N_40592);
or U42687 (N_42687,N_40945,N_40696);
and U42688 (N_42688,N_41722,N_40561);
nand U42689 (N_42689,N_41745,N_40024);
or U42690 (N_42690,N_40873,N_41142);
nand U42691 (N_42691,N_40425,N_40408);
xnor U42692 (N_42692,N_41367,N_40311);
nor U42693 (N_42693,N_40355,N_41494);
and U42694 (N_42694,N_40734,N_40057);
nand U42695 (N_42695,N_41444,N_41931);
and U42696 (N_42696,N_41792,N_40749);
nand U42697 (N_42697,N_40385,N_41240);
and U42698 (N_42698,N_40236,N_41377);
nor U42699 (N_42699,N_41696,N_40446);
nand U42700 (N_42700,N_40200,N_41803);
xor U42701 (N_42701,N_41263,N_40458);
or U42702 (N_42702,N_40083,N_40750);
and U42703 (N_42703,N_41521,N_40996);
xnor U42704 (N_42704,N_41515,N_41318);
and U42705 (N_42705,N_40937,N_41473);
and U42706 (N_42706,N_41885,N_40847);
nand U42707 (N_42707,N_40975,N_41158);
xnor U42708 (N_42708,N_41616,N_41063);
nand U42709 (N_42709,N_41864,N_41949);
nor U42710 (N_42710,N_41513,N_41953);
nand U42711 (N_42711,N_40346,N_41203);
or U42712 (N_42712,N_41704,N_41822);
nand U42713 (N_42713,N_40949,N_41637);
nand U42714 (N_42714,N_41645,N_40841);
or U42715 (N_42715,N_40924,N_41041);
xor U42716 (N_42716,N_40264,N_41698);
xnor U42717 (N_42717,N_41502,N_41674);
nand U42718 (N_42718,N_40986,N_41003);
xnor U42719 (N_42719,N_40121,N_41346);
and U42720 (N_42720,N_40839,N_41319);
xor U42721 (N_42721,N_40344,N_41743);
and U42722 (N_42722,N_41607,N_41118);
nor U42723 (N_42723,N_40233,N_40198);
nor U42724 (N_42724,N_40431,N_41055);
xnor U42725 (N_42725,N_40087,N_41214);
or U42726 (N_42726,N_40151,N_40881);
nand U42727 (N_42727,N_40558,N_41125);
xnor U42728 (N_42728,N_40744,N_40602);
nand U42729 (N_42729,N_41724,N_40234);
or U42730 (N_42730,N_41193,N_41983);
or U42731 (N_42731,N_41602,N_40032);
xnor U42732 (N_42732,N_41084,N_41580);
or U42733 (N_42733,N_41879,N_40310);
and U42734 (N_42734,N_40819,N_41459);
nor U42735 (N_42735,N_41666,N_40025);
or U42736 (N_42736,N_40582,N_40226);
or U42737 (N_42737,N_41254,N_40472);
nor U42738 (N_42738,N_41337,N_40348);
xor U42739 (N_42739,N_40676,N_40395);
and U42740 (N_42740,N_41441,N_41206);
or U42741 (N_42741,N_41347,N_40669);
and U42742 (N_42742,N_40775,N_40587);
and U42743 (N_42743,N_40168,N_40284);
nor U42744 (N_42744,N_40146,N_40660);
or U42745 (N_42745,N_41641,N_41117);
xnor U42746 (N_42746,N_41511,N_41035);
nand U42747 (N_42747,N_40138,N_40089);
and U42748 (N_42748,N_40807,N_40060);
xor U42749 (N_42749,N_41824,N_40705);
nand U42750 (N_42750,N_41883,N_41285);
nand U42751 (N_42751,N_40513,N_41257);
or U42752 (N_42752,N_40801,N_41324);
nor U42753 (N_42753,N_41077,N_41823);
nor U42754 (N_42754,N_41909,N_41115);
nand U42755 (N_42755,N_41130,N_40709);
nand U42756 (N_42756,N_40361,N_41171);
and U42757 (N_42757,N_40922,N_40469);
and U42758 (N_42758,N_41358,N_40476);
nor U42759 (N_42759,N_41819,N_41788);
and U42760 (N_42760,N_40691,N_41971);
and U42761 (N_42761,N_41093,N_41085);
xor U42762 (N_42762,N_40907,N_41017);
and U42763 (N_42763,N_41439,N_40914);
and U42764 (N_42764,N_40599,N_40163);
nor U42765 (N_42765,N_41961,N_40056);
or U42766 (N_42766,N_40463,N_41552);
or U42767 (N_42767,N_40837,N_41555);
xor U42768 (N_42768,N_40268,N_40619);
or U42769 (N_42769,N_40071,N_40918);
and U42770 (N_42770,N_41276,N_40950);
nor U42771 (N_42771,N_40008,N_40601);
and U42772 (N_42772,N_40338,N_41300);
or U42773 (N_42773,N_40445,N_40915);
or U42774 (N_42774,N_40932,N_40142);
or U42775 (N_42775,N_41934,N_40465);
and U42776 (N_42776,N_40097,N_40470);
and U42777 (N_42777,N_41849,N_41429);
xnor U42778 (N_42778,N_40989,N_41913);
nor U42779 (N_42779,N_41540,N_40580);
nor U42780 (N_42780,N_40358,N_41710);
or U42781 (N_42781,N_41016,N_40386);
or U42782 (N_42782,N_40160,N_41785);
xnor U42783 (N_42783,N_41611,N_40059);
xor U42784 (N_42784,N_40882,N_41915);
xor U42785 (N_42785,N_40248,N_41464);
nor U42786 (N_42786,N_40280,N_41215);
nand U42787 (N_42787,N_41466,N_41149);
nand U42788 (N_42788,N_40777,N_41262);
or U42789 (N_42789,N_41062,N_41454);
nand U42790 (N_42790,N_41136,N_40717);
and U42791 (N_42791,N_41461,N_40783);
xnor U42792 (N_42792,N_40547,N_41729);
nor U42793 (N_42793,N_40629,N_41844);
xor U42794 (N_42794,N_40811,N_41784);
nor U42795 (N_42795,N_40081,N_41851);
xor U42796 (N_42796,N_40093,N_40805);
and U42797 (N_42797,N_41156,N_40126);
xor U42798 (N_42798,N_41378,N_41395);
and U42799 (N_42799,N_41065,N_40449);
nand U42800 (N_42800,N_41195,N_40433);
or U42801 (N_42801,N_41375,N_41284);
xnor U42802 (N_42802,N_40840,N_41568);
xnor U42803 (N_42803,N_40724,N_41688);
xnor U42804 (N_42804,N_40507,N_41228);
nor U42805 (N_42805,N_41304,N_41201);
nor U42806 (N_42806,N_40537,N_41105);
xor U42807 (N_42807,N_40506,N_40763);
and U42808 (N_42808,N_41204,N_41121);
and U42809 (N_42809,N_40844,N_40867);
and U42810 (N_42810,N_40595,N_41579);
nand U42811 (N_42811,N_40257,N_40426);
xnor U42812 (N_42812,N_41112,N_40757);
nor U42813 (N_42813,N_40654,N_41443);
or U42814 (N_42814,N_40963,N_40374);
nor U42815 (N_42815,N_41164,N_41216);
xor U42816 (N_42816,N_41058,N_41890);
and U42817 (N_42817,N_40738,N_40678);
or U42818 (N_42818,N_41309,N_41101);
and U42819 (N_42819,N_41557,N_41748);
or U42820 (N_42820,N_40846,N_40100);
and U42821 (N_42821,N_41831,N_40373);
xnor U42822 (N_42822,N_41243,N_41020);
and U42823 (N_42823,N_40642,N_40178);
nor U42824 (N_42824,N_41755,N_41079);
and U42825 (N_42825,N_41259,N_40870);
nor U42826 (N_42826,N_41001,N_40102);
or U42827 (N_42827,N_41417,N_40668);
xnor U42828 (N_42828,N_40708,N_41128);
nor U42829 (N_42829,N_40341,N_41807);
and U42830 (N_42830,N_40605,N_41272);
nor U42831 (N_42831,N_41977,N_41589);
and U42832 (N_42832,N_40265,N_40191);
nor U42833 (N_42833,N_41250,N_40650);
nor U42834 (N_42834,N_41208,N_41475);
and U42835 (N_42835,N_40725,N_41458);
or U42836 (N_42836,N_41157,N_40515);
xor U42837 (N_42837,N_40640,N_40860);
or U42838 (N_42838,N_41870,N_40769);
and U42839 (N_42839,N_40597,N_40345);
nor U42840 (N_42840,N_41271,N_40052);
nand U42841 (N_42841,N_41192,N_41881);
nor U42842 (N_42842,N_41942,N_40266);
nor U42843 (N_42843,N_40917,N_40868);
xnor U42844 (N_42844,N_40790,N_41435);
and U42845 (N_42845,N_40101,N_41211);
nor U42846 (N_42846,N_41599,N_40002);
xnor U42847 (N_42847,N_41132,N_40565);
nand U42848 (N_42848,N_41042,N_41622);
xor U42849 (N_42849,N_40437,N_41941);
or U42850 (N_42850,N_41876,N_41472);
nor U42851 (N_42851,N_41389,N_40269);
xor U42852 (N_42852,N_41025,N_40622);
xor U42853 (N_42853,N_40866,N_41964);
xor U42854 (N_42854,N_40277,N_40328);
or U42855 (N_42855,N_41593,N_40970);
xnor U42856 (N_42856,N_41027,N_40401);
nor U42857 (N_42857,N_40630,N_41007);
and U42858 (N_42858,N_40133,N_41731);
and U42859 (N_42859,N_41143,N_40721);
or U42860 (N_42860,N_41131,N_41361);
xor U42861 (N_42861,N_41590,N_40973);
and U42862 (N_42862,N_40365,N_41230);
and U42863 (N_42863,N_40424,N_41669);
or U42864 (N_42864,N_40028,N_40030);
nand U42865 (N_42865,N_40312,N_41083);
nand U42866 (N_42866,N_41708,N_40808);
nand U42867 (N_42867,N_41119,N_40851);
xnor U42868 (N_42868,N_40684,N_41972);
and U42869 (N_42869,N_40186,N_40495);
or U42870 (N_42870,N_40791,N_41873);
nand U42871 (N_42871,N_41268,N_41670);
and U42872 (N_42872,N_41457,N_41733);
or U42873 (N_42873,N_41774,N_41390);
or U42874 (N_42874,N_41716,N_41097);
or U42875 (N_42875,N_40516,N_40609);
or U42876 (N_42876,N_41910,N_41470);
xor U42877 (N_42877,N_41618,N_41497);
nor U42878 (N_42878,N_40887,N_41293);
nor U42879 (N_42879,N_40143,N_41282);
nor U42880 (N_42880,N_41974,N_41231);
or U42881 (N_42881,N_40359,N_41952);
or U42882 (N_42882,N_40011,N_40187);
nor U42883 (N_42883,N_41239,N_41392);
and U42884 (N_42884,N_40332,N_41664);
xor U42885 (N_42885,N_41330,N_41799);
nand U42886 (N_42886,N_41642,N_41553);
nand U42887 (N_42887,N_40806,N_41846);
or U42888 (N_42888,N_40290,N_41837);
nand U42889 (N_42889,N_40898,N_40330);
nor U42890 (N_42890,N_41024,N_41298);
xnor U42891 (N_42891,N_40334,N_41013);
and U42892 (N_42892,N_40948,N_40697);
and U42893 (N_42893,N_41279,N_40214);
or U42894 (N_42894,N_41707,N_41834);
or U42895 (N_42895,N_40999,N_41106);
nand U42896 (N_42896,N_40523,N_41546);
nand U42897 (N_42897,N_40732,N_40833);
and U42898 (N_42898,N_41144,N_41857);
nor U42899 (N_42899,N_40347,N_41753);
xnor U42900 (N_42900,N_40185,N_41778);
and U42901 (N_42901,N_40407,N_41996);
and U42902 (N_42902,N_41332,N_41320);
and U42903 (N_42903,N_41342,N_41040);
xnor U42904 (N_42904,N_40267,N_40611);
and U42905 (N_42905,N_41904,N_40078);
nand U42906 (N_42906,N_40680,N_40225);
nand U42907 (N_42907,N_40711,N_40303);
xor U42908 (N_42908,N_40339,N_41423);
or U42909 (N_42909,N_40646,N_40301);
nor U42910 (N_42910,N_40990,N_41402);
nand U42911 (N_42911,N_40004,N_40181);
or U42912 (N_42912,N_40012,N_41725);
or U42913 (N_42913,N_41487,N_40514);
nor U42914 (N_42914,N_41574,N_41653);
xor U42915 (N_42915,N_40620,N_41336);
nand U42916 (N_42916,N_40812,N_41989);
or U42917 (N_42917,N_40238,N_40455);
or U42918 (N_42918,N_40658,N_40015);
or U42919 (N_42919,N_41999,N_41019);
nor U42920 (N_42920,N_41751,N_40079);
nand U42921 (N_42921,N_40020,N_40325);
and U42922 (N_42922,N_40383,N_40553);
xor U42923 (N_42923,N_40411,N_40891);
nand U42924 (N_42924,N_41418,N_41388);
and U42925 (N_42925,N_40205,N_40664);
and U42926 (N_42926,N_41921,N_40871);
nand U42927 (N_42927,N_41258,N_40628);
and U42928 (N_42928,N_40413,N_40771);
or U42929 (N_42929,N_40533,N_40159);
and U42930 (N_42930,N_41812,N_40202);
nor U42931 (N_42931,N_40627,N_40354);
or U42932 (N_42932,N_41297,N_40462);
or U42933 (N_42933,N_41684,N_40477);
and U42934 (N_42934,N_40036,N_40244);
or U42935 (N_42935,N_40356,N_41168);
xnor U42936 (N_42936,N_40481,N_41838);
nor U42937 (N_42937,N_41210,N_41159);
xnor U42938 (N_42938,N_40239,N_41775);
nor U42939 (N_42939,N_41369,N_40023);
or U42940 (N_42940,N_41770,N_41884);
nor U42941 (N_42941,N_41982,N_40103);
and U42942 (N_42942,N_41973,N_40132);
xnor U42943 (N_42943,N_41415,N_41307);
or U42944 (N_42944,N_41229,N_40755);
nand U42945 (N_42945,N_41406,N_40606);
nand U42946 (N_42946,N_41226,N_40636);
nor U42947 (N_42947,N_40053,N_41327);
and U42948 (N_42948,N_40743,N_41340);
or U42949 (N_42949,N_41255,N_41223);
and U42950 (N_42950,N_41056,N_40417);
nand U42951 (N_42951,N_40050,N_41266);
and U42952 (N_42952,N_40615,N_40797);
nand U42953 (N_42953,N_41556,N_40828);
nand U42954 (N_42954,N_41154,N_41532);
and U42955 (N_42955,N_41789,N_41145);
xnor U42956 (N_42956,N_41928,N_41661);
and U42957 (N_42957,N_40995,N_40935);
and U42958 (N_42958,N_41726,N_40194);
nand U42959 (N_42959,N_41478,N_41817);
and U42960 (N_42960,N_40529,N_41080);
nand U42961 (N_42961,N_40038,N_41234);
xnor U42962 (N_42962,N_41202,N_41182);
xnor U42963 (N_42963,N_40457,N_40227);
or U42964 (N_42964,N_41919,N_40475);
and U42965 (N_42965,N_41345,N_41028);
xor U42966 (N_42966,N_41539,N_40534);
nand U42967 (N_42967,N_40742,N_40730);
and U42968 (N_42968,N_40764,N_40471);
and U42969 (N_42969,N_40987,N_40329);
and U42970 (N_42970,N_41245,N_40855);
nor U42971 (N_42971,N_41492,N_40707);
nor U42972 (N_42972,N_40082,N_40309);
nand U42973 (N_42973,N_40522,N_40435);
or U42974 (N_42974,N_41779,N_41104);
or U42975 (N_42975,N_40139,N_41917);
or U42976 (N_42976,N_40106,N_41765);
xor U42977 (N_42977,N_41650,N_40337);
or U42978 (N_42978,N_41232,N_40467);
or U42979 (N_42979,N_40375,N_41365);
and U42980 (N_42980,N_40681,N_40183);
and U42981 (N_42981,N_40501,N_41486);
xor U42982 (N_42982,N_40521,N_40809);
nand U42983 (N_42983,N_40498,N_41867);
or U42984 (N_42984,N_41946,N_40639);
or U42985 (N_42985,N_40333,N_40010);
nor U42986 (N_42986,N_41907,N_40933);
and U42987 (N_42987,N_41137,N_40754);
and U42988 (N_42988,N_41363,N_41236);
nor U42989 (N_42989,N_40129,N_40088);
nor U42990 (N_42990,N_41408,N_40591);
nand U42991 (N_42991,N_41421,N_41043);
and U42992 (N_42992,N_40270,N_40869);
nor U42993 (N_42993,N_40215,N_41256);
or U42994 (N_42994,N_41205,N_40564);
and U42995 (N_42995,N_40823,N_40596);
nor U42996 (N_42996,N_40510,N_40271);
nand U42997 (N_42997,N_40557,N_41975);
or U42998 (N_42998,N_40041,N_40575);
and U42999 (N_42999,N_41512,N_41008);
or U43000 (N_43000,N_40887,N_40361);
nand U43001 (N_43001,N_40730,N_41839);
and U43002 (N_43002,N_40442,N_41156);
nand U43003 (N_43003,N_40091,N_40547);
xnor U43004 (N_43004,N_41080,N_40258);
and U43005 (N_43005,N_40519,N_40781);
or U43006 (N_43006,N_40154,N_40256);
or U43007 (N_43007,N_40892,N_40012);
xor U43008 (N_43008,N_40120,N_41065);
nand U43009 (N_43009,N_41156,N_40201);
xor U43010 (N_43010,N_40650,N_40758);
xnor U43011 (N_43011,N_41183,N_41943);
nand U43012 (N_43012,N_40241,N_40161);
or U43013 (N_43013,N_41272,N_41314);
nand U43014 (N_43014,N_41814,N_40116);
xnor U43015 (N_43015,N_40536,N_41194);
nor U43016 (N_43016,N_40246,N_40257);
or U43017 (N_43017,N_40790,N_41741);
and U43018 (N_43018,N_41204,N_40268);
nand U43019 (N_43019,N_40638,N_40161);
nand U43020 (N_43020,N_41684,N_41553);
xor U43021 (N_43021,N_40633,N_40928);
or U43022 (N_43022,N_41601,N_40355);
nor U43023 (N_43023,N_41119,N_40390);
nand U43024 (N_43024,N_41643,N_40926);
nand U43025 (N_43025,N_40467,N_40776);
xnor U43026 (N_43026,N_40435,N_41721);
nand U43027 (N_43027,N_40690,N_41947);
or U43028 (N_43028,N_41303,N_40351);
nor U43029 (N_43029,N_40509,N_41788);
xor U43030 (N_43030,N_40582,N_41706);
and U43031 (N_43031,N_41729,N_41035);
and U43032 (N_43032,N_41430,N_41257);
and U43033 (N_43033,N_40283,N_40287);
xor U43034 (N_43034,N_41823,N_41686);
xor U43035 (N_43035,N_40748,N_41387);
xnor U43036 (N_43036,N_41608,N_41400);
or U43037 (N_43037,N_41183,N_41708);
or U43038 (N_43038,N_40236,N_40070);
and U43039 (N_43039,N_41952,N_40478);
xnor U43040 (N_43040,N_40953,N_41020);
xnor U43041 (N_43041,N_41597,N_41481);
nand U43042 (N_43042,N_41417,N_41991);
and U43043 (N_43043,N_41172,N_41402);
and U43044 (N_43044,N_40694,N_41254);
xor U43045 (N_43045,N_40061,N_41300);
nor U43046 (N_43046,N_40612,N_40532);
nand U43047 (N_43047,N_40270,N_40132);
nand U43048 (N_43048,N_40946,N_41809);
or U43049 (N_43049,N_41482,N_40517);
and U43050 (N_43050,N_41576,N_40727);
and U43051 (N_43051,N_41651,N_40062);
xor U43052 (N_43052,N_41656,N_40043);
nor U43053 (N_43053,N_41234,N_41255);
nor U43054 (N_43054,N_41211,N_41815);
xor U43055 (N_43055,N_40618,N_41577);
or U43056 (N_43056,N_40590,N_41972);
and U43057 (N_43057,N_41473,N_41397);
or U43058 (N_43058,N_40622,N_41921);
and U43059 (N_43059,N_40022,N_40512);
nor U43060 (N_43060,N_40348,N_40693);
nor U43061 (N_43061,N_40720,N_40894);
and U43062 (N_43062,N_40728,N_40080);
nand U43063 (N_43063,N_40326,N_40387);
xor U43064 (N_43064,N_40534,N_41744);
or U43065 (N_43065,N_40211,N_41587);
nand U43066 (N_43066,N_41089,N_41993);
nor U43067 (N_43067,N_41989,N_40127);
and U43068 (N_43068,N_40647,N_40778);
nor U43069 (N_43069,N_40538,N_41313);
or U43070 (N_43070,N_40144,N_41160);
nor U43071 (N_43071,N_40507,N_40021);
xnor U43072 (N_43072,N_40152,N_40157);
xor U43073 (N_43073,N_41857,N_41326);
and U43074 (N_43074,N_41587,N_41512);
and U43075 (N_43075,N_40399,N_41373);
nor U43076 (N_43076,N_40652,N_41682);
or U43077 (N_43077,N_41623,N_40788);
or U43078 (N_43078,N_40819,N_40906);
or U43079 (N_43079,N_40583,N_41756);
xnor U43080 (N_43080,N_41067,N_41358);
nor U43081 (N_43081,N_41302,N_41304);
or U43082 (N_43082,N_41634,N_40847);
and U43083 (N_43083,N_41195,N_40799);
nor U43084 (N_43084,N_40493,N_40252);
xnor U43085 (N_43085,N_41505,N_40134);
and U43086 (N_43086,N_40479,N_40456);
nor U43087 (N_43087,N_41725,N_41422);
nand U43088 (N_43088,N_41414,N_40671);
and U43089 (N_43089,N_40093,N_40053);
nand U43090 (N_43090,N_40750,N_40788);
xor U43091 (N_43091,N_41947,N_40624);
or U43092 (N_43092,N_41268,N_40839);
and U43093 (N_43093,N_40559,N_41609);
xor U43094 (N_43094,N_40155,N_41288);
nor U43095 (N_43095,N_40171,N_40096);
or U43096 (N_43096,N_41114,N_40558);
nor U43097 (N_43097,N_40474,N_41295);
nand U43098 (N_43098,N_41438,N_40279);
nand U43099 (N_43099,N_40232,N_40151);
or U43100 (N_43100,N_41610,N_40125);
xor U43101 (N_43101,N_40581,N_41288);
and U43102 (N_43102,N_41093,N_41646);
nor U43103 (N_43103,N_40342,N_41340);
and U43104 (N_43104,N_41581,N_40963);
and U43105 (N_43105,N_40770,N_40847);
nand U43106 (N_43106,N_41343,N_40472);
and U43107 (N_43107,N_40673,N_41690);
or U43108 (N_43108,N_40250,N_41386);
nor U43109 (N_43109,N_40811,N_40377);
xnor U43110 (N_43110,N_41231,N_40147);
nand U43111 (N_43111,N_40624,N_40720);
and U43112 (N_43112,N_40112,N_41377);
nor U43113 (N_43113,N_41992,N_41784);
nor U43114 (N_43114,N_41244,N_40670);
xnor U43115 (N_43115,N_40199,N_41256);
xor U43116 (N_43116,N_41730,N_41882);
nor U43117 (N_43117,N_40258,N_41348);
and U43118 (N_43118,N_41520,N_40752);
or U43119 (N_43119,N_40622,N_41792);
nand U43120 (N_43120,N_41467,N_40375);
nor U43121 (N_43121,N_41869,N_40631);
nand U43122 (N_43122,N_41313,N_40884);
and U43123 (N_43123,N_40902,N_41414);
xor U43124 (N_43124,N_40548,N_40378);
and U43125 (N_43125,N_40839,N_41287);
and U43126 (N_43126,N_41343,N_40913);
and U43127 (N_43127,N_41952,N_41730);
nor U43128 (N_43128,N_41273,N_41517);
nand U43129 (N_43129,N_40444,N_40280);
nor U43130 (N_43130,N_41723,N_40604);
nand U43131 (N_43131,N_41788,N_40196);
nor U43132 (N_43132,N_41023,N_40696);
nand U43133 (N_43133,N_40939,N_41453);
nand U43134 (N_43134,N_41383,N_41503);
nand U43135 (N_43135,N_40148,N_40312);
xnor U43136 (N_43136,N_40348,N_41494);
and U43137 (N_43137,N_41283,N_40206);
xnor U43138 (N_43138,N_41696,N_41708);
or U43139 (N_43139,N_41377,N_41467);
xor U43140 (N_43140,N_41960,N_40803);
or U43141 (N_43141,N_40694,N_41732);
nand U43142 (N_43142,N_41668,N_41655);
nor U43143 (N_43143,N_40039,N_41985);
or U43144 (N_43144,N_41053,N_41773);
nand U43145 (N_43145,N_41272,N_41335);
and U43146 (N_43146,N_40209,N_41927);
xnor U43147 (N_43147,N_41474,N_41523);
nand U43148 (N_43148,N_41677,N_40606);
nor U43149 (N_43149,N_41063,N_41047);
and U43150 (N_43150,N_40911,N_41960);
nand U43151 (N_43151,N_41733,N_40089);
or U43152 (N_43152,N_41473,N_40516);
and U43153 (N_43153,N_40435,N_41924);
and U43154 (N_43154,N_41275,N_41112);
or U43155 (N_43155,N_41783,N_40628);
xnor U43156 (N_43156,N_41142,N_41521);
nand U43157 (N_43157,N_41986,N_41874);
and U43158 (N_43158,N_41834,N_41132);
or U43159 (N_43159,N_40826,N_40058);
nand U43160 (N_43160,N_41956,N_41902);
or U43161 (N_43161,N_41525,N_40207);
nand U43162 (N_43162,N_40651,N_41889);
or U43163 (N_43163,N_41328,N_40994);
nor U43164 (N_43164,N_40965,N_40714);
or U43165 (N_43165,N_40129,N_40474);
nand U43166 (N_43166,N_40622,N_41225);
or U43167 (N_43167,N_40702,N_41304);
nor U43168 (N_43168,N_40439,N_41030);
xnor U43169 (N_43169,N_40176,N_41290);
or U43170 (N_43170,N_41432,N_41245);
nand U43171 (N_43171,N_41496,N_41537);
nor U43172 (N_43172,N_41524,N_40055);
xnor U43173 (N_43173,N_41987,N_40291);
nor U43174 (N_43174,N_41481,N_41537);
and U43175 (N_43175,N_40063,N_41180);
xor U43176 (N_43176,N_41703,N_41479);
xor U43177 (N_43177,N_40889,N_40858);
nor U43178 (N_43178,N_41561,N_40142);
xnor U43179 (N_43179,N_41464,N_40143);
or U43180 (N_43180,N_41066,N_40889);
and U43181 (N_43181,N_41220,N_41123);
xor U43182 (N_43182,N_40430,N_40125);
or U43183 (N_43183,N_41526,N_40193);
or U43184 (N_43184,N_40919,N_40315);
xnor U43185 (N_43185,N_41487,N_41733);
nor U43186 (N_43186,N_41380,N_40006);
or U43187 (N_43187,N_41242,N_41437);
or U43188 (N_43188,N_40849,N_41823);
nor U43189 (N_43189,N_41418,N_41718);
nand U43190 (N_43190,N_40657,N_41979);
or U43191 (N_43191,N_41855,N_41129);
or U43192 (N_43192,N_41270,N_40001);
nand U43193 (N_43193,N_40149,N_40416);
or U43194 (N_43194,N_41724,N_41714);
nor U43195 (N_43195,N_41814,N_40535);
and U43196 (N_43196,N_40917,N_40908);
and U43197 (N_43197,N_40693,N_41117);
or U43198 (N_43198,N_41902,N_40054);
and U43199 (N_43199,N_40111,N_40187);
nor U43200 (N_43200,N_41819,N_41107);
xor U43201 (N_43201,N_40962,N_40692);
and U43202 (N_43202,N_40268,N_41967);
xnor U43203 (N_43203,N_40813,N_41752);
xor U43204 (N_43204,N_40977,N_40338);
xnor U43205 (N_43205,N_40851,N_41222);
xor U43206 (N_43206,N_40372,N_40744);
or U43207 (N_43207,N_40858,N_40264);
or U43208 (N_43208,N_40107,N_40714);
xor U43209 (N_43209,N_41799,N_41107);
and U43210 (N_43210,N_40838,N_40328);
and U43211 (N_43211,N_41858,N_41904);
nor U43212 (N_43212,N_40984,N_40222);
and U43213 (N_43213,N_41791,N_40267);
nor U43214 (N_43214,N_41219,N_41375);
or U43215 (N_43215,N_41294,N_40874);
nand U43216 (N_43216,N_41967,N_41444);
or U43217 (N_43217,N_41228,N_41455);
nor U43218 (N_43218,N_40558,N_40211);
xnor U43219 (N_43219,N_40688,N_40749);
and U43220 (N_43220,N_40833,N_40174);
and U43221 (N_43221,N_41508,N_41944);
or U43222 (N_43222,N_41214,N_40960);
or U43223 (N_43223,N_40507,N_40939);
and U43224 (N_43224,N_40600,N_40532);
nand U43225 (N_43225,N_41603,N_40929);
nor U43226 (N_43226,N_40344,N_41000);
or U43227 (N_43227,N_40611,N_41122);
nor U43228 (N_43228,N_40273,N_40395);
nand U43229 (N_43229,N_40736,N_41553);
nand U43230 (N_43230,N_41816,N_41583);
and U43231 (N_43231,N_40785,N_40440);
or U43232 (N_43232,N_41667,N_40319);
nor U43233 (N_43233,N_40455,N_41245);
nand U43234 (N_43234,N_40484,N_41684);
or U43235 (N_43235,N_40340,N_40056);
nor U43236 (N_43236,N_40805,N_41945);
and U43237 (N_43237,N_40865,N_40227);
nand U43238 (N_43238,N_40999,N_40051);
nor U43239 (N_43239,N_40036,N_41672);
or U43240 (N_43240,N_40745,N_40353);
and U43241 (N_43241,N_40321,N_40436);
nand U43242 (N_43242,N_40113,N_41822);
and U43243 (N_43243,N_41103,N_41390);
and U43244 (N_43244,N_41875,N_41794);
and U43245 (N_43245,N_41181,N_40528);
nor U43246 (N_43246,N_41065,N_41743);
and U43247 (N_43247,N_41324,N_40552);
nand U43248 (N_43248,N_40742,N_40906);
or U43249 (N_43249,N_40929,N_41087);
xor U43250 (N_43250,N_40599,N_40856);
xnor U43251 (N_43251,N_41286,N_41395);
or U43252 (N_43252,N_40020,N_40894);
xor U43253 (N_43253,N_41924,N_41532);
nand U43254 (N_43254,N_41216,N_41158);
and U43255 (N_43255,N_40284,N_40326);
or U43256 (N_43256,N_40143,N_40545);
xnor U43257 (N_43257,N_40913,N_40295);
or U43258 (N_43258,N_41219,N_40873);
xor U43259 (N_43259,N_41453,N_41519);
nand U43260 (N_43260,N_40358,N_40485);
nor U43261 (N_43261,N_40322,N_41610);
xor U43262 (N_43262,N_40439,N_40368);
and U43263 (N_43263,N_40216,N_40219);
nor U43264 (N_43264,N_41381,N_40526);
and U43265 (N_43265,N_40061,N_40484);
or U43266 (N_43266,N_41403,N_40659);
nand U43267 (N_43267,N_40706,N_40548);
or U43268 (N_43268,N_40685,N_41046);
nand U43269 (N_43269,N_40812,N_41099);
and U43270 (N_43270,N_41243,N_40041);
nor U43271 (N_43271,N_40468,N_40528);
and U43272 (N_43272,N_40087,N_40494);
or U43273 (N_43273,N_40293,N_41294);
and U43274 (N_43274,N_40995,N_41510);
nand U43275 (N_43275,N_40167,N_41178);
nand U43276 (N_43276,N_40309,N_40728);
and U43277 (N_43277,N_40263,N_40578);
xnor U43278 (N_43278,N_41629,N_41956);
nand U43279 (N_43279,N_40670,N_41017);
and U43280 (N_43280,N_40619,N_41777);
and U43281 (N_43281,N_41887,N_41074);
nor U43282 (N_43282,N_40080,N_40913);
and U43283 (N_43283,N_41538,N_40282);
nor U43284 (N_43284,N_40295,N_40542);
and U43285 (N_43285,N_40309,N_40026);
and U43286 (N_43286,N_40836,N_40791);
xor U43287 (N_43287,N_41539,N_41638);
nor U43288 (N_43288,N_40721,N_41161);
nor U43289 (N_43289,N_40138,N_40267);
nand U43290 (N_43290,N_40008,N_40037);
or U43291 (N_43291,N_40379,N_40529);
xnor U43292 (N_43292,N_40458,N_40152);
xor U43293 (N_43293,N_40756,N_40984);
nor U43294 (N_43294,N_40837,N_40018);
or U43295 (N_43295,N_41899,N_40898);
xnor U43296 (N_43296,N_41065,N_41900);
and U43297 (N_43297,N_40576,N_40412);
and U43298 (N_43298,N_41136,N_41677);
or U43299 (N_43299,N_40683,N_40057);
nor U43300 (N_43300,N_41827,N_41550);
nand U43301 (N_43301,N_40566,N_40279);
or U43302 (N_43302,N_40023,N_41041);
nor U43303 (N_43303,N_40491,N_41559);
and U43304 (N_43304,N_40091,N_40997);
or U43305 (N_43305,N_40398,N_40948);
nor U43306 (N_43306,N_41482,N_40173);
or U43307 (N_43307,N_40721,N_41767);
nand U43308 (N_43308,N_40386,N_40516);
nand U43309 (N_43309,N_40696,N_41593);
and U43310 (N_43310,N_40338,N_41144);
and U43311 (N_43311,N_40453,N_40152);
nor U43312 (N_43312,N_40699,N_40729);
xor U43313 (N_43313,N_40867,N_40091);
nand U43314 (N_43314,N_41912,N_41449);
nor U43315 (N_43315,N_40659,N_40203);
nand U43316 (N_43316,N_40581,N_40373);
nand U43317 (N_43317,N_40725,N_41153);
and U43318 (N_43318,N_41540,N_40059);
or U43319 (N_43319,N_40543,N_40629);
and U43320 (N_43320,N_40031,N_40226);
and U43321 (N_43321,N_40107,N_40127);
nand U43322 (N_43322,N_41759,N_41858);
xor U43323 (N_43323,N_40342,N_40812);
xnor U43324 (N_43324,N_41402,N_41122);
and U43325 (N_43325,N_40763,N_40168);
and U43326 (N_43326,N_40210,N_40229);
nor U43327 (N_43327,N_41455,N_40564);
xnor U43328 (N_43328,N_41665,N_40933);
or U43329 (N_43329,N_41733,N_41039);
nand U43330 (N_43330,N_41967,N_41422);
or U43331 (N_43331,N_40707,N_40480);
and U43332 (N_43332,N_41376,N_40227);
and U43333 (N_43333,N_41472,N_41357);
nor U43334 (N_43334,N_41429,N_40623);
or U43335 (N_43335,N_40325,N_41085);
xor U43336 (N_43336,N_40965,N_41718);
nand U43337 (N_43337,N_41559,N_41913);
nor U43338 (N_43338,N_40305,N_40175);
or U43339 (N_43339,N_40335,N_40697);
nor U43340 (N_43340,N_40295,N_41970);
and U43341 (N_43341,N_40159,N_41463);
xor U43342 (N_43342,N_41371,N_41490);
nand U43343 (N_43343,N_41421,N_41144);
nand U43344 (N_43344,N_41098,N_41960);
and U43345 (N_43345,N_40054,N_41197);
xnor U43346 (N_43346,N_41520,N_41474);
or U43347 (N_43347,N_41683,N_41817);
or U43348 (N_43348,N_40527,N_40841);
or U43349 (N_43349,N_40443,N_41286);
xor U43350 (N_43350,N_40813,N_41385);
nor U43351 (N_43351,N_40856,N_40633);
nand U43352 (N_43352,N_40723,N_40868);
xor U43353 (N_43353,N_40902,N_40492);
nor U43354 (N_43354,N_40326,N_41466);
xnor U43355 (N_43355,N_40988,N_40482);
nand U43356 (N_43356,N_40855,N_40538);
or U43357 (N_43357,N_41012,N_41341);
and U43358 (N_43358,N_40555,N_41932);
nor U43359 (N_43359,N_40745,N_40747);
nor U43360 (N_43360,N_40019,N_41027);
xnor U43361 (N_43361,N_40221,N_40126);
xnor U43362 (N_43362,N_40323,N_40459);
or U43363 (N_43363,N_41453,N_41128);
or U43364 (N_43364,N_40674,N_40149);
nor U43365 (N_43365,N_40661,N_41349);
nor U43366 (N_43366,N_41346,N_41166);
and U43367 (N_43367,N_41056,N_40302);
nor U43368 (N_43368,N_41429,N_40256);
nor U43369 (N_43369,N_41204,N_41616);
nor U43370 (N_43370,N_41061,N_41252);
nor U43371 (N_43371,N_40959,N_40123);
nand U43372 (N_43372,N_41590,N_40028);
nor U43373 (N_43373,N_40780,N_40494);
or U43374 (N_43374,N_40024,N_40870);
xor U43375 (N_43375,N_41579,N_41881);
xnor U43376 (N_43376,N_40625,N_40231);
xnor U43377 (N_43377,N_40325,N_40752);
xor U43378 (N_43378,N_40083,N_40074);
or U43379 (N_43379,N_40388,N_40782);
xor U43380 (N_43380,N_41578,N_41476);
nand U43381 (N_43381,N_41266,N_40666);
xnor U43382 (N_43382,N_41580,N_41099);
and U43383 (N_43383,N_41927,N_40367);
or U43384 (N_43384,N_41597,N_41874);
and U43385 (N_43385,N_41533,N_41801);
nand U43386 (N_43386,N_41468,N_41828);
nand U43387 (N_43387,N_40845,N_41866);
nor U43388 (N_43388,N_40856,N_40646);
nor U43389 (N_43389,N_40732,N_40832);
nor U43390 (N_43390,N_41087,N_41275);
and U43391 (N_43391,N_41784,N_40521);
and U43392 (N_43392,N_41980,N_40982);
xor U43393 (N_43393,N_40639,N_40327);
or U43394 (N_43394,N_40726,N_41517);
and U43395 (N_43395,N_40495,N_40674);
nand U43396 (N_43396,N_41661,N_41321);
xnor U43397 (N_43397,N_40294,N_41549);
nand U43398 (N_43398,N_41693,N_41031);
and U43399 (N_43399,N_40786,N_40262);
and U43400 (N_43400,N_40882,N_40357);
xor U43401 (N_43401,N_41409,N_40188);
xor U43402 (N_43402,N_41063,N_40509);
or U43403 (N_43403,N_40971,N_41256);
xor U43404 (N_43404,N_40418,N_40018);
or U43405 (N_43405,N_41972,N_41820);
xor U43406 (N_43406,N_40010,N_41850);
xnor U43407 (N_43407,N_40133,N_40961);
and U43408 (N_43408,N_40598,N_41794);
nand U43409 (N_43409,N_40433,N_41907);
nor U43410 (N_43410,N_40570,N_40554);
nor U43411 (N_43411,N_41743,N_40743);
nand U43412 (N_43412,N_41260,N_41039);
nand U43413 (N_43413,N_41212,N_41621);
xnor U43414 (N_43414,N_41240,N_40572);
nor U43415 (N_43415,N_41092,N_40067);
nor U43416 (N_43416,N_40039,N_40091);
xnor U43417 (N_43417,N_41852,N_40550);
nor U43418 (N_43418,N_40142,N_41399);
or U43419 (N_43419,N_40407,N_40013);
nand U43420 (N_43420,N_41773,N_40664);
and U43421 (N_43421,N_40469,N_40241);
or U43422 (N_43422,N_40356,N_41799);
nor U43423 (N_43423,N_41345,N_40675);
or U43424 (N_43424,N_40501,N_41064);
or U43425 (N_43425,N_40402,N_41133);
xor U43426 (N_43426,N_41130,N_40150);
nand U43427 (N_43427,N_41785,N_41437);
nand U43428 (N_43428,N_41415,N_41155);
or U43429 (N_43429,N_41562,N_41820);
xor U43430 (N_43430,N_40903,N_40114);
and U43431 (N_43431,N_40193,N_41949);
and U43432 (N_43432,N_40859,N_40114);
nor U43433 (N_43433,N_40359,N_40418);
nor U43434 (N_43434,N_40003,N_40238);
or U43435 (N_43435,N_41154,N_41215);
or U43436 (N_43436,N_41585,N_40065);
xor U43437 (N_43437,N_41076,N_40480);
or U43438 (N_43438,N_40842,N_41833);
xnor U43439 (N_43439,N_41827,N_40627);
and U43440 (N_43440,N_41608,N_40642);
and U43441 (N_43441,N_41558,N_40911);
nand U43442 (N_43442,N_40351,N_40743);
xor U43443 (N_43443,N_41060,N_40753);
nor U43444 (N_43444,N_40361,N_40454);
and U43445 (N_43445,N_40732,N_41828);
nand U43446 (N_43446,N_40181,N_40571);
or U43447 (N_43447,N_41511,N_40900);
or U43448 (N_43448,N_41031,N_41568);
or U43449 (N_43449,N_40359,N_40688);
xor U43450 (N_43450,N_41734,N_40722);
nor U43451 (N_43451,N_41970,N_41850);
and U43452 (N_43452,N_41177,N_40703);
xor U43453 (N_43453,N_41097,N_40501);
nand U43454 (N_43454,N_41413,N_41130);
and U43455 (N_43455,N_40506,N_41754);
nand U43456 (N_43456,N_41632,N_41125);
or U43457 (N_43457,N_40536,N_41849);
or U43458 (N_43458,N_41634,N_40720);
or U43459 (N_43459,N_41724,N_40096);
xor U43460 (N_43460,N_40307,N_40887);
nor U43461 (N_43461,N_41945,N_40392);
or U43462 (N_43462,N_41398,N_40305);
or U43463 (N_43463,N_40018,N_41315);
and U43464 (N_43464,N_40894,N_41736);
xor U43465 (N_43465,N_40748,N_40239);
and U43466 (N_43466,N_41252,N_40809);
xnor U43467 (N_43467,N_41958,N_40956);
and U43468 (N_43468,N_40947,N_41245);
nor U43469 (N_43469,N_40777,N_40934);
or U43470 (N_43470,N_41104,N_41755);
and U43471 (N_43471,N_40180,N_41055);
and U43472 (N_43472,N_41396,N_40802);
nand U43473 (N_43473,N_40339,N_40083);
and U43474 (N_43474,N_40708,N_40039);
or U43475 (N_43475,N_40878,N_41911);
nor U43476 (N_43476,N_40058,N_40202);
xor U43477 (N_43477,N_41733,N_40547);
nand U43478 (N_43478,N_41600,N_41237);
and U43479 (N_43479,N_40948,N_40035);
nand U43480 (N_43480,N_41526,N_41989);
nand U43481 (N_43481,N_41273,N_41437);
nand U43482 (N_43482,N_40049,N_40690);
nand U43483 (N_43483,N_40420,N_40376);
nor U43484 (N_43484,N_41678,N_41979);
nor U43485 (N_43485,N_40756,N_40742);
or U43486 (N_43486,N_41667,N_40955);
or U43487 (N_43487,N_40171,N_41623);
nor U43488 (N_43488,N_40889,N_40023);
xor U43489 (N_43489,N_40898,N_41123);
and U43490 (N_43490,N_41718,N_40746);
xnor U43491 (N_43491,N_41550,N_40347);
nor U43492 (N_43492,N_40946,N_40124);
or U43493 (N_43493,N_41618,N_41282);
or U43494 (N_43494,N_40597,N_41861);
or U43495 (N_43495,N_41578,N_41134);
xnor U43496 (N_43496,N_41736,N_41309);
nor U43497 (N_43497,N_40443,N_40020);
nand U43498 (N_43498,N_40829,N_41295);
or U43499 (N_43499,N_40238,N_41989);
and U43500 (N_43500,N_41262,N_41490);
or U43501 (N_43501,N_40641,N_40699);
nor U43502 (N_43502,N_41327,N_41116);
and U43503 (N_43503,N_41290,N_41460);
or U43504 (N_43504,N_40019,N_40129);
xnor U43505 (N_43505,N_40590,N_41557);
or U43506 (N_43506,N_41046,N_40835);
and U43507 (N_43507,N_40264,N_40271);
nor U43508 (N_43508,N_41085,N_41119);
xor U43509 (N_43509,N_41686,N_41995);
nor U43510 (N_43510,N_40613,N_41877);
and U43511 (N_43511,N_40386,N_41088);
and U43512 (N_43512,N_40430,N_41880);
or U43513 (N_43513,N_41102,N_40884);
nand U43514 (N_43514,N_40460,N_40236);
and U43515 (N_43515,N_40746,N_41902);
xnor U43516 (N_43516,N_40134,N_41815);
and U43517 (N_43517,N_41702,N_40991);
nand U43518 (N_43518,N_40600,N_40816);
and U43519 (N_43519,N_41069,N_41870);
nand U43520 (N_43520,N_40178,N_41279);
nand U43521 (N_43521,N_41277,N_41961);
and U43522 (N_43522,N_40740,N_41451);
xor U43523 (N_43523,N_41159,N_40476);
xnor U43524 (N_43524,N_40110,N_40607);
and U43525 (N_43525,N_40683,N_40164);
nor U43526 (N_43526,N_40896,N_41592);
or U43527 (N_43527,N_40868,N_41104);
or U43528 (N_43528,N_40194,N_41421);
nand U43529 (N_43529,N_41822,N_40174);
or U43530 (N_43530,N_40416,N_40401);
or U43531 (N_43531,N_40278,N_40144);
or U43532 (N_43532,N_41233,N_40455);
or U43533 (N_43533,N_40920,N_41763);
and U43534 (N_43534,N_40531,N_40419);
or U43535 (N_43535,N_41458,N_41038);
and U43536 (N_43536,N_41765,N_40279);
xnor U43537 (N_43537,N_40561,N_40777);
and U43538 (N_43538,N_40056,N_40003);
nor U43539 (N_43539,N_40800,N_40979);
and U43540 (N_43540,N_41350,N_40059);
nand U43541 (N_43541,N_40544,N_41289);
and U43542 (N_43542,N_41239,N_40228);
or U43543 (N_43543,N_41642,N_40327);
nand U43544 (N_43544,N_41546,N_40265);
or U43545 (N_43545,N_40890,N_41478);
nand U43546 (N_43546,N_41239,N_41583);
nor U43547 (N_43547,N_40265,N_41399);
or U43548 (N_43548,N_40846,N_41848);
or U43549 (N_43549,N_41111,N_41972);
nand U43550 (N_43550,N_40266,N_40492);
xor U43551 (N_43551,N_41886,N_40127);
nand U43552 (N_43552,N_40311,N_41848);
nand U43553 (N_43553,N_41353,N_41337);
or U43554 (N_43554,N_40313,N_41715);
nand U43555 (N_43555,N_40912,N_41034);
xor U43556 (N_43556,N_40988,N_41959);
nand U43557 (N_43557,N_40749,N_41755);
or U43558 (N_43558,N_40700,N_41535);
xor U43559 (N_43559,N_40402,N_41044);
nor U43560 (N_43560,N_41937,N_41417);
and U43561 (N_43561,N_41613,N_40267);
and U43562 (N_43562,N_41601,N_40603);
and U43563 (N_43563,N_40855,N_40366);
xor U43564 (N_43564,N_41540,N_40206);
and U43565 (N_43565,N_40250,N_41980);
nor U43566 (N_43566,N_41309,N_40628);
and U43567 (N_43567,N_40638,N_40203);
xnor U43568 (N_43568,N_41890,N_40578);
xnor U43569 (N_43569,N_40966,N_41225);
or U43570 (N_43570,N_41031,N_41139);
nor U43571 (N_43571,N_41640,N_40024);
or U43572 (N_43572,N_40962,N_41020);
or U43573 (N_43573,N_40508,N_40089);
and U43574 (N_43574,N_40424,N_41145);
nand U43575 (N_43575,N_41409,N_40938);
and U43576 (N_43576,N_41315,N_41675);
nor U43577 (N_43577,N_41023,N_40855);
xor U43578 (N_43578,N_41854,N_41183);
xor U43579 (N_43579,N_40093,N_41693);
xnor U43580 (N_43580,N_41454,N_41904);
xor U43581 (N_43581,N_40974,N_40498);
nor U43582 (N_43582,N_41481,N_41621);
or U43583 (N_43583,N_40087,N_40869);
xnor U43584 (N_43584,N_40336,N_40299);
or U43585 (N_43585,N_40698,N_41020);
xnor U43586 (N_43586,N_41543,N_41049);
and U43587 (N_43587,N_41643,N_40633);
xor U43588 (N_43588,N_41553,N_40386);
or U43589 (N_43589,N_40773,N_41410);
nor U43590 (N_43590,N_40359,N_41846);
nand U43591 (N_43591,N_40545,N_41604);
nand U43592 (N_43592,N_41749,N_40995);
nor U43593 (N_43593,N_41663,N_41675);
xor U43594 (N_43594,N_41202,N_41983);
xor U43595 (N_43595,N_40215,N_40651);
nor U43596 (N_43596,N_41190,N_41648);
or U43597 (N_43597,N_41713,N_41949);
or U43598 (N_43598,N_40516,N_41067);
nor U43599 (N_43599,N_40228,N_41505);
and U43600 (N_43600,N_41923,N_40459);
and U43601 (N_43601,N_41358,N_40533);
and U43602 (N_43602,N_41734,N_41561);
nor U43603 (N_43603,N_41916,N_40627);
nand U43604 (N_43604,N_40924,N_40162);
xnor U43605 (N_43605,N_40375,N_41283);
or U43606 (N_43606,N_41964,N_40798);
xnor U43607 (N_43607,N_41065,N_41984);
nand U43608 (N_43608,N_40791,N_40642);
or U43609 (N_43609,N_41694,N_40993);
or U43610 (N_43610,N_41051,N_41348);
nand U43611 (N_43611,N_41918,N_41180);
xnor U43612 (N_43612,N_41265,N_40296);
nand U43613 (N_43613,N_40169,N_40988);
nor U43614 (N_43614,N_41875,N_40644);
and U43615 (N_43615,N_41676,N_40858);
and U43616 (N_43616,N_41737,N_40755);
xnor U43617 (N_43617,N_40858,N_40106);
or U43618 (N_43618,N_40788,N_40122);
and U43619 (N_43619,N_41487,N_40191);
xor U43620 (N_43620,N_40911,N_41542);
or U43621 (N_43621,N_40339,N_40023);
xor U43622 (N_43622,N_40724,N_41296);
nor U43623 (N_43623,N_40115,N_41075);
xnor U43624 (N_43624,N_40374,N_41765);
and U43625 (N_43625,N_40595,N_41045);
nand U43626 (N_43626,N_40107,N_41786);
nor U43627 (N_43627,N_41241,N_41392);
or U43628 (N_43628,N_40111,N_41602);
nand U43629 (N_43629,N_41323,N_41100);
nor U43630 (N_43630,N_41331,N_40897);
nor U43631 (N_43631,N_40760,N_41479);
or U43632 (N_43632,N_41763,N_40811);
or U43633 (N_43633,N_41436,N_41804);
or U43634 (N_43634,N_40784,N_41966);
nor U43635 (N_43635,N_40120,N_41568);
or U43636 (N_43636,N_41414,N_40662);
xor U43637 (N_43637,N_40554,N_40919);
or U43638 (N_43638,N_41261,N_40890);
and U43639 (N_43639,N_40316,N_41209);
xor U43640 (N_43640,N_41151,N_40674);
xnor U43641 (N_43641,N_41950,N_41567);
xnor U43642 (N_43642,N_40317,N_40446);
and U43643 (N_43643,N_41978,N_41533);
and U43644 (N_43644,N_40202,N_40455);
and U43645 (N_43645,N_40637,N_40942);
nand U43646 (N_43646,N_40125,N_41158);
or U43647 (N_43647,N_41877,N_40677);
nand U43648 (N_43648,N_41568,N_41087);
and U43649 (N_43649,N_41131,N_40590);
xnor U43650 (N_43650,N_40506,N_41951);
nor U43651 (N_43651,N_40917,N_41567);
nand U43652 (N_43652,N_41946,N_41669);
or U43653 (N_43653,N_40066,N_41066);
xnor U43654 (N_43654,N_40473,N_41355);
or U43655 (N_43655,N_40836,N_40313);
nand U43656 (N_43656,N_40521,N_40501);
nor U43657 (N_43657,N_41066,N_40160);
or U43658 (N_43658,N_40857,N_41916);
nand U43659 (N_43659,N_41679,N_40476);
and U43660 (N_43660,N_41149,N_40620);
nand U43661 (N_43661,N_41180,N_40656);
xnor U43662 (N_43662,N_40625,N_40822);
or U43663 (N_43663,N_40071,N_41004);
or U43664 (N_43664,N_40238,N_40291);
xnor U43665 (N_43665,N_41940,N_41021);
or U43666 (N_43666,N_41591,N_40056);
xor U43667 (N_43667,N_40444,N_40980);
and U43668 (N_43668,N_41455,N_40328);
nor U43669 (N_43669,N_40735,N_41055);
xor U43670 (N_43670,N_41244,N_40734);
and U43671 (N_43671,N_41001,N_40200);
or U43672 (N_43672,N_41329,N_40107);
nand U43673 (N_43673,N_41750,N_40521);
and U43674 (N_43674,N_41869,N_40087);
xor U43675 (N_43675,N_40171,N_40134);
and U43676 (N_43676,N_40594,N_40144);
or U43677 (N_43677,N_40235,N_40541);
xor U43678 (N_43678,N_41139,N_41070);
xor U43679 (N_43679,N_41329,N_41946);
xor U43680 (N_43680,N_40341,N_41193);
nand U43681 (N_43681,N_41498,N_41351);
and U43682 (N_43682,N_40147,N_40951);
nand U43683 (N_43683,N_41527,N_41442);
xor U43684 (N_43684,N_40041,N_41333);
nor U43685 (N_43685,N_40915,N_41777);
nor U43686 (N_43686,N_41900,N_40456);
nand U43687 (N_43687,N_40678,N_40799);
and U43688 (N_43688,N_41513,N_41924);
or U43689 (N_43689,N_40137,N_41459);
and U43690 (N_43690,N_41949,N_41830);
xnor U43691 (N_43691,N_41897,N_41121);
nand U43692 (N_43692,N_40077,N_41059);
nand U43693 (N_43693,N_41886,N_40696);
and U43694 (N_43694,N_40097,N_40980);
or U43695 (N_43695,N_40709,N_41365);
nor U43696 (N_43696,N_40798,N_40073);
xnor U43697 (N_43697,N_41159,N_40321);
nor U43698 (N_43698,N_40851,N_40782);
or U43699 (N_43699,N_41858,N_40710);
nand U43700 (N_43700,N_41342,N_40046);
xnor U43701 (N_43701,N_40911,N_41231);
or U43702 (N_43702,N_41101,N_40664);
or U43703 (N_43703,N_40248,N_40956);
or U43704 (N_43704,N_40808,N_40015);
or U43705 (N_43705,N_40209,N_41943);
nor U43706 (N_43706,N_41975,N_41791);
nand U43707 (N_43707,N_40192,N_40215);
xnor U43708 (N_43708,N_41557,N_41528);
and U43709 (N_43709,N_40414,N_41023);
or U43710 (N_43710,N_41777,N_41697);
and U43711 (N_43711,N_40380,N_41664);
nand U43712 (N_43712,N_40457,N_41206);
nor U43713 (N_43713,N_41728,N_40648);
nor U43714 (N_43714,N_41640,N_41677);
nor U43715 (N_43715,N_41767,N_40598);
and U43716 (N_43716,N_41487,N_41241);
xor U43717 (N_43717,N_40401,N_41846);
or U43718 (N_43718,N_41100,N_41592);
xor U43719 (N_43719,N_41778,N_40899);
or U43720 (N_43720,N_40069,N_41800);
xnor U43721 (N_43721,N_40921,N_40803);
nor U43722 (N_43722,N_41239,N_40954);
and U43723 (N_43723,N_40802,N_40270);
nand U43724 (N_43724,N_40897,N_40439);
and U43725 (N_43725,N_41211,N_40327);
nand U43726 (N_43726,N_41494,N_40036);
or U43727 (N_43727,N_40996,N_40729);
nor U43728 (N_43728,N_41403,N_41215);
nor U43729 (N_43729,N_41551,N_40020);
nand U43730 (N_43730,N_40701,N_40859);
xor U43731 (N_43731,N_40894,N_40537);
or U43732 (N_43732,N_40115,N_41371);
or U43733 (N_43733,N_41533,N_40477);
or U43734 (N_43734,N_40009,N_41748);
nand U43735 (N_43735,N_40643,N_41438);
nor U43736 (N_43736,N_41034,N_40310);
xnor U43737 (N_43737,N_40721,N_41522);
nor U43738 (N_43738,N_40338,N_41431);
and U43739 (N_43739,N_41004,N_41209);
nand U43740 (N_43740,N_40181,N_40659);
and U43741 (N_43741,N_41574,N_40130);
nand U43742 (N_43742,N_40514,N_41935);
and U43743 (N_43743,N_41659,N_40739);
nor U43744 (N_43744,N_41080,N_41795);
xnor U43745 (N_43745,N_40741,N_40464);
xnor U43746 (N_43746,N_40594,N_41730);
xnor U43747 (N_43747,N_41762,N_40061);
xnor U43748 (N_43748,N_41890,N_41139);
and U43749 (N_43749,N_41508,N_41438);
nor U43750 (N_43750,N_41562,N_40478);
nand U43751 (N_43751,N_41127,N_40747);
nand U43752 (N_43752,N_41794,N_40933);
and U43753 (N_43753,N_40829,N_41282);
nor U43754 (N_43754,N_41515,N_41768);
or U43755 (N_43755,N_40593,N_40886);
nor U43756 (N_43756,N_41295,N_41555);
xor U43757 (N_43757,N_41317,N_40912);
nand U43758 (N_43758,N_41293,N_41218);
nor U43759 (N_43759,N_41693,N_40828);
nor U43760 (N_43760,N_41638,N_40045);
xor U43761 (N_43761,N_41370,N_40462);
nor U43762 (N_43762,N_40548,N_40159);
nand U43763 (N_43763,N_40500,N_41899);
or U43764 (N_43764,N_40443,N_41938);
xnor U43765 (N_43765,N_40366,N_41009);
nand U43766 (N_43766,N_40357,N_41323);
or U43767 (N_43767,N_40894,N_40757);
xnor U43768 (N_43768,N_41052,N_40913);
or U43769 (N_43769,N_40296,N_41262);
nor U43770 (N_43770,N_40013,N_40582);
and U43771 (N_43771,N_40484,N_41996);
and U43772 (N_43772,N_41346,N_41435);
nor U43773 (N_43773,N_40492,N_40694);
xor U43774 (N_43774,N_40458,N_40608);
and U43775 (N_43775,N_41101,N_40616);
and U43776 (N_43776,N_41863,N_41123);
nand U43777 (N_43777,N_40916,N_41882);
nor U43778 (N_43778,N_40977,N_41988);
and U43779 (N_43779,N_41254,N_40879);
nor U43780 (N_43780,N_41516,N_41547);
or U43781 (N_43781,N_40303,N_41528);
and U43782 (N_43782,N_41551,N_40210);
or U43783 (N_43783,N_41145,N_40929);
nor U43784 (N_43784,N_41272,N_41244);
or U43785 (N_43785,N_41804,N_40276);
nand U43786 (N_43786,N_40837,N_41142);
and U43787 (N_43787,N_41751,N_40663);
nand U43788 (N_43788,N_41396,N_40933);
nor U43789 (N_43789,N_41082,N_40961);
nor U43790 (N_43790,N_41992,N_41592);
and U43791 (N_43791,N_41974,N_40723);
or U43792 (N_43792,N_41812,N_41379);
nand U43793 (N_43793,N_40506,N_40949);
or U43794 (N_43794,N_41347,N_41056);
or U43795 (N_43795,N_41199,N_40507);
and U43796 (N_43796,N_41555,N_41122);
or U43797 (N_43797,N_40805,N_40916);
nand U43798 (N_43798,N_40797,N_41426);
or U43799 (N_43799,N_41906,N_41563);
nor U43800 (N_43800,N_40324,N_40340);
xor U43801 (N_43801,N_41121,N_41786);
and U43802 (N_43802,N_40242,N_41445);
and U43803 (N_43803,N_41611,N_41401);
or U43804 (N_43804,N_40862,N_40894);
nor U43805 (N_43805,N_40012,N_40580);
and U43806 (N_43806,N_40510,N_40405);
nand U43807 (N_43807,N_40420,N_40444);
or U43808 (N_43808,N_41365,N_41202);
and U43809 (N_43809,N_41691,N_40058);
nor U43810 (N_43810,N_40391,N_40936);
xnor U43811 (N_43811,N_41778,N_41185);
and U43812 (N_43812,N_41200,N_41442);
or U43813 (N_43813,N_41543,N_40595);
or U43814 (N_43814,N_40148,N_40197);
nor U43815 (N_43815,N_41538,N_41701);
nor U43816 (N_43816,N_40119,N_40551);
or U43817 (N_43817,N_41756,N_41797);
nor U43818 (N_43818,N_41253,N_41408);
nand U43819 (N_43819,N_41078,N_41406);
xor U43820 (N_43820,N_40988,N_41919);
nor U43821 (N_43821,N_41858,N_40701);
xor U43822 (N_43822,N_41241,N_41976);
nand U43823 (N_43823,N_40299,N_41445);
nor U43824 (N_43824,N_40338,N_41232);
nand U43825 (N_43825,N_40424,N_40112);
xor U43826 (N_43826,N_41653,N_40962);
nand U43827 (N_43827,N_40549,N_40851);
and U43828 (N_43828,N_41589,N_41849);
nand U43829 (N_43829,N_40261,N_41031);
and U43830 (N_43830,N_40962,N_41749);
nor U43831 (N_43831,N_40528,N_41732);
xor U43832 (N_43832,N_41874,N_40409);
nor U43833 (N_43833,N_40227,N_40281);
nor U43834 (N_43834,N_40545,N_41996);
and U43835 (N_43835,N_41109,N_41205);
nor U43836 (N_43836,N_40422,N_41455);
nor U43837 (N_43837,N_41879,N_41292);
xnor U43838 (N_43838,N_40372,N_41017);
nand U43839 (N_43839,N_41920,N_40718);
and U43840 (N_43840,N_41615,N_40174);
and U43841 (N_43841,N_40010,N_41602);
xnor U43842 (N_43842,N_40268,N_41736);
xnor U43843 (N_43843,N_40437,N_41955);
nor U43844 (N_43844,N_40777,N_40877);
or U43845 (N_43845,N_40726,N_40090);
or U43846 (N_43846,N_41882,N_40191);
and U43847 (N_43847,N_40796,N_40032);
nor U43848 (N_43848,N_40503,N_40614);
and U43849 (N_43849,N_40352,N_40206);
or U43850 (N_43850,N_40443,N_40862);
nor U43851 (N_43851,N_40003,N_40409);
or U43852 (N_43852,N_41436,N_41454);
and U43853 (N_43853,N_41933,N_40758);
xor U43854 (N_43854,N_41486,N_41809);
xnor U43855 (N_43855,N_40414,N_40747);
nand U43856 (N_43856,N_40465,N_41037);
nor U43857 (N_43857,N_41676,N_40215);
nand U43858 (N_43858,N_40692,N_41885);
nor U43859 (N_43859,N_40469,N_40957);
nand U43860 (N_43860,N_40305,N_41529);
nand U43861 (N_43861,N_40153,N_40998);
or U43862 (N_43862,N_41323,N_41310);
nand U43863 (N_43863,N_41327,N_40867);
and U43864 (N_43864,N_40585,N_40243);
nand U43865 (N_43865,N_41098,N_40697);
xnor U43866 (N_43866,N_41965,N_40844);
xnor U43867 (N_43867,N_41103,N_40494);
and U43868 (N_43868,N_41602,N_40565);
nor U43869 (N_43869,N_41856,N_40170);
and U43870 (N_43870,N_40709,N_40882);
xnor U43871 (N_43871,N_41881,N_41629);
or U43872 (N_43872,N_41179,N_40505);
or U43873 (N_43873,N_40075,N_41402);
nor U43874 (N_43874,N_40578,N_41355);
nor U43875 (N_43875,N_40120,N_40784);
or U43876 (N_43876,N_40748,N_40141);
or U43877 (N_43877,N_40951,N_41493);
nor U43878 (N_43878,N_41536,N_40201);
and U43879 (N_43879,N_40113,N_41611);
xnor U43880 (N_43880,N_40070,N_40728);
nand U43881 (N_43881,N_40204,N_40103);
or U43882 (N_43882,N_40209,N_40915);
xor U43883 (N_43883,N_40765,N_41865);
xnor U43884 (N_43884,N_41482,N_40299);
or U43885 (N_43885,N_40722,N_41522);
xnor U43886 (N_43886,N_41290,N_41865);
or U43887 (N_43887,N_41560,N_40633);
or U43888 (N_43888,N_41834,N_40500);
and U43889 (N_43889,N_41075,N_41790);
and U43890 (N_43890,N_40536,N_40723);
xor U43891 (N_43891,N_40555,N_40770);
or U43892 (N_43892,N_40577,N_40399);
and U43893 (N_43893,N_41877,N_40398);
and U43894 (N_43894,N_40329,N_40861);
and U43895 (N_43895,N_41120,N_40239);
nand U43896 (N_43896,N_41232,N_40539);
and U43897 (N_43897,N_40995,N_40259);
xnor U43898 (N_43898,N_41195,N_41810);
or U43899 (N_43899,N_40002,N_40887);
xor U43900 (N_43900,N_40852,N_40129);
nor U43901 (N_43901,N_40458,N_41803);
xor U43902 (N_43902,N_40677,N_41865);
nand U43903 (N_43903,N_40134,N_41870);
or U43904 (N_43904,N_41033,N_41543);
and U43905 (N_43905,N_40222,N_40277);
nand U43906 (N_43906,N_40763,N_41395);
and U43907 (N_43907,N_41590,N_40760);
and U43908 (N_43908,N_41306,N_41968);
xor U43909 (N_43909,N_41546,N_40134);
nor U43910 (N_43910,N_41260,N_41253);
nand U43911 (N_43911,N_41328,N_40377);
nand U43912 (N_43912,N_40440,N_40628);
nand U43913 (N_43913,N_41620,N_41887);
or U43914 (N_43914,N_41038,N_41109);
nand U43915 (N_43915,N_41782,N_40122);
or U43916 (N_43916,N_41154,N_40259);
or U43917 (N_43917,N_41891,N_40355);
nand U43918 (N_43918,N_41013,N_41118);
xnor U43919 (N_43919,N_40061,N_40597);
nor U43920 (N_43920,N_40942,N_40348);
and U43921 (N_43921,N_41968,N_40186);
or U43922 (N_43922,N_40546,N_41096);
nand U43923 (N_43923,N_40851,N_40840);
nor U43924 (N_43924,N_40179,N_41550);
xor U43925 (N_43925,N_40289,N_41029);
xor U43926 (N_43926,N_41851,N_41957);
nand U43927 (N_43927,N_40572,N_40086);
and U43928 (N_43928,N_41750,N_40977);
nand U43929 (N_43929,N_40866,N_40882);
nor U43930 (N_43930,N_41118,N_40470);
xnor U43931 (N_43931,N_40050,N_40613);
or U43932 (N_43932,N_40032,N_41623);
nor U43933 (N_43933,N_40796,N_40950);
xnor U43934 (N_43934,N_40498,N_41200);
nand U43935 (N_43935,N_41486,N_41631);
or U43936 (N_43936,N_41628,N_41860);
nor U43937 (N_43937,N_40038,N_41786);
or U43938 (N_43938,N_41437,N_40734);
nor U43939 (N_43939,N_41641,N_41948);
xnor U43940 (N_43940,N_41296,N_41574);
or U43941 (N_43941,N_40465,N_41328);
nor U43942 (N_43942,N_40443,N_40101);
nand U43943 (N_43943,N_40804,N_41148);
xor U43944 (N_43944,N_41977,N_41316);
and U43945 (N_43945,N_41206,N_40348);
and U43946 (N_43946,N_40952,N_41603);
xnor U43947 (N_43947,N_41611,N_40361);
nor U43948 (N_43948,N_41313,N_40816);
and U43949 (N_43949,N_41096,N_41361);
nand U43950 (N_43950,N_40452,N_41490);
or U43951 (N_43951,N_41634,N_41426);
and U43952 (N_43952,N_41064,N_40258);
nand U43953 (N_43953,N_40711,N_40733);
xor U43954 (N_43954,N_41298,N_41232);
xnor U43955 (N_43955,N_41439,N_40601);
nor U43956 (N_43956,N_40273,N_40463);
and U43957 (N_43957,N_40210,N_40658);
or U43958 (N_43958,N_40726,N_40228);
or U43959 (N_43959,N_40023,N_41467);
nor U43960 (N_43960,N_41323,N_40343);
nand U43961 (N_43961,N_41577,N_41250);
or U43962 (N_43962,N_40748,N_41332);
or U43963 (N_43963,N_41819,N_40172);
or U43964 (N_43964,N_41000,N_41776);
and U43965 (N_43965,N_41504,N_40917);
xor U43966 (N_43966,N_40404,N_40182);
nand U43967 (N_43967,N_40304,N_41866);
or U43968 (N_43968,N_41775,N_41305);
xnor U43969 (N_43969,N_40857,N_41062);
or U43970 (N_43970,N_40159,N_41079);
nand U43971 (N_43971,N_41551,N_41250);
nor U43972 (N_43972,N_41959,N_40800);
and U43973 (N_43973,N_41475,N_41494);
nand U43974 (N_43974,N_40246,N_41202);
nand U43975 (N_43975,N_40968,N_41588);
or U43976 (N_43976,N_41453,N_41849);
nand U43977 (N_43977,N_40587,N_40912);
or U43978 (N_43978,N_40576,N_41846);
xnor U43979 (N_43979,N_41773,N_40392);
and U43980 (N_43980,N_40114,N_41933);
nand U43981 (N_43981,N_40115,N_40973);
and U43982 (N_43982,N_41396,N_41249);
nor U43983 (N_43983,N_41538,N_41910);
nor U43984 (N_43984,N_40859,N_40620);
nor U43985 (N_43985,N_40211,N_41920);
and U43986 (N_43986,N_41210,N_40276);
xnor U43987 (N_43987,N_40454,N_40778);
nand U43988 (N_43988,N_41155,N_40610);
nor U43989 (N_43989,N_41639,N_41444);
or U43990 (N_43990,N_40919,N_40869);
xor U43991 (N_43991,N_40060,N_41646);
and U43992 (N_43992,N_41700,N_40232);
nor U43993 (N_43993,N_40590,N_41187);
or U43994 (N_43994,N_41865,N_40832);
nand U43995 (N_43995,N_41332,N_40434);
and U43996 (N_43996,N_40950,N_41044);
nor U43997 (N_43997,N_41232,N_41825);
or U43998 (N_43998,N_40391,N_41719);
or U43999 (N_43999,N_41056,N_41266);
xor U44000 (N_44000,N_42265,N_43426);
xor U44001 (N_44001,N_42975,N_42856);
nor U44002 (N_44002,N_43532,N_42101);
nor U44003 (N_44003,N_42325,N_43933);
nand U44004 (N_44004,N_42873,N_42755);
nand U44005 (N_44005,N_43405,N_42296);
xnor U44006 (N_44006,N_42528,N_43095);
or U44007 (N_44007,N_43615,N_43288);
nor U44008 (N_44008,N_42716,N_42200);
and U44009 (N_44009,N_43300,N_42159);
or U44010 (N_44010,N_43268,N_43726);
or U44011 (N_44011,N_42480,N_42401);
and U44012 (N_44012,N_42494,N_43780);
nand U44013 (N_44013,N_42854,N_42525);
nand U44014 (N_44014,N_43092,N_43454);
xnor U44015 (N_44015,N_42710,N_43896);
nand U44016 (N_44016,N_43675,N_43919);
xor U44017 (N_44017,N_42523,N_42366);
nor U44018 (N_44018,N_43473,N_42505);
and U44019 (N_44019,N_42536,N_42396);
nor U44020 (N_44020,N_43635,N_43321);
xnor U44021 (N_44021,N_42133,N_43330);
and U44022 (N_44022,N_43350,N_42051);
nor U44023 (N_44023,N_42287,N_43659);
xor U44024 (N_44024,N_43966,N_43328);
and U44025 (N_44025,N_43179,N_42823);
and U44026 (N_44026,N_42979,N_43612);
nor U44027 (N_44027,N_43723,N_43779);
nand U44028 (N_44028,N_42499,N_43510);
nand U44029 (N_44029,N_42583,N_42461);
nand U44030 (N_44030,N_42920,N_43741);
or U44031 (N_44031,N_43442,N_43724);
nand U44032 (N_44032,N_42228,N_42564);
or U44033 (N_44033,N_42596,N_43422);
nor U44034 (N_44034,N_42207,N_42286);
or U44035 (N_44035,N_43519,N_42990);
and U44036 (N_44036,N_42481,N_42758);
and U44037 (N_44037,N_42273,N_42322);
nand U44038 (N_44038,N_42683,N_42381);
or U44039 (N_44039,N_43208,N_43381);
nand U44040 (N_44040,N_43900,N_43667);
and U44041 (N_44041,N_43834,N_43359);
or U44042 (N_44042,N_43531,N_43158);
or U44043 (N_44043,N_43607,N_43941);
nor U44044 (N_44044,N_43589,N_43820);
or U44045 (N_44045,N_42341,N_42654);
nor U44046 (N_44046,N_43694,N_43545);
nor U44047 (N_44047,N_43560,N_42387);
xor U44048 (N_44048,N_43989,N_42967);
xor U44049 (N_44049,N_42139,N_43187);
or U44050 (N_44050,N_43700,N_42037);
nor U44051 (N_44051,N_42509,N_42684);
xor U44052 (N_44052,N_43656,N_42947);
nor U44053 (N_44053,N_42548,N_43790);
nand U44054 (N_44054,N_43879,N_42867);
nor U44055 (N_44055,N_43735,N_43356);
and U44056 (N_44056,N_43807,N_43235);
xnor U44057 (N_44057,N_43291,N_42250);
xnor U44058 (N_44058,N_42812,N_42246);
xnor U44059 (N_44059,N_42306,N_42877);
nand U44060 (N_44060,N_42456,N_43445);
nand U44061 (N_44061,N_42348,N_42451);
xnor U44062 (N_44062,N_42060,N_42665);
nand U44063 (N_44063,N_42066,N_43410);
and U44064 (N_44064,N_43468,N_43903);
and U44065 (N_44065,N_42421,N_42516);
nand U44066 (N_44066,N_43523,N_43110);
nor U44067 (N_44067,N_42188,N_42019);
xor U44068 (N_44068,N_43222,N_42978);
nand U44069 (N_44069,N_43928,N_43809);
xnor U44070 (N_44070,N_43249,N_42989);
and U44071 (N_44071,N_43793,N_43492);
or U44072 (N_44072,N_42770,N_42988);
nor U44073 (N_44073,N_42468,N_42087);
nand U44074 (N_44074,N_43768,N_42125);
xor U44075 (N_44075,N_42760,N_42734);
xor U44076 (N_44076,N_42879,N_42437);
and U44077 (N_44077,N_42913,N_43916);
xnor U44078 (N_44078,N_43509,N_42476);
xnor U44079 (N_44079,N_43609,N_42206);
xor U44080 (N_44080,N_43574,N_43148);
nor U44081 (N_44081,N_42094,N_42722);
xnor U44082 (N_44082,N_42418,N_43645);
xnor U44083 (N_44083,N_43096,N_43565);
xnor U44084 (N_44084,N_42930,N_43155);
xor U44085 (N_44085,N_42490,N_43596);
nor U44086 (N_44086,N_43011,N_43149);
xor U44087 (N_44087,N_43870,N_42338);
xor U44088 (N_44088,N_43296,N_43844);
and U44089 (N_44089,N_42120,N_43062);
and U44090 (N_44090,N_42268,N_42283);
or U44091 (N_44091,N_42068,N_42891);
xor U44092 (N_44092,N_42906,N_43009);
nand U44093 (N_44093,N_43570,N_43542);
nand U44094 (N_44094,N_43465,N_43230);
nand U44095 (N_44095,N_43353,N_43976);
and U44096 (N_44096,N_42141,N_43457);
nor U44097 (N_44097,N_42969,N_42820);
nor U44098 (N_44098,N_43681,N_43898);
and U44099 (N_44099,N_43354,N_43854);
nor U44100 (N_44100,N_42416,N_42460);
nand U44101 (N_44101,N_43950,N_42897);
xnor U44102 (N_44102,N_42963,N_43205);
xor U44103 (N_44103,N_42715,N_42303);
xnor U44104 (N_44104,N_43083,N_42669);
xor U44105 (N_44105,N_43070,N_42714);
nand U44106 (N_44106,N_42189,N_43335);
nor U44107 (N_44107,N_42049,N_42732);
or U44108 (N_44108,N_42332,N_42771);
xnor U44109 (N_44109,N_43924,N_42956);
xnor U44110 (N_44110,N_43974,N_42233);
and U44111 (N_44111,N_42796,N_42953);
or U44112 (N_44112,N_42198,N_42545);
and U44113 (N_44113,N_43409,N_42199);
or U44114 (N_44114,N_43370,N_42067);
and U44115 (N_44115,N_42522,N_43622);
or U44116 (N_44116,N_43676,N_42267);
nand U44117 (N_44117,N_43481,N_42748);
or U44118 (N_44118,N_43555,N_42933);
or U44119 (N_44119,N_43057,N_43623);
or U44120 (N_44120,N_42290,N_42939);
or U44121 (N_44121,N_42797,N_42475);
nor U44122 (N_44122,N_42254,N_42258);
xor U44123 (N_44123,N_43411,N_42831);
or U44124 (N_44124,N_43026,N_43526);
and U44125 (N_44125,N_43434,N_42380);
nor U44126 (N_44126,N_43297,N_43628);
nor U44127 (N_44127,N_43708,N_43392);
or U44128 (N_44128,N_42036,N_42657);
nor U44129 (N_44129,N_42833,N_43818);
nand U44130 (N_44130,N_42343,N_42680);
nor U44131 (N_44131,N_42048,N_42574);
or U44132 (N_44132,N_43488,N_43241);
nand U44133 (N_44133,N_43051,N_43355);
nor U44134 (N_44134,N_43416,N_43498);
xnor U44135 (N_44135,N_42183,N_42486);
or U44136 (N_44136,N_43730,N_42663);
xor U44137 (N_44137,N_42294,N_42611);
and U44138 (N_44138,N_42845,N_43455);
or U44139 (N_44139,N_43716,N_42603);
and U44140 (N_44140,N_42768,N_42088);
nor U44141 (N_44141,N_42358,N_43649);
and U44142 (N_44142,N_43247,N_43922);
nor U44143 (N_44143,N_43368,N_43143);
xor U44144 (N_44144,N_43415,N_43069);
xnor U44145 (N_44145,N_42726,N_43431);
nand U44146 (N_44146,N_42135,N_42488);
or U44147 (N_44147,N_42085,N_42422);
and U44148 (N_44148,N_42737,N_42610);
nand U44149 (N_44149,N_43734,N_43064);
or U44150 (N_44150,N_42888,N_43859);
or U44151 (N_44151,N_43207,N_42001);
and U44152 (N_44152,N_42373,N_42558);
nand U44153 (N_44153,N_43054,N_42081);
and U44154 (N_44154,N_42644,N_42617);
or U44155 (N_44155,N_43094,N_42292);
or U44156 (N_44156,N_42744,N_43315);
nor U44157 (N_44157,N_42701,N_43319);
nor U44158 (N_44158,N_42407,N_43124);
or U44159 (N_44159,N_42600,N_43944);
nand U44160 (N_44160,N_43866,N_42613);
nor U44161 (N_44161,N_42500,N_42559);
xor U44162 (N_44162,N_42450,N_42328);
xnor U44163 (N_44163,N_43672,N_42858);
and U44164 (N_44164,N_43243,N_42289);
and U44165 (N_44165,N_43078,N_42720);
or U44166 (N_44166,N_43202,N_42997);
xnor U44167 (N_44167,N_43638,N_42666);
xor U44168 (N_44168,N_43458,N_42474);
xnor U44169 (N_44169,N_43799,N_42569);
nor U44170 (N_44170,N_43657,N_42910);
and U44171 (N_44171,N_42570,N_43801);
xor U44172 (N_44172,N_43237,N_42918);
or U44173 (N_44173,N_43508,N_42115);
nor U44174 (N_44174,N_43142,N_42314);
or U44175 (N_44175,N_43290,N_42792);
xor U44176 (N_44176,N_42646,N_42083);
xor U44177 (N_44177,N_42080,N_42752);
or U44178 (N_44178,N_42109,N_43037);
nor U44179 (N_44179,N_43246,N_43863);
nor U44180 (N_44180,N_42908,N_43908);
or U44181 (N_44181,N_42255,N_42593);
nand U44182 (N_44182,N_43378,N_42923);
nor U44183 (N_44183,N_42590,N_42517);
nor U44184 (N_44184,N_42262,N_43192);
nand U44185 (N_44185,N_42712,N_42467);
or U44186 (N_44186,N_42021,N_42998);
or U44187 (N_44187,N_42044,N_42899);
nor U44188 (N_44188,N_43206,N_42973);
or U44189 (N_44189,N_43892,N_42059);
nor U44190 (N_44190,N_43324,N_42544);
or U44191 (N_44191,N_42130,N_43753);
nand U44192 (N_44192,N_42194,N_42148);
nor U44193 (N_44193,N_42581,N_43952);
or U44194 (N_44194,N_42546,N_43891);
xnor U44195 (N_44195,N_42575,N_43275);
nand U44196 (N_44196,N_42632,N_43851);
and U44197 (N_44197,N_43500,N_43188);
nor U44198 (N_44198,N_43418,N_43169);
or U44199 (N_44199,N_43389,N_42635);
and U44200 (N_44200,N_43788,N_42190);
nand U44201 (N_44201,N_42986,N_43402);
nand U44202 (N_44202,N_43758,N_43384);
or U44203 (N_44203,N_42673,N_43137);
nand U44204 (N_44204,N_42731,N_43270);
nor U44205 (N_44205,N_42946,N_42203);
xor U44206 (N_44206,N_42595,N_43079);
or U44207 (N_44207,N_42093,N_42230);
nor U44208 (N_44208,N_43619,N_42038);
or U44209 (N_44209,N_42645,N_42420);
nor U44210 (N_44210,N_42129,N_42608);
or U44211 (N_44211,N_43929,N_42782);
or U44212 (N_44212,N_42822,N_42786);
nor U44213 (N_44213,N_43115,N_42165);
nor U44214 (N_44214,N_43541,N_42064);
or U44215 (N_44215,N_42662,N_42761);
or U44216 (N_44216,N_43374,N_42697);
nor U44217 (N_44217,N_42402,N_42929);
or U44218 (N_44218,N_42876,N_43761);
xor U44219 (N_44219,N_43244,N_43386);
or U44220 (N_44220,N_42372,N_42333);
and U44221 (N_44221,N_42878,N_43164);
xor U44222 (N_44222,N_43191,N_43961);
and U44223 (N_44223,N_42153,N_43817);
nand U44224 (N_44224,N_43477,N_43698);
xor U44225 (N_44225,N_43212,N_42285);
nand U44226 (N_44226,N_43447,N_42394);
nand U44227 (N_44227,N_42449,N_43387);
nor U44228 (N_44228,N_43086,N_43170);
or U44229 (N_44229,N_43639,N_43475);
nor U44230 (N_44230,N_42735,N_42851);
or U44231 (N_44231,N_42312,N_42147);
nor U44232 (N_44232,N_43015,N_42553);
xor U44233 (N_44233,N_42390,N_42506);
or U44234 (N_44234,N_42146,N_43616);
nor U44235 (N_44235,N_43577,N_43990);
xnor U44236 (N_44236,N_42024,N_43152);
xor U44237 (N_44237,N_42301,N_43334);
and U44238 (N_44238,N_43647,N_42084);
or U44239 (N_44239,N_43583,N_42244);
xor U44240 (N_44240,N_42004,N_42917);
or U44241 (N_44241,N_42234,N_42524);
nand U44242 (N_44242,N_43603,N_42927);
or U44243 (N_44243,N_43154,N_42779);
nor U44244 (N_44244,N_43112,N_42648);
or U44245 (N_44245,N_42784,N_43162);
and U44246 (N_44246,N_42948,N_43595);
xnor U44247 (N_44247,N_42007,N_42497);
xnor U44248 (N_44248,N_42193,N_43636);
or U44249 (N_44249,N_42844,N_42905);
and U44250 (N_44250,N_43413,N_42540);
xnor U44251 (N_44251,N_43449,N_42766);
nor U44252 (N_44252,N_43665,N_43762);
nor U44253 (N_44253,N_42945,N_43914);
nand U44254 (N_44254,N_43918,N_43407);
and U44255 (N_44255,N_43128,N_42994);
xor U44256 (N_44256,N_43557,N_42925);
nand U44257 (N_44257,N_42547,N_43253);
and U44258 (N_44258,N_42607,N_42470);
nor U44259 (N_44259,N_42614,N_42346);
or U44260 (N_44260,N_43783,N_42937);
xor U44261 (N_44261,N_43283,N_42363);
xnor U44262 (N_44262,N_42113,N_43401);
nor U44263 (N_44263,N_43678,N_42668);
nand U44264 (N_44264,N_42803,N_42477);
and U44265 (N_44265,N_43361,N_42859);
or U44266 (N_44266,N_42916,N_42638);
nand U44267 (N_44267,N_42043,N_43050);
nor U44268 (N_44268,N_43610,N_42386);
xnor U44269 (N_44269,N_42526,N_42238);
or U44270 (N_44270,N_43752,N_42172);
nand U44271 (N_44271,N_43585,N_42335);
or U44272 (N_44272,N_43175,N_43505);
and U44273 (N_44273,N_43289,N_42368);
or U44274 (N_44274,N_43940,N_43204);
and U44275 (N_44275,N_43403,N_42733);
and U44276 (N_44276,N_42349,N_42119);
or U44277 (N_44277,N_42056,N_43857);
and U44278 (N_44278,N_43232,N_42054);
and U44279 (N_44279,N_43931,N_42252);
nand U44280 (N_44280,N_42826,N_43608);
nor U44281 (N_44281,N_42580,N_42058);
nor U44282 (N_44282,N_43061,N_43751);
xor U44283 (N_44283,N_42724,N_42950);
nor U44284 (N_44284,N_42411,N_42802);
xnor U44285 (N_44285,N_43215,N_43141);
nand U44286 (N_44286,N_42185,N_42417);
nand U44287 (N_44287,N_42445,N_43814);
nor U44288 (N_44288,N_43016,N_42098);
nand U44289 (N_44289,N_43067,N_42655);
nor U44290 (N_44290,N_42209,N_42033);
nand U44291 (N_44291,N_43282,N_42319);
or U44292 (N_44292,N_43703,N_42708);
nand U44293 (N_44293,N_42299,N_43731);
nand U44294 (N_44294,N_42729,N_43058);
nand U44295 (N_44295,N_43456,N_42414);
xor U44296 (N_44296,N_43960,N_42839);
nor U44297 (N_44297,N_42212,N_42819);
and U44298 (N_44298,N_42884,N_43781);
or U44299 (N_44299,N_43875,N_42894);
nand U44300 (N_44300,N_43145,N_43874);
nand U44301 (N_44301,N_42848,N_42985);
nor U44302 (N_44302,N_43005,N_43433);
xnor U44303 (N_44303,N_42483,N_42686);
or U44304 (N_44304,N_43512,N_43298);
xor U44305 (N_44305,N_43994,N_42378);
xnor U44306 (N_44306,N_43320,N_42723);
and U44307 (N_44307,N_43867,N_43065);
nand U44308 (N_44308,N_43840,N_42754);
or U44309 (N_44309,N_42487,N_42079);
xor U44310 (N_44310,N_42073,N_42459);
or U44311 (N_44311,N_42857,N_42482);
and U44312 (N_44312,N_43849,N_43209);
nor U44313 (N_44313,N_42126,N_43059);
and U44314 (N_44314,N_43294,N_43709);
xor U44315 (N_44315,N_42798,N_43177);
nand U44316 (N_44316,N_43261,N_43800);
nand U44317 (N_44317,N_42764,N_43024);
or U44318 (N_44318,N_42305,N_43651);
xor U44319 (N_44319,N_43032,N_42187);
nor U44320 (N_44320,N_42895,N_43216);
or U44321 (N_44321,N_42790,N_42075);
xor U44322 (N_44322,N_42242,N_43028);
and U44323 (N_44323,N_43652,N_43114);
or U44324 (N_44324,N_43895,N_42365);
nand U44325 (N_44325,N_42659,N_42624);
nor U44326 (N_44326,N_42072,N_42495);
nand U44327 (N_44327,N_42743,N_43076);
nor U44328 (N_44328,N_42154,N_43642);
nand U44329 (N_44329,N_43196,N_43920);
or U44330 (N_44330,N_42337,N_42571);
and U44331 (N_44331,N_42114,N_43968);
or U44332 (N_44332,N_43868,N_43889);
xor U44333 (N_44333,N_43673,N_43101);
xnor U44334 (N_44334,N_43038,N_42436);
and U44335 (N_44335,N_43306,N_43880);
xnor U44336 (N_44336,N_42807,N_43970);
and U44337 (N_44337,N_43347,N_43075);
and U44338 (N_44338,N_43325,N_42280);
nor U44339 (N_44339,N_43591,N_42818);
and U44340 (N_44340,N_42216,N_42862);
nand U44341 (N_44341,N_43372,N_43313);
nand U44342 (N_44342,N_42248,N_42281);
xor U44343 (N_44343,N_42713,N_43487);
nand U44344 (N_44344,N_43602,N_43000);
xnor U44345 (N_44345,N_43576,N_42377);
or U44346 (N_44346,N_43474,N_42229);
or U44347 (N_44347,N_42279,N_42621);
or U44348 (N_44348,N_43553,N_42220);
nand U44349 (N_44349,N_43269,N_42788);
nand U44350 (N_44350,N_42828,N_43072);
xor U44351 (N_44351,N_42965,N_43293);
or U44352 (N_44352,N_42406,N_42275);
nor U44353 (N_44353,N_43327,N_43018);
xnor U44354 (N_44354,N_43424,N_42618);
nor U44355 (N_44355,N_42881,N_43138);
xor U44356 (N_44356,N_42040,N_43262);
nor U44357 (N_44357,N_42016,N_43496);
or U44358 (N_44358,N_43025,N_43251);
nand U44359 (N_44359,N_42589,N_43967);
and U44360 (N_44360,N_43766,N_43331);
or U44361 (N_44361,N_42022,N_42582);
and U44362 (N_44362,N_42308,N_42074);
or U44363 (N_44363,N_42814,N_42893);
or U44364 (N_44364,N_42237,N_42205);
and U44365 (N_44365,N_42222,N_43443);
xnor U44366 (N_44366,N_42327,N_43287);
nor U44367 (N_44367,N_43732,N_43634);
and U44368 (N_44368,N_43625,N_43841);
nand U44369 (N_44369,N_42170,N_43157);
nor U44370 (N_44370,N_42940,N_42840);
xor U44371 (N_44371,N_42435,N_42959);
or U44372 (N_44372,N_43692,N_42560);
xnor U44373 (N_44373,N_43071,N_43947);
and U44374 (N_44374,N_42800,N_42805);
and U44375 (N_44375,N_42011,N_43238);
or U44376 (N_44376,N_42543,N_42124);
xnor U44377 (N_44377,N_42431,N_43343);
or U44378 (N_44378,N_43821,N_43108);
nand U44379 (N_44379,N_43661,N_43684);
or U44380 (N_44380,N_42993,N_42682);
nand U44381 (N_44381,N_43943,N_43997);
nor U44382 (N_44382,N_42046,N_42443);
nand U44383 (N_44383,N_43004,N_43184);
and U44384 (N_44384,N_42849,N_43862);
and U44385 (N_44385,N_43013,N_43575);
xor U44386 (N_44386,N_42442,N_43160);
nor U44387 (N_44387,N_42503,N_43836);
and U44388 (N_44388,N_42453,N_42750);
or U44389 (N_44389,N_42599,N_43877);
or U44390 (N_44390,N_43795,N_43664);
or U44391 (N_44391,N_42999,N_43563);
and U44392 (N_44392,N_42020,N_42323);
and U44393 (N_44393,N_43530,N_42128);
nand U44394 (N_44394,N_43146,N_42441);
nand U44395 (N_44395,N_42465,N_42834);
nand U44396 (N_44396,N_43687,N_42112);
and U44397 (N_44397,N_42772,N_42433);
and U44398 (N_44398,N_42954,N_43539);
nand U44399 (N_44399,N_43459,N_43771);
and U44400 (N_44400,N_42935,N_43686);
or U44401 (N_44401,N_43236,N_43740);
nand U44402 (N_44402,N_43257,N_43631);
nand U44403 (N_44403,N_43643,N_43827);
xor U44404 (N_44404,N_43792,N_43121);
and U44405 (N_44405,N_43521,N_43632);
or U44406 (N_44406,N_42552,N_43176);
or U44407 (N_44407,N_42169,N_42756);
xor U44408 (N_44408,N_43364,N_42271);
and U44409 (N_44409,N_43562,N_42972);
and U44410 (N_44410,N_42374,N_43345);
nand U44411 (N_44411,N_43586,N_42002);
or U44412 (N_44412,N_42423,N_42239);
and U44413 (N_44413,N_42132,N_43648);
nand U44414 (N_44414,N_42392,N_43581);
nand U44415 (N_44415,N_42535,N_42097);
nor U44416 (N_44416,N_43936,N_43670);
or U44417 (N_44417,N_42099,N_43520);
or U44418 (N_44418,N_43010,N_42631);
nand U44419 (N_44419,N_42180,N_42871);
nor U44420 (N_44420,N_42951,N_43339);
xor U44421 (N_44421,N_43436,N_42371);
or U44422 (N_44422,N_43566,N_42000);
xnor U44423 (N_44423,N_43173,N_42177);
nand U44424 (N_44424,N_43118,N_43470);
or U44425 (N_44425,N_42149,N_42957);
and U44426 (N_44426,N_42588,N_42577);
and U44427 (N_44427,N_42429,N_42780);
nand U44428 (N_44428,N_43946,N_43178);
or U44429 (N_44429,N_43199,N_43464);
xnor U44430 (N_44430,N_43116,N_43939);
and U44431 (N_44431,N_43839,N_43958);
nor U44432 (N_44432,N_42091,N_43653);
nand U44433 (N_44433,N_43316,N_42685);
xnor U44434 (N_44434,N_43150,N_42838);
xnor U44435 (N_44435,N_42316,N_43461);
or U44436 (N_44436,N_42410,N_43400);
nand U44437 (N_44437,N_42911,N_42711);
and U44438 (N_44438,N_43346,N_42984);
or U44439 (N_44439,N_42376,N_43002);
and U44440 (N_44440,N_42507,N_43996);
xnor U44441 (N_44441,N_42721,N_43739);
and U44442 (N_44442,N_43524,N_42136);
and U44443 (N_44443,N_42650,N_42042);
or U44444 (N_44444,N_43856,N_43008);
nor U44445 (N_44445,N_42747,N_42360);
xnor U44446 (N_44446,N_42329,N_42887);
or U44447 (N_44447,N_43301,N_42783);
and U44448 (N_44448,N_43425,N_42705);
or U44449 (N_44449,N_43646,N_42739);
or U44450 (N_44450,N_42869,N_42105);
nand U44451 (N_44451,N_42027,N_42594);
nand U44452 (N_44452,N_42354,N_43637);
or U44453 (N_44453,N_43971,N_42412);
or U44454 (N_44454,N_42257,N_42245);
or U44455 (N_44455,N_43310,N_43240);
or U44456 (N_44456,N_43564,N_43308);
xor U44457 (N_44457,N_43229,N_42241);
nand U44458 (N_44458,N_42479,N_43323);
nor U44459 (N_44459,N_42472,N_43992);
xnor U44460 (N_44460,N_43802,N_43161);
or U44461 (N_44461,N_43884,N_42642);
nand U44462 (N_44462,N_43810,N_43926);
or U44463 (N_44463,N_43778,N_42942);
nand U44464 (N_44464,N_43446,N_43782);
or U44465 (N_44465,N_43953,N_42478);
xnor U44466 (N_44466,N_42107,N_42649);
nand U44467 (N_44467,N_43549,N_43039);
xnor U44468 (N_44468,N_42519,N_42359);
or U44469 (N_44469,N_42639,N_43451);
or U44470 (N_44470,N_43963,N_43699);
nor U44471 (N_44471,N_43969,N_43536);
and U44472 (N_44472,N_42566,N_42415);
nand U44473 (N_44473,N_43544,N_42227);
nand U44474 (N_44474,N_43180,N_43853);
xor U44475 (N_44475,N_42513,N_43683);
nor U44476 (N_44476,N_43182,N_42510);
nor U44477 (N_44477,N_42320,N_42003);
xnor U44478 (N_44478,N_42740,N_43427);
nor U44479 (N_44479,N_43878,N_42061);
or U44480 (N_44480,N_42484,N_43909);
xnor U44481 (N_44481,N_42466,N_42585);
xor U44482 (N_44482,N_42041,N_43630);
xnor U44483 (N_44483,N_43406,N_43421);
or U44484 (N_44484,N_42164,N_43453);
nor U44485 (N_44485,N_43340,N_43080);
and U44486 (N_44486,N_42336,N_42231);
nor U44487 (N_44487,N_42841,N_42157);
or U44488 (N_44488,N_42898,N_43304);
nor U44489 (N_44489,N_43399,N_42738);
nand U44490 (N_44490,N_43813,N_43535);
nor U44491 (N_44491,N_43975,N_42679);
or U44492 (N_44492,N_42342,N_43045);
and U44493 (N_44493,N_43561,N_42537);
xor U44494 (N_44494,N_43088,N_43869);
nand U44495 (N_44495,N_42439,N_43842);
nand U44496 (N_44496,N_42604,N_42270);
nand U44497 (N_44497,N_43412,N_42630);
and U44498 (N_44498,N_42196,N_42932);
nand U44499 (N_44499,N_42949,N_42530);
or U44500 (N_44500,N_43558,N_42078);
or U44501 (N_44501,N_43483,N_42127);
or U44502 (N_44502,N_42055,N_42471);
and U44503 (N_44503,N_42602,N_42902);
xnor U44504 (N_44504,N_43597,N_43104);
and U44505 (N_44505,N_43255,N_43713);
and U44506 (N_44506,N_42514,N_42214);
or U44507 (N_44507,N_42432,N_42176);
and U44508 (N_44508,N_42627,N_42077);
and U44509 (N_44509,N_43093,N_43838);
nor U44510 (N_44510,N_43765,N_43794);
or U44511 (N_44511,N_43671,N_43362);
nor U44512 (N_44512,N_42689,N_42086);
or U44513 (N_44513,N_42527,N_43266);
and U44514 (N_44514,N_42964,N_42794);
or U44515 (N_44515,N_42634,N_43972);
xnor U44516 (N_44516,N_43942,N_42647);
xnor U44517 (N_44517,N_43482,N_43166);
nor U44518 (N_44518,N_43336,N_42226);
nor U44519 (N_44519,N_42936,N_42695);
nor U44520 (N_44520,N_42824,N_43174);
nand U44521 (N_44521,N_42551,N_43956);
or U44522 (N_44522,N_43654,N_42492);
xnor U44523 (N_44523,N_43624,N_43501);
and U44524 (N_44524,N_42440,N_42926);
xnor U44525 (N_44525,N_43302,N_42017);
and U44526 (N_44526,N_42026,N_42508);
or U44527 (N_44527,N_43134,N_43034);
xor U44528 (N_44528,N_43830,N_42504);
and U44529 (N_44529,N_42904,N_43949);
nand U44530 (N_44530,N_43998,N_43991);
xnor U44531 (N_44531,N_42746,N_42829);
xor U44532 (N_44532,N_42704,N_43770);
or U44533 (N_44533,N_43886,N_43745);
xor U44534 (N_44534,N_42347,N_43627);
xnor U44535 (N_44535,N_43662,N_43264);
or U44536 (N_44536,N_43396,N_42025);
nor U44537 (N_44537,N_42868,N_43201);
xor U44538 (N_44538,N_42717,N_43186);
or U44539 (N_44539,N_43733,N_43084);
or U44540 (N_44540,N_42702,N_43882);
nand U44541 (N_44541,N_42369,N_43438);
or U44542 (N_44542,N_42298,N_43806);
nor U44543 (N_44543,N_43132,N_42676);
or U44544 (N_44544,N_42511,N_43021);
or U44545 (N_44545,N_43516,N_43254);
xnor U44546 (N_44546,N_43620,N_43567);
xor U44547 (N_44547,N_43515,N_43633);
nand U44548 (N_44548,N_42789,N_42762);
or U44549 (N_44549,N_42616,N_43213);
xor U44550 (N_44550,N_43507,N_43123);
nor U44551 (N_44551,N_42554,N_42864);
nor U44552 (N_44552,N_43358,N_42277);
nor U44553 (N_44553,N_42162,N_43897);
nand U44554 (N_44554,N_43395,N_42350);
xor U44555 (N_44555,N_43312,N_43522);
nand U44556 (N_44556,N_43278,N_42974);
or U44557 (N_44557,N_42550,N_43193);
nor U44558 (N_44558,N_42643,N_42063);
and U44559 (N_44559,N_43450,N_43604);
xor U44560 (N_44560,N_43214,N_43168);
nand U44561 (N_44561,N_42757,N_43448);
xnor U44562 (N_44562,N_43718,N_43349);
and U44563 (N_44563,N_43973,N_43106);
and U44564 (N_44564,N_43326,N_43641);
nor U44565 (N_44565,N_42977,N_43550);
and U44566 (N_44566,N_42438,N_43573);
nand U44567 (N_44567,N_42123,N_42145);
nor U44568 (N_44568,N_43518,N_42300);
nor U44569 (N_44569,N_42140,N_43452);
nand U44570 (N_44570,N_42455,N_42591);
nor U44571 (N_44571,N_42243,N_43749);
nor U44572 (N_44572,N_42232,N_43951);
and U44573 (N_44573,N_43832,N_42491);
nand U44574 (N_44574,N_42870,N_43398);
xor U44575 (N_44575,N_43463,N_43476);
and U44576 (N_44576,N_43728,N_43663);
or U44577 (N_44577,N_43218,N_43824);
or U44578 (N_44578,N_42221,N_42633);
or U44579 (N_44579,N_42090,N_43383);
nand U44580 (N_44580,N_43881,N_42907);
nand U44581 (N_44581,N_42515,N_42843);
or U44582 (N_44582,N_42652,N_43147);
nand U44583 (N_44583,N_42311,N_43677);
and U44584 (N_44584,N_43815,N_42256);
nand U44585 (N_44585,N_42391,N_42076);
nor U44586 (N_44586,N_43819,N_42096);
or U44587 (N_44587,N_43375,N_43200);
nor U44588 (N_44588,N_43435,N_43587);
and U44589 (N_44589,N_42691,N_42446);
nor U44590 (N_44590,N_42192,N_42028);
nand U44591 (N_44591,N_42736,N_42557);
and U44592 (N_44592,N_43714,N_43621);
nand U44593 (N_44593,N_42875,N_43538);
xnor U44594 (N_44594,N_43905,N_43685);
and U44595 (N_44595,N_42053,N_42403);
or U44596 (N_44596,N_43333,N_43747);
and U44597 (N_44597,N_43760,N_42938);
and U44598 (N_44598,N_43466,N_43082);
and U44599 (N_44599,N_43462,N_43036);
nand U44600 (N_44600,N_42727,N_42121);
and U44601 (N_44601,N_42493,N_43429);
nor U44602 (N_44602,N_42623,N_43529);
or U44603 (N_44603,N_43493,N_42409);
nand U44604 (N_44604,N_42675,N_42151);
or U44605 (N_44605,N_43777,N_42161);
xnor U44606 (N_44606,N_43183,N_43357);
nand U44607 (N_44607,N_43408,N_42882);
and U44608 (N_44608,N_43710,N_42393);
or U44609 (N_44609,N_43224,N_43210);
nand U44610 (N_44610,N_43414,N_42572);
or U44611 (N_44611,N_42413,N_43893);
nor U44612 (N_44612,N_42035,N_42259);
nand U44613 (N_44613,N_43285,N_43171);
nand U44614 (N_44614,N_43031,N_42690);
xnor U44615 (N_44615,N_43056,N_43317);
or U44616 (N_44616,N_43272,N_43485);
or U44617 (N_44617,N_43367,N_43125);
nand U44618 (N_44618,N_43495,N_43221);
or U44619 (N_44619,N_42719,N_43548);
or U44620 (N_44620,N_43784,N_42785);
nor U44621 (N_44621,N_43776,N_42383);
nand U44622 (N_44622,N_43618,N_43126);
or U44623 (N_44623,N_42251,N_43769);
and U44624 (N_44624,N_43717,N_43682);
xor U44625 (N_44625,N_42134,N_43774);
xnor U44626 (N_44626,N_43796,N_42464);
or U44627 (N_44627,N_42223,N_43292);
and U44628 (N_44628,N_42131,N_43706);
or U44629 (N_44629,N_42208,N_42573);
or U44630 (N_44630,N_43729,N_42218);
and U44631 (N_44631,N_43767,N_42806);
nor U44632 (N_44632,N_43592,N_42102);
xnor U44633 (N_44633,N_43484,N_43130);
or U44634 (N_44634,N_43030,N_43260);
nand U44635 (N_44635,N_42352,N_42009);
or U44636 (N_44636,N_43195,N_43363);
xor U44637 (N_44637,N_43365,N_43601);
nor U44638 (N_44638,N_42264,N_43371);
or U44639 (N_44639,N_43502,N_43910);
nor U44640 (N_44640,N_43923,N_43379);
and U44641 (N_44641,N_42670,N_43883);
nor U44642 (N_44642,N_43514,N_43309);
nor U44643 (N_44643,N_43578,N_43074);
nand U44644 (N_44644,N_42776,N_42071);
and U44645 (N_44645,N_42832,N_42331);
nand U44646 (N_44646,N_43828,N_42728);
and U44647 (N_44647,N_43829,N_42458);
or U44648 (N_44648,N_42397,N_42533);
nor U44649 (N_44649,N_42430,N_42751);
or U44650 (N_44650,N_42047,N_42781);
xnor U44651 (N_44651,N_42837,N_43003);
and U44652 (N_44652,N_43393,N_42357);
xor U44653 (N_44653,N_43478,N_42677);
or U44654 (N_44654,N_43099,N_43593);
xnor U44655 (N_44655,N_42883,N_42775);
xor U44656 (N_44656,N_42191,N_42778);
nor U44657 (N_44657,N_42317,N_42156);
nand U44658 (N_44658,N_43369,N_43650);
or U44659 (N_44659,N_43808,N_43668);
nand U44660 (N_44660,N_43499,N_43419);
xnor U44661 (N_44661,N_42057,N_43917);
or U44662 (N_44662,N_42971,N_42263);
xnor U44663 (N_44663,N_43303,N_43007);
xor U44664 (N_44664,N_43263,N_43680);
nand U44665 (N_44665,N_43720,N_42693);
and U44666 (N_44666,N_42835,N_43140);
and U44667 (N_44667,N_43722,N_42454);
and U44668 (N_44668,N_42339,N_43227);
and U44669 (N_44669,N_42315,N_42641);
nor U44670 (N_44670,N_43833,N_42619);
nor U44671 (N_44671,N_42167,N_43228);
xnor U44672 (N_44672,N_43023,N_43727);
or U44673 (N_44673,N_42195,N_43197);
nor U44674 (N_44674,N_42344,N_42749);
or U44675 (N_44675,N_43773,N_42579);
nor U44676 (N_44676,N_42601,N_42759);
or U44677 (N_44677,N_42008,N_43131);
and U44678 (N_44678,N_42830,N_43077);
xnor U44679 (N_44679,N_42240,N_43721);
xor U44680 (N_44680,N_43705,N_42725);
and U44681 (N_44681,N_43139,N_43391);
nor U44682 (N_44682,N_42774,N_42922);
and U44683 (N_44683,N_43165,N_42168);
nor U44684 (N_44684,N_42900,N_43085);
nand U44685 (N_44685,N_42178,N_42542);
nor U44686 (N_44686,N_42106,N_43534);
and U44687 (N_44687,N_42626,N_43725);
nor U44688 (N_44688,N_42291,N_42225);
and U44689 (N_44689,N_43525,N_42235);
or U44690 (N_44690,N_42034,N_42295);
xnor U44691 (N_44691,N_42817,N_43554);
nor U44692 (N_44692,N_42448,N_43234);
nor U44693 (N_44693,N_43469,N_43081);
xor U44694 (N_44694,N_43113,N_43764);
nand U44695 (N_44695,N_43019,N_42116);
or U44696 (N_44696,N_42023,N_42353);
or U44697 (N_44697,N_43252,N_42658);
or U44698 (N_44698,N_42427,N_42903);
nand U44699 (N_44699,N_42293,N_43988);
xnor U44700 (N_44700,N_42815,N_42269);
or U44701 (N_44701,N_43480,N_42987);
or U44702 (N_44702,N_43156,N_42667);
and U44703 (N_44703,N_42866,N_42555);
xor U44704 (N_44704,N_42549,N_43690);
nor U44705 (N_44705,N_43540,N_43904);
or U44706 (N_44706,N_43219,N_42598);
nor U44707 (N_44707,N_43122,N_42801);
and U44708 (N_44708,N_43644,N_43280);
and U44709 (N_44709,N_43423,N_42674);
nor U44710 (N_44710,N_42521,N_42816);
nor U44711 (N_44711,N_43744,N_43927);
xor U44712 (N_44712,N_43388,N_42142);
xnor U44713 (N_44713,N_42100,N_43506);
nor U44714 (N_44714,N_42889,N_43259);
and U44715 (N_44715,N_43719,N_43811);
nor U44716 (N_44716,N_42825,N_42408);
nor U44717 (N_44717,N_43437,N_42605);
nor U44718 (N_44718,N_42567,N_43376);
and U44719 (N_44719,N_43763,N_42861);
nor U44720 (N_44720,N_43097,N_42108);
nor U44721 (N_44721,N_43755,N_43812);
nand U44722 (N_44722,N_43479,N_42388);
and U44723 (N_44723,N_42718,N_42541);
xor U44724 (N_44724,N_42586,N_43925);
xnor U44725 (N_44725,N_42171,N_43858);
nor U44726 (N_44726,N_43102,N_43341);
nand U44727 (N_44727,N_43250,N_42672);
and U44728 (N_44728,N_42584,N_42874);
xnor U44729 (N_44729,N_42062,N_42795);
xor U44730 (N_44730,N_43144,N_43660);
and U44731 (N_44731,N_42653,N_43552);
xnor U44732 (N_44732,N_43281,N_43352);
nand U44733 (N_44733,N_43100,N_43772);
and U44734 (N_44734,N_42609,N_42664);
or U44735 (N_44735,N_42943,N_43098);
or U44736 (N_44736,N_43825,N_43020);
nor U44737 (N_44737,N_43605,N_43276);
xor U44738 (N_44738,N_43861,N_42224);
nor U44739 (N_44739,N_42958,N_43504);
nand U44740 (N_44740,N_43119,N_42846);
and U44741 (N_44741,N_42769,N_43979);
or U44742 (N_44742,N_42629,N_42092);
or U44743 (N_44743,N_43787,N_42745);
nor U44744 (N_44744,N_43876,N_43052);
xor U44745 (N_44745,N_43190,N_43899);
nand U44746 (N_44746,N_43993,N_42821);
or U44747 (N_44747,N_43711,N_42952);
and U44748 (N_44748,N_42330,N_43850);
nor U44749 (N_44749,N_43959,N_42996);
nor U44750 (N_44750,N_43404,N_42010);
nand U44751 (N_44751,N_42118,N_42181);
or U44752 (N_44752,N_42274,N_42561);
nand U44753 (N_44753,N_42260,N_43329);
nor U44754 (N_44754,N_42612,N_42914);
nor U44755 (N_44755,N_42694,N_42361);
nor U44756 (N_44756,N_43256,N_43962);
nor U44757 (N_44757,N_42651,N_43852);
nand U44758 (N_44758,N_43105,N_42110);
xnor U44759 (N_44759,N_43360,N_43584);
nand U44760 (N_44760,N_43517,N_42981);
nand U44761 (N_44761,N_42030,N_43894);
and U44762 (N_44762,N_43277,N_43885);
nand U44763 (N_44763,N_43053,N_43211);
nor U44764 (N_44764,N_42787,N_43040);
and U44765 (N_44765,N_43513,N_43865);
xor U44766 (N_44766,N_42031,N_43757);
or U44767 (N_44767,N_42452,N_42029);
xnor U44768 (N_44768,N_42976,N_42700);
nor U44769 (N_44769,N_43497,N_43117);
or U44770 (N_44770,N_42150,N_42276);
nand U44771 (N_44771,N_42400,N_43695);
xnor U44772 (N_44772,N_43432,N_43981);
xor U44773 (N_44773,N_42763,N_42249);
nand U44774 (N_44774,N_43912,N_43033);
nor U44775 (N_44775,N_42144,N_43977);
and U44776 (N_44776,N_42529,N_43233);
or U44777 (N_44777,N_43688,N_43674);
or U44778 (N_44778,N_43527,N_43954);
and U44779 (N_44779,N_43528,N_43629);
or U44780 (N_44780,N_42032,N_43533);
nand U44781 (N_44781,N_42919,N_43932);
and U44782 (N_44782,N_43847,N_42356);
nand U44783 (N_44783,N_42405,N_43985);
nand U44784 (N_44784,N_43580,N_43344);
nor U44785 (N_44785,N_43579,N_42272);
nand U44786 (N_44786,N_42419,N_42345);
or U44787 (N_44787,N_43696,N_42069);
nor U44788 (N_44788,N_43440,N_43906);
xnor U44789 (N_44789,N_42597,N_42399);
and U44790 (N_44790,N_43789,N_43494);
or U44791 (N_44791,N_42219,N_43697);
xnor U44792 (N_44792,N_42213,N_43373);
and U44793 (N_44793,N_42095,N_43945);
or U44794 (N_44794,N_42173,N_42236);
or U44795 (N_44795,N_42912,N_43701);
nor U44796 (N_44796,N_42706,N_42186);
xor U44797 (N_44797,N_42703,N_43047);
or U44798 (N_44798,N_43394,N_42777);
nand U44799 (N_44799,N_42065,N_42155);
nand U44800 (N_44800,N_42850,N_42182);
xnor U44801 (N_44801,N_43265,N_43307);
or U44802 (N_44802,N_42628,N_42791);
nand U44803 (N_44803,N_43153,N_43006);
xor U44804 (N_44804,N_42852,N_43743);
and U44805 (N_44805,N_42473,N_43305);
xnor U44806 (N_44806,N_43348,N_43135);
nor U44807 (N_44807,N_42809,N_43198);
and U44808 (N_44808,N_42428,N_42699);
or U44809 (N_44809,N_43258,N_42885);
and U44810 (N_44810,N_43055,N_43888);
or U44811 (N_44811,N_43707,N_42367);
nor U44812 (N_44812,N_42520,N_43689);
or U44813 (N_44813,N_42375,N_43913);
or U44814 (N_44814,N_42288,N_43921);
and U44815 (N_44815,N_42793,N_42578);
xnor U44816 (N_44816,N_43775,N_43311);
nor U44817 (N_44817,N_43380,N_43655);
nor U44818 (N_44818,N_42532,N_42808);
nor U44819 (N_44819,N_43239,N_42362);
xnor U44820 (N_44820,N_42678,N_43823);
or U44821 (N_44821,N_43582,N_43822);
nor U44822 (N_44822,N_43569,N_42266);
and U44823 (N_44823,N_43556,N_42556);
nor U44824 (N_44824,N_43746,N_43890);
and U44825 (N_44825,N_43491,N_43136);
nor U44826 (N_44826,N_43614,N_42014);
nand U44827 (N_44827,N_42982,N_43872);
nor U44828 (N_44828,N_43127,N_43172);
nor U44829 (N_44829,N_43299,N_42447);
nand U44830 (N_44830,N_42568,N_43543);
and U44831 (N_44831,N_42174,N_43750);
nand U44832 (N_44832,N_42143,N_43983);
nand U44833 (N_44833,N_42204,N_43163);
or U44834 (N_44834,N_42321,N_42742);
nor U44835 (N_44835,N_43286,N_43245);
nand U44836 (N_44836,N_42640,N_42966);
nand U44837 (N_44837,N_43231,N_42842);
nor U44838 (N_44838,N_43295,N_43472);
nand U44839 (N_44839,N_43066,N_42163);
and U44840 (N_44840,N_43658,N_42215);
nand U44841 (N_44841,N_42804,N_42810);
or U44842 (N_44842,N_43742,N_43980);
nand U44843 (N_44843,N_42995,N_43754);
or U44844 (N_44844,N_43843,N_43803);
nand U44845 (N_44845,N_42992,N_42425);
nand U44846 (N_44846,N_42395,N_43428);
and U44847 (N_44847,N_43797,N_43786);
or U44848 (N_44848,N_43274,N_42606);
nor U44849 (N_44849,N_43044,N_42434);
or U44850 (N_44850,N_42382,N_43444);
xor U44851 (N_44851,N_43617,N_42955);
and U44852 (N_44852,N_42896,N_42302);
and U44853 (N_44853,N_42364,N_42827);
xnor U44854 (N_44854,N_43559,N_43873);
or U44855 (N_44855,N_43600,N_42636);
and U44856 (N_44856,N_43551,N_43611);
nand U44857 (N_44857,N_43978,N_43738);
nand U44858 (N_44858,N_43167,N_42687);
nor U44859 (N_44859,N_42531,N_43109);
xor U44860 (N_44860,N_42324,N_42211);
nand U44861 (N_44861,N_42671,N_43915);
nor U44862 (N_44862,N_42853,N_43107);
or U44863 (N_44863,N_43322,N_43855);
and U44864 (N_44864,N_43043,N_43737);
nor U44865 (N_44865,N_43948,N_43490);
nand U44866 (N_44866,N_43835,N_42404);
or U44867 (N_44867,N_42799,N_43986);
nand U44868 (N_44868,N_43022,N_43831);
xnor U44869 (N_44869,N_43223,N_42013);
xnor U44870 (N_44870,N_42039,N_42313);
nand U44871 (N_44871,N_43090,N_43957);
xor U44872 (N_44872,N_42384,N_42282);
nor U44873 (N_44873,N_42498,N_43046);
and U44874 (N_44874,N_43471,N_43901);
or U44875 (N_44875,N_42538,N_42563);
nor U44876 (N_44876,N_43068,N_42622);
nor U44877 (N_44877,N_43103,N_43702);
or U44878 (N_44878,N_42501,N_42765);
nand U44879 (N_44879,N_43087,N_42620);
nor U44880 (N_44880,N_42909,N_43571);
xnor U44881 (N_44881,N_42179,N_43511);
nand U44882 (N_44882,N_43666,N_42901);
nand U44883 (N_44883,N_43382,N_43460);
or U44884 (N_44884,N_43151,N_42688);
or U44885 (N_44885,N_43042,N_42625);
and U44886 (N_44886,N_43017,N_43804);
xor U44887 (N_44887,N_43995,N_43679);
xnor U44888 (N_44888,N_42890,N_43273);
xnor U44889 (N_44889,N_43189,N_43805);
nand U44890 (N_44890,N_43366,N_43041);
or U44891 (N_44891,N_43217,N_43284);
or U44892 (N_44892,N_43704,N_43712);
nand U44893 (N_44893,N_43640,N_43606);
nor U44894 (N_44894,N_42692,N_42297);
nor U44895 (N_44895,N_42166,N_42351);
nand U44896 (N_44896,N_42462,N_43248);
xor U44897 (N_44897,N_42424,N_42355);
nand U44898 (N_44898,N_43871,N_42880);
and U44899 (N_44899,N_42082,N_43503);
and U44900 (N_44900,N_42104,N_42444);
and U44901 (N_44901,N_43332,N_42012);
nor U44902 (N_44902,N_42847,N_43934);
xor U44903 (N_44903,N_42045,N_42122);
nor U44904 (N_44904,N_42915,N_42117);
nor U44905 (N_44905,N_42539,N_42006);
nand U44906 (N_44906,N_43014,N_43048);
nand U44907 (N_44907,N_42962,N_42534);
and U44908 (N_44908,N_42576,N_42980);
or U44909 (N_44909,N_43930,N_42389);
xnor U44910 (N_44910,N_43027,N_42592);
nand U44911 (N_44911,N_43826,N_43691);
nand U44912 (N_44912,N_43314,N_43489);
and U44913 (N_44913,N_42615,N_43271);
or U44914 (N_44914,N_43279,N_43756);
nor U44915 (N_44915,N_42070,N_42991);
or U44916 (N_44916,N_42152,N_42924);
xor U44917 (N_44917,N_43785,N_43669);
xnor U44918 (N_44918,N_43185,N_42587);
nor U44919 (N_44919,N_43351,N_42865);
and U44920 (N_44920,N_43035,N_43846);
and U44921 (N_44921,N_43439,N_43547);
nor U44922 (N_44922,N_43420,N_43441);
nand U44923 (N_44923,N_43377,N_43907);
or U44924 (N_44924,N_42928,N_43568);
nor U44925 (N_44925,N_42340,N_43430);
nand U44926 (N_44926,N_42707,N_42197);
xnor U44927 (N_44927,N_43337,N_42730);
xnor U44928 (N_44928,N_43111,N_43572);
and U44929 (N_44929,N_42562,N_42175);
or U44930 (N_44930,N_43626,N_43133);
and U44931 (N_44931,N_42217,N_43964);
nor U44932 (N_44932,N_42565,N_42767);
nor U44933 (N_44933,N_42284,N_43759);
and U44934 (N_44934,N_42934,N_42656);
and U44935 (N_44935,N_42138,N_42334);
nand U44936 (N_44936,N_42426,N_43613);
or U44937 (N_44937,N_43537,N_42158);
xnor U44938 (N_44938,N_43486,N_42457);
and U44939 (N_44939,N_42201,N_43935);
and U44940 (N_44940,N_42469,N_42278);
nand U44941 (N_44941,N_42518,N_42202);
nand U44942 (N_44942,N_42379,N_42696);
nor U44943 (N_44943,N_43267,N_43338);
nor U44944 (N_44944,N_42050,N_43999);
or U44945 (N_44945,N_42310,N_42018);
and U44946 (N_44946,N_42637,N_43599);
or U44947 (N_44947,N_42892,N_42811);
or U44948 (N_44948,N_42489,N_43791);
nand U44949 (N_44949,N_42660,N_43049);
nand U44950 (N_44950,N_43226,N_43012);
and U44951 (N_44951,N_42941,N_43816);
and U44952 (N_44952,N_42960,N_42944);
or U44953 (N_44953,N_43060,N_42137);
nand U44954 (N_44954,N_43837,N_43860);
and U44955 (N_44955,N_43965,N_43588);
xor U44956 (N_44956,N_42111,N_43029);
nand U44957 (N_44957,N_42886,N_43467);
and U44958 (N_44958,N_42005,N_43955);
nand U44959 (N_44959,N_42921,N_42261);
xnor U44960 (N_44960,N_43937,N_42318);
and U44961 (N_44961,N_42160,N_42968);
nand U44962 (N_44962,N_43194,N_42931);
nor U44963 (N_44963,N_43848,N_42253);
and U44964 (N_44964,N_43736,N_43987);
nor U44965 (N_44965,N_43887,N_43225);
and U44966 (N_44966,N_43911,N_42983);
nand U44967 (N_44967,N_42753,N_42326);
and U44968 (N_44968,N_43546,N_43242);
xor U44969 (N_44969,N_42661,N_42813);
nor U44970 (N_44970,N_43748,N_42385);
nor U44971 (N_44971,N_43089,N_42247);
nor U44972 (N_44972,N_42860,N_43203);
and U44973 (N_44973,N_43594,N_43342);
nand U44974 (N_44974,N_43938,N_42496);
and U44975 (N_44975,N_42304,N_42307);
or U44976 (N_44976,N_42089,N_43181);
xnor U44977 (N_44977,N_42370,N_42052);
and U44978 (N_44978,N_42709,N_42970);
and U44979 (N_44979,N_42485,N_42872);
nand U44980 (N_44980,N_43120,N_42512);
and U44981 (N_44981,N_43984,N_42103);
or U44982 (N_44982,N_42398,N_43091);
and U44983 (N_44983,N_43982,N_43063);
nand U44984 (N_44984,N_42961,N_42015);
nor U44985 (N_44985,N_43397,N_43385);
nor U44986 (N_44986,N_43159,N_43864);
nor U44987 (N_44987,N_42836,N_43693);
nand U44988 (N_44988,N_42309,N_43798);
or U44989 (N_44989,N_43001,N_42855);
or U44990 (N_44990,N_43318,N_43715);
nor U44991 (N_44991,N_42863,N_42773);
or U44992 (N_44992,N_43220,N_43845);
or U44993 (N_44993,N_43590,N_42698);
and U44994 (N_44994,N_43598,N_42463);
or U44995 (N_44995,N_42741,N_42184);
nor U44996 (N_44996,N_43129,N_42210);
nand U44997 (N_44997,N_43902,N_42502);
or U44998 (N_44998,N_43417,N_43390);
nand U44999 (N_44999,N_42681,N_43073);
nor U45000 (N_45000,N_42106,N_42540);
xnor U45001 (N_45001,N_43158,N_42545);
or U45002 (N_45002,N_42670,N_42383);
nand U45003 (N_45003,N_42734,N_42820);
nor U45004 (N_45004,N_43832,N_43013);
and U45005 (N_45005,N_43652,N_42593);
and U45006 (N_45006,N_43919,N_43798);
nor U45007 (N_45007,N_42305,N_42898);
nor U45008 (N_45008,N_43264,N_43046);
nand U45009 (N_45009,N_43449,N_42426);
xor U45010 (N_45010,N_42254,N_43537);
nand U45011 (N_45011,N_43021,N_42199);
and U45012 (N_45012,N_42488,N_42097);
and U45013 (N_45013,N_43965,N_43418);
nand U45014 (N_45014,N_43217,N_42047);
and U45015 (N_45015,N_43967,N_42586);
or U45016 (N_45016,N_42400,N_42523);
or U45017 (N_45017,N_43763,N_43058);
nand U45018 (N_45018,N_43932,N_43748);
or U45019 (N_45019,N_43584,N_42519);
or U45020 (N_45020,N_43597,N_42684);
nand U45021 (N_45021,N_43993,N_42993);
nor U45022 (N_45022,N_43701,N_43252);
or U45023 (N_45023,N_43965,N_42697);
or U45024 (N_45024,N_42752,N_43909);
nand U45025 (N_45025,N_42618,N_43827);
nor U45026 (N_45026,N_42619,N_42883);
and U45027 (N_45027,N_43064,N_43477);
or U45028 (N_45028,N_42677,N_42869);
and U45029 (N_45029,N_43802,N_42279);
nand U45030 (N_45030,N_42209,N_43651);
xor U45031 (N_45031,N_43718,N_42563);
and U45032 (N_45032,N_43556,N_42143);
and U45033 (N_45033,N_43689,N_43099);
or U45034 (N_45034,N_43399,N_43683);
xor U45035 (N_45035,N_42018,N_43497);
xnor U45036 (N_45036,N_43489,N_43611);
nor U45037 (N_45037,N_42548,N_43069);
nor U45038 (N_45038,N_42963,N_42900);
and U45039 (N_45039,N_43120,N_43835);
nand U45040 (N_45040,N_43100,N_42308);
and U45041 (N_45041,N_42374,N_43882);
nor U45042 (N_45042,N_43189,N_43483);
and U45043 (N_45043,N_42382,N_42855);
nor U45044 (N_45044,N_43760,N_43851);
nand U45045 (N_45045,N_43578,N_43158);
xnor U45046 (N_45046,N_42539,N_43419);
and U45047 (N_45047,N_43755,N_43765);
or U45048 (N_45048,N_42678,N_43608);
and U45049 (N_45049,N_43934,N_42592);
xor U45050 (N_45050,N_43251,N_43312);
nor U45051 (N_45051,N_43453,N_43608);
nand U45052 (N_45052,N_43183,N_42666);
or U45053 (N_45053,N_43682,N_42953);
and U45054 (N_45054,N_42545,N_42495);
nor U45055 (N_45055,N_43084,N_42275);
xnor U45056 (N_45056,N_42200,N_43514);
nand U45057 (N_45057,N_43674,N_43320);
and U45058 (N_45058,N_43767,N_42427);
nand U45059 (N_45059,N_43829,N_42855);
nand U45060 (N_45060,N_43783,N_42182);
xor U45061 (N_45061,N_43035,N_42866);
or U45062 (N_45062,N_42224,N_43885);
xnor U45063 (N_45063,N_42182,N_43306);
and U45064 (N_45064,N_42385,N_43138);
and U45065 (N_45065,N_43420,N_43281);
nor U45066 (N_45066,N_43792,N_42247);
xnor U45067 (N_45067,N_42900,N_42796);
and U45068 (N_45068,N_43471,N_42381);
and U45069 (N_45069,N_42385,N_43130);
nor U45070 (N_45070,N_43248,N_43250);
nand U45071 (N_45071,N_43357,N_43715);
nor U45072 (N_45072,N_42727,N_43693);
nor U45073 (N_45073,N_42819,N_43247);
nor U45074 (N_45074,N_43185,N_43602);
xor U45075 (N_45075,N_43399,N_42240);
nor U45076 (N_45076,N_42436,N_43074);
nand U45077 (N_45077,N_42066,N_43923);
xor U45078 (N_45078,N_43388,N_43586);
xor U45079 (N_45079,N_42381,N_42197);
nor U45080 (N_45080,N_42623,N_42492);
xor U45081 (N_45081,N_42335,N_43241);
nand U45082 (N_45082,N_43123,N_42144);
and U45083 (N_45083,N_42577,N_42416);
nor U45084 (N_45084,N_42259,N_43634);
nor U45085 (N_45085,N_42068,N_43953);
or U45086 (N_45086,N_42871,N_42950);
and U45087 (N_45087,N_43591,N_43026);
or U45088 (N_45088,N_43597,N_42990);
and U45089 (N_45089,N_43901,N_43539);
or U45090 (N_45090,N_42733,N_43742);
nand U45091 (N_45091,N_42186,N_42162);
nand U45092 (N_45092,N_43624,N_42989);
and U45093 (N_45093,N_43055,N_42389);
or U45094 (N_45094,N_42096,N_43074);
nand U45095 (N_45095,N_42872,N_43852);
nand U45096 (N_45096,N_43795,N_43389);
and U45097 (N_45097,N_43875,N_42878);
nor U45098 (N_45098,N_42886,N_43540);
and U45099 (N_45099,N_43338,N_43623);
and U45100 (N_45100,N_43270,N_43311);
or U45101 (N_45101,N_43821,N_43526);
and U45102 (N_45102,N_43491,N_42236);
nor U45103 (N_45103,N_42718,N_42725);
nor U45104 (N_45104,N_43786,N_42796);
nor U45105 (N_45105,N_43614,N_42654);
nand U45106 (N_45106,N_42828,N_43750);
xnor U45107 (N_45107,N_43788,N_42121);
and U45108 (N_45108,N_43512,N_42020);
and U45109 (N_45109,N_42465,N_42857);
nor U45110 (N_45110,N_43083,N_42425);
and U45111 (N_45111,N_43061,N_43703);
nor U45112 (N_45112,N_43078,N_43265);
and U45113 (N_45113,N_42360,N_43512);
and U45114 (N_45114,N_42527,N_43182);
nor U45115 (N_45115,N_43256,N_43191);
xnor U45116 (N_45116,N_42947,N_42845);
xnor U45117 (N_45117,N_43167,N_43969);
nand U45118 (N_45118,N_43619,N_42203);
nand U45119 (N_45119,N_42821,N_42307);
or U45120 (N_45120,N_43375,N_43877);
and U45121 (N_45121,N_43877,N_43106);
or U45122 (N_45122,N_42822,N_43078);
nor U45123 (N_45123,N_42860,N_43474);
or U45124 (N_45124,N_42937,N_43507);
and U45125 (N_45125,N_43116,N_43563);
nand U45126 (N_45126,N_42266,N_42732);
nand U45127 (N_45127,N_43496,N_42804);
nand U45128 (N_45128,N_42213,N_43325);
xnor U45129 (N_45129,N_42875,N_43814);
and U45130 (N_45130,N_43866,N_43284);
or U45131 (N_45131,N_43224,N_42700);
nor U45132 (N_45132,N_43332,N_43680);
nand U45133 (N_45133,N_42211,N_43009);
or U45134 (N_45134,N_43818,N_43469);
nand U45135 (N_45135,N_42788,N_43757);
and U45136 (N_45136,N_42599,N_42693);
nor U45137 (N_45137,N_43845,N_42199);
nor U45138 (N_45138,N_42409,N_43958);
or U45139 (N_45139,N_43320,N_43198);
xnor U45140 (N_45140,N_42716,N_43140);
xor U45141 (N_45141,N_42505,N_43739);
and U45142 (N_45142,N_43797,N_42690);
and U45143 (N_45143,N_42884,N_43490);
nor U45144 (N_45144,N_42668,N_42046);
nor U45145 (N_45145,N_42580,N_43955);
or U45146 (N_45146,N_42535,N_42079);
and U45147 (N_45147,N_43577,N_42256);
nor U45148 (N_45148,N_43407,N_43390);
or U45149 (N_45149,N_43951,N_42927);
nand U45150 (N_45150,N_43988,N_42239);
or U45151 (N_45151,N_42958,N_42806);
or U45152 (N_45152,N_42693,N_43546);
or U45153 (N_45153,N_42077,N_42087);
or U45154 (N_45154,N_43150,N_43257);
nand U45155 (N_45155,N_43526,N_43580);
and U45156 (N_45156,N_43690,N_42004);
xnor U45157 (N_45157,N_42373,N_42107);
or U45158 (N_45158,N_42426,N_42674);
or U45159 (N_45159,N_43876,N_42178);
nor U45160 (N_45160,N_42218,N_43235);
nand U45161 (N_45161,N_43385,N_43010);
or U45162 (N_45162,N_43047,N_42515);
nor U45163 (N_45163,N_42808,N_42998);
nand U45164 (N_45164,N_43603,N_43080);
and U45165 (N_45165,N_42905,N_43906);
xor U45166 (N_45166,N_43857,N_42855);
or U45167 (N_45167,N_43429,N_42348);
nor U45168 (N_45168,N_43115,N_43228);
and U45169 (N_45169,N_42740,N_42293);
and U45170 (N_45170,N_42100,N_43238);
xnor U45171 (N_45171,N_43166,N_43349);
and U45172 (N_45172,N_43294,N_42877);
and U45173 (N_45173,N_42299,N_42620);
xor U45174 (N_45174,N_42849,N_43794);
or U45175 (N_45175,N_42605,N_42026);
xor U45176 (N_45176,N_43963,N_42554);
or U45177 (N_45177,N_43388,N_43420);
or U45178 (N_45178,N_43725,N_42480);
and U45179 (N_45179,N_43540,N_43452);
nor U45180 (N_45180,N_43178,N_42444);
nor U45181 (N_45181,N_42959,N_43799);
and U45182 (N_45182,N_43388,N_42257);
or U45183 (N_45183,N_43255,N_43320);
nor U45184 (N_45184,N_43117,N_42470);
or U45185 (N_45185,N_42513,N_42538);
nor U45186 (N_45186,N_43472,N_42337);
and U45187 (N_45187,N_42728,N_43402);
nor U45188 (N_45188,N_43633,N_42266);
and U45189 (N_45189,N_43253,N_42758);
and U45190 (N_45190,N_42006,N_43106);
nand U45191 (N_45191,N_42565,N_43271);
nor U45192 (N_45192,N_43453,N_42726);
or U45193 (N_45193,N_42506,N_42048);
nor U45194 (N_45194,N_43633,N_43072);
or U45195 (N_45195,N_43803,N_42058);
nand U45196 (N_45196,N_42692,N_43595);
or U45197 (N_45197,N_43128,N_43743);
or U45198 (N_45198,N_43956,N_43859);
xor U45199 (N_45199,N_43938,N_42815);
and U45200 (N_45200,N_42887,N_42978);
nand U45201 (N_45201,N_42874,N_42084);
or U45202 (N_45202,N_42638,N_42469);
nor U45203 (N_45203,N_42423,N_42286);
nand U45204 (N_45204,N_43095,N_42481);
nand U45205 (N_45205,N_43854,N_42133);
xnor U45206 (N_45206,N_42100,N_42793);
and U45207 (N_45207,N_43039,N_43439);
and U45208 (N_45208,N_43512,N_43750);
xor U45209 (N_45209,N_42118,N_43638);
nand U45210 (N_45210,N_42790,N_43624);
nand U45211 (N_45211,N_42174,N_43447);
nand U45212 (N_45212,N_42176,N_43696);
nand U45213 (N_45213,N_42205,N_42776);
nor U45214 (N_45214,N_43518,N_43605);
and U45215 (N_45215,N_43720,N_42564);
xor U45216 (N_45216,N_43466,N_43628);
and U45217 (N_45217,N_42192,N_42260);
and U45218 (N_45218,N_43790,N_43156);
nand U45219 (N_45219,N_42824,N_43285);
nor U45220 (N_45220,N_42499,N_42694);
nor U45221 (N_45221,N_43067,N_42597);
nand U45222 (N_45222,N_42820,N_42904);
and U45223 (N_45223,N_42386,N_43196);
nor U45224 (N_45224,N_42325,N_42327);
xor U45225 (N_45225,N_43422,N_42104);
xnor U45226 (N_45226,N_42536,N_42222);
xor U45227 (N_45227,N_42039,N_42544);
nor U45228 (N_45228,N_42954,N_43128);
nor U45229 (N_45229,N_42500,N_42466);
or U45230 (N_45230,N_43506,N_42410);
xor U45231 (N_45231,N_43967,N_42393);
and U45232 (N_45232,N_43084,N_42552);
or U45233 (N_45233,N_43754,N_42932);
and U45234 (N_45234,N_43915,N_43962);
xor U45235 (N_45235,N_43894,N_42351);
or U45236 (N_45236,N_43978,N_42349);
xnor U45237 (N_45237,N_43368,N_42831);
nand U45238 (N_45238,N_43580,N_43617);
or U45239 (N_45239,N_43568,N_43947);
nand U45240 (N_45240,N_43771,N_43717);
and U45241 (N_45241,N_43086,N_43449);
xor U45242 (N_45242,N_42321,N_43638);
or U45243 (N_45243,N_42054,N_42992);
xor U45244 (N_45244,N_42955,N_43295);
or U45245 (N_45245,N_42951,N_42518);
nor U45246 (N_45246,N_43021,N_42761);
nor U45247 (N_45247,N_43338,N_42474);
or U45248 (N_45248,N_43125,N_42609);
nand U45249 (N_45249,N_43216,N_43813);
nor U45250 (N_45250,N_42151,N_43858);
and U45251 (N_45251,N_42882,N_43450);
nand U45252 (N_45252,N_42887,N_43350);
and U45253 (N_45253,N_43473,N_42733);
or U45254 (N_45254,N_43647,N_42681);
xnor U45255 (N_45255,N_42721,N_43723);
and U45256 (N_45256,N_43424,N_42152);
and U45257 (N_45257,N_43602,N_43061);
or U45258 (N_45258,N_42650,N_43762);
xnor U45259 (N_45259,N_42746,N_42952);
or U45260 (N_45260,N_42709,N_43454);
xor U45261 (N_45261,N_43265,N_42824);
nand U45262 (N_45262,N_43559,N_43803);
xnor U45263 (N_45263,N_42839,N_43951);
or U45264 (N_45264,N_43070,N_43952);
nand U45265 (N_45265,N_42475,N_43562);
xnor U45266 (N_45266,N_43915,N_43577);
xor U45267 (N_45267,N_42239,N_43606);
nor U45268 (N_45268,N_43832,N_43745);
nor U45269 (N_45269,N_42958,N_43446);
nand U45270 (N_45270,N_43006,N_42981);
or U45271 (N_45271,N_42954,N_43140);
and U45272 (N_45272,N_43321,N_43714);
xor U45273 (N_45273,N_43826,N_42305);
and U45274 (N_45274,N_42900,N_42154);
and U45275 (N_45275,N_43672,N_42205);
xor U45276 (N_45276,N_43062,N_42534);
nand U45277 (N_45277,N_43414,N_43958);
nand U45278 (N_45278,N_42036,N_43037);
xor U45279 (N_45279,N_43644,N_43710);
xnor U45280 (N_45280,N_42396,N_43574);
or U45281 (N_45281,N_42705,N_42577);
or U45282 (N_45282,N_42456,N_43165);
nor U45283 (N_45283,N_42423,N_42771);
nor U45284 (N_45284,N_42187,N_42308);
and U45285 (N_45285,N_43747,N_43051);
xnor U45286 (N_45286,N_43298,N_42829);
nor U45287 (N_45287,N_42818,N_42104);
nand U45288 (N_45288,N_42062,N_42269);
nand U45289 (N_45289,N_42954,N_43149);
or U45290 (N_45290,N_43079,N_42362);
or U45291 (N_45291,N_43074,N_42474);
and U45292 (N_45292,N_42992,N_43374);
xnor U45293 (N_45293,N_43202,N_43495);
xor U45294 (N_45294,N_43007,N_42592);
nor U45295 (N_45295,N_43735,N_42135);
nand U45296 (N_45296,N_43507,N_42773);
nand U45297 (N_45297,N_43777,N_43283);
xor U45298 (N_45298,N_42393,N_42610);
nand U45299 (N_45299,N_43175,N_43804);
or U45300 (N_45300,N_43093,N_42635);
or U45301 (N_45301,N_43642,N_42409);
or U45302 (N_45302,N_43794,N_42836);
nor U45303 (N_45303,N_42298,N_43014);
xnor U45304 (N_45304,N_42068,N_42218);
or U45305 (N_45305,N_43132,N_42146);
nor U45306 (N_45306,N_43578,N_42780);
nand U45307 (N_45307,N_42920,N_43208);
xor U45308 (N_45308,N_43336,N_42746);
xnor U45309 (N_45309,N_42977,N_42347);
or U45310 (N_45310,N_42318,N_42279);
and U45311 (N_45311,N_43236,N_43843);
xor U45312 (N_45312,N_43193,N_42477);
and U45313 (N_45313,N_43200,N_43303);
nand U45314 (N_45314,N_43740,N_42782);
nand U45315 (N_45315,N_42525,N_42789);
xnor U45316 (N_45316,N_43529,N_42245);
nand U45317 (N_45317,N_43060,N_43204);
nand U45318 (N_45318,N_43568,N_42050);
and U45319 (N_45319,N_42769,N_43994);
nand U45320 (N_45320,N_43605,N_43187);
nor U45321 (N_45321,N_42269,N_42750);
nand U45322 (N_45322,N_43941,N_43038);
nand U45323 (N_45323,N_42041,N_43183);
or U45324 (N_45324,N_43659,N_42373);
and U45325 (N_45325,N_42299,N_42400);
nand U45326 (N_45326,N_43261,N_43069);
xnor U45327 (N_45327,N_43208,N_42157);
or U45328 (N_45328,N_42541,N_43806);
and U45329 (N_45329,N_42966,N_42833);
nand U45330 (N_45330,N_42802,N_42046);
nor U45331 (N_45331,N_43480,N_42590);
xnor U45332 (N_45332,N_42764,N_42960);
nand U45333 (N_45333,N_42024,N_42457);
or U45334 (N_45334,N_42718,N_43567);
or U45335 (N_45335,N_43090,N_43893);
nor U45336 (N_45336,N_42037,N_42922);
and U45337 (N_45337,N_43131,N_43844);
nor U45338 (N_45338,N_42167,N_43639);
or U45339 (N_45339,N_43942,N_43781);
nor U45340 (N_45340,N_42314,N_43249);
xor U45341 (N_45341,N_43961,N_42655);
and U45342 (N_45342,N_42434,N_42983);
and U45343 (N_45343,N_42140,N_43169);
and U45344 (N_45344,N_42471,N_42673);
nor U45345 (N_45345,N_43682,N_42296);
and U45346 (N_45346,N_43953,N_42521);
nand U45347 (N_45347,N_42714,N_42653);
nor U45348 (N_45348,N_43191,N_43876);
nor U45349 (N_45349,N_43777,N_42610);
nor U45350 (N_45350,N_43042,N_43810);
xnor U45351 (N_45351,N_43210,N_43999);
and U45352 (N_45352,N_43449,N_42069);
nor U45353 (N_45353,N_42036,N_42041);
xor U45354 (N_45354,N_43705,N_42452);
and U45355 (N_45355,N_43314,N_43307);
nor U45356 (N_45356,N_42815,N_43013);
and U45357 (N_45357,N_42021,N_42172);
and U45358 (N_45358,N_42707,N_42442);
and U45359 (N_45359,N_42860,N_43353);
xnor U45360 (N_45360,N_43570,N_42361);
xnor U45361 (N_45361,N_43470,N_42058);
xor U45362 (N_45362,N_42991,N_43385);
or U45363 (N_45363,N_42360,N_42851);
xor U45364 (N_45364,N_42342,N_43296);
nand U45365 (N_45365,N_43528,N_43075);
xor U45366 (N_45366,N_42957,N_43360);
or U45367 (N_45367,N_42315,N_43896);
nand U45368 (N_45368,N_43739,N_43861);
and U45369 (N_45369,N_42860,N_43780);
xor U45370 (N_45370,N_42055,N_42934);
nor U45371 (N_45371,N_43315,N_42451);
or U45372 (N_45372,N_43820,N_43504);
nand U45373 (N_45373,N_42929,N_43836);
or U45374 (N_45374,N_42683,N_42262);
nor U45375 (N_45375,N_43323,N_43267);
nor U45376 (N_45376,N_42928,N_43249);
nor U45377 (N_45377,N_42121,N_42638);
and U45378 (N_45378,N_42567,N_42757);
and U45379 (N_45379,N_43272,N_42976);
xor U45380 (N_45380,N_42677,N_43583);
xnor U45381 (N_45381,N_42763,N_43177);
and U45382 (N_45382,N_42971,N_43231);
nand U45383 (N_45383,N_43337,N_43566);
nand U45384 (N_45384,N_43538,N_42853);
nand U45385 (N_45385,N_43539,N_42255);
or U45386 (N_45386,N_43075,N_42861);
nor U45387 (N_45387,N_42432,N_43351);
nor U45388 (N_45388,N_43376,N_43247);
xnor U45389 (N_45389,N_43718,N_43575);
or U45390 (N_45390,N_42470,N_42629);
nor U45391 (N_45391,N_43583,N_43255);
or U45392 (N_45392,N_42625,N_42367);
nand U45393 (N_45393,N_42097,N_42850);
nor U45394 (N_45394,N_43538,N_42310);
nand U45395 (N_45395,N_42182,N_43237);
nand U45396 (N_45396,N_43692,N_43827);
nor U45397 (N_45397,N_43716,N_43116);
nand U45398 (N_45398,N_43907,N_43817);
or U45399 (N_45399,N_42841,N_42876);
or U45400 (N_45400,N_43794,N_43527);
and U45401 (N_45401,N_43862,N_43938);
nand U45402 (N_45402,N_43659,N_43473);
or U45403 (N_45403,N_42002,N_43313);
nand U45404 (N_45404,N_42283,N_43256);
nand U45405 (N_45405,N_43643,N_42141);
or U45406 (N_45406,N_43715,N_43392);
and U45407 (N_45407,N_42752,N_43784);
xor U45408 (N_45408,N_42171,N_42253);
nor U45409 (N_45409,N_42026,N_43062);
and U45410 (N_45410,N_42795,N_42052);
nor U45411 (N_45411,N_42710,N_42579);
nor U45412 (N_45412,N_43863,N_43017);
xnor U45413 (N_45413,N_42319,N_42665);
or U45414 (N_45414,N_42184,N_43091);
xor U45415 (N_45415,N_42381,N_42830);
nor U45416 (N_45416,N_42138,N_42499);
or U45417 (N_45417,N_42124,N_42609);
xor U45418 (N_45418,N_43590,N_42060);
xor U45419 (N_45419,N_43366,N_42910);
and U45420 (N_45420,N_43618,N_43148);
nor U45421 (N_45421,N_42292,N_43470);
and U45422 (N_45422,N_43251,N_43405);
nor U45423 (N_45423,N_42556,N_43177);
or U45424 (N_45424,N_43748,N_43791);
and U45425 (N_45425,N_42349,N_43635);
xor U45426 (N_45426,N_43470,N_43567);
and U45427 (N_45427,N_42688,N_42866);
or U45428 (N_45428,N_43198,N_43307);
xnor U45429 (N_45429,N_42444,N_42299);
or U45430 (N_45430,N_42870,N_42280);
nand U45431 (N_45431,N_42849,N_43490);
and U45432 (N_45432,N_43915,N_42405);
xnor U45433 (N_45433,N_43786,N_42941);
or U45434 (N_45434,N_43926,N_43195);
nand U45435 (N_45435,N_43366,N_42004);
or U45436 (N_45436,N_42608,N_42241);
or U45437 (N_45437,N_43289,N_42504);
xnor U45438 (N_45438,N_43564,N_43476);
or U45439 (N_45439,N_43783,N_42952);
and U45440 (N_45440,N_43987,N_42111);
xnor U45441 (N_45441,N_43942,N_43868);
nand U45442 (N_45442,N_42414,N_43056);
nand U45443 (N_45443,N_43492,N_43062);
nor U45444 (N_45444,N_43789,N_43350);
or U45445 (N_45445,N_43252,N_42081);
and U45446 (N_45446,N_43618,N_43487);
nor U45447 (N_45447,N_42915,N_42672);
and U45448 (N_45448,N_42009,N_43289);
nor U45449 (N_45449,N_42012,N_42883);
nand U45450 (N_45450,N_42626,N_42549);
xnor U45451 (N_45451,N_42022,N_42560);
nor U45452 (N_45452,N_42600,N_42708);
and U45453 (N_45453,N_42547,N_43788);
nand U45454 (N_45454,N_43431,N_42301);
nand U45455 (N_45455,N_42534,N_42836);
nor U45456 (N_45456,N_43838,N_42426);
nand U45457 (N_45457,N_43481,N_42838);
nand U45458 (N_45458,N_42312,N_42752);
nand U45459 (N_45459,N_43888,N_43952);
and U45460 (N_45460,N_42958,N_43644);
and U45461 (N_45461,N_42339,N_42689);
xnor U45462 (N_45462,N_43469,N_42256);
and U45463 (N_45463,N_43445,N_43805);
nand U45464 (N_45464,N_42704,N_42138);
nor U45465 (N_45465,N_42574,N_43210);
and U45466 (N_45466,N_42518,N_42595);
nand U45467 (N_45467,N_42055,N_42716);
xnor U45468 (N_45468,N_43559,N_42619);
xor U45469 (N_45469,N_43981,N_43109);
and U45470 (N_45470,N_43332,N_43120);
nand U45471 (N_45471,N_43262,N_43151);
or U45472 (N_45472,N_42449,N_42139);
nand U45473 (N_45473,N_42681,N_43343);
and U45474 (N_45474,N_42808,N_43001);
and U45475 (N_45475,N_43173,N_43817);
and U45476 (N_45476,N_43483,N_43121);
or U45477 (N_45477,N_43839,N_43686);
nand U45478 (N_45478,N_42287,N_42475);
nand U45479 (N_45479,N_42675,N_43168);
xor U45480 (N_45480,N_43739,N_42357);
or U45481 (N_45481,N_43009,N_43116);
and U45482 (N_45482,N_42072,N_43349);
and U45483 (N_45483,N_43534,N_42367);
and U45484 (N_45484,N_43320,N_43099);
xor U45485 (N_45485,N_42857,N_43455);
and U45486 (N_45486,N_42072,N_43256);
or U45487 (N_45487,N_42195,N_43294);
and U45488 (N_45488,N_42253,N_43295);
xor U45489 (N_45489,N_42153,N_43467);
nand U45490 (N_45490,N_42488,N_42547);
nand U45491 (N_45491,N_43879,N_43312);
and U45492 (N_45492,N_42918,N_43998);
or U45493 (N_45493,N_42071,N_42372);
or U45494 (N_45494,N_43857,N_43100);
or U45495 (N_45495,N_43672,N_43247);
xor U45496 (N_45496,N_42782,N_42446);
nand U45497 (N_45497,N_43396,N_43378);
xor U45498 (N_45498,N_43847,N_43098);
xnor U45499 (N_45499,N_42557,N_43843);
and U45500 (N_45500,N_43430,N_42634);
nor U45501 (N_45501,N_42333,N_43771);
and U45502 (N_45502,N_43492,N_42098);
and U45503 (N_45503,N_43698,N_42998);
nor U45504 (N_45504,N_43947,N_42975);
xor U45505 (N_45505,N_42822,N_43784);
and U45506 (N_45506,N_43278,N_43632);
xor U45507 (N_45507,N_42909,N_43476);
nor U45508 (N_45508,N_42779,N_43372);
or U45509 (N_45509,N_42066,N_42385);
nor U45510 (N_45510,N_43193,N_42604);
xnor U45511 (N_45511,N_43352,N_43819);
nand U45512 (N_45512,N_42187,N_43299);
or U45513 (N_45513,N_43483,N_43165);
xor U45514 (N_45514,N_42150,N_42336);
nand U45515 (N_45515,N_43996,N_43706);
and U45516 (N_45516,N_42705,N_42718);
and U45517 (N_45517,N_43468,N_43001);
or U45518 (N_45518,N_43685,N_42903);
and U45519 (N_45519,N_43381,N_42087);
nand U45520 (N_45520,N_42346,N_42546);
or U45521 (N_45521,N_43941,N_42525);
nor U45522 (N_45522,N_42824,N_42346);
and U45523 (N_45523,N_43007,N_43349);
xor U45524 (N_45524,N_42189,N_43482);
and U45525 (N_45525,N_42466,N_42573);
and U45526 (N_45526,N_43184,N_43250);
nand U45527 (N_45527,N_43785,N_42030);
and U45528 (N_45528,N_43521,N_43194);
nor U45529 (N_45529,N_42260,N_43726);
nor U45530 (N_45530,N_42095,N_42122);
xor U45531 (N_45531,N_42943,N_42383);
nor U45532 (N_45532,N_43321,N_42370);
nand U45533 (N_45533,N_43008,N_43697);
nand U45534 (N_45534,N_43024,N_43872);
or U45535 (N_45535,N_42683,N_43351);
nor U45536 (N_45536,N_42632,N_42041);
nor U45537 (N_45537,N_43439,N_42626);
nand U45538 (N_45538,N_42449,N_43364);
and U45539 (N_45539,N_42794,N_42978);
nand U45540 (N_45540,N_43639,N_43673);
and U45541 (N_45541,N_42350,N_43563);
and U45542 (N_45542,N_42213,N_43316);
xnor U45543 (N_45543,N_42338,N_42916);
xnor U45544 (N_45544,N_42896,N_42348);
and U45545 (N_45545,N_43655,N_43172);
nand U45546 (N_45546,N_42939,N_42092);
and U45547 (N_45547,N_42713,N_42134);
and U45548 (N_45548,N_43918,N_42803);
xor U45549 (N_45549,N_42768,N_42609);
nor U45550 (N_45550,N_43301,N_43762);
nor U45551 (N_45551,N_42395,N_43062);
nor U45552 (N_45552,N_42448,N_42402);
nand U45553 (N_45553,N_42665,N_42430);
nand U45554 (N_45554,N_43016,N_42431);
nand U45555 (N_45555,N_42531,N_43283);
or U45556 (N_45556,N_43071,N_42374);
or U45557 (N_45557,N_43470,N_42483);
and U45558 (N_45558,N_43779,N_43143);
nand U45559 (N_45559,N_42299,N_43613);
xor U45560 (N_45560,N_43139,N_43055);
and U45561 (N_45561,N_43773,N_42127);
xnor U45562 (N_45562,N_42565,N_42172);
and U45563 (N_45563,N_42366,N_43755);
and U45564 (N_45564,N_42481,N_42235);
or U45565 (N_45565,N_42557,N_42241);
and U45566 (N_45566,N_42445,N_42193);
xnor U45567 (N_45567,N_42851,N_43319);
nand U45568 (N_45568,N_43088,N_43359);
nor U45569 (N_45569,N_42618,N_43318);
or U45570 (N_45570,N_43354,N_42450);
nand U45571 (N_45571,N_43222,N_42846);
xnor U45572 (N_45572,N_42803,N_42481);
and U45573 (N_45573,N_43157,N_43071);
xor U45574 (N_45574,N_42111,N_43810);
nand U45575 (N_45575,N_42609,N_42890);
nand U45576 (N_45576,N_43578,N_42038);
nand U45577 (N_45577,N_43891,N_43902);
and U45578 (N_45578,N_42765,N_43261);
and U45579 (N_45579,N_43277,N_42769);
xor U45580 (N_45580,N_42961,N_42941);
nand U45581 (N_45581,N_43757,N_43891);
xnor U45582 (N_45582,N_43199,N_43035);
xor U45583 (N_45583,N_43764,N_43876);
xor U45584 (N_45584,N_42787,N_42290);
and U45585 (N_45585,N_42923,N_42401);
or U45586 (N_45586,N_42858,N_42626);
nand U45587 (N_45587,N_43610,N_42874);
nand U45588 (N_45588,N_43348,N_42845);
nand U45589 (N_45589,N_43636,N_43291);
nor U45590 (N_45590,N_42569,N_42032);
nor U45591 (N_45591,N_43905,N_42548);
and U45592 (N_45592,N_43094,N_42129);
nor U45593 (N_45593,N_43972,N_43791);
or U45594 (N_45594,N_43413,N_43211);
xnor U45595 (N_45595,N_43258,N_43768);
nor U45596 (N_45596,N_42778,N_42160);
and U45597 (N_45597,N_42845,N_43242);
nor U45598 (N_45598,N_42959,N_43205);
and U45599 (N_45599,N_42089,N_43351);
nand U45600 (N_45600,N_43967,N_43409);
or U45601 (N_45601,N_42488,N_42523);
or U45602 (N_45602,N_42316,N_42421);
nand U45603 (N_45603,N_42574,N_42855);
nand U45604 (N_45604,N_42686,N_43276);
and U45605 (N_45605,N_42635,N_43698);
nor U45606 (N_45606,N_42214,N_43818);
or U45607 (N_45607,N_43873,N_43019);
nand U45608 (N_45608,N_43642,N_43515);
xor U45609 (N_45609,N_43206,N_43529);
nand U45610 (N_45610,N_43274,N_43734);
nor U45611 (N_45611,N_43103,N_43723);
and U45612 (N_45612,N_42002,N_43496);
and U45613 (N_45613,N_43907,N_42044);
xor U45614 (N_45614,N_42521,N_42360);
nand U45615 (N_45615,N_42194,N_42405);
and U45616 (N_45616,N_43527,N_42239);
or U45617 (N_45617,N_42107,N_42423);
xnor U45618 (N_45618,N_43256,N_42857);
nand U45619 (N_45619,N_43242,N_43041);
or U45620 (N_45620,N_42268,N_43994);
or U45621 (N_45621,N_42631,N_43972);
nor U45622 (N_45622,N_42726,N_42117);
nor U45623 (N_45623,N_42734,N_43810);
and U45624 (N_45624,N_42244,N_43859);
or U45625 (N_45625,N_42446,N_43981);
nor U45626 (N_45626,N_43668,N_42633);
nand U45627 (N_45627,N_43663,N_42769);
and U45628 (N_45628,N_43073,N_42338);
and U45629 (N_45629,N_43366,N_43062);
xnor U45630 (N_45630,N_43649,N_43176);
or U45631 (N_45631,N_42061,N_43608);
nor U45632 (N_45632,N_42315,N_43784);
or U45633 (N_45633,N_43743,N_43479);
and U45634 (N_45634,N_42648,N_43097);
nor U45635 (N_45635,N_43529,N_42024);
nand U45636 (N_45636,N_43886,N_42048);
or U45637 (N_45637,N_43948,N_42133);
and U45638 (N_45638,N_42346,N_42158);
nand U45639 (N_45639,N_42602,N_42852);
nor U45640 (N_45640,N_43886,N_43691);
nand U45641 (N_45641,N_43469,N_43573);
nor U45642 (N_45642,N_43528,N_42292);
xor U45643 (N_45643,N_42938,N_42345);
and U45644 (N_45644,N_43984,N_43171);
and U45645 (N_45645,N_42090,N_43188);
xor U45646 (N_45646,N_42659,N_42145);
xnor U45647 (N_45647,N_42577,N_42935);
nand U45648 (N_45648,N_43575,N_43129);
nand U45649 (N_45649,N_42106,N_43169);
xnor U45650 (N_45650,N_42390,N_43785);
nor U45651 (N_45651,N_42696,N_43477);
and U45652 (N_45652,N_43601,N_42463);
nand U45653 (N_45653,N_42312,N_42136);
nor U45654 (N_45654,N_42381,N_42784);
xnor U45655 (N_45655,N_42847,N_43717);
or U45656 (N_45656,N_43299,N_42371);
and U45657 (N_45657,N_42959,N_42730);
nand U45658 (N_45658,N_42435,N_43819);
or U45659 (N_45659,N_42730,N_43668);
and U45660 (N_45660,N_42717,N_43808);
nand U45661 (N_45661,N_42983,N_42134);
nand U45662 (N_45662,N_43935,N_42610);
xor U45663 (N_45663,N_43772,N_43769);
nor U45664 (N_45664,N_43809,N_43977);
nor U45665 (N_45665,N_42999,N_42044);
xor U45666 (N_45666,N_42624,N_43902);
and U45667 (N_45667,N_43995,N_43232);
or U45668 (N_45668,N_42389,N_42843);
nor U45669 (N_45669,N_42938,N_43529);
xnor U45670 (N_45670,N_43022,N_42444);
xor U45671 (N_45671,N_43075,N_43572);
nand U45672 (N_45672,N_42496,N_42173);
xnor U45673 (N_45673,N_43714,N_42865);
nor U45674 (N_45674,N_42994,N_42087);
or U45675 (N_45675,N_43486,N_42834);
nand U45676 (N_45676,N_43467,N_43694);
and U45677 (N_45677,N_42176,N_42178);
nor U45678 (N_45678,N_42996,N_42870);
nand U45679 (N_45679,N_42843,N_42895);
and U45680 (N_45680,N_43618,N_43250);
or U45681 (N_45681,N_43304,N_42081);
and U45682 (N_45682,N_43116,N_42021);
nand U45683 (N_45683,N_42139,N_42735);
nor U45684 (N_45684,N_42142,N_43717);
nand U45685 (N_45685,N_42350,N_43547);
xnor U45686 (N_45686,N_42535,N_43006);
xnor U45687 (N_45687,N_42505,N_43683);
or U45688 (N_45688,N_42612,N_43464);
and U45689 (N_45689,N_43632,N_43960);
xnor U45690 (N_45690,N_42477,N_43281);
and U45691 (N_45691,N_43680,N_42280);
and U45692 (N_45692,N_43121,N_42134);
or U45693 (N_45693,N_42118,N_43566);
nand U45694 (N_45694,N_42929,N_42330);
xor U45695 (N_45695,N_42163,N_42551);
nor U45696 (N_45696,N_42859,N_43145);
xnor U45697 (N_45697,N_43780,N_43814);
and U45698 (N_45698,N_43622,N_43866);
or U45699 (N_45699,N_43190,N_42452);
nand U45700 (N_45700,N_42959,N_42590);
or U45701 (N_45701,N_42939,N_43518);
and U45702 (N_45702,N_43613,N_42476);
xor U45703 (N_45703,N_43773,N_43761);
nor U45704 (N_45704,N_42592,N_42751);
or U45705 (N_45705,N_43443,N_42550);
xnor U45706 (N_45706,N_42948,N_42302);
and U45707 (N_45707,N_42491,N_42878);
and U45708 (N_45708,N_43469,N_43975);
xnor U45709 (N_45709,N_43487,N_42988);
or U45710 (N_45710,N_42015,N_43710);
xnor U45711 (N_45711,N_43220,N_43964);
xor U45712 (N_45712,N_43845,N_43570);
or U45713 (N_45713,N_43499,N_43342);
xnor U45714 (N_45714,N_42477,N_43072);
nor U45715 (N_45715,N_42979,N_43419);
or U45716 (N_45716,N_43437,N_43115);
or U45717 (N_45717,N_42739,N_43161);
and U45718 (N_45718,N_42172,N_42268);
xnor U45719 (N_45719,N_42407,N_43760);
xor U45720 (N_45720,N_42489,N_43172);
nor U45721 (N_45721,N_42407,N_42134);
nor U45722 (N_45722,N_42353,N_43303);
or U45723 (N_45723,N_42616,N_43680);
nand U45724 (N_45724,N_42835,N_43158);
and U45725 (N_45725,N_42591,N_43060);
and U45726 (N_45726,N_42768,N_43580);
and U45727 (N_45727,N_42916,N_42223);
or U45728 (N_45728,N_43927,N_43537);
nand U45729 (N_45729,N_43795,N_42970);
or U45730 (N_45730,N_43177,N_42326);
nor U45731 (N_45731,N_42065,N_43293);
or U45732 (N_45732,N_42693,N_42475);
or U45733 (N_45733,N_42115,N_42901);
nand U45734 (N_45734,N_43974,N_43548);
nand U45735 (N_45735,N_43186,N_43476);
xor U45736 (N_45736,N_42349,N_42983);
xnor U45737 (N_45737,N_43844,N_42567);
nor U45738 (N_45738,N_43124,N_43468);
nor U45739 (N_45739,N_43322,N_43208);
and U45740 (N_45740,N_42646,N_43529);
xor U45741 (N_45741,N_43500,N_43119);
and U45742 (N_45742,N_43796,N_43359);
nand U45743 (N_45743,N_42454,N_43304);
xnor U45744 (N_45744,N_43733,N_43358);
and U45745 (N_45745,N_43720,N_43349);
nand U45746 (N_45746,N_43479,N_42097);
nand U45747 (N_45747,N_43599,N_43892);
xnor U45748 (N_45748,N_43320,N_43526);
nand U45749 (N_45749,N_43384,N_43289);
xnor U45750 (N_45750,N_42808,N_42798);
or U45751 (N_45751,N_42200,N_42655);
or U45752 (N_45752,N_43997,N_43875);
and U45753 (N_45753,N_42699,N_42159);
nand U45754 (N_45754,N_42095,N_42429);
nand U45755 (N_45755,N_42954,N_42501);
and U45756 (N_45756,N_42652,N_43563);
nor U45757 (N_45757,N_43047,N_43792);
nor U45758 (N_45758,N_42340,N_42514);
or U45759 (N_45759,N_43033,N_42370);
nor U45760 (N_45760,N_43001,N_43411);
nand U45761 (N_45761,N_43895,N_43764);
or U45762 (N_45762,N_43971,N_42994);
nor U45763 (N_45763,N_43580,N_43220);
nand U45764 (N_45764,N_43151,N_42400);
and U45765 (N_45765,N_42113,N_43743);
xnor U45766 (N_45766,N_43153,N_42187);
nand U45767 (N_45767,N_43021,N_42336);
xnor U45768 (N_45768,N_43278,N_42007);
nor U45769 (N_45769,N_43305,N_42319);
nor U45770 (N_45770,N_42609,N_43830);
and U45771 (N_45771,N_42743,N_42943);
or U45772 (N_45772,N_43614,N_43606);
xnor U45773 (N_45773,N_42790,N_42058);
and U45774 (N_45774,N_42756,N_42546);
and U45775 (N_45775,N_42919,N_43025);
and U45776 (N_45776,N_43186,N_42894);
and U45777 (N_45777,N_42418,N_42103);
or U45778 (N_45778,N_42790,N_43370);
nor U45779 (N_45779,N_42857,N_43980);
and U45780 (N_45780,N_43917,N_43566);
nand U45781 (N_45781,N_43436,N_43780);
nand U45782 (N_45782,N_42529,N_42455);
xor U45783 (N_45783,N_43147,N_42015);
and U45784 (N_45784,N_42397,N_43739);
nand U45785 (N_45785,N_43682,N_43059);
nor U45786 (N_45786,N_42066,N_42299);
nor U45787 (N_45787,N_42961,N_43334);
or U45788 (N_45788,N_43832,N_42912);
or U45789 (N_45789,N_43074,N_42782);
xnor U45790 (N_45790,N_43775,N_43987);
nand U45791 (N_45791,N_42502,N_42030);
nor U45792 (N_45792,N_43025,N_43571);
nor U45793 (N_45793,N_43097,N_43026);
or U45794 (N_45794,N_42243,N_42654);
or U45795 (N_45795,N_43685,N_43491);
nor U45796 (N_45796,N_42639,N_43660);
and U45797 (N_45797,N_42108,N_42242);
and U45798 (N_45798,N_43896,N_42769);
xor U45799 (N_45799,N_43139,N_43543);
and U45800 (N_45800,N_43905,N_42043);
nor U45801 (N_45801,N_43697,N_42097);
or U45802 (N_45802,N_42002,N_42870);
xor U45803 (N_45803,N_43174,N_42487);
nand U45804 (N_45804,N_43630,N_43556);
nor U45805 (N_45805,N_43421,N_43973);
or U45806 (N_45806,N_42255,N_42912);
or U45807 (N_45807,N_43575,N_42372);
nor U45808 (N_45808,N_42597,N_43653);
nor U45809 (N_45809,N_43768,N_43465);
nor U45810 (N_45810,N_42531,N_43769);
nand U45811 (N_45811,N_42349,N_43484);
xnor U45812 (N_45812,N_42638,N_42733);
xor U45813 (N_45813,N_42110,N_43187);
and U45814 (N_45814,N_42533,N_42009);
or U45815 (N_45815,N_43374,N_43393);
and U45816 (N_45816,N_42471,N_42150);
xor U45817 (N_45817,N_42076,N_43714);
and U45818 (N_45818,N_43611,N_42569);
nor U45819 (N_45819,N_43261,N_43205);
nor U45820 (N_45820,N_43886,N_43393);
xnor U45821 (N_45821,N_42581,N_42215);
nor U45822 (N_45822,N_43052,N_43140);
nor U45823 (N_45823,N_43901,N_43306);
nand U45824 (N_45824,N_43397,N_42551);
and U45825 (N_45825,N_43627,N_42045);
and U45826 (N_45826,N_43675,N_42355);
or U45827 (N_45827,N_43432,N_42966);
nor U45828 (N_45828,N_43135,N_42460);
nand U45829 (N_45829,N_43653,N_42238);
nand U45830 (N_45830,N_43180,N_42154);
xor U45831 (N_45831,N_42030,N_42962);
and U45832 (N_45832,N_43548,N_43137);
or U45833 (N_45833,N_42706,N_43947);
nand U45834 (N_45834,N_43767,N_42211);
and U45835 (N_45835,N_43724,N_42420);
nor U45836 (N_45836,N_43110,N_42860);
or U45837 (N_45837,N_42592,N_42787);
nor U45838 (N_45838,N_43623,N_42293);
or U45839 (N_45839,N_42650,N_43337);
or U45840 (N_45840,N_43071,N_42818);
nor U45841 (N_45841,N_42016,N_43258);
and U45842 (N_45842,N_43947,N_42688);
xor U45843 (N_45843,N_42110,N_42146);
xor U45844 (N_45844,N_43600,N_42154);
nand U45845 (N_45845,N_43755,N_43544);
nor U45846 (N_45846,N_43873,N_43631);
nand U45847 (N_45847,N_42713,N_42952);
xor U45848 (N_45848,N_42471,N_43557);
xnor U45849 (N_45849,N_43107,N_42307);
nand U45850 (N_45850,N_42700,N_42366);
nor U45851 (N_45851,N_42806,N_43078);
and U45852 (N_45852,N_43028,N_42968);
xnor U45853 (N_45853,N_42142,N_42181);
nand U45854 (N_45854,N_42473,N_43045);
nor U45855 (N_45855,N_42927,N_42770);
or U45856 (N_45856,N_43494,N_42338);
or U45857 (N_45857,N_42290,N_42486);
and U45858 (N_45858,N_43502,N_43352);
xor U45859 (N_45859,N_42011,N_43431);
nor U45860 (N_45860,N_42306,N_42769);
nand U45861 (N_45861,N_43980,N_43832);
nor U45862 (N_45862,N_42359,N_42706);
nand U45863 (N_45863,N_42322,N_43886);
xnor U45864 (N_45864,N_43023,N_42528);
or U45865 (N_45865,N_42105,N_43203);
nor U45866 (N_45866,N_42290,N_43937);
nand U45867 (N_45867,N_43079,N_42348);
or U45868 (N_45868,N_42005,N_43411);
nor U45869 (N_45869,N_43871,N_42488);
nor U45870 (N_45870,N_43757,N_43523);
nor U45871 (N_45871,N_42980,N_43549);
nand U45872 (N_45872,N_42084,N_43100);
or U45873 (N_45873,N_43716,N_43779);
nand U45874 (N_45874,N_42379,N_42899);
nand U45875 (N_45875,N_42005,N_42818);
nand U45876 (N_45876,N_42645,N_43300);
xnor U45877 (N_45877,N_43755,N_42093);
xnor U45878 (N_45878,N_43028,N_42749);
nand U45879 (N_45879,N_42763,N_42792);
or U45880 (N_45880,N_43446,N_43552);
nand U45881 (N_45881,N_42253,N_43538);
and U45882 (N_45882,N_43034,N_42612);
nand U45883 (N_45883,N_43819,N_43980);
or U45884 (N_45884,N_43421,N_42914);
and U45885 (N_45885,N_43380,N_43347);
xor U45886 (N_45886,N_42423,N_42784);
xnor U45887 (N_45887,N_43378,N_42904);
nand U45888 (N_45888,N_42744,N_42234);
or U45889 (N_45889,N_43877,N_43039);
and U45890 (N_45890,N_42673,N_43166);
nand U45891 (N_45891,N_43675,N_43011);
or U45892 (N_45892,N_43080,N_42917);
nor U45893 (N_45893,N_43048,N_43597);
xor U45894 (N_45894,N_42061,N_43693);
or U45895 (N_45895,N_43947,N_43986);
nor U45896 (N_45896,N_42932,N_43321);
nand U45897 (N_45897,N_43012,N_43219);
nor U45898 (N_45898,N_42450,N_42872);
xor U45899 (N_45899,N_43234,N_42537);
or U45900 (N_45900,N_43531,N_42443);
and U45901 (N_45901,N_43993,N_43686);
or U45902 (N_45902,N_42155,N_42425);
or U45903 (N_45903,N_42035,N_42528);
and U45904 (N_45904,N_42209,N_42655);
or U45905 (N_45905,N_43287,N_42527);
and U45906 (N_45906,N_42807,N_43488);
or U45907 (N_45907,N_43668,N_43869);
nor U45908 (N_45908,N_43286,N_42866);
nand U45909 (N_45909,N_43731,N_43979);
xor U45910 (N_45910,N_43591,N_42341);
nor U45911 (N_45911,N_43167,N_43550);
nor U45912 (N_45912,N_43566,N_43657);
nand U45913 (N_45913,N_43404,N_42485);
and U45914 (N_45914,N_42631,N_43271);
or U45915 (N_45915,N_42689,N_43244);
or U45916 (N_45916,N_42490,N_42012);
nor U45917 (N_45917,N_43868,N_43588);
and U45918 (N_45918,N_43671,N_43989);
xnor U45919 (N_45919,N_43869,N_43378);
nand U45920 (N_45920,N_42409,N_43896);
or U45921 (N_45921,N_42208,N_43060);
nand U45922 (N_45922,N_42722,N_43136);
nand U45923 (N_45923,N_43099,N_42528);
nor U45924 (N_45924,N_43543,N_42186);
nand U45925 (N_45925,N_42292,N_42257);
or U45926 (N_45926,N_43630,N_43961);
nand U45927 (N_45927,N_43503,N_43972);
or U45928 (N_45928,N_42830,N_42059);
nand U45929 (N_45929,N_42156,N_43149);
xnor U45930 (N_45930,N_42901,N_43612);
xnor U45931 (N_45931,N_43789,N_42088);
or U45932 (N_45932,N_43805,N_43857);
nor U45933 (N_45933,N_43429,N_42484);
or U45934 (N_45934,N_43557,N_42196);
nor U45935 (N_45935,N_42784,N_42890);
nand U45936 (N_45936,N_43222,N_43396);
or U45937 (N_45937,N_42000,N_42777);
and U45938 (N_45938,N_43391,N_43870);
and U45939 (N_45939,N_43883,N_43432);
nor U45940 (N_45940,N_43832,N_43487);
nor U45941 (N_45941,N_42500,N_43656);
and U45942 (N_45942,N_42168,N_42214);
or U45943 (N_45943,N_43826,N_43673);
nand U45944 (N_45944,N_42570,N_43031);
and U45945 (N_45945,N_42668,N_42816);
or U45946 (N_45946,N_42725,N_42182);
nor U45947 (N_45947,N_43951,N_43338);
or U45948 (N_45948,N_42012,N_43854);
nand U45949 (N_45949,N_43727,N_43932);
or U45950 (N_45950,N_43786,N_42497);
nand U45951 (N_45951,N_43391,N_42592);
nor U45952 (N_45952,N_43341,N_42993);
nand U45953 (N_45953,N_43233,N_42471);
nor U45954 (N_45954,N_43512,N_43909);
or U45955 (N_45955,N_43307,N_43194);
xnor U45956 (N_45956,N_43693,N_42498);
nand U45957 (N_45957,N_43270,N_43768);
nand U45958 (N_45958,N_42490,N_43959);
and U45959 (N_45959,N_42611,N_42357);
xnor U45960 (N_45960,N_43383,N_43341);
xor U45961 (N_45961,N_43211,N_43838);
or U45962 (N_45962,N_43118,N_42227);
and U45963 (N_45963,N_43481,N_43503);
nand U45964 (N_45964,N_43328,N_42056);
or U45965 (N_45965,N_42020,N_43422);
xor U45966 (N_45966,N_43158,N_42997);
and U45967 (N_45967,N_43594,N_43856);
xor U45968 (N_45968,N_43311,N_42858);
nand U45969 (N_45969,N_43156,N_43116);
or U45970 (N_45970,N_42903,N_43628);
nor U45971 (N_45971,N_42744,N_43306);
or U45972 (N_45972,N_43789,N_43553);
or U45973 (N_45973,N_42837,N_42893);
nor U45974 (N_45974,N_43416,N_42906);
or U45975 (N_45975,N_43318,N_42537);
xor U45976 (N_45976,N_42416,N_43659);
and U45977 (N_45977,N_43882,N_43343);
and U45978 (N_45978,N_42669,N_43872);
and U45979 (N_45979,N_42074,N_42921);
xnor U45980 (N_45980,N_42335,N_43433);
nor U45981 (N_45981,N_43213,N_43620);
nor U45982 (N_45982,N_42115,N_42983);
or U45983 (N_45983,N_43848,N_42180);
or U45984 (N_45984,N_43848,N_42514);
xnor U45985 (N_45985,N_43526,N_42746);
and U45986 (N_45986,N_42122,N_42199);
nor U45987 (N_45987,N_43871,N_42111);
and U45988 (N_45988,N_43016,N_42785);
and U45989 (N_45989,N_42255,N_42885);
nand U45990 (N_45990,N_42522,N_43460);
xnor U45991 (N_45991,N_42889,N_42042);
and U45992 (N_45992,N_42273,N_43060);
nor U45993 (N_45993,N_42888,N_42407);
xor U45994 (N_45994,N_43892,N_42816);
nor U45995 (N_45995,N_42747,N_43646);
nand U45996 (N_45996,N_43445,N_43943);
or U45997 (N_45997,N_43110,N_43951);
or U45998 (N_45998,N_43471,N_43948);
or U45999 (N_45999,N_43907,N_43475);
xnor U46000 (N_46000,N_44135,N_45374);
xor U46001 (N_46001,N_45214,N_44763);
or U46002 (N_46002,N_45538,N_45697);
and U46003 (N_46003,N_44397,N_44557);
nor U46004 (N_46004,N_45689,N_44857);
nor U46005 (N_46005,N_45714,N_45163);
nor U46006 (N_46006,N_44113,N_44509);
and U46007 (N_46007,N_45941,N_44726);
and U46008 (N_46008,N_44388,N_44988);
nand U46009 (N_46009,N_45099,N_45720);
xnor U46010 (N_46010,N_45742,N_44665);
and U46011 (N_46011,N_44972,N_45853);
nor U46012 (N_46012,N_45082,N_44915);
nor U46013 (N_46013,N_45023,N_45961);
nor U46014 (N_46014,N_45121,N_44204);
or U46015 (N_46015,N_44682,N_45037);
nor U46016 (N_46016,N_45621,N_44872);
nand U46017 (N_46017,N_45244,N_44712);
and U46018 (N_46018,N_45314,N_44986);
nor U46019 (N_46019,N_44463,N_44057);
xnor U46020 (N_46020,N_44883,N_45945);
nand U46021 (N_46021,N_44183,N_45187);
xnor U46022 (N_46022,N_44875,N_45827);
nand U46023 (N_46023,N_44950,N_45886);
nand U46024 (N_46024,N_45691,N_45390);
or U46025 (N_46025,N_44770,N_45957);
and U46026 (N_46026,N_45043,N_44862);
xor U46027 (N_46027,N_44871,N_44010);
nand U46028 (N_46028,N_44394,N_44497);
or U46029 (N_46029,N_45539,N_44744);
nand U46030 (N_46030,N_44107,N_44534);
nand U46031 (N_46031,N_45597,N_44808);
nor U46032 (N_46032,N_45553,N_45052);
nand U46033 (N_46033,N_45094,N_44533);
or U46034 (N_46034,N_44620,N_44047);
and U46035 (N_46035,N_44052,N_45382);
or U46036 (N_46036,N_44468,N_44622);
nand U46037 (N_46037,N_45171,N_44322);
and U46038 (N_46038,N_44079,N_45372);
and U46039 (N_46039,N_44266,N_44541);
nor U46040 (N_46040,N_44009,N_45457);
nand U46041 (N_46041,N_45406,N_44191);
or U46042 (N_46042,N_44237,N_44403);
and U46043 (N_46043,N_45350,N_44980);
or U46044 (N_46044,N_45473,N_44589);
nor U46045 (N_46045,N_44663,N_44318);
xor U46046 (N_46046,N_45563,N_44908);
xor U46047 (N_46047,N_44676,N_44678);
or U46048 (N_46048,N_44898,N_45832);
or U46049 (N_46049,N_45748,N_44299);
nand U46050 (N_46050,N_44870,N_45152);
xor U46051 (N_46051,N_44496,N_45825);
nor U46052 (N_46052,N_45859,N_44874);
nor U46053 (N_46053,N_45062,N_44361);
or U46054 (N_46054,N_44615,N_45786);
or U46055 (N_46055,N_45041,N_45826);
nor U46056 (N_46056,N_45419,N_45070);
nor U46057 (N_46057,N_45633,N_44163);
xor U46058 (N_46058,N_44903,N_45366);
nand U46059 (N_46059,N_44005,N_45225);
xnor U46060 (N_46060,N_45224,N_44034);
or U46061 (N_46061,N_44947,N_44918);
or U46062 (N_46062,N_45236,N_44913);
xnor U46063 (N_46063,N_45282,N_45210);
xor U46064 (N_46064,N_44020,N_44181);
and U46065 (N_46065,N_44085,N_44131);
nor U46066 (N_46066,N_44768,N_44041);
nand U46067 (N_46067,N_44840,N_44490);
nor U46068 (N_46068,N_45974,N_44152);
or U46069 (N_46069,N_44006,N_45617);
nor U46070 (N_46070,N_44088,N_45493);
or U46071 (N_46071,N_44687,N_45164);
xor U46072 (N_46072,N_45324,N_45577);
nand U46073 (N_46073,N_45085,N_44619);
and U46074 (N_46074,N_45892,N_44485);
nand U46075 (N_46075,N_44479,N_44143);
and U46076 (N_46076,N_45531,N_44441);
or U46077 (N_46077,N_44545,N_45894);
and U46078 (N_46078,N_45663,N_44424);
nor U46079 (N_46079,N_44936,N_44758);
nand U46080 (N_46080,N_45294,N_45959);
xor U46081 (N_46081,N_45669,N_44562);
nor U46082 (N_46082,N_45556,N_44836);
and U46083 (N_46083,N_44944,N_45025);
xnor U46084 (N_46084,N_44911,N_44314);
and U46085 (N_46085,N_45927,N_45769);
and U46086 (N_46086,N_44084,N_45931);
xnor U46087 (N_46087,N_44724,N_45511);
or U46088 (N_46088,N_45205,N_44411);
and U46089 (N_46089,N_45463,N_45309);
xor U46090 (N_46090,N_45862,N_44408);
and U46091 (N_46091,N_45650,N_45370);
nor U46092 (N_46092,N_44607,N_44218);
or U46093 (N_46093,N_45346,N_44339);
and U46094 (N_46094,N_45271,N_45734);
nor U46095 (N_46095,N_44037,N_44332);
and U46096 (N_46096,N_45492,N_45222);
and U46097 (N_46097,N_45676,N_44654);
nor U46098 (N_46098,N_44952,N_44605);
or U46099 (N_46099,N_45719,N_45943);
xnor U46100 (N_46100,N_44777,N_44550);
nand U46101 (N_46101,N_44839,N_44074);
and U46102 (N_46102,N_45740,N_45264);
or U46103 (N_46103,N_45836,N_45280);
nand U46104 (N_46104,N_44112,N_45807);
xor U46105 (N_46105,N_44159,N_44737);
and U46106 (N_46106,N_44285,N_45606);
nor U46107 (N_46107,N_44505,N_45850);
xnor U46108 (N_46108,N_45747,N_44951);
and U46109 (N_46109,N_44161,N_45662);
or U46110 (N_46110,N_45149,N_44896);
and U46111 (N_46111,N_44157,N_44506);
nand U46112 (N_46112,N_44308,N_44454);
nor U46113 (N_46113,N_45129,N_45991);
xnor U46114 (N_46114,N_45332,N_44273);
nand U46115 (N_46115,N_44484,N_45865);
xnor U46116 (N_46116,N_44739,N_44795);
or U46117 (N_46117,N_45487,N_44070);
or U46118 (N_46118,N_44643,N_44141);
or U46119 (N_46119,N_45933,N_45458);
and U46120 (N_46120,N_44150,N_44588);
nand U46121 (N_46121,N_45453,N_44887);
xor U46122 (N_46122,N_44234,N_44595);
and U46123 (N_46123,N_44969,N_44032);
nor U46124 (N_46124,N_44312,N_44548);
or U46125 (N_46125,N_44031,N_45202);
or U46126 (N_46126,N_44279,N_45508);
or U46127 (N_46127,N_44306,N_45576);
nand U46128 (N_46128,N_45460,N_45808);
nand U46129 (N_46129,N_44766,N_44476);
and U46130 (N_46130,N_44679,N_44136);
xor U46131 (N_46131,N_44478,N_44120);
or U46132 (N_46132,N_45920,N_44649);
nand U46133 (N_46133,N_44783,N_45188);
xnor U46134 (N_46134,N_45535,N_44169);
nor U46135 (N_46135,N_45316,N_45976);
xnor U46136 (N_46136,N_45201,N_45980);
or U46137 (N_46137,N_45495,N_45821);
or U46138 (N_46138,N_45569,N_45496);
xnor U46139 (N_46139,N_45966,N_45878);
nand U46140 (N_46140,N_44193,N_44945);
nand U46141 (N_46141,N_45422,N_45902);
nand U46142 (N_46142,N_44501,N_44603);
nand U46143 (N_46143,N_45359,N_44330);
nand U46144 (N_46144,N_44417,N_44221);
xnor U46145 (N_46145,N_44699,N_44069);
xnor U46146 (N_46146,N_44097,N_45756);
or U46147 (N_46147,N_44636,N_44166);
and U46148 (N_46148,N_44559,N_44801);
nor U46149 (N_46149,N_45263,N_44924);
nand U46150 (N_46150,N_44053,N_45512);
xnor U46151 (N_46151,N_44717,N_45051);
or U46152 (N_46152,N_45660,N_45634);
nand U46153 (N_46153,N_45186,N_44540);
nor U46154 (N_46154,N_45643,N_44953);
and U46155 (N_46155,N_45770,N_44943);
and U46156 (N_46156,N_45628,N_45695);
or U46157 (N_46157,N_45234,N_44511);
and U46158 (N_46158,N_44657,N_45678);
nor U46159 (N_46159,N_44409,N_44902);
or U46160 (N_46160,N_45701,N_44613);
or U46161 (N_46161,N_44334,N_44216);
xor U46162 (N_46162,N_45404,N_45958);
or U46163 (N_46163,N_45513,N_45746);
nand U46164 (N_46164,N_45640,N_45603);
xnor U46165 (N_46165,N_44384,N_44797);
nor U46166 (N_46166,N_45955,N_45226);
nand U46167 (N_46167,N_44232,N_44873);
and U46168 (N_46168,N_45532,N_44283);
xnor U46169 (N_46169,N_45415,N_44743);
and U46170 (N_46170,N_45433,N_44223);
nor U46171 (N_46171,N_44055,N_45609);
nand U46172 (N_46172,N_44539,N_45174);
xnor U46173 (N_46173,N_45279,N_44922);
and U46174 (N_46174,N_45743,N_45065);
nand U46175 (N_46175,N_44342,N_44442);
xor U46176 (N_46176,N_45593,N_44729);
nand U46177 (N_46177,N_44775,N_44133);
xor U46178 (N_46178,N_44486,N_45083);
nand U46179 (N_46179,N_44503,N_45349);
and U46180 (N_46180,N_45856,N_44247);
nand U46181 (N_46181,N_45774,N_44933);
nor U46182 (N_46182,N_45954,N_45586);
or U46183 (N_46183,N_44522,N_44660);
nor U46184 (N_46184,N_44741,N_45622);
and U46185 (N_46185,N_44610,N_44267);
nand U46186 (N_46186,N_45694,N_44985);
and U46187 (N_46187,N_45510,N_44659);
or U46188 (N_46188,N_44211,N_44023);
or U46189 (N_46189,N_44348,N_44290);
nand U46190 (N_46190,N_44740,N_44959);
nor U46191 (N_46191,N_45292,N_44907);
and U46192 (N_46192,N_45520,N_45269);
nor U46193 (N_46193,N_44720,N_45339);
nor U46194 (N_46194,N_45034,N_45962);
nor U46195 (N_46195,N_44859,N_45753);
and U46196 (N_46196,N_45078,N_45028);
and U46197 (N_46197,N_44570,N_45930);
or U46198 (N_46198,N_44086,N_44481);
nand U46199 (N_46199,N_45792,N_44482);
and U46200 (N_46200,N_45968,N_45267);
nand U46201 (N_46201,N_45744,N_45494);
xor U46202 (N_46202,N_44921,N_45548);
nor U46203 (N_46203,N_44272,N_45373);
and U46204 (N_46204,N_44528,N_45076);
xnor U46205 (N_46205,N_44822,N_45053);
xnor U46206 (N_46206,N_45820,N_44329);
or U46207 (N_46207,N_45286,N_44058);
and U46208 (N_46208,N_45448,N_45542);
and U46209 (N_46209,N_45754,N_45154);
or U46210 (N_46210,N_45815,N_45302);
and U46211 (N_46211,N_44958,N_45388);
and U46212 (N_46212,N_44674,N_45138);
xor U46213 (N_46213,N_44640,N_44270);
xor U46214 (N_46214,N_45275,N_45858);
and U46215 (N_46215,N_45912,N_44168);
or U46216 (N_46216,N_44456,N_44328);
nor U46217 (N_46217,N_44300,N_45241);
and U46218 (N_46218,N_44920,N_44251);
and U46219 (N_46219,N_44868,N_44160);
and U46220 (N_46220,N_45331,N_45323);
and U46221 (N_46221,N_45408,N_44154);
nor U46222 (N_46222,N_44071,N_44721);
and U46223 (N_46223,N_44170,N_45905);
nand U46224 (N_46224,N_45762,N_45342);
nand U46225 (N_46225,N_45001,N_44791);
nor U46226 (N_46226,N_45502,N_45247);
nor U46227 (N_46227,N_44225,N_44530);
and U46228 (N_46228,N_44851,N_44416);
nand U46229 (N_46229,N_45897,N_44618);
nand U46230 (N_46230,N_44782,N_44723);
or U46231 (N_46231,N_44434,N_45861);
nand U46232 (N_46232,N_44208,N_45300);
or U46233 (N_46233,N_45805,N_45117);
or U46234 (N_46234,N_44414,N_45570);
xor U46235 (N_46235,N_44672,N_45984);
nor U46236 (N_46236,N_44294,N_45200);
nand U46237 (N_46237,N_45871,N_45467);
and U46238 (N_46238,N_44087,N_44437);
or U46239 (N_46239,N_44310,N_44098);
or U46240 (N_46240,N_45822,N_45946);
nand U46241 (N_46241,N_45904,N_44100);
and U46242 (N_46242,N_45184,N_44536);
and U46243 (N_46243,N_45107,N_44241);
nor U46244 (N_46244,N_44359,N_44419);
nand U46245 (N_46245,N_45327,N_44016);
nand U46246 (N_46246,N_44799,N_44994);
and U46247 (N_46247,N_45291,N_45360);
and U46248 (N_46248,N_45900,N_44623);
xnor U46249 (N_46249,N_44828,N_44563);
and U46250 (N_46250,N_45898,N_44675);
or U46251 (N_46251,N_45153,N_45155);
nor U46252 (N_46252,N_44718,N_44923);
nor U46253 (N_46253,N_44691,N_45591);
or U46254 (N_46254,N_44658,N_45702);
nand U46255 (N_46255,N_44428,N_45838);
or U46256 (N_46256,N_45290,N_44527);
nand U46257 (N_46257,N_45104,N_44807);
and U46258 (N_46258,N_45345,N_45722);
or U46259 (N_46259,N_45673,N_45518);
or U46260 (N_46260,N_44116,N_44909);
nand U46261 (N_46261,N_45347,N_44398);
and U46262 (N_46262,N_45783,N_45208);
or U46263 (N_46263,N_45427,N_45883);
nor U46264 (N_46264,N_44171,N_45935);
and U46265 (N_46265,N_45568,N_44044);
and U46266 (N_46266,N_44917,N_44313);
nor U46267 (N_46267,N_44608,N_45560);
or U46268 (N_46268,N_45238,N_44022);
xnor U46269 (N_46269,N_45914,N_45340);
nand U46270 (N_46270,N_45687,N_44750);
nand U46271 (N_46271,N_44700,N_45006);
xnor U46272 (N_46272,N_44573,N_45891);
nand U46273 (N_46273,N_44982,N_44002);
and U46274 (N_46274,N_44863,N_45150);
nor U46275 (N_46275,N_45533,N_45489);
xnor U46276 (N_46276,N_45110,N_45320);
or U46277 (N_46277,N_45135,N_44080);
nor U46278 (N_46278,N_45004,N_44549);
nand U46279 (N_46279,N_44473,N_45362);
nand U46280 (N_46280,N_44593,N_44582);
or U46281 (N_46281,N_44867,N_45075);
nor U46282 (N_46282,N_45194,N_45266);
xnor U46283 (N_46283,N_44803,N_45369);
or U46284 (N_46284,N_45212,N_45377);
or U46285 (N_46285,N_45637,N_45343);
xor U46286 (N_46286,N_45937,N_45461);
or U46287 (N_46287,N_44488,N_45018);
nand U46288 (N_46288,N_45218,N_45315);
xnor U46289 (N_46289,N_45679,N_44324);
or U46290 (N_46290,N_44819,N_45887);
and U46291 (N_46291,N_44829,N_44612);
or U46292 (N_46292,N_45172,N_45215);
xnor U46293 (N_46293,N_45585,N_45772);
nor U46294 (N_46294,N_45398,N_44462);
nor U46295 (N_46295,N_45501,N_44302);
xnor U46296 (N_46296,N_44004,N_45969);
nand U46297 (N_46297,N_44440,N_45718);
and U46298 (N_46298,N_44716,N_44860);
xnor U46299 (N_46299,N_44537,N_44435);
xnor U46300 (N_46300,N_44039,N_44470);
xor U46301 (N_46301,N_44402,N_45181);
xor U46302 (N_46302,N_45704,N_44229);
and U46303 (N_46303,N_45009,N_45642);
nand U46304 (N_46304,N_45242,N_45007);
nor U46305 (N_46305,N_45964,N_45465);
or U46306 (N_46306,N_44200,N_44964);
or U46307 (N_46307,N_44759,N_45411);
nand U46308 (N_46308,N_45823,N_44275);
or U46309 (N_46309,N_44063,N_44162);
or U46310 (N_46310,N_44110,N_44260);
nand U46311 (N_46311,N_45651,N_44962);
or U46312 (N_46312,N_45040,N_44629);
or U46313 (N_46313,N_45375,N_45909);
nor U46314 (N_46314,N_45896,N_44628);
nor U46315 (N_46315,N_45947,N_44802);
nor U46316 (N_46316,N_44927,N_44786);
nor U46317 (N_46317,N_44710,N_44790);
nor U46318 (N_46318,N_44752,N_45641);
and U46319 (N_46319,N_44206,N_45063);
or U46320 (N_46320,N_45466,N_44987);
xor U46321 (N_46321,N_45574,N_44895);
and U46322 (N_46322,N_45700,N_45627);
or U46323 (N_46323,N_45341,N_45417);
nand U46324 (N_46324,N_45013,N_45594);
nand U46325 (N_46325,N_45992,N_44841);
or U46326 (N_46326,N_44578,N_45519);
nand U46327 (N_46327,N_45470,N_45889);
nor U46328 (N_46328,N_45793,N_45401);
and U46329 (N_46329,N_44554,N_44568);
xnor U46330 (N_46330,N_44126,N_45449);
and U46331 (N_46331,N_44114,N_45221);
or U46332 (N_46332,N_44469,N_45410);
nor U46333 (N_46333,N_44475,N_45491);
nand U46334 (N_46334,N_44349,N_45298);
and U46335 (N_46335,N_44391,N_44467);
and U46336 (N_46336,N_45400,N_45630);
and U46337 (N_46337,N_44970,N_44850);
xnor U46338 (N_46338,N_44714,N_45088);
nor U46339 (N_46339,N_44794,N_45472);
nor U46340 (N_46340,N_44626,N_44543);
nor U46341 (N_46341,N_45777,N_45177);
nand U46342 (N_46342,N_45682,N_45840);
or U46343 (N_46343,N_44246,N_44600);
nor U46344 (N_46344,N_44708,N_44066);
xnor U46345 (N_46345,N_45189,N_44552);
or U46346 (N_46346,N_44728,N_45423);
nor U46347 (N_46347,N_44878,N_44180);
nor U46348 (N_46348,N_45624,N_45002);
or U46349 (N_46349,N_44585,N_44938);
nand U46350 (N_46350,N_44239,N_44771);
nor U46351 (N_46351,N_44753,N_45197);
nor U46352 (N_46352,N_44974,N_44912);
nand U46353 (N_46353,N_45060,N_44774);
xor U46354 (N_46354,N_45635,N_45103);
and U46355 (N_46355,N_44577,N_45612);
nor U46356 (N_46356,N_45297,N_45301);
nor U46357 (N_46357,N_44195,N_44443);
and U46358 (N_46358,N_45058,N_44689);
nor U46359 (N_46359,N_44189,N_45385);
nand U46360 (N_46360,N_44880,N_44781);
or U46361 (N_46361,N_44445,N_44635);
nand U46362 (N_46362,N_44624,N_44215);
xor U46363 (N_46363,N_44321,N_45745);
nand U46364 (N_46364,N_44104,N_45333);
xor U46365 (N_46365,N_45045,N_44683);
nor U46366 (N_46366,N_45686,N_44495);
nand U46367 (N_46367,N_44033,N_45581);
nand U46368 (N_46368,N_44356,N_45668);
nand U46369 (N_46369,N_44115,N_45273);
nor U46370 (N_46370,N_45038,N_45875);
nor U46371 (N_46371,N_44165,N_44413);
nor U46372 (N_46372,N_44081,N_45287);
xor U46373 (N_46373,N_45183,N_45477);
or U46374 (N_46374,N_45050,N_45371);
nand U46375 (N_46375,N_44590,N_45671);
nor U46376 (N_46376,N_45599,N_45313);
nor U46377 (N_46377,N_44351,N_44655);
xnor U46378 (N_46378,N_45995,N_44210);
or U46379 (N_46379,N_44276,N_44638);
and U46380 (N_46380,N_45386,N_45381);
nor U46381 (N_46381,N_44845,N_45357);
or U46382 (N_46382,N_44190,N_44282);
xor U46383 (N_46383,N_44788,N_44499);
or U46384 (N_46384,N_44957,N_44778);
xor U46385 (N_46385,N_45860,N_44664);
xor U46386 (N_46386,N_45717,N_45384);
and U46387 (N_46387,N_44932,N_44274);
and U46388 (N_46388,N_45451,N_44949);
xnor U46389 (N_46389,N_45317,N_44438);
nor U46390 (N_46390,N_45596,N_45337);
or U46391 (N_46391,N_44265,N_44426);
nor U46392 (N_46392,N_44137,N_44231);
nand U46393 (N_46393,N_45924,N_44401);
nor U46394 (N_46394,N_44854,N_44119);
nand U46395 (N_46395,N_44754,N_45546);
xor U46396 (N_46396,N_45140,N_45464);
or U46397 (N_46397,N_45178,N_44560);
nor U46398 (N_46398,N_45391,N_44681);
nor U46399 (N_46399,N_44914,N_45664);
xnor U46400 (N_46400,N_45182,N_45054);
nor U46401 (N_46401,N_44331,N_45849);
nand U46402 (N_46402,N_44571,N_45265);
nor U46403 (N_46403,N_45874,N_44027);
nor U46404 (N_46404,N_45893,N_44931);
xor U46405 (N_46405,N_44993,N_44036);
xor U46406 (N_46406,N_45289,N_45737);
nand U46407 (N_46407,N_45270,N_45550);
nor U46408 (N_46408,N_44926,N_44466);
or U46409 (N_46409,N_45245,N_45873);
xor U46410 (N_46410,N_45170,N_44301);
or U46411 (N_46411,N_44688,N_44965);
and U46412 (N_46412,N_44813,N_45755);
or U46413 (N_46413,N_45575,N_44500);
and U46414 (N_46414,N_44824,N_44960);
nor U46415 (N_46415,N_44392,N_45973);
nand U46416 (N_46416,N_45365,N_44971);
or U46417 (N_46417,N_44298,N_45926);
nand U46418 (N_46418,N_45979,N_45424);
or U46419 (N_46419,N_45235,N_44789);
nor U46420 (N_46420,N_44293,N_44864);
nor U46421 (N_46421,N_45476,N_44125);
and U46422 (N_46422,N_45312,N_45420);
xor U46423 (N_46423,N_44187,N_44186);
nor U46424 (N_46424,N_45814,N_45810);
and U46425 (N_46425,N_45598,N_45529);
xor U46426 (N_46426,N_45250,N_44167);
nor U46427 (N_46427,N_44142,N_45403);
nand U46428 (N_46428,N_44386,N_44706);
or U46429 (N_46429,N_44458,N_44652);
xor U46430 (N_46430,N_44519,N_44630);
or U46431 (N_46431,N_45142,N_45817);
or U46432 (N_46432,N_45975,N_45260);
nand U46433 (N_46433,N_44518,N_45851);
nor U46434 (N_46434,N_45728,N_44042);
xnor U46435 (N_46435,N_44606,N_45950);
and U46436 (N_46436,N_45207,N_44345);
xor U46437 (N_46437,N_44212,N_45151);
nor U46438 (N_46438,N_45281,N_45363);
nor U46439 (N_46439,N_45750,N_44694);
xnor U46440 (N_46440,N_44019,N_45443);
xor U46441 (N_46441,N_45852,N_45092);
nor U46442 (N_46442,N_44427,N_45899);
nor U46443 (N_46443,N_44433,N_44461);
or U46444 (N_46444,N_44399,N_44271);
and U46445 (N_46445,N_45418,N_44257);
or U46446 (N_46446,N_45126,N_45024);
or U46447 (N_46447,N_45960,N_45738);
nand U46448 (N_46448,N_44641,N_44963);
nor U46449 (N_46449,N_44217,N_44996);
and U46450 (N_46450,N_45936,N_45674);
and U46451 (N_46451,N_45394,N_44722);
and U46452 (N_46452,N_45049,N_45983);
xnor U46453 (N_46453,N_45989,N_45087);
and U46454 (N_46454,N_44051,N_45452);
and U46455 (N_46455,N_44747,N_45649);
nand U46456 (N_46456,N_45632,N_45032);
nand U46457 (N_46457,N_45779,N_44973);
nand U46458 (N_46458,N_44396,N_45921);
and U46459 (N_46459,N_44000,N_44644);
and U46460 (N_46460,N_44881,N_44444);
or U46461 (N_46461,N_45191,N_45106);
nand U46462 (N_46462,N_44684,N_44303);
xnor U46463 (N_46463,N_45086,N_44059);
nor U46464 (N_46464,N_44378,N_45499);
xor U46465 (N_46465,N_44226,N_44404);
and U46466 (N_46466,N_44637,N_44734);
nor U46467 (N_46467,N_44955,N_44227);
nor U46468 (N_46468,N_44814,N_44833);
xnor U46469 (N_46469,N_44625,N_44147);
nand U46470 (N_46470,N_44904,N_44551);
or U46471 (N_46471,N_44669,N_44925);
xnor U46472 (N_46472,N_45308,N_44385);
nand U46473 (N_46473,N_44148,N_44838);
nor U46474 (N_46474,N_44579,N_45438);
nor U46475 (N_46475,N_44288,N_45412);
xnor U46476 (N_46476,N_45967,N_44474);
nor U46477 (N_46477,N_44072,N_44291);
nand U46478 (N_46478,N_45399,N_44253);
or U46479 (N_46479,N_45407,N_44455);
or U46480 (N_46480,N_45173,N_45685);
and U46481 (N_46481,N_45667,N_45061);
nand U46482 (N_46482,N_45219,N_45030);
and U46483 (N_46483,N_45986,N_45509);
nand U46484 (N_46484,N_45102,N_44961);
nor U46485 (N_46485,N_45982,N_45435);
xor U46486 (N_46486,N_45439,N_44235);
and U46487 (N_46487,N_44352,N_44842);
or U46488 (N_46488,N_44263,N_44255);
nand U46489 (N_46489,N_44611,N_44172);
nor U46490 (N_46490,N_45798,N_44292);
or U46491 (N_46491,N_45733,N_45877);
nor U46492 (N_46492,N_45485,N_45338);
nand U46493 (N_46493,N_45732,N_44719);
xor U46494 (N_46494,N_45048,N_44363);
nand U46495 (N_46495,N_45789,N_45486);
xor U46496 (N_46496,N_44315,N_45620);
nand U46497 (N_46497,N_44151,N_45284);
and U46498 (N_46498,N_45021,N_44028);
and U46499 (N_46499,N_45652,N_44203);
nor U46500 (N_46500,N_44156,N_44192);
xor U46501 (N_46501,N_44677,N_44449);
and U46502 (N_46502,N_44531,N_45834);
and U46503 (N_46503,N_44866,N_44757);
or U46504 (N_46504,N_44939,N_45118);
nor U46505 (N_46505,N_45185,N_45578);
nand U46506 (N_46506,N_45796,N_44566);
nor U46507 (N_46507,N_45253,N_45376);
and U46508 (N_46508,N_45882,N_44800);
xnor U46509 (N_46509,N_45133,N_45758);
nand U46510 (N_46510,N_44976,N_44897);
and U46511 (N_46511,N_44093,N_45128);
and U46512 (N_46512,N_44756,N_45527);
nand U46513 (N_46513,N_44564,N_44284);
and U46514 (N_46514,N_44343,N_45305);
nand U46515 (N_46515,N_44240,N_44040);
or U46516 (N_46516,N_44806,N_45478);
or U46517 (N_46517,N_45547,N_44983);
and U46518 (N_46518,N_45444,N_45739);
xor U46519 (N_46519,N_44858,N_44410);
or U46520 (N_46520,N_44899,N_45631);
xnor U46521 (N_46521,N_44844,N_44632);
nor U46522 (N_46522,N_44375,N_45517);
nand U46523 (N_46523,N_45469,N_44893);
nand U46524 (N_46524,N_45646,N_45409);
or U46525 (N_46525,N_44553,N_44647);
xnor U46526 (N_46526,N_45657,N_45644);
and U46527 (N_46527,N_45525,N_45368);
and U46528 (N_46528,N_44121,N_44346);
and U46529 (N_46529,N_45056,N_45693);
nand U46530 (N_46530,N_44056,N_44197);
nand U46531 (N_46531,N_44614,N_44264);
and U46532 (N_46532,N_45903,N_45175);
nand U46533 (N_46533,N_45232,N_44289);
nand U46534 (N_46534,N_44111,N_45356);
xnor U46535 (N_46535,N_45097,N_45095);
or U46536 (N_46536,N_45776,N_45582);
xnor U46537 (N_46537,N_45837,N_45690);
nor U46538 (N_46538,N_45276,N_45167);
xor U46539 (N_46539,N_45616,N_45071);
and U46540 (N_46540,N_44432,N_45811);
nand U46541 (N_46541,N_44158,N_44017);
nand U46542 (N_46542,N_45067,N_45285);
xor U46543 (N_46543,N_45648,N_44507);
xor U46544 (N_46544,N_45785,N_45699);
nand U46545 (N_46545,N_44592,N_45545);
xor U46546 (N_46546,N_44262,N_45012);
and U46547 (N_46547,N_44995,N_45141);
or U46548 (N_46548,N_45680,N_44230);
nand U46549 (N_46549,N_45348,N_45240);
xor U46550 (N_46550,N_45829,N_45925);
xnor U46551 (N_46551,N_45918,N_44146);
and U46552 (N_46552,N_44024,N_44929);
or U46553 (N_46553,N_44731,N_44320);
nand U46554 (N_46554,N_45441,N_45206);
or U46555 (N_46555,N_44662,N_45146);
and U46556 (N_46556,N_45601,N_45364);
and U46557 (N_46557,N_45421,N_44556);
nand U46558 (N_46558,N_44011,N_45911);
nand U46559 (N_46559,N_44817,N_45072);
nand U46560 (N_46560,N_45551,N_44572);
or U46561 (N_46561,N_45334,N_45354);
nor U46562 (N_46562,N_45555,N_44650);
or U46563 (N_46563,N_45672,N_45254);
or U46564 (N_46564,N_45725,N_45389);
nor U46565 (N_46565,N_45572,N_45318);
xor U46566 (N_46566,N_44502,N_45119);
xor U46567 (N_46567,N_45046,N_44544);
nand U46568 (N_46568,N_45600,N_44894);
nand U46569 (N_46569,N_45778,N_44574);
nand U46570 (N_46570,N_44984,N_44835);
nor U46571 (N_46571,N_44374,N_45766);
nor U46572 (N_46572,N_44425,N_45257);
nor U46573 (N_46573,N_45447,N_45255);
nor U46574 (N_46574,N_45507,N_44576);
nor U46575 (N_46575,N_44524,N_44295);
and U46576 (N_46576,N_45405,N_44003);
xnor U46577 (N_46577,N_44884,N_44882);
or U46578 (N_46578,N_45895,N_45537);
nor U46579 (N_46579,N_45698,N_45658);
nand U46580 (N_46580,N_45352,N_45554);
nor U46581 (N_46581,N_44380,N_44892);
nand U46582 (N_46582,N_45831,N_45993);
and U46583 (N_46583,N_44395,N_45251);
nand U46584 (N_46584,N_44287,N_44709);
nor U46585 (N_46585,N_44450,N_44335);
and U46586 (N_46586,N_45521,N_45870);
or U46587 (N_46587,N_45145,N_44105);
xor U46588 (N_46588,N_44992,N_44853);
or U46589 (N_46589,N_45736,N_45806);
nand U46590 (N_46590,N_44280,N_45784);
xnor U46591 (N_46591,N_45951,N_44693);
and U46592 (N_46592,N_45797,N_45198);
xnor U46593 (N_46593,N_45474,N_45397);
xor U46594 (N_46594,N_44068,N_44268);
nand U46595 (N_46595,N_44372,N_44304);
nand U46596 (N_46596,N_45116,N_44307);
xnor U46597 (N_46597,N_45064,N_44847);
and U46598 (N_46598,N_44812,N_45763);
and U46599 (N_46599,N_45353,N_44516);
nor U46600 (N_46600,N_45351,N_44935);
nor U46601 (N_46601,N_44062,N_44843);
and U46602 (N_46602,N_45812,N_44823);
nand U46603 (N_46603,N_44178,N_45130);
and U46604 (N_46604,N_44376,N_45761);
and U46605 (N_46605,N_44686,N_45454);
or U46606 (N_46606,N_45425,N_44406);
nand U46607 (N_46607,N_45080,N_44018);
nand U46608 (N_46608,N_44326,N_45835);
xor U46609 (N_46609,N_45217,N_45272);
nand U46610 (N_46610,N_45213,N_45842);
nor U46611 (N_46611,N_44793,N_45209);
nand U46612 (N_46612,N_45055,N_44742);
or U46613 (N_46613,N_45000,N_44222);
and U46614 (N_46614,N_44928,N_45735);
or U46615 (N_46615,N_44008,N_45923);
nor U46616 (N_46616,N_45246,N_45203);
nor U46617 (N_46617,N_45115,N_44670);
xnor U46618 (N_46618,N_44617,N_45869);
nor U46619 (N_46619,N_44480,N_44692);
or U46620 (N_46620,N_44095,N_44007);
nand U46621 (N_46621,N_44364,N_45136);
nor U46622 (N_46622,N_45432,N_44736);
or U46623 (N_46623,N_44591,N_44333);
and U46624 (N_46624,N_44666,N_44680);
and U46625 (N_46625,N_45614,N_45830);
and U46626 (N_46626,N_44368,N_44269);
nand U46627 (N_46627,N_44220,N_45876);
or U46628 (N_46628,N_45639,N_44746);
nand U46629 (N_46629,N_44277,N_45122);
xnor U46630 (N_46630,N_45019,N_44515);
or U46631 (N_46631,N_45355,N_44138);
xnor U46632 (N_46632,N_44890,N_44811);
and U46633 (N_46633,N_44244,N_45490);
and U46634 (N_46634,N_45482,N_44685);
or U46635 (N_46635,N_45319,N_44733);
nor U46636 (N_46636,N_44598,N_44575);
nand U46637 (N_46637,N_45033,N_45462);
xnor U46638 (N_46638,N_45204,N_44645);
and U46639 (N_46639,N_45500,N_44772);
nor U46640 (N_46640,N_45727,N_45752);
or U46641 (N_46641,N_45999,N_44639);
and U46642 (N_46642,N_45442,N_45330);
or U46643 (N_46643,N_44013,N_44459);
xnor U46644 (N_46644,N_44050,N_44900);
nand U46645 (N_46645,N_45402,N_44809);
nand U46646 (N_46646,N_45677,N_45166);
nand U46647 (N_46647,N_45843,N_45505);
or U46648 (N_46648,N_45994,N_45039);
nand U46649 (N_46649,N_44798,N_44785);
or U46650 (N_46650,N_45710,N_45380);
xnor U46651 (N_46651,N_45655,N_45031);
nor U46652 (N_46652,N_44583,N_44360);
nand U46653 (N_46653,N_45775,N_44948);
and U46654 (N_46654,N_45703,N_44471);
nand U46655 (N_46655,N_44014,N_44132);
and U46656 (N_46656,N_45261,N_45712);
and U46657 (N_46657,N_44096,N_45296);
and U46658 (N_46658,N_45195,N_44855);
and U46659 (N_46659,N_44997,N_45258);
nand U46660 (N_46660,N_44219,N_44642);
xor U46661 (N_46661,N_45636,N_45216);
or U46662 (N_46662,N_44705,N_44510);
and U46663 (N_46663,N_45378,N_44344);
or U46664 (N_46664,N_44730,N_44916);
xnor U46665 (N_46665,N_45647,N_44365);
or U46666 (N_46666,N_44646,N_44453);
and U46667 (N_46667,N_44094,N_44472);
nand U46668 (N_46668,N_45395,N_44587);
xnor U46669 (N_46669,N_45262,N_45864);
nor U46670 (N_46670,N_45387,N_44127);
nor U46671 (N_46671,N_45638,N_45988);
nand U46672 (N_46672,N_45716,N_44930);
nand U46673 (N_46673,N_44889,N_45977);
nor U46674 (N_46674,N_44238,N_44377);
and U46675 (N_46675,N_44383,N_45675);
xor U46676 (N_46676,N_45607,N_45611);
or U46677 (N_46677,N_45844,N_45863);
nand U46678 (N_46678,N_44370,N_45998);
nand U46679 (N_46679,N_44555,N_44586);
nand U46680 (N_46680,N_45970,N_44517);
nand U46681 (N_46681,N_45559,N_45158);
and U46682 (N_46682,N_45125,N_45430);
and U46683 (N_46683,N_44787,N_44029);
and U46684 (N_46684,N_45259,N_44532);
nand U46685 (N_46685,N_45881,N_44357);
xor U46686 (N_46686,N_45868,N_45450);
nor U46687 (N_46687,N_45583,N_44140);
and U46688 (N_46688,N_44604,N_45584);
and U46689 (N_46689,N_45344,N_44358);
and U46690 (N_46690,N_45828,N_44707);
nand U46691 (N_46691,N_45137,N_44184);
and U46692 (N_46692,N_44249,N_45307);
xnor U46693 (N_46693,N_45940,N_45692);
xnor U46694 (N_46694,N_44077,N_44735);
nor U46695 (N_46695,N_45751,N_45566);
or U46696 (N_46696,N_44538,N_45741);
and U46697 (N_46697,N_45613,N_44422);
nor U46698 (N_46698,N_44128,N_45587);
nand U46699 (N_46699,N_44337,N_45066);
xnor U46700 (N_46700,N_44174,N_44745);
and U46701 (N_46701,N_45956,N_44999);
xor U46702 (N_46702,N_44201,N_45580);
nor U46703 (N_46703,N_45764,N_44477);
nand U46704 (N_46704,N_45211,N_45456);
and U46705 (N_46705,N_45413,N_45654);
nand U46706 (N_46706,N_45483,N_44810);
xnor U46707 (N_46707,N_44245,N_45179);
nor U46708 (N_46708,N_44910,N_45625);
xor U46709 (N_46709,N_45949,N_45917);
nand U46710 (N_46710,N_45608,N_44651);
xor U46711 (N_46711,N_45922,N_44954);
or U46712 (N_46712,N_44012,N_44494);
xnor U46713 (N_46713,N_44751,N_45656);
nor U46714 (N_46714,N_44382,N_45480);
xor U46715 (N_46715,N_44108,N_45857);
nor U46716 (N_46716,N_45708,N_44861);
or U46717 (N_46717,N_45709,N_44489);
nor U46718 (N_46718,N_45096,N_44341);
and U46719 (N_46719,N_44760,N_44767);
xor U46720 (N_46720,N_44418,N_44423);
nor U46721 (N_46721,N_44015,N_45729);
and U46722 (N_46722,N_45475,N_45367);
or U46723 (N_46723,N_44305,N_45801);
xor U46724 (N_46724,N_45468,N_44565);
xor U46725 (N_46725,N_45091,N_45228);
or U46726 (N_46726,N_45972,N_44196);
or U46727 (N_46727,N_44149,N_44580);
or U46728 (N_46728,N_44256,N_44355);
and U46729 (N_46729,N_45759,N_45552);
and U46730 (N_46730,N_45928,N_45017);
xnor U46731 (N_46731,N_44317,N_45003);
xnor U46732 (N_46732,N_44837,N_45929);
nor U46733 (N_46733,N_45268,N_45997);
xnor U46734 (N_46734,N_44199,N_44431);
nor U46735 (N_46735,N_45605,N_44597);
nor U46736 (N_46736,N_45132,N_44325);
nand U46737 (N_46737,N_45256,N_45011);
nand U46738 (N_46738,N_45392,N_44956);
nor U46739 (N_46739,N_45794,N_44940);
nor U46740 (N_46740,N_44134,N_45223);
nand U46741 (N_46741,N_44493,N_44885);
or U46742 (N_46742,N_44026,N_45446);
nand U46743 (N_46743,N_45093,N_44547);
nor U46744 (N_46744,N_45721,N_44998);
and U46745 (N_46745,N_44968,N_44164);
nand U46746 (N_46746,N_44671,N_45645);
nand U46747 (N_46747,N_44129,N_45015);
nand U46748 (N_46748,N_44046,N_45782);
nand U46749 (N_46749,N_44083,N_45230);
xnor U46750 (N_46750,N_45278,N_44323);
or U46751 (N_46751,N_44701,N_45996);
xor U46752 (N_46752,N_45426,N_45787);
nor U46753 (N_46753,N_45014,N_45239);
and U46754 (N_46754,N_44073,N_44690);
xnor U46755 (N_46755,N_45180,N_44393);
and U46756 (N_46756,N_45610,N_44762);
and U46757 (N_46757,N_44173,N_45534);
and U46758 (N_46758,N_45565,N_44354);
or U46759 (N_46759,N_44001,N_44830);
xor U46760 (N_46760,N_45488,N_45229);
or U46761 (N_46761,N_44448,N_44067);
or U46762 (N_46762,N_44021,N_45978);
or U46763 (N_46763,N_44297,N_44905);
nor U46764 (N_46764,N_44048,N_44460);
or U46765 (N_46765,N_44124,N_45987);
nand U46766 (N_46766,N_45530,N_45558);
nand U46767 (N_46767,N_44103,N_44869);
nand U46768 (N_46768,N_45321,N_44436);
nand U46769 (N_46769,N_44340,N_44627);
xor U46770 (N_46770,N_45383,N_45027);
and U46771 (N_46771,N_45431,N_45090);
nor U46772 (N_46772,N_44064,N_45567);
or U46773 (N_46773,N_45653,N_44102);
nand U46774 (N_46774,N_45965,N_45953);
or U46775 (N_46775,N_44248,N_44465);
or U46776 (N_46776,N_45791,N_44233);
nor U46777 (N_46777,N_44038,N_44697);
nand U46778 (N_46778,N_45549,N_45802);
nor U46779 (N_46779,N_45176,N_44609);
xor U46780 (N_46780,N_44713,N_45564);
xor U46781 (N_46781,N_45114,N_44834);
and U46782 (N_46782,N_45059,N_45629);
or U46783 (N_46783,N_44569,N_44941);
or U46784 (N_46784,N_44525,N_45523);
xor U46785 (N_46785,N_44286,N_44153);
nand U46786 (N_46786,N_44091,N_45939);
and U46787 (N_46787,N_45073,N_45277);
nor U46788 (N_46788,N_45615,N_44919);
xor U46789 (N_46789,N_45068,N_44430);
xnor U46790 (N_46790,N_45227,N_45757);
xor U46791 (N_46791,N_45803,N_45196);
xor U46792 (N_46792,N_44089,N_44703);
nand U46793 (N_46793,N_45005,N_44827);
nand U46794 (N_46794,N_45681,N_44661);
nand U46795 (N_46795,N_45765,N_45109);
or U46796 (N_46796,N_45771,N_45618);
nand U46797 (N_46797,N_45872,N_44526);
nand U46798 (N_46798,N_44065,N_44738);
and U46799 (N_46799,N_44452,N_45790);
or U46800 (N_46800,N_44182,N_45788);
nand U46801 (N_46801,N_45839,N_45516);
nor U46802 (N_46802,N_44243,N_44601);
nand U46803 (N_46803,N_45169,N_44846);
xnor U46804 (N_46804,N_44258,N_45479);
and U46805 (N_46805,N_45022,N_44535);
nor U46806 (N_46806,N_45846,N_45026);
or U46807 (N_46807,N_45528,N_45833);
and U46808 (N_46808,N_44512,N_44373);
nand U46809 (N_46809,N_44177,N_45471);
nand U46810 (N_46810,N_45819,N_44784);
and U46811 (N_46811,N_44209,N_44621);
xnor U46812 (N_46812,N_44139,N_44732);
nor U46813 (N_46813,N_45436,N_45105);
or U46814 (N_46814,N_44888,N_45619);
and U46815 (N_46815,N_45124,N_45243);
and U46816 (N_46816,N_44748,N_44176);
nor U46817 (N_46817,N_44978,N_45901);
or U46818 (N_46818,N_45880,N_45595);
xor U46819 (N_46819,N_44420,N_45885);
nand U46820 (N_46820,N_44967,N_44698);
xnor U46821 (N_46821,N_45981,N_44906);
nand U46822 (N_46822,N_44076,N_44049);
or U46823 (N_46823,N_44099,N_45157);
or U46824 (N_46824,N_44491,N_44155);
and U46825 (N_46825,N_45147,N_45329);
and U46826 (N_46826,N_44296,N_44979);
or U46827 (N_46827,N_44749,N_44224);
and U46828 (N_46828,N_44977,N_45866);
nand U46829 (N_46829,N_44213,N_44106);
and U46830 (N_46830,N_44876,N_45526);
and U46831 (N_46831,N_45799,N_44379);
nand U46832 (N_46832,N_44558,N_45010);
and U46833 (N_46833,N_45156,N_44075);
nor U46834 (N_46834,N_45161,N_44702);
and U46835 (N_46835,N_44514,N_45544);
xnor U46836 (N_46836,N_44879,N_45768);
or U46837 (N_46837,N_45711,N_45506);
nand U46838 (N_46838,N_44371,N_44891);
xnor U46839 (N_46839,N_45306,N_45131);
nor U46840 (N_46840,N_45057,N_45325);
or U46841 (N_46841,N_44336,N_45414);
and U46842 (N_46842,N_45481,N_44122);
xor U46843 (N_46843,N_44390,N_44725);
nor U46844 (N_46844,N_44796,N_44901);
or U46845 (N_46845,N_45543,N_45809);
nand U46846 (N_46846,N_45942,N_45910);
and U46847 (N_46847,N_44508,N_44769);
xor U46848 (N_46848,N_44228,N_44369);
nand U46849 (N_46849,N_45437,N_44561);
xor U46850 (N_46850,N_44185,N_45688);
or U46851 (N_46851,N_44596,N_45162);
or U46852 (N_46852,N_45592,N_44145);
or U46853 (N_46853,N_44761,N_44205);
xor U46854 (N_46854,N_44567,N_44309);
xor U46855 (N_46855,N_45589,N_44242);
and U46856 (N_46856,N_45659,N_44523);
or U46857 (N_46857,N_44092,N_45288);
nor U46858 (N_46858,N_45336,N_44780);
xnor U46859 (N_46859,N_44381,N_44942);
and U46860 (N_46860,N_44865,N_44188);
and U46861 (N_46861,N_45042,N_45867);
nor U46862 (N_46862,N_44101,N_45938);
xnor U46863 (N_46863,N_44281,N_44877);
or U46864 (N_46864,N_45602,N_45715);
and U46865 (N_46865,N_44025,N_44804);
nor U46866 (N_46866,N_45948,N_45706);
nand U46867 (N_46867,N_44054,N_44429);
nor U46868 (N_46868,N_44175,N_44695);
or U46869 (N_46869,N_44792,N_44856);
xnor U46870 (N_46870,N_44194,N_45670);
nand U46871 (N_46871,N_45579,N_44631);
or U46872 (N_46872,N_44989,N_45089);
and U46873 (N_46873,N_44776,N_45879);
nand U46874 (N_46874,N_45252,N_45100);
nor U46875 (N_46875,N_45841,N_44389);
xnor U46876 (N_46876,N_45079,N_44130);
and U46877 (N_46877,N_45168,N_45561);
or U46878 (N_46878,N_45913,N_45074);
or U46879 (N_46879,N_45963,N_45029);
and U46880 (N_46880,N_45160,N_45726);
nand U46881 (N_46881,N_45588,N_45335);
or U46882 (N_46882,N_45934,N_44118);
nor U46883 (N_46883,N_45626,N_44937);
nor U46884 (N_46884,N_45192,N_44981);
xor U46885 (N_46885,N_45113,N_45919);
and U46886 (N_46886,N_45795,N_45445);
or U46887 (N_46887,N_45816,N_45623);
and U46888 (N_46888,N_45854,N_45190);
nand U46889 (N_46889,N_44250,N_44831);
xor U46890 (N_46890,N_44816,N_45148);
and U46891 (N_46891,N_44711,N_45522);
or U46892 (N_46892,N_44633,N_45393);
or U46893 (N_46893,N_45248,N_44765);
xnor U46894 (N_46894,N_45035,N_44815);
xnor U46895 (N_46895,N_44821,N_45661);
xor U46896 (N_46896,N_45781,N_44236);
and U46897 (N_46897,N_45036,N_44090);
xor U46898 (N_46898,N_44826,N_44198);
nor U46899 (N_46899,N_44362,N_44668);
and U46900 (N_46900,N_45193,N_44043);
xnor U46901 (N_46901,N_45731,N_45112);
nand U46902 (N_46902,N_45804,N_44773);
and U46903 (N_46903,N_45249,N_44207);
and U46904 (N_46904,N_44446,N_45081);
or U46905 (N_46905,N_45429,N_45199);
xor U46906 (N_46906,N_44634,N_44520);
nor U46907 (N_46907,N_45990,N_45684);
or U46908 (N_46908,N_45730,N_45514);
nor U46909 (N_46909,N_45666,N_45293);
or U46910 (N_46910,N_45295,N_45541);
nor U46911 (N_46911,N_45434,N_44412);
nor U46912 (N_46912,N_44673,N_45044);
nand U46913 (N_46913,N_45604,N_45139);
and U46914 (N_46914,N_44991,N_45890);
and U46915 (N_46915,N_44109,N_44082);
nand U46916 (N_46916,N_45237,N_44616);
nand U46917 (N_46917,N_44366,N_44832);
or U46918 (N_46918,N_45665,N_45760);
nor U46919 (N_46919,N_45134,N_45773);
or U46920 (N_46920,N_45127,N_45503);
or U46921 (N_46921,N_44447,N_44779);
xor U46922 (N_46922,N_44316,N_45971);
and U46923 (N_46923,N_45540,N_45707);
or U46924 (N_46924,N_44820,N_44602);
nand U46925 (N_46925,N_45705,N_44078);
nor U46926 (N_46926,N_45944,N_45515);
or U46927 (N_46927,N_44400,N_44347);
xor U46928 (N_46928,N_45952,N_44327);
nand U46929 (N_46929,N_45020,N_45274);
xor U46930 (N_46930,N_45907,N_45123);
or U46931 (N_46931,N_44990,N_44045);
nand U46932 (N_46932,N_44755,N_44849);
nor U46933 (N_46933,N_45932,N_44439);
nand U46934 (N_46934,N_45683,N_44353);
nor U46935 (N_46935,N_45428,N_45455);
or U46936 (N_46936,N_45884,N_44656);
or U46937 (N_46937,N_45855,N_44584);
nand U46938 (N_46938,N_45696,N_45985);
or U46939 (N_46939,N_44648,N_44311);
xnor U46940 (N_46940,N_44259,N_44261);
or U46941 (N_46941,N_45159,N_44594);
nor U46942 (N_46942,N_44696,N_45818);
and U46943 (N_46943,N_44704,N_45016);
xor U46944 (N_46944,N_45915,N_45299);
xor U46945 (N_46945,N_44946,N_45524);
and U46946 (N_46946,N_44030,N_45847);
xnor U46947 (N_46947,N_45848,N_44852);
nor U46948 (N_46948,N_45713,N_44487);
or U46949 (N_46949,N_45723,N_44387);
and U46950 (N_46950,N_45322,N_44504);
xor U46951 (N_46951,N_45916,N_45311);
or U46952 (N_46952,N_45767,N_45047);
or U46953 (N_46953,N_44975,N_45220);
and U46954 (N_46954,N_45231,N_44653);
xor U46955 (N_46955,N_44179,N_45165);
or U46956 (N_46956,N_44825,N_45283);
or U46957 (N_46957,N_44254,N_45361);
nand U46958 (N_46958,N_44599,N_45143);
nor U46959 (N_46959,N_44966,N_44667);
and U46960 (N_46960,N_45077,N_44035);
xnor U46961 (N_46961,N_45557,N_44405);
nand U46962 (N_46962,N_45571,N_44818);
nand U46963 (N_46963,N_45120,N_44581);
or U46964 (N_46964,N_44727,N_44457);
xor U46965 (N_46965,N_45824,N_45396);
nand U46966 (N_46966,N_44415,N_45440);
nor U46967 (N_46967,N_45108,N_45536);
or U46968 (N_46968,N_44202,N_44513);
nor U46969 (N_46969,N_44542,N_45498);
nand U46970 (N_46970,N_45358,N_45303);
nor U46971 (N_46971,N_44805,N_45144);
or U46972 (N_46972,N_44123,N_45800);
nand U46973 (N_46973,N_44214,N_44061);
xor U46974 (N_46974,N_44546,N_44886);
nor U46975 (N_46975,N_44483,N_45328);
xor U46976 (N_46976,N_45484,N_45233);
nand U46977 (N_46977,N_44764,N_45888);
and U46978 (N_46978,N_44144,N_45101);
xnor U46979 (N_46979,N_44464,N_45749);
nand U46980 (N_46980,N_45008,N_45111);
and U46981 (N_46981,N_45590,N_44252);
nand U46982 (N_46982,N_44117,N_45845);
nor U46983 (N_46983,N_44060,N_44350);
nand U46984 (N_46984,N_45084,N_45813);
nand U46985 (N_46985,N_44848,N_44421);
xor U46986 (N_46986,N_45497,N_45906);
xnor U46987 (N_46987,N_45416,N_44498);
or U46988 (N_46988,N_44278,N_44934);
xnor U46989 (N_46989,N_45310,N_44451);
xnor U46990 (N_46990,N_44715,N_45304);
and U46991 (N_46991,N_45724,N_45908);
xor U46992 (N_46992,N_45069,N_45459);
or U46993 (N_46993,N_45780,N_45573);
nor U46994 (N_46994,N_44529,N_45098);
xnor U46995 (N_46995,N_45379,N_44492);
and U46996 (N_46996,N_45326,N_44319);
nor U46997 (N_46997,N_44338,N_44521);
nor U46998 (N_46998,N_44367,N_45562);
nor U46999 (N_46999,N_44407,N_45504);
nand U47000 (N_47000,N_45856,N_44309);
and U47001 (N_47001,N_44914,N_45885);
nand U47002 (N_47002,N_44683,N_45033);
or U47003 (N_47003,N_44898,N_44759);
and U47004 (N_47004,N_45928,N_45900);
and U47005 (N_47005,N_45786,N_44233);
nand U47006 (N_47006,N_45766,N_44711);
and U47007 (N_47007,N_45879,N_45214);
nand U47008 (N_47008,N_44483,N_44149);
and U47009 (N_47009,N_45655,N_44202);
nand U47010 (N_47010,N_45980,N_45584);
nand U47011 (N_47011,N_44081,N_44970);
nand U47012 (N_47012,N_44899,N_44402);
nand U47013 (N_47013,N_45577,N_45522);
nand U47014 (N_47014,N_45329,N_44489);
nand U47015 (N_47015,N_44143,N_44042);
xnor U47016 (N_47016,N_44372,N_45983);
nor U47017 (N_47017,N_45878,N_44164);
and U47018 (N_47018,N_44944,N_44538);
or U47019 (N_47019,N_45792,N_45206);
xor U47020 (N_47020,N_44311,N_44945);
and U47021 (N_47021,N_45004,N_45447);
and U47022 (N_47022,N_45974,N_45786);
xor U47023 (N_47023,N_45290,N_44861);
or U47024 (N_47024,N_44965,N_45467);
nand U47025 (N_47025,N_44978,N_45190);
and U47026 (N_47026,N_44295,N_45434);
nor U47027 (N_47027,N_45852,N_45531);
or U47028 (N_47028,N_44688,N_45911);
and U47029 (N_47029,N_45125,N_45278);
nor U47030 (N_47030,N_45874,N_45987);
nand U47031 (N_47031,N_45053,N_44961);
nor U47032 (N_47032,N_45777,N_45478);
xor U47033 (N_47033,N_44219,N_44536);
xor U47034 (N_47034,N_44019,N_44858);
or U47035 (N_47035,N_45183,N_45502);
nand U47036 (N_47036,N_44581,N_44915);
nor U47037 (N_47037,N_45391,N_45530);
and U47038 (N_47038,N_45210,N_45843);
and U47039 (N_47039,N_45797,N_45465);
xnor U47040 (N_47040,N_45800,N_44581);
nand U47041 (N_47041,N_45193,N_45656);
and U47042 (N_47042,N_44392,N_44473);
nand U47043 (N_47043,N_44165,N_45399);
xnor U47044 (N_47044,N_44913,N_45388);
and U47045 (N_47045,N_44559,N_44223);
nand U47046 (N_47046,N_44607,N_45116);
nand U47047 (N_47047,N_44447,N_45970);
nand U47048 (N_47048,N_44507,N_45948);
nand U47049 (N_47049,N_44319,N_45361);
or U47050 (N_47050,N_45857,N_44807);
or U47051 (N_47051,N_45545,N_44768);
nor U47052 (N_47052,N_44844,N_44386);
nor U47053 (N_47053,N_44198,N_45756);
and U47054 (N_47054,N_45866,N_44483);
xor U47055 (N_47055,N_44509,N_44619);
and U47056 (N_47056,N_45293,N_44482);
nand U47057 (N_47057,N_45726,N_45952);
and U47058 (N_47058,N_44070,N_44524);
or U47059 (N_47059,N_44432,N_45360);
xor U47060 (N_47060,N_45331,N_44563);
and U47061 (N_47061,N_45809,N_45853);
and U47062 (N_47062,N_45242,N_44867);
and U47063 (N_47063,N_44688,N_44099);
nand U47064 (N_47064,N_44266,N_44743);
nor U47065 (N_47065,N_45473,N_45853);
and U47066 (N_47066,N_45818,N_45259);
and U47067 (N_47067,N_44537,N_45963);
nor U47068 (N_47068,N_44666,N_45717);
nor U47069 (N_47069,N_44107,N_44728);
and U47070 (N_47070,N_45487,N_44860);
or U47071 (N_47071,N_45417,N_44782);
or U47072 (N_47072,N_44117,N_44006);
xor U47073 (N_47073,N_45567,N_44419);
xor U47074 (N_47074,N_44318,N_44732);
xnor U47075 (N_47075,N_45649,N_44595);
xnor U47076 (N_47076,N_44774,N_45398);
or U47077 (N_47077,N_45614,N_44280);
and U47078 (N_47078,N_45838,N_45752);
nand U47079 (N_47079,N_44593,N_45850);
xnor U47080 (N_47080,N_44923,N_45314);
xnor U47081 (N_47081,N_44187,N_45034);
xnor U47082 (N_47082,N_44973,N_44959);
and U47083 (N_47083,N_45541,N_45717);
or U47084 (N_47084,N_45964,N_44536);
or U47085 (N_47085,N_44705,N_44265);
nand U47086 (N_47086,N_44424,N_45288);
xnor U47087 (N_47087,N_45724,N_44773);
and U47088 (N_47088,N_45468,N_45808);
or U47089 (N_47089,N_44852,N_44292);
nand U47090 (N_47090,N_45425,N_44262);
nand U47091 (N_47091,N_45279,N_45626);
and U47092 (N_47092,N_44600,N_44934);
nand U47093 (N_47093,N_44707,N_45960);
and U47094 (N_47094,N_45440,N_45105);
nand U47095 (N_47095,N_44347,N_45213);
or U47096 (N_47096,N_44799,N_44250);
xor U47097 (N_47097,N_45531,N_45881);
nor U47098 (N_47098,N_45752,N_45900);
or U47099 (N_47099,N_45730,N_45121);
xor U47100 (N_47100,N_45886,N_44010);
nor U47101 (N_47101,N_45782,N_45569);
nand U47102 (N_47102,N_45638,N_45551);
xnor U47103 (N_47103,N_45599,N_45337);
nor U47104 (N_47104,N_45555,N_45022);
and U47105 (N_47105,N_44974,N_45162);
xnor U47106 (N_47106,N_45314,N_44203);
xor U47107 (N_47107,N_45440,N_44259);
nor U47108 (N_47108,N_45289,N_44494);
xnor U47109 (N_47109,N_44665,N_45058);
or U47110 (N_47110,N_44586,N_45479);
xnor U47111 (N_47111,N_45044,N_45414);
nor U47112 (N_47112,N_44515,N_44511);
xor U47113 (N_47113,N_44778,N_44801);
or U47114 (N_47114,N_44606,N_45354);
nand U47115 (N_47115,N_45206,N_44929);
and U47116 (N_47116,N_44993,N_45553);
and U47117 (N_47117,N_45448,N_44711);
and U47118 (N_47118,N_44442,N_44973);
nand U47119 (N_47119,N_44719,N_45449);
or U47120 (N_47120,N_45746,N_45852);
and U47121 (N_47121,N_44726,N_44700);
nor U47122 (N_47122,N_45695,N_44137);
xor U47123 (N_47123,N_45965,N_45047);
nor U47124 (N_47124,N_44441,N_44838);
and U47125 (N_47125,N_45725,N_44381);
nand U47126 (N_47126,N_45568,N_44641);
xor U47127 (N_47127,N_45205,N_45584);
nor U47128 (N_47128,N_44984,N_45488);
nand U47129 (N_47129,N_44817,N_44343);
or U47130 (N_47130,N_45343,N_44930);
nor U47131 (N_47131,N_45165,N_45504);
xnor U47132 (N_47132,N_45088,N_45778);
and U47133 (N_47133,N_45903,N_45880);
xor U47134 (N_47134,N_45711,N_44196);
or U47135 (N_47135,N_45116,N_45935);
xnor U47136 (N_47136,N_44971,N_45116);
or U47137 (N_47137,N_45704,N_45715);
xnor U47138 (N_47138,N_45978,N_45958);
or U47139 (N_47139,N_45008,N_44094);
and U47140 (N_47140,N_44843,N_45691);
nand U47141 (N_47141,N_45853,N_45427);
or U47142 (N_47142,N_44326,N_45410);
and U47143 (N_47143,N_44280,N_45908);
nand U47144 (N_47144,N_45519,N_45354);
nand U47145 (N_47145,N_45742,N_44149);
nand U47146 (N_47146,N_45671,N_44544);
or U47147 (N_47147,N_44327,N_45618);
and U47148 (N_47148,N_44964,N_45284);
nand U47149 (N_47149,N_45316,N_44284);
nand U47150 (N_47150,N_45203,N_45534);
or U47151 (N_47151,N_45992,N_45854);
and U47152 (N_47152,N_44984,N_44087);
nand U47153 (N_47153,N_45123,N_44286);
nor U47154 (N_47154,N_45044,N_45229);
and U47155 (N_47155,N_44972,N_45600);
or U47156 (N_47156,N_44568,N_45318);
nor U47157 (N_47157,N_44187,N_45041);
or U47158 (N_47158,N_45398,N_44545);
nand U47159 (N_47159,N_45834,N_45149);
and U47160 (N_47160,N_44952,N_44564);
xnor U47161 (N_47161,N_44822,N_44140);
nand U47162 (N_47162,N_45149,N_45048);
or U47163 (N_47163,N_44327,N_44256);
nor U47164 (N_47164,N_44238,N_44865);
xor U47165 (N_47165,N_45322,N_45302);
or U47166 (N_47166,N_44977,N_45032);
nor U47167 (N_47167,N_45966,N_45964);
or U47168 (N_47168,N_45435,N_45826);
and U47169 (N_47169,N_45436,N_44941);
and U47170 (N_47170,N_44668,N_44461);
nand U47171 (N_47171,N_44191,N_44021);
or U47172 (N_47172,N_44425,N_44578);
nor U47173 (N_47173,N_45731,N_44898);
nand U47174 (N_47174,N_45906,N_44333);
nand U47175 (N_47175,N_45680,N_45623);
nor U47176 (N_47176,N_44613,N_44191);
nor U47177 (N_47177,N_45252,N_44218);
and U47178 (N_47178,N_44157,N_45607);
nor U47179 (N_47179,N_44030,N_45467);
or U47180 (N_47180,N_44527,N_45245);
or U47181 (N_47181,N_44170,N_44444);
and U47182 (N_47182,N_44025,N_44834);
nor U47183 (N_47183,N_45460,N_44611);
nand U47184 (N_47184,N_45162,N_45234);
nand U47185 (N_47185,N_44575,N_45853);
nor U47186 (N_47186,N_45911,N_45201);
and U47187 (N_47187,N_45198,N_44971);
nor U47188 (N_47188,N_44163,N_45655);
nand U47189 (N_47189,N_44790,N_44923);
nor U47190 (N_47190,N_44068,N_45316);
or U47191 (N_47191,N_45269,N_44089);
xor U47192 (N_47192,N_44860,N_44183);
and U47193 (N_47193,N_45047,N_44701);
and U47194 (N_47194,N_45677,N_44109);
and U47195 (N_47195,N_44102,N_44166);
xor U47196 (N_47196,N_44499,N_44021);
xor U47197 (N_47197,N_44802,N_44193);
and U47198 (N_47198,N_45990,N_44410);
xor U47199 (N_47199,N_44955,N_44425);
or U47200 (N_47200,N_45454,N_44454);
xnor U47201 (N_47201,N_45278,N_45995);
or U47202 (N_47202,N_45317,N_44005);
xnor U47203 (N_47203,N_44316,N_45629);
or U47204 (N_47204,N_44072,N_45967);
or U47205 (N_47205,N_44321,N_45517);
and U47206 (N_47206,N_44929,N_44778);
or U47207 (N_47207,N_45362,N_44150);
xor U47208 (N_47208,N_44937,N_44250);
xnor U47209 (N_47209,N_44962,N_44867);
nor U47210 (N_47210,N_45239,N_45797);
or U47211 (N_47211,N_44525,N_45227);
nor U47212 (N_47212,N_45581,N_44325);
nor U47213 (N_47213,N_44614,N_45990);
nand U47214 (N_47214,N_45055,N_45447);
or U47215 (N_47215,N_45223,N_45907);
nor U47216 (N_47216,N_45641,N_45799);
or U47217 (N_47217,N_44248,N_44948);
nor U47218 (N_47218,N_44419,N_44701);
nor U47219 (N_47219,N_44120,N_45673);
and U47220 (N_47220,N_44793,N_45600);
or U47221 (N_47221,N_44314,N_45861);
nor U47222 (N_47222,N_44882,N_44478);
nor U47223 (N_47223,N_44418,N_45961);
nor U47224 (N_47224,N_45666,N_44804);
nand U47225 (N_47225,N_44606,N_44795);
or U47226 (N_47226,N_45028,N_44766);
nand U47227 (N_47227,N_44041,N_44107);
xnor U47228 (N_47228,N_44730,N_44901);
or U47229 (N_47229,N_44562,N_45765);
xnor U47230 (N_47230,N_45412,N_44026);
xnor U47231 (N_47231,N_45511,N_44265);
and U47232 (N_47232,N_45586,N_44605);
xor U47233 (N_47233,N_44481,N_44691);
nor U47234 (N_47234,N_45130,N_45979);
or U47235 (N_47235,N_45039,N_44764);
xor U47236 (N_47236,N_45247,N_45651);
nor U47237 (N_47237,N_45135,N_45979);
or U47238 (N_47238,N_45851,N_45068);
nand U47239 (N_47239,N_45161,N_44201);
nand U47240 (N_47240,N_45650,N_44101);
nor U47241 (N_47241,N_45224,N_45683);
or U47242 (N_47242,N_45328,N_44590);
xnor U47243 (N_47243,N_45261,N_44974);
nor U47244 (N_47244,N_44745,N_44220);
xor U47245 (N_47245,N_45673,N_44436);
and U47246 (N_47246,N_45061,N_44298);
nand U47247 (N_47247,N_44612,N_44486);
nand U47248 (N_47248,N_45316,N_44550);
and U47249 (N_47249,N_45793,N_44446);
and U47250 (N_47250,N_44241,N_45101);
and U47251 (N_47251,N_45587,N_44573);
or U47252 (N_47252,N_45903,N_45236);
and U47253 (N_47253,N_44879,N_44912);
and U47254 (N_47254,N_44809,N_45795);
nand U47255 (N_47255,N_44760,N_44853);
nand U47256 (N_47256,N_45823,N_45715);
and U47257 (N_47257,N_44165,N_44135);
nand U47258 (N_47258,N_45674,N_44077);
xnor U47259 (N_47259,N_44586,N_45384);
and U47260 (N_47260,N_44659,N_44591);
nand U47261 (N_47261,N_44024,N_44690);
nor U47262 (N_47262,N_45396,N_45167);
and U47263 (N_47263,N_44335,N_45429);
nand U47264 (N_47264,N_44175,N_44096);
and U47265 (N_47265,N_45657,N_45034);
or U47266 (N_47266,N_45166,N_45956);
or U47267 (N_47267,N_45539,N_45404);
xnor U47268 (N_47268,N_44232,N_44239);
nor U47269 (N_47269,N_45085,N_44527);
nor U47270 (N_47270,N_44497,N_45712);
nor U47271 (N_47271,N_44041,N_45194);
xnor U47272 (N_47272,N_44789,N_45744);
and U47273 (N_47273,N_45862,N_44943);
nand U47274 (N_47274,N_44363,N_45737);
and U47275 (N_47275,N_44756,N_44777);
and U47276 (N_47276,N_44312,N_45497);
xor U47277 (N_47277,N_44622,N_45208);
and U47278 (N_47278,N_44788,N_44298);
and U47279 (N_47279,N_45056,N_45553);
xor U47280 (N_47280,N_44942,N_44275);
and U47281 (N_47281,N_44184,N_45038);
and U47282 (N_47282,N_44094,N_44039);
or U47283 (N_47283,N_45878,N_45417);
or U47284 (N_47284,N_44572,N_45064);
nor U47285 (N_47285,N_45090,N_44103);
and U47286 (N_47286,N_44117,N_45684);
or U47287 (N_47287,N_45985,N_44870);
nor U47288 (N_47288,N_45987,N_44231);
nor U47289 (N_47289,N_45395,N_45518);
nor U47290 (N_47290,N_45747,N_45171);
xor U47291 (N_47291,N_45918,N_45737);
xor U47292 (N_47292,N_44972,N_44790);
or U47293 (N_47293,N_44161,N_45794);
nor U47294 (N_47294,N_44814,N_44020);
and U47295 (N_47295,N_44121,N_44089);
nand U47296 (N_47296,N_45924,N_45357);
or U47297 (N_47297,N_44187,N_45830);
nand U47298 (N_47298,N_45586,N_45230);
xor U47299 (N_47299,N_45336,N_45732);
xnor U47300 (N_47300,N_45075,N_45232);
xnor U47301 (N_47301,N_45507,N_44950);
xor U47302 (N_47302,N_45410,N_44431);
and U47303 (N_47303,N_45669,N_44823);
nor U47304 (N_47304,N_45089,N_45643);
nand U47305 (N_47305,N_44570,N_45403);
xor U47306 (N_47306,N_44048,N_44141);
xor U47307 (N_47307,N_44418,N_44946);
or U47308 (N_47308,N_44533,N_45217);
xnor U47309 (N_47309,N_44399,N_45707);
and U47310 (N_47310,N_45307,N_44490);
nand U47311 (N_47311,N_44282,N_45372);
nor U47312 (N_47312,N_45362,N_45590);
xor U47313 (N_47313,N_44783,N_45597);
and U47314 (N_47314,N_44807,N_45932);
nand U47315 (N_47315,N_45188,N_44934);
and U47316 (N_47316,N_44488,N_45263);
and U47317 (N_47317,N_44464,N_44099);
nor U47318 (N_47318,N_45856,N_45197);
xor U47319 (N_47319,N_45030,N_44690);
and U47320 (N_47320,N_45926,N_45618);
nand U47321 (N_47321,N_44673,N_45944);
nand U47322 (N_47322,N_44857,N_44040);
and U47323 (N_47323,N_45876,N_44301);
xnor U47324 (N_47324,N_45200,N_45347);
or U47325 (N_47325,N_44879,N_44759);
xnor U47326 (N_47326,N_44264,N_45781);
nand U47327 (N_47327,N_45659,N_44905);
and U47328 (N_47328,N_45706,N_44606);
or U47329 (N_47329,N_45766,N_45506);
nand U47330 (N_47330,N_44678,N_45474);
nor U47331 (N_47331,N_44643,N_44185);
xor U47332 (N_47332,N_44084,N_45897);
nor U47333 (N_47333,N_45770,N_45495);
nand U47334 (N_47334,N_45890,N_45802);
xor U47335 (N_47335,N_45096,N_45525);
and U47336 (N_47336,N_44350,N_45919);
xor U47337 (N_47337,N_45219,N_44271);
xnor U47338 (N_47338,N_44709,N_44213);
nor U47339 (N_47339,N_44244,N_44140);
xor U47340 (N_47340,N_44158,N_45546);
xor U47341 (N_47341,N_45197,N_45403);
xor U47342 (N_47342,N_44244,N_45244);
or U47343 (N_47343,N_44674,N_45252);
nand U47344 (N_47344,N_44844,N_44188);
and U47345 (N_47345,N_45705,N_45365);
nor U47346 (N_47346,N_44584,N_44616);
or U47347 (N_47347,N_45425,N_44984);
and U47348 (N_47348,N_44836,N_44393);
nor U47349 (N_47349,N_44558,N_44713);
and U47350 (N_47350,N_44963,N_44622);
nor U47351 (N_47351,N_45823,N_44638);
nand U47352 (N_47352,N_45894,N_44683);
nand U47353 (N_47353,N_45936,N_45004);
nand U47354 (N_47354,N_44264,N_44863);
nand U47355 (N_47355,N_44298,N_45034);
nor U47356 (N_47356,N_45345,N_45299);
nand U47357 (N_47357,N_45986,N_44107);
and U47358 (N_47358,N_45184,N_44662);
nand U47359 (N_47359,N_45665,N_44008);
nand U47360 (N_47360,N_44287,N_45991);
nor U47361 (N_47361,N_45327,N_44977);
and U47362 (N_47362,N_45066,N_44969);
xor U47363 (N_47363,N_45299,N_44112);
nor U47364 (N_47364,N_44221,N_44667);
nand U47365 (N_47365,N_45966,N_44603);
or U47366 (N_47366,N_44131,N_44967);
nor U47367 (N_47367,N_44941,N_44759);
or U47368 (N_47368,N_44744,N_44341);
and U47369 (N_47369,N_45836,N_45530);
and U47370 (N_47370,N_45975,N_44880);
xnor U47371 (N_47371,N_44359,N_44073);
and U47372 (N_47372,N_44336,N_45052);
nand U47373 (N_47373,N_44965,N_44609);
xnor U47374 (N_47374,N_45195,N_44869);
or U47375 (N_47375,N_44891,N_45518);
and U47376 (N_47376,N_44923,N_45925);
xor U47377 (N_47377,N_45256,N_44515);
and U47378 (N_47378,N_45943,N_44814);
nand U47379 (N_47379,N_44024,N_44307);
or U47380 (N_47380,N_44898,N_45763);
nor U47381 (N_47381,N_44207,N_44598);
or U47382 (N_47382,N_44649,N_44473);
xor U47383 (N_47383,N_44957,N_44185);
nand U47384 (N_47384,N_45818,N_44101);
nand U47385 (N_47385,N_45726,N_45056);
nand U47386 (N_47386,N_44492,N_45277);
or U47387 (N_47387,N_44214,N_44763);
nand U47388 (N_47388,N_44329,N_44764);
xor U47389 (N_47389,N_45178,N_45359);
or U47390 (N_47390,N_45765,N_45523);
xnor U47391 (N_47391,N_44352,N_44311);
nand U47392 (N_47392,N_45531,N_45304);
or U47393 (N_47393,N_45344,N_45470);
and U47394 (N_47394,N_44105,N_44175);
or U47395 (N_47395,N_44493,N_44285);
nand U47396 (N_47396,N_44589,N_44391);
and U47397 (N_47397,N_45819,N_45956);
nand U47398 (N_47398,N_45490,N_45030);
and U47399 (N_47399,N_45577,N_44724);
nand U47400 (N_47400,N_45169,N_44964);
or U47401 (N_47401,N_44640,N_44918);
xor U47402 (N_47402,N_44759,N_45432);
xor U47403 (N_47403,N_45786,N_45815);
nor U47404 (N_47404,N_44466,N_45772);
xnor U47405 (N_47405,N_45286,N_44673);
and U47406 (N_47406,N_44848,N_44566);
and U47407 (N_47407,N_44192,N_44460);
xnor U47408 (N_47408,N_45271,N_44742);
or U47409 (N_47409,N_44051,N_45611);
nand U47410 (N_47410,N_45576,N_44738);
nor U47411 (N_47411,N_44372,N_45057);
and U47412 (N_47412,N_45459,N_45461);
xor U47413 (N_47413,N_44398,N_45225);
or U47414 (N_47414,N_44322,N_44140);
nand U47415 (N_47415,N_45875,N_44975);
and U47416 (N_47416,N_44335,N_45981);
nor U47417 (N_47417,N_45134,N_45528);
xor U47418 (N_47418,N_45405,N_44632);
nand U47419 (N_47419,N_45024,N_45116);
xnor U47420 (N_47420,N_45163,N_44530);
nand U47421 (N_47421,N_44181,N_44150);
or U47422 (N_47422,N_45311,N_45770);
xor U47423 (N_47423,N_44303,N_45358);
and U47424 (N_47424,N_44462,N_44803);
and U47425 (N_47425,N_45927,N_45259);
or U47426 (N_47426,N_44280,N_44101);
or U47427 (N_47427,N_44020,N_44119);
nand U47428 (N_47428,N_44836,N_44856);
nand U47429 (N_47429,N_45839,N_45436);
xor U47430 (N_47430,N_44323,N_45242);
nor U47431 (N_47431,N_44489,N_44031);
nand U47432 (N_47432,N_45961,N_45640);
xor U47433 (N_47433,N_45238,N_44051);
nor U47434 (N_47434,N_45783,N_44116);
nand U47435 (N_47435,N_45140,N_44689);
nand U47436 (N_47436,N_45875,N_45280);
nor U47437 (N_47437,N_45001,N_45293);
or U47438 (N_47438,N_44771,N_44367);
and U47439 (N_47439,N_44231,N_45909);
or U47440 (N_47440,N_45898,N_44993);
nor U47441 (N_47441,N_45125,N_44073);
xor U47442 (N_47442,N_45727,N_44011);
or U47443 (N_47443,N_44160,N_44753);
xor U47444 (N_47444,N_45490,N_45602);
nor U47445 (N_47445,N_44437,N_44959);
nor U47446 (N_47446,N_45566,N_45164);
and U47447 (N_47447,N_45431,N_44772);
or U47448 (N_47448,N_44208,N_44434);
xor U47449 (N_47449,N_45271,N_45759);
xor U47450 (N_47450,N_44294,N_45143);
nand U47451 (N_47451,N_45177,N_44044);
nor U47452 (N_47452,N_44161,N_45896);
nor U47453 (N_47453,N_45013,N_45511);
nor U47454 (N_47454,N_45470,N_44985);
nor U47455 (N_47455,N_44095,N_44586);
xor U47456 (N_47456,N_44818,N_44310);
and U47457 (N_47457,N_44966,N_45550);
and U47458 (N_47458,N_44369,N_45033);
xor U47459 (N_47459,N_44299,N_45703);
or U47460 (N_47460,N_45997,N_44639);
or U47461 (N_47461,N_44275,N_44502);
xnor U47462 (N_47462,N_45580,N_44328);
nand U47463 (N_47463,N_45985,N_45631);
and U47464 (N_47464,N_45614,N_45169);
xor U47465 (N_47465,N_44833,N_44832);
nor U47466 (N_47466,N_44743,N_44438);
xor U47467 (N_47467,N_44526,N_45773);
or U47468 (N_47468,N_44427,N_45250);
nand U47469 (N_47469,N_45465,N_45206);
nor U47470 (N_47470,N_44630,N_45627);
or U47471 (N_47471,N_44631,N_45144);
and U47472 (N_47472,N_45549,N_44213);
xor U47473 (N_47473,N_45192,N_44714);
nor U47474 (N_47474,N_45519,N_44087);
or U47475 (N_47475,N_44074,N_44186);
nand U47476 (N_47476,N_44832,N_44175);
xor U47477 (N_47477,N_45001,N_45094);
nor U47478 (N_47478,N_45613,N_44454);
nand U47479 (N_47479,N_44735,N_45765);
or U47480 (N_47480,N_44277,N_44115);
nor U47481 (N_47481,N_44700,N_44542);
xor U47482 (N_47482,N_45637,N_45250);
nor U47483 (N_47483,N_45380,N_44181);
and U47484 (N_47484,N_44003,N_45261);
nor U47485 (N_47485,N_45050,N_44129);
nand U47486 (N_47486,N_44684,N_45149);
nor U47487 (N_47487,N_45328,N_45507);
nor U47488 (N_47488,N_44135,N_45224);
or U47489 (N_47489,N_45847,N_44527);
nor U47490 (N_47490,N_45269,N_45637);
and U47491 (N_47491,N_45282,N_44501);
nor U47492 (N_47492,N_45335,N_44244);
or U47493 (N_47493,N_45270,N_44342);
xor U47494 (N_47494,N_45607,N_44736);
and U47495 (N_47495,N_44643,N_45806);
and U47496 (N_47496,N_45056,N_44002);
nand U47497 (N_47497,N_44971,N_45861);
or U47498 (N_47498,N_45201,N_45463);
and U47499 (N_47499,N_45766,N_44066);
nand U47500 (N_47500,N_44374,N_44974);
nor U47501 (N_47501,N_45040,N_44547);
and U47502 (N_47502,N_45530,N_45178);
and U47503 (N_47503,N_45891,N_44322);
and U47504 (N_47504,N_45136,N_45453);
or U47505 (N_47505,N_44062,N_45773);
nor U47506 (N_47506,N_45985,N_44045);
nor U47507 (N_47507,N_45012,N_44715);
or U47508 (N_47508,N_44662,N_45990);
nor U47509 (N_47509,N_45994,N_45473);
or U47510 (N_47510,N_45543,N_44148);
nor U47511 (N_47511,N_44163,N_44861);
and U47512 (N_47512,N_44867,N_45130);
nor U47513 (N_47513,N_44304,N_45498);
or U47514 (N_47514,N_45463,N_45125);
xnor U47515 (N_47515,N_45784,N_45887);
nand U47516 (N_47516,N_44707,N_44710);
or U47517 (N_47517,N_45519,N_45415);
and U47518 (N_47518,N_45192,N_45703);
nand U47519 (N_47519,N_44143,N_44442);
or U47520 (N_47520,N_44023,N_45699);
nand U47521 (N_47521,N_45356,N_45024);
nand U47522 (N_47522,N_44485,N_44940);
xnor U47523 (N_47523,N_45400,N_45779);
and U47524 (N_47524,N_45674,N_44406);
and U47525 (N_47525,N_44551,N_45190);
xor U47526 (N_47526,N_45896,N_45230);
nor U47527 (N_47527,N_45687,N_45070);
and U47528 (N_47528,N_45170,N_45076);
nor U47529 (N_47529,N_45508,N_44895);
xor U47530 (N_47530,N_45075,N_44776);
nand U47531 (N_47531,N_45484,N_44435);
and U47532 (N_47532,N_45656,N_44325);
nand U47533 (N_47533,N_45494,N_45117);
and U47534 (N_47534,N_45109,N_44601);
nand U47535 (N_47535,N_44442,N_44397);
nor U47536 (N_47536,N_44434,N_44599);
or U47537 (N_47537,N_45930,N_45798);
nand U47538 (N_47538,N_45129,N_44094);
and U47539 (N_47539,N_45346,N_45777);
and U47540 (N_47540,N_45382,N_45830);
nand U47541 (N_47541,N_44226,N_44824);
xor U47542 (N_47542,N_45461,N_44478);
nor U47543 (N_47543,N_44390,N_44112);
nand U47544 (N_47544,N_44061,N_45333);
nand U47545 (N_47545,N_45464,N_45290);
xnor U47546 (N_47546,N_45832,N_44832);
or U47547 (N_47547,N_44400,N_45435);
nand U47548 (N_47548,N_45096,N_45115);
or U47549 (N_47549,N_45323,N_45804);
nor U47550 (N_47550,N_45743,N_44460);
or U47551 (N_47551,N_44578,N_45430);
and U47552 (N_47552,N_45540,N_44268);
or U47553 (N_47553,N_44409,N_45593);
nand U47554 (N_47554,N_44011,N_44166);
and U47555 (N_47555,N_45997,N_45260);
or U47556 (N_47556,N_45276,N_45125);
nor U47557 (N_47557,N_45048,N_44589);
xor U47558 (N_47558,N_45852,N_44291);
and U47559 (N_47559,N_44415,N_44697);
nand U47560 (N_47560,N_44768,N_44820);
or U47561 (N_47561,N_44648,N_44895);
nor U47562 (N_47562,N_45963,N_44321);
and U47563 (N_47563,N_45637,N_44231);
nand U47564 (N_47564,N_45348,N_45778);
or U47565 (N_47565,N_45260,N_44168);
and U47566 (N_47566,N_44756,N_44633);
nand U47567 (N_47567,N_45066,N_44354);
nand U47568 (N_47568,N_44128,N_45716);
xor U47569 (N_47569,N_45538,N_45138);
nor U47570 (N_47570,N_44191,N_45512);
nor U47571 (N_47571,N_45610,N_44515);
or U47572 (N_47572,N_45266,N_44478);
or U47573 (N_47573,N_45831,N_45285);
xnor U47574 (N_47574,N_44185,N_45190);
nand U47575 (N_47575,N_44491,N_44007);
and U47576 (N_47576,N_44248,N_44722);
nand U47577 (N_47577,N_44292,N_45237);
or U47578 (N_47578,N_44183,N_44603);
xnor U47579 (N_47579,N_45431,N_44609);
and U47580 (N_47580,N_44093,N_44972);
and U47581 (N_47581,N_45459,N_45049);
nor U47582 (N_47582,N_45196,N_45788);
nor U47583 (N_47583,N_45760,N_44137);
nand U47584 (N_47584,N_44979,N_45340);
nor U47585 (N_47585,N_45171,N_44975);
nand U47586 (N_47586,N_45382,N_44142);
and U47587 (N_47587,N_45055,N_45356);
nor U47588 (N_47588,N_44136,N_44688);
nor U47589 (N_47589,N_45620,N_44043);
xor U47590 (N_47590,N_45610,N_45085);
nor U47591 (N_47591,N_45539,N_45693);
or U47592 (N_47592,N_45952,N_44943);
or U47593 (N_47593,N_45592,N_45791);
nand U47594 (N_47594,N_44261,N_44574);
nor U47595 (N_47595,N_44332,N_45784);
and U47596 (N_47596,N_44068,N_44115);
or U47597 (N_47597,N_44462,N_45951);
nor U47598 (N_47598,N_45588,N_45861);
or U47599 (N_47599,N_45483,N_44490);
nand U47600 (N_47600,N_44914,N_44182);
nand U47601 (N_47601,N_45730,N_44440);
nand U47602 (N_47602,N_45757,N_44859);
xor U47603 (N_47603,N_44630,N_45922);
nand U47604 (N_47604,N_44750,N_45645);
xor U47605 (N_47605,N_45251,N_44595);
nor U47606 (N_47606,N_44050,N_44764);
xnor U47607 (N_47607,N_45708,N_45030);
xor U47608 (N_47608,N_45141,N_44003);
xnor U47609 (N_47609,N_44578,N_45934);
nand U47610 (N_47610,N_44192,N_44937);
nor U47611 (N_47611,N_45674,N_45285);
nand U47612 (N_47612,N_44730,N_45172);
or U47613 (N_47613,N_45454,N_44695);
nand U47614 (N_47614,N_45786,N_44708);
nor U47615 (N_47615,N_45069,N_44333);
xor U47616 (N_47616,N_44399,N_44446);
nor U47617 (N_47617,N_45592,N_44526);
xor U47618 (N_47618,N_44371,N_44639);
nand U47619 (N_47619,N_45124,N_44964);
nor U47620 (N_47620,N_44894,N_45423);
xor U47621 (N_47621,N_45276,N_44574);
or U47622 (N_47622,N_44861,N_45256);
nand U47623 (N_47623,N_44258,N_44456);
xnor U47624 (N_47624,N_44653,N_44931);
and U47625 (N_47625,N_45585,N_45010);
nor U47626 (N_47626,N_44001,N_45814);
or U47627 (N_47627,N_44681,N_44161);
xor U47628 (N_47628,N_45570,N_44895);
or U47629 (N_47629,N_45065,N_44491);
nor U47630 (N_47630,N_45786,N_44701);
nand U47631 (N_47631,N_45657,N_45445);
and U47632 (N_47632,N_44538,N_44519);
or U47633 (N_47633,N_44946,N_44558);
nor U47634 (N_47634,N_44292,N_44456);
xnor U47635 (N_47635,N_45021,N_45295);
and U47636 (N_47636,N_44364,N_44975);
nor U47637 (N_47637,N_45300,N_45168);
nand U47638 (N_47638,N_44790,N_44014);
nor U47639 (N_47639,N_45019,N_44813);
or U47640 (N_47640,N_45951,N_44631);
xnor U47641 (N_47641,N_45723,N_45675);
xor U47642 (N_47642,N_44647,N_44358);
and U47643 (N_47643,N_44113,N_44762);
nand U47644 (N_47644,N_45151,N_44575);
xnor U47645 (N_47645,N_45634,N_44933);
nor U47646 (N_47646,N_45967,N_44304);
and U47647 (N_47647,N_44889,N_44485);
or U47648 (N_47648,N_44466,N_44070);
nand U47649 (N_47649,N_44934,N_45884);
or U47650 (N_47650,N_44138,N_44943);
or U47651 (N_47651,N_45669,N_45087);
xnor U47652 (N_47652,N_45884,N_45248);
xor U47653 (N_47653,N_44021,N_44655);
xor U47654 (N_47654,N_45900,N_44907);
xnor U47655 (N_47655,N_44082,N_44872);
nand U47656 (N_47656,N_44796,N_44498);
and U47657 (N_47657,N_44775,N_45403);
and U47658 (N_47658,N_45948,N_44338);
or U47659 (N_47659,N_45463,N_45931);
or U47660 (N_47660,N_45224,N_45080);
nor U47661 (N_47661,N_45531,N_45481);
or U47662 (N_47662,N_44757,N_45747);
and U47663 (N_47663,N_44138,N_45922);
nor U47664 (N_47664,N_44341,N_45098);
xnor U47665 (N_47665,N_45184,N_45234);
and U47666 (N_47666,N_45805,N_44851);
nor U47667 (N_47667,N_45931,N_44190);
nor U47668 (N_47668,N_44557,N_45386);
or U47669 (N_47669,N_45107,N_45250);
or U47670 (N_47670,N_45964,N_45822);
nor U47671 (N_47671,N_45265,N_44998);
xor U47672 (N_47672,N_45746,N_44540);
nor U47673 (N_47673,N_44224,N_45392);
nor U47674 (N_47674,N_44159,N_44224);
nor U47675 (N_47675,N_45493,N_45769);
nand U47676 (N_47676,N_44781,N_44941);
and U47677 (N_47677,N_45547,N_44482);
xor U47678 (N_47678,N_45388,N_44540);
nand U47679 (N_47679,N_44056,N_45666);
xnor U47680 (N_47680,N_44056,N_45566);
nand U47681 (N_47681,N_45919,N_45518);
nand U47682 (N_47682,N_44427,N_45193);
or U47683 (N_47683,N_44908,N_45265);
nand U47684 (N_47684,N_44034,N_45802);
or U47685 (N_47685,N_45045,N_45563);
and U47686 (N_47686,N_45857,N_45263);
xor U47687 (N_47687,N_45456,N_45405);
xor U47688 (N_47688,N_45854,N_45201);
nor U47689 (N_47689,N_45364,N_45653);
nand U47690 (N_47690,N_45200,N_45000);
xor U47691 (N_47691,N_45250,N_44724);
and U47692 (N_47692,N_45527,N_45526);
and U47693 (N_47693,N_45835,N_45227);
and U47694 (N_47694,N_44356,N_44964);
nand U47695 (N_47695,N_45226,N_45729);
or U47696 (N_47696,N_44288,N_44808);
xnor U47697 (N_47697,N_45296,N_45495);
nand U47698 (N_47698,N_45396,N_44727);
and U47699 (N_47699,N_44170,N_44575);
nor U47700 (N_47700,N_45849,N_45052);
or U47701 (N_47701,N_45613,N_45630);
nor U47702 (N_47702,N_45517,N_45547);
nor U47703 (N_47703,N_44201,N_44876);
xor U47704 (N_47704,N_45990,N_44041);
nor U47705 (N_47705,N_44271,N_44798);
and U47706 (N_47706,N_45536,N_44986);
and U47707 (N_47707,N_44801,N_45039);
or U47708 (N_47708,N_45814,N_45607);
or U47709 (N_47709,N_45234,N_45256);
nand U47710 (N_47710,N_45206,N_45854);
and U47711 (N_47711,N_44868,N_44119);
or U47712 (N_47712,N_45977,N_45767);
nor U47713 (N_47713,N_45101,N_44310);
xor U47714 (N_47714,N_45772,N_44434);
nor U47715 (N_47715,N_45942,N_44641);
xor U47716 (N_47716,N_45110,N_44126);
and U47717 (N_47717,N_44862,N_44998);
nor U47718 (N_47718,N_45008,N_45863);
and U47719 (N_47719,N_44845,N_44257);
and U47720 (N_47720,N_44562,N_45801);
and U47721 (N_47721,N_44468,N_45729);
xor U47722 (N_47722,N_44068,N_44083);
xnor U47723 (N_47723,N_45601,N_45398);
nand U47724 (N_47724,N_44944,N_45730);
nand U47725 (N_47725,N_45131,N_45620);
or U47726 (N_47726,N_45005,N_44184);
nand U47727 (N_47727,N_44825,N_45278);
xor U47728 (N_47728,N_44027,N_45291);
nand U47729 (N_47729,N_45565,N_44654);
nor U47730 (N_47730,N_45500,N_45640);
or U47731 (N_47731,N_45183,N_44097);
or U47732 (N_47732,N_44424,N_44221);
nand U47733 (N_47733,N_44235,N_44893);
or U47734 (N_47734,N_45384,N_44205);
and U47735 (N_47735,N_45770,N_45422);
and U47736 (N_47736,N_44731,N_45345);
and U47737 (N_47737,N_45003,N_45009);
and U47738 (N_47738,N_44853,N_44342);
or U47739 (N_47739,N_44154,N_44567);
xnor U47740 (N_47740,N_45257,N_45854);
nor U47741 (N_47741,N_45049,N_45926);
nor U47742 (N_47742,N_44479,N_44977);
xor U47743 (N_47743,N_45973,N_44407);
nor U47744 (N_47744,N_45962,N_45751);
nor U47745 (N_47745,N_45174,N_44604);
nor U47746 (N_47746,N_44034,N_44757);
or U47747 (N_47747,N_45360,N_45318);
or U47748 (N_47748,N_44758,N_44404);
or U47749 (N_47749,N_45644,N_45336);
nand U47750 (N_47750,N_45476,N_45857);
and U47751 (N_47751,N_45103,N_45167);
nor U47752 (N_47752,N_45086,N_45003);
or U47753 (N_47753,N_44571,N_45288);
xor U47754 (N_47754,N_44208,N_44025);
xor U47755 (N_47755,N_44065,N_44846);
nor U47756 (N_47756,N_45330,N_44198);
xnor U47757 (N_47757,N_44499,N_45920);
or U47758 (N_47758,N_45263,N_45355);
nand U47759 (N_47759,N_45816,N_44333);
and U47760 (N_47760,N_44451,N_44047);
nor U47761 (N_47761,N_45102,N_44233);
xor U47762 (N_47762,N_44799,N_45084);
and U47763 (N_47763,N_45359,N_44616);
nor U47764 (N_47764,N_45982,N_44541);
and U47765 (N_47765,N_44730,N_44833);
or U47766 (N_47766,N_44660,N_45301);
nand U47767 (N_47767,N_44948,N_45482);
nor U47768 (N_47768,N_44203,N_45567);
or U47769 (N_47769,N_45479,N_44825);
and U47770 (N_47770,N_44731,N_44107);
nor U47771 (N_47771,N_45939,N_45437);
nand U47772 (N_47772,N_45405,N_44982);
nor U47773 (N_47773,N_44202,N_45479);
and U47774 (N_47774,N_44917,N_44000);
xor U47775 (N_47775,N_45056,N_45716);
nor U47776 (N_47776,N_45041,N_45259);
xnor U47777 (N_47777,N_45986,N_45037);
or U47778 (N_47778,N_45028,N_44702);
nor U47779 (N_47779,N_44371,N_44252);
nor U47780 (N_47780,N_45228,N_44428);
and U47781 (N_47781,N_45317,N_44657);
nor U47782 (N_47782,N_44560,N_45790);
and U47783 (N_47783,N_45608,N_45880);
and U47784 (N_47784,N_44147,N_45492);
and U47785 (N_47785,N_44536,N_45962);
nor U47786 (N_47786,N_44582,N_44335);
nand U47787 (N_47787,N_44270,N_45396);
nor U47788 (N_47788,N_45533,N_45275);
and U47789 (N_47789,N_45429,N_44189);
nor U47790 (N_47790,N_45494,N_44490);
nand U47791 (N_47791,N_45577,N_44381);
nor U47792 (N_47792,N_45648,N_45219);
xnor U47793 (N_47793,N_45178,N_45364);
or U47794 (N_47794,N_44656,N_44110);
nand U47795 (N_47795,N_44080,N_44541);
and U47796 (N_47796,N_44322,N_44189);
or U47797 (N_47797,N_44386,N_44104);
xor U47798 (N_47798,N_45906,N_44014);
nor U47799 (N_47799,N_45934,N_44837);
xnor U47800 (N_47800,N_44094,N_44449);
xnor U47801 (N_47801,N_45444,N_45979);
and U47802 (N_47802,N_45179,N_44340);
and U47803 (N_47803,N_44643,N_44676);
or U47804 (N_47804,N_44393,N_45960);
xor U47805 (N_47805,N_45951,N_44644);
and U47806 (N_47806,N_44859,N_44475);
nor U47807 (N_47807,N_45992,N_44326);
nand U47808 (N_47808,N_44817,N_44570);
nand U47809 (N_47809,N_45204,N_44665);
nand U47810 (N_47810,N_45024,N_44019);
nand U47811 (N_47811,N_44575,N_45139);
or U47812 (N_47812,N_44985,N_45434);
and U47813 (N_47813,N_45561,N_45889);
or U47814 (N_47814,N_44587,N_44034);
xor U47815 (N_47815,N_44618,N_44290);
xnor U47816 (N_47816,N_45140,N_44463);
or U47817 (N_47817,N_45793,N_45261);
nand U47818 (N_47818,N_44694,N_45822);
or U47819 (N_47819,N_44032,N_45511);
nor U47820 (N_47820,N_45718,N_44279);
nor U47821 (N_47821,N_44824,N_44091);
or U47822 (N_47822,N_44350,N_44461);
and U47823 (N_47823,N_44626,N_44477);
or U47824 (N_47824,N_45275,N_45913);
and U47825 (N_47825,N_45942,N_45442);
nand U47826 (N_47826,N_44751,N_45804);
xnor U47827 (N_47827,N_45669,N_45411);
or U47828 (N_47828,N_44916,N_45182);
nand U47829 (N_47829,N_45560,N_44703);
nand U47830 (N_47830,N_44913,N_44004);
xnor U47831 (N_47831,N_45628,N_45045);
xnor U47832 (N_47832,N_44924,N_44408);
xor U47833 (N_47833,N_44125,N_44762);
nor U47834 (N_47834,N_45091,N_45256);
nor U47835 (N_47835,N_45068,N_45452);
xor U47836 (N_47836,N_45690,N_45892);
or U47837 (N_47837,N_45588,N_45361);
xor U47838 (N_47838,N_44587,N_44366);
nor U47839 (N_47839,N_44034,N_45561);
xor U47840 (N_47840,N_45105,N_45529);
xnor U47841 (N_47841,N_44873,N_44242);
nor U47842 (N_47842,N_44501,N_45677);
or U47843 (N_47843,N_45562,N_45756);
xor U47844 (N_47844,N_44725,N_44640);
xor U47845 (N_47845,N_44830,N_44296);
and U47846 (N_47846,N_44551,N_44193);
xor U47847 (N_47847,N_44937,N_45392);
and U47848 (N_47848,N_45012,N_44432);
nand U47849 (N_47849,N_44502,N_44054);
or U47850 (N_47850,N_45214,N_45911);
nand U47851 (N_47851,N_44527,N_45362);
nand U47852 (N_47852,N_44208,N_45850);
or U47853 (N_47853,N_45100,N_45264);
and U47854 (N_47854,N_44605,N_44741);
nor U47855 (N_47855,N_44049,N_44969);
xnor U47856 (N_47856,N_45006,N_44628);
nor U47857 (N_47857,N_44677,N_45901);
nand U47858 (N_47858,N_44820,N_44785);
or U47859 (N_47859,N_45537,N_44101);
nor U47860 (N_47860,N_45925,N_45119);
nand U47861 (N_47861,N_45255,N_44296);
and U47862 (N_47862,N_45629,N_44352);
and U47863 (N_47863,N_45334,N_44695);
nor U47864 (N_47864,N_44554,N_45936);
nor U47865 (N_47865,N_45520,N_44246);
or U47866 (N_47866,N_44978,N_45522);
nor U47867 (N_47867,N_44867,N_45415);
nor U47868 (N_47868,N_45982,N_45914);
nor U47869 (N_47869,N_44479,N_45427);
nor U47870 (N_47870,N_45961,N_45393);
xnor U47871 (N_47871,N_45033,N_44176);
or U47872 (N_47872,N_44037,N_44171);
or U47873 (N_47873,N_44026,N_45509);
nor U47874 (N_47874,N_45677,N_44673);
xnor U47875 (N_47875,N_44919,N_45398);
nor U47876 (N_47876,N_45028,N_44450);
nand U47877 (N_47877,N_44138,N_45213);
nand U47878 (N_47878,N_45834,N_44860);
xnor U47879 (N_47879,N_44388,N_45234);
nand U47880 (N_47880,N_45407,N_45392);
xnor U47881 (N_47881,N_44086,N_45424);
or U47882 (N_47882,N_44893,N_44535);
nor U47883 (N_47883,N_44975,N_44626);
xnor U47884 (N_47884,N_45423,N_44815);
and U47885 (N_47885,N_44063,N_44442);
nor U47886 (N_47886,N_45997,N_45062);
nand U47887 (N_47887,N_44642,N_45603);
nand U47888 (N_47888,N_44939,N_45102);
and U47889 (N_47889,N_45457,N_45169);
nand U47890 (N_47890,N_44546,N_45248);
nand U47891 (N_47891,N_45766,N_44408);
nor U47892 (N_47892,N_45214,N_44313);
and U47893 (N_47893,N_45614,N_45150);
and U47894 (N_47894,N_44900,N_44830);
nor U47895 (N_47895,N_44698,N_45113);
xnor U47896 (N_47896,N_45619,N_44205);
or U47897 (N_47897,N_44960,N_45190);
and U47898 (N_47898,N_45719,N_44027);
nor U47899 (N_47899,N_44897,N_44296);
or U47900 (N_47900,N_44148,N_45571);
and U47901 (N_47901,N_44218,N_45170);
nand U47902 (N_47902,N_44895,N_45053);
or U47903 (N_47903,N_44624,N_44764);
xor U47904 (N_47904,N_44828,N_44892);
nand U47905 (N_47905,N_44984,N_45519);
and U47906 (N_47906,N_44628,N_44497);
xnor U47907 (N_47907,N_45680,N_44427);
nor U47908 (N_47908,N_45841,N_45074);
nand U47909 (N_47909,N_44869,N_44457);
and U47910 (N_47910,N_45767,N_44436);
nand U47911 (N_47911,N_44139,N_45859);
nand U47912 (N_47912,N_44235,N_45232);
and U47913 (N_47913,N_44095,N_45971);
nor U47914 (N_47914,N_45211,N_45559);
and U47915 (N_47915,N_44670,N_45835);
or U47916 (N_47916,N_44352,N_44910);
nand U47917 (N_47917,N_44927,N_45366);
and U47918 (N_47918,N_44057,N_45963);
nand U47919 (N_47919,N_44783,N_45065);
xor U47920 (N_47920,N_45888,N_45159);
nand U47921 (N_47921,N_45673,N_45217);
xor U47922 (N_47922,N_45987,N_44715);
nand U47923 (N_47923,N_45572,N_45734);
and U47924 (N_47924,N_45303,N_44254);
or U47925 (N_47925,N_44212,N_44805);
or U47926 (N_47926,N_45613,N_45770);
or U47927 (N_47927,N_45528,N_45333);
nor U47928 (N_47928,N_45218,N_44511);
or U47929 (N_47929,N_44072,N_45111);
nor U47930 (N_47930,N_44184,N_44707);
xor U47931 (N_47931,N_44142,N_45356);
or U47932 (N_47932,N_44019,N_45915);
and U47933 (N_47933,N_45292,N_44804);
or U47934 (N_47934,N_44329,N_44266);
nand U47935 (N_47935,N_45444,N_45438);
nand U47936 (N_47936,N_44550,N_45077);
nor U47937 (N_47937,N_45437,N_44543);
nor U47938 (N_47938,N_44351,N_45897);
xnor U47939 (N_47939,N_44318,N_44198);
and U47940 (N_47940,N_45247,N_45253);
or U47941 (N_47941,N_45102,N_45311);
or U47942 (N_47942,N_45903,N_45027);
nor U47943 (N_47943,N_44413,N_44685);
nor U47944 (N_47944,N_45323,N_44627);
xor U47945 (N_47945,N_44100,N_45264);
xnor U47946 (N_47946,N_44547,N_45981);
nand U47947 (N_47947,N_45101,N_45903);
or U47948 (N_47948,N_45486,N_44134);
nand U47949 (N_47949,N_44790,N_45161);
and U47950 (N_47950,N_44365,N_44113);
or U47951 (N_47951,N_44016,N_45295);
nand U47952 (N_47952,N_45134,N_45196);
nor U47953 (N_47953,N_45546,N_44248);
nand U47954 (N_47954,N_45986,N_44116);
and U47955 (N_47955,N_45243,N_44485);
xor U47956 (N_47956,N_44737,N_45539);
nand U47957 (N_47957,N_45041,N_45815);
or U47958 (N_47958,N_44117,N_45166);
xnor U47959 (N_47959,N_45890,N_45004);
xor U47960 (N_47960,N_44494,N_44193);
nand U47961 (N_47961,N_44049,N_45007);
and U47962 (N_47962,N_44451,N_45455);
nor U47963 (N_47963,N_44079,N_45368);
nand U47964 (N_47964,N_44335,N_44391);
and U47965 (N_47965,N_45687,N_45093);
xnor U47966 (N_47966,N_45036,N_44087);
and U47967 (N_47967,N_44355,N_45927);
nand U47968 (N_47968,N_44609,N_45897);
and U47969 (N_47969,N_45846,N_45880);
nand U47970 (N_47970,N_45864,N_44883);
nand U47971 (N_47971,N_44659,N_45053);
or U47972 (N_47972,N_44025,N_44180);
or U47973 (N_47973,N_44833,N_44243);
or U47974 (N_47974,N_44038,N_45255);
nand U47975 (N_47975,N_45824,N_44443);
and U47976 (N_47976,N_45822,N_44995);
xnor U47977 (N_47977,N_44152,N_44162);
nand U47978 (N_47978,N_45435,N_45026);
nor U47979 (N_47979,N_44707,N_44726);
and U47980 (N_47980,N_44481,N_44556);
nor U47981 (N_47981,N_45609,N_44528);
nor U47982 (N_47982,N_45998,N_44105);
or U47983 (N_47983,N_44793,N_44534);
nand U47984 (N_47984,N_45186,N_45427);
and U47985 (N_47985,N_44361,N_45956);
xnor U47986 (N_47986,N_45529,N_44564);
xnor U47987 (N_47987,N_45135,N_44833);
nand U47988 (N_47988,N_44833,N_44088);
nor U47989 (N_47989,N_44473,N_44751);
xor U47990 (N_47990,N_45559,N_45610);
nor U47991 (N_47991,N_44389,N_45616);
and U47992 (N_47992,N_45400,N_45951);
nor U47993 (N_47993,N_44700,N_44032);
and U47994 (N_47994,N_44554,N_44009);
xor U47995 (N_47995,N_44424,N_45652);
nand U47996 (N_47996,N_45212,N_44356);
nand U47997 (N_47997,N_44165,N_44229);
nor U47998 (N_47998,N_44663,N_44226);
xnor U47999 (N_47999,N_44031,N_44825);
or U48000 (N_48000,N_46307,N_47182);
nand U48001 (N_48001,N_46829,N_46702);
nor U48002 (N_48002,N_47265,N_46860);
nand U48003 (N_48003,N_47143,N_46556);
and U48004 (N_48004,N_46792,N_46077);
and U48005 (N_48005,N_46318,N_47199);
xor U48006 (N_48006,N_46636,N_46946);
nor U48007 (N_48007,N_47363,N_47141);
nand U48008 (N_48008,N_47628,N_47658);
xnor U48009 (N_48009,N_47942,N_47772);
nand U48010 (N_48010,N_47682,N_46156);
and U48011 (N_48011,N_47513,N_47410);
xor U48012 (N_48012,N_46424,N_46930);
and U48013 (N_48013,N_47538,N_46907);
or U48014 (N_48014,N_47178,N_47024);
nor U48015 (N_48015,N_47999,N_47471);
nand U48016 (N_48016,N_47689,N_47277);
or U48017 (N_48017,N_46580,N_47960);
and U48018 (N_48018,N_46087,N_47381);
and U48019 (N_48019,N_47710,N_46145);
nor U48020 (N_48020,N_47519,N_47261);
xnor U48021 (N_48021,N_47493,N_47430);
and U48022 (N_48022,N_46102,N_47859);
and U48023 (N_48023,N_46836,N_47864);
xnor U48024 (N_48024,N_47762,N_47070);
and U48025 (N_48025,N_47729,N_46088);
nand U48026 (N_48026,N_46328,N_46004);
or U48027 (N_48027,N_47985,N_46308);
or U48028 (N_48028,N_47019,N_46669);
and U48029 (N_48029,N_47338,N_47606);
nand U48030 (N_48030,N_47631,N_46058);
nand U48031 (N_48031,N_47703,N_46412);
and U48032 (N_48032,N_46182,N_47723);
nand U48033 (N_48033,N_47680,N_46996);
xor U48034 (N_48034,N_46014,N_46715);
xor U48035 (N_48035,N_46039,N_47695);
xnor U48036 (N_48036,N_46271,N_47622);
or U48037 (N_48037,N_47986,N_47262);
nor U48038 (N_48038,N_47115,N_46713);
nand U48039 (N_48039,N_46236,N_46413);
or U48040 (N_48040,N_46332,N_47624);
nand U48041 (N_48041,N_47349,N_47755);
xor U48042 (N_48042,N_46223,N_47328);
and U48043 (N_48043,N_46148,N_47061);
nand U48044 (N_48044,N_46871,N_46176);
or U48045 (N_48045,N_46422,N_46588);
xnor U48046 (N_48046,N_47207,N_46289);
xnor U48047 (N_48047,N_47092,N_47874);
and U48048 (N_48048,N_47260,N_46602);
or U48049 (N_48049,N_46681,N_47868);
nor U48050 (N_48050,N_47116,N_46431);
and U48051 (N_48051,N_46734,N_47078);
and U48052 (N_48052,N_46514,N_47018);
nand U48053 (N_48053,N_46352,N_47322);
and U48054 (N_48054,N_47768,N_46870);
and U48055 (N_48055,N_46754,N_47004);
nor U48056 (N_48056,N_47201,N_46900);
or U48057 (N_48057,N_46915,N_47975);
and U48058 (N_48058,N_46293,N_46187);
nor U48059 (N_48059,N_46017,N_46130);
xor U48060 (N_48060,N_47095,N_47733);
xnor U48061 (N_48061,N_47777,N_47648);
and U48062 (N_48062,N_46587,N_46643);
xor U48063 (N_48063,N_47066,N_47692);
xnor U48064 (N_48064,N_46274,N_46408);
xor U48065 (N_48065,N_46692,N_46767);
xor U48066 (N_48066,N_47323,N_47367);
nor U48067 (N_48067,N_47039,N_47884);
nand U48068 (N_48068,N_47020,N_47091);
nand U48069 (N_48069,N_46095,N_47717);
nand U48070 (N_48070,N_47104,N_47219);
nor U48071 (N_48071,N_47094,N_46158);
or U48072 (N_48072,N_46262,N_46582);
nor U48073 (N_48073,N_46801,N_46820);
or U48074 (N_48074,N_46344,N_46482);
nand U48075 (N_48075,N_47973,N_47785);
and U48076 (N_48076,N_46208,N_46876);
nand U48077 (N_48077,N_46195,N_46065);
or U48078 (N_48078,N_46761,N_47077);
and U48079 (N_48079,N_46106,N_46673);
or U48080 (N_48080,N_46697,N_46638);
nand U48081 (N_48081,N_47337,N_46265);
nor U48082 (N_48082,N_46085,N_46654);
nor U48083 (N_48083,N_46722,N_47280);
nand U48084 (N_48084,N_47734,N_46656);
and U48085 (N_48085,N_46938,N_47279);
or U48086 (N_48086,N_46320,N_47840);
or U48087 (N_48087,N_47636,N_47394);
nor U48088 (N_48088,N_47283,N_46802);
nor U48089 (N_48089,N_46567,N_46611);
and U48090 (N_48090,N_47368,N_47882);
nor U48091 (N_48091,N_47854,N_47064);
and U48092 (N_48092,N_47467,N_46120);
and U48093 (N_48093,N_47657,N_46239);
nor U48094 (N_48094,N_46585,N_46159);
or U48095 (N_48095,N_46943,N_46969);
nor U48096 (N_48096,N_46126,N_47312);
or U48097 (N_48097,N_47997,N_47102);
xnor U48098 (N_48098,N_46841,N_46407);
xor U48099 (N_48099,N_46859,N_47415);
and U48100 (N_48100,N_47005,N_46693);
nand U48101 (N_48101,N_46502,N_47883);
nand U48102 (N_48102,N_47525,N_47751);
nor U48103 (N_48103,N_46748,N_46746);
nor U48104 (N_48104,N_46132,N_47998);
and U48105 (N_48105,N_46745,N_46062);
nor U48106 (N_48106,N_47915,N_47118);
or U48107 (N_48107,N_46140,N_47305);
xor U48108 (N_48108,N_47914,N_47294);
or U48109 (N_48109,N_46434,N_47730);
xnor U48110 (N_48110,N_47351,N_47111);
xor U48111 (N_48111,N_47902,N_47093);
xor U48112 (N_48112,N_47870,N_46224);
or U48113 (N_48113,N_46565,N_47524);
nand U48114 (N_48114,N_47907,N_46649);
nand U48115 (N_48115,N_46546,N_47802);
xnor U48116 (N_48116,N_46566,N_47107);
xor U48117 (N_48117,N_47167,N_47575);
nor U48118 (N_48118,N_47954,N_47520);
nor U48119 (N_48119,N_47809,N_47523);
and U48120 (N_48120,N_47278,N_47567);
nor U48121 (N_48121,N_47925,N_46368);
nor U48122 (N_48122,N_46980,N_47983);
and U48123 (N_48123,N_46939,N_46389);
or U48124 (N_48124,N_47849,N_46618);
nor U48125 (N_48125,N_47675,N_46338);
or U48126 (N_48126,N_47736,N_46861);
nand U48127 (N_48127,N_47812,N_47900);
or U48128 (N_48128,N_46789,N_46916);
nor U48129 (N_48129,N_46622,N_47617);
nor U48130 (N_48130,N_46286,N_46315);
nand U48131 (N_48131,N_46612,N_46167);
nand U48132 (N_48132,N_47568,N_47041);
and U48133 (N_48133,N_46460,N_46592);
and U48134 (N_48134,N_46682,N_47597);
or U48135 (N_48135,N_47741,N_47379);
nor U48136 (N_48136,N_47578,N_46282);
nor U48137 (N_48137,N_46506,N_46775);
xnor U48138 (N_48138,N_46849,N_46152);
nor U48139 (N_48139,N_46272,N_47805);
xor U48140 (N_48140,N_47535,N_47784);
nor U48141 (N_48141,N_47579,N_47159);
and U48142 (N_48142,N_46312,N_46259);
nor U48143 (N_48143,N_46735,N_46909);
or U48144 (N_48144,N_46207,N_47258);
nor U48145 (N_48145,N_46816,N_46326);
or U48146 (N_48146,N_46908,N_46512);
and U48147 (N_48147,N_47359,N_46711);
nand U48148 (N_48148,N_46586,N_46114);
or U48149 (N_48149,N_46363,N_47635);
and U48150 (N_48150,N_46350,N_46658);
xnor U48151 (N_48151,N_47711,N_47639);
and U48152 (N_48152,N_47724,N_46927);
nor U48153 (N_48153,N_47477,N_47487);
or U48154 (N_48154,N_47296,N_46401);
nor U48155 (N_48155,N_46015,N_47082);
nor U48156 (N_48156,N_46064,N_46013);
nand U48157 (N_48157,N_47853,N_46942);
xnor U48158 (N_48158,N_46978,N_46624);
and U48159 (N_48159,N_47715,N_46743);
xor U48160 (N_48160,N_47508,N_46881);
nand U48161 (N_48161,N_46610,N_46022);
xor U48162 (N_48162,N_47042,N_46241);
and U48163 (N_48163,N_46222,N_47652);
and U48164 (N_48164,N_46299,N_46552);
or U48165 (N_48165,N_47592,N_47456);
nor U48166 (N_48166,N_47509,N_46304);
nor U48167 (N_48167,N_47128,N_46897);
nand U48168 (N_48168,N_46119,N_47079);
xor U48169 (N_48169,N_47289,N_47681);
nand U48170 (N_48170,N_46772,N_47901);
and U48171 (N_48171,N_47310,N_47284);
nor U48172 (N_48172,N_47282,N_47946);
xnor U48173 (N_48173,N_46008,N_47129);
and U48174 (N_48174,N_47320,N_47237);
nand U48175 (N_48175,N_46548,N_46477);
or U48176 (N_48176,N_46986,N_46420);
or U48177 (N_48177,N_47259,N_46827);
or U48178 (N_48178,N_46740,N_46979);
or U48179 (N_48179,N_47881,N_47684);
xnor U48180 (N_48180,N_46832,N_47197);
or U48181 (N_48181,N_47439,N_47669);
nor U48182 (N_48182,N_47123,N_46717);
and U48183 (N_48183,N_47164,N_47062);
xnor U48184 (N_48184,N_46519,N_46281);
or U48185 (N_48185,N_46472,N_47132);
and U48186 (N_48186,N_46071,N_46079);
nor U48187 (N_48187,N_46024,N_47562);
and U48188 (N_48188,N_46788,N_46601);
xnor U48189 (N_48189,N_46887,N_46052);
or U48190 (N_48190,N_47352,N_46982);
xnor U48191 (N_48191,N_47887,N_47056);
or U48192 (N_48192,N_47268,N_46616);
or U48193 (N_48193,N_46518,N_46003);
or U48194 (N_48194,N_46410,N_47555);
nor U48195 (N_48195,N_46822,N_46421);
nor U48196 (N_48196,N_46497,N_47701);
and U48197 (N_48197,N_46254,N_46992);
or U48198 (N_48198,N_47945,N_46009);
nand U48199 (N_48199,N_47676,N_47748);
nor U48200 (N_48200,N_46521,N_46354);
or U48201 (N_48201,N_47651,N_47926);
xor U48202 (N_48202,N_46409,N_46342);
and U48203 (N_48203,N_46764,N_46090);
nor U48204 (N_48204,N_46296,N_47503);
and U48205 (N_48205,N_46139,N_46560);
nor U48206 (N_48206,N_46288,N_47440);
nor U48207 (N_48207,N_46457,N_46233);
nor U48208 (N_48208,N_47226,N_46183);
xor U48209 (N_48209,N_46667,N_47697);
or U48210 (N_48210,N_47362,N_46971);
and U48211 (N_48211,N_46781,N_46771);
and U48212 (N_48212,N_47889,N_46988);
and U48213 (N_48213,N_47667,N_47099);
xor U48214 (N_48214,N_47817,N_47637);
nor U48215 (N_48215,N_46203,N_46995);
or U48216 (N_48216,N_47895,N_46112);
xor U48217 (N_48217,N_47489,N_47463);
and U48218 (N_48218,N_46796,N_46600);
or U48219 (N_48219,N_47964,N_47690);
and U48220 (N_48220,N_47671,N_47819);
nor U48221 (N_48221,N_46301,N_47534);
nor U48222 (N_48222,N_47632,N_47458);
and U48223 (N_48223,N_46426,N_46813);
xor U48224 (N_48224,N_47878,N_46495);
nor U48225 (N_48225,N_46154,N_46739);
nand U48226 (N_48226,N_46977,N_47787);
or U48227 (N_48227,N_47659,N_46689);
and U48228 (N_48228,N_47786,N_46498);
and U48229 (N_48229,N_46635,N_47836);
and U48230 (N_48230,N_47827,N_47021);
or U48231 (N_48231,N_47416,N_47893);
or U48232 (N_48232,N_47758,N_46303);
nor U48233 (N_48233,N_46773,N_46337);
nand U48234 (N_48234,N_47443,N_46345);
or U48235 (N_48235,N_46261,N_47030);
nand U48236 (N_48236,N_47344,N_46068);
or U48237 (N_48237,N_47529,N_46736);
and U48238 (N_48238,N_46642,N_47700);
nand U48239 (N_48239,N_47557,N_46517);
nand U48240 (N_48240,N_47332,N_46650);
xnor U48241 (N_48241,N_47756,N_46554);
xor U48242 (N_48242,N_47565,N_47105);
xnor U48243 (N_48243,N_46089,N_46379);
xor U48244 (N_48244,N_47574,N_46672);
nand U48245 (N_48245,N_46808,N_46830);
xor U48246 (N_48246,N_47623,N_47331);
or U48247 (N_48247,N_47838,N_46339);
nor U48248 (N_48248,N_47497,N_46800);
and U48249 (N_48249,N_47502,N_47314);
and U48250 (N_48250,N_46553,N_47488);
xnor U48251 (N_48251,N_46425,N_46873);
and U48252 (N_48252,N_46967,N_46248);
nor U48253 (N_48253,N_47761,N_47453);
xor U48254 (N_48254,N_47372,N_46968);
nor U48255 (N_48255,N_46151,N_47913);
xor U48256 (N_48256,N_46049,N_47776);
xnor U48257 (N_48257,N_47770,N_46583);
nor U48258 (N_48258,N_46718,N_47022);
and U48259 (N_48259,N_46917,N_47273);
nor U48260 (N_48260,N_46509,N_47791);
nand U48261 (N_48261,N_47186,N_47297);
xnor U48262 (N_48262,N_47252,N_47457);
or U48263 (N_48263,N_46858,N_46851);
nor U48264 (N_48264,N_47494,N_47125);
xnor U48265 (N_48265,N_46125,N_46903);
nand U48266 (N_48266,N_46640,N_46284);
nor U48267 (N_48267,N_47154,N_47144);
xor U48268 (N_48268,N_46629,N_47820);
xnor U48269 (N_48269,N_46668,N_47345);
and U48270 (N_48270,N_46885,N_46507);
xnor U48271 (N_48271,N_47603,N_46061);
nand U48272 (N_48272,N_46442,N_47448);
nor U48273 (N_48273,N_46879,N_46138);
nor U48274 (N_48274,N_47974,N_47088);
xor U48275 (N_48275,N_47807,N_47798);
and U48276 (N_48276,N_47923,N_46235);
nand U48277 (N_48277,N_47293,N_46042);
and U48278 (N_48278,N_47605,N_46868);
nand U48279 (N_48279,N_47580,N_47043);
xnor U48280 (N_48280,N_47003,N_46486);
xor U48281 (N_48281,N_47561,N_47200);
nor U48282 (N_48282,N_46365,N_47090);
xor U48283 (N_48283,N_46824,N_46230);
nand U48284 (N_48284,N_47747,N_47187);
xnor U48285 (N_48285,N_47549,N_47403);
xor U48286 (N_48286,N_47988,N_47560);
nand U48287 (N_48287,N_46007,N_46795);
nor U48288 (N_48288,N_47384,N_46411);
nor U48289 (N_48289,N_46378,N_47743);
nand U48290 (N_48290,N_46807,N_46825);
or U48291 (N_48291,N_47364,N_46200);
and U48292 (N_48292,N_46291,N_46229);
and U48293 (N_48293,N_46645,N_47204);
and U48294 (N_48294,N_47609,N_46314);
nor U48295 (N_48295,N_46755,N_47444);
and U48296 (N_48296,N_46277,N_46021);
or U48297 (N_48297,N_47135,N_47928);
and U48298 (N_48298,N_46057,N_46309);
nand U48299 (N_48299,N_47220,N_46446);
nor U48300 (N_48300,N_47546,N_47202);
and U48301 (N_48301,N_47190,N_47112);
nor U48302 (N_48302,N_47388,N_46972);
nor U48303 (N_48303,N_46921,N_47131);
nand U48304 (N_48304,N_47335,N_46295);
xnor U48305 (N_48305,N_46720,N_46137);
or U48306 (N_48306,N_47140,N_46104);
nand U48307 (N_48307,N_47959,N_47674);
xor U48308 (N_48308,N_46542,N_47234);
nand U48309 (N_48309,N_47542,N_47499);
nand U48310 (N_48310,N_46578,N_47387);
or U48311 (N_48311,N_47963,N_46330);
xor U48312 (N_48312,N_47891,N_46465);
and U48313 (N_48313,N_47516,N_46430);
or U48314 (N_48314,N_46564,N_47894);
nand U48315 (N_48315,N_47012,N_46853);
and U48316 (N_48316,N_47506,N_46310);
or U48317 (N_48317,N_46956,N_47006);
xor U48318 (N_48318,N_46346,N_47712);
nand U48319 (N_48319,N_47446,N_46540);
nand U48320 (N_48320,N_46703,N_46780);
xnor U48321 (N_48321,N_46516,N_47475);
nor U48322 (N_48322,N_47414,N_46627);
xnor U48323 (N_48323,N_46931,N_47081);
and U48324 (N_48324,N_47057,N_46854);
nand U48325 (N_48325,N_46439,N_47570);
and U48326 (N_48326,N_46957,N_47653);
and U48327 (N_48327,N_47539,N_46249);
nor U48328 (N_48328,N_47627,N_46247);
or U48329 (N_48329,N_46467,N_46144);
or U48330 (N_48330,N_47452,N_47984);
nor U48331 (N_48331,N_47841,N_46628);
nor U48332 (N_48332,N_47833,N_47530);
nor U48333 (N_48333,N_47329,N_47354);
nor U48334 (N_48334,N_46835,N_47350);
nand U48335 (N_48335,N_46597,N_46016);
nand U48336 (N_48336,N_47319,N_47302);
or U48337 (N_48337,N_46856,N_46489);
and U48338 (N_48338,N_46614,N_46245);
or U48339 (N_48339,N_46877,N_46768);
and U48340 (N_48340,N_46894,N_46710);
nand U48341 (N_48341,N_46663,N_46226);
or U48342 (N_48342,N_47767,N_46698);
nand U48343 (N_48343,N_46402,N_47334);
or U48344 (N_48344,N_47716,N_47011);
nand U48345 (N_48345,N_47968,N_46466);
xnor U48346 (N_48346,N_47573,N_46216);
xor U48347 (N_48347,N_47391,N_46581);
or U48348 (N_48348,N_47917,N_46406);
nand U48349 (N_48349,N_46899,N_46384);
and U48350 (N_48350,N_46175,N_46505);
nand U48351 (N_48351,N_46633,N_47994);
xnor U48352 (N_48352,N_47462,N_46347);
nand U48353 (N_48353,N_46846,N_47673);
or U48354 (N_48354,N_47205,N_47233);
nor U48355 (N_48355,N_46108,N_47848);
nand U48356 (N_48356,N_47466,N_47225);
and U48357 (N_48357,N_46960,N_46081);
nor U48358 (N_48358,N_46129,N_47735);
xnor U48359 (N_48359,N_47348,N_46092);
or U48360 (N_48360,N_47427,N_47356);
nor U48361 (N_48361,N_47947,N_46059);
or U48362 (N_48362,N_47906,N_46018);
xnor U48363 (N_48363,N_46043,N_47792);
nor U48364 (N_48364,N_47537,N_47185);
and U48365 (N_48365,N_47569,N_47972);
and U48366 (N_48366,N_47825,N_47879);
nand U48367 (N_48367,N_46173,N_47655);
or U48368 (N_48368,N_47342,N_47179);
and U48369 (N_48369,N_47377,N_47438);
and U48370 (N_48370,N_47548,N_46741);
nand U48371 (N_48371,N_47275,N_47707);
nand U48372 (N_48372,N_47604,N_46926);
and U48373 (N_48373,N_47801,N_47845);
nor U48374 (N_48374,N_46932,N_46515);
or U48375 (N_48375,N_46591,N_47670);
nor U48376 (N_48376,N_46723,N_47993);
nand U48377 (N_48377,N_47980,N_46237);
nor U48378 (N_48378,N_47068,N_46532);
or U48379 (N_48379,N_47382,N_47905);
nand U48380 (N_48380,N_47424,N_46026);
xor U48381 (N_48381,N_47656,N_46607);
or U48382 (N_48382,N_47232,N_46372);
or U48383 (N_48383,N_47647,N_46452);
or U48384 (N_48384,N_47392,N_47922);
and U48385 (N_48385,N_46010,N_47428);
xnor U48386 (N_48386,N_47961,N_46811);
nand U48387 (N_48387,N_47484,N_46561);
nand U48388 (N_48388,N_47654,N_47436);
nand U48389 (N_48389,N_46044,N_47230);
nand U48390 (N_48390,N_47396,N_46950);
xor U48391 (N_48391,N_47754,N_46527);
or U48392 (N_48392,N_46302,N_47120);
xnor U48393 (N_48393,N_46762,N_46273);
nor U48394 (N_48394,N_47732,N_47031);
xnor U48395 (N_48395,N_47029,N_46766);
or U48396 (N_48396,N_47445,N_47970);
and U48397 (N_48397,N_47113,N_46845);
or U48398 (N_48398,N_46965,N_46122);
and U48399 (N_48399,N_46370,N_47704);
or U48400 (N_48400,N_47270,N_46324);
nor U48401 (N_48401,N_46544,N_47172);
and U48402 (N_48402,N_46604,N_47492);
or U48403 (N_48403,N_47939,N_46572);
and U48404 (N_48404,N_46250,N_47110);
nand U48405 (N_48405,N_47799,N_47844);
and U48406 (N_48406,N_46925,N_47165);
nor U48407 (N_48407,N_47087,N_47152);
nor U48408 (N_48408,N_46695,N_46278);
or U48409 (N_48409,N_46691,N_46983);
xnor U48410 (N_48410,N_47324,N_47393);
xnor U48411 (N_48411,N_47927,N_47124);
xnor U48412 (N_48412,N_47249,N_46797);
or U48413 (N_48413,N_47325,N_46889);
or U48414 (N_48414,N_47369,N_47666);
nand U48415 (N_48415,N_46919,N_47221);
and U48416 (N_48416,N_47137,N_46367);
xnor U48417 (N_48417,N_47514,N_47935);
nor U48418 (N_48418,N_46810,N_47979);
nor U48419 (N_48419,N_46360,N_46400);
nor U48420 (N_48420,N_47346,N_47757);
nor U48421 (N_48421,N_47480,N_47683);
xor U48422 (N_48422,N_46419,N_47134);
nor U48423 (N_48423,N_46625,N_47694);
nand U48424 (N_48424,N_46630,N_47083);
xor U48425 (N_48425,N_47114,N_47739);
nand U48426 (N_48426,N_46869,N_47050);
xor U48427 (N_48427,N_46989,N_46571);
nor U48428 (N_48428,N_47290,N_46082);
or U48429 (N_48429,N_47281,N_46670);
nor U48430 (N_48430,N_46666,N_46496);
and U48431 (N_48431,N_46416,N_46392);
and U48432 (N_48432,N_47048,N_47130);
or U48433 (N_48433,N_47545,N_47584);
and U48434 (N_48434,N_47184,N_47254);
nor U48435 (N_48435,N_47815,N_47912);
nand U48436 (N_48436,N_47442,N_46415);
nor U48437 (N_48437,N_46317,N_47419);
xnor U48438 (N_48438,N_46644,N_46492);
and U48439 (N_48439,N_46074,N_46714);
nand U48440 (N_48440,N_46776,N_47371);
nand U48441 (N_48441,N_46242,N_47850);
nand U48442 (N_48442,N_47175,N_46892);
xnor U48443 (N_48443,N_46169,N_46511);
nand U48444 (N_48444,N_47663,N_46657);
and U48445 (N_48445,N_47528,N_47872);
or U48446 (N_48446,N_46923,N_47903);
nor U48447 (N_48447,N_46481,N_47242);
or U48448 (N_48448,N_47588,N_46440);
and U48449 (N_48449,N_46056,N_46450);
nor U48450 (N_48450,N_47067,N_47223);
or U48451 (N_48451,N_46298,N_46751);
and U48452 (N_48452,N_46047,N_47714);
or U48453 (N_48453,N_46852,N_47981);
or U48454 (N_48454,N_47846,N_47750);
or U48455 (N_48455,N_46471,N_47407);
xor U48456 (N_48456,N_46866,N_46545);
nor U48457 (N_48457,N_46549,N_47978);
nand U48458 (N_48458,N_46355,N_47507);
and U48459 (N_48459,N_46403,N_47842);
nand U48460 (N_48460,N_46744,N_47089);
and U48461 (N_48461,N_46435,N_47235);
xor U48462 (N_48462,N_46316,N_47992);
xor U48463 (N_48463,N_46478,N_47590);
nor U48464 (N_48464,N_46340,N_46508);
and U48465 (N_48465,N_47619,N_47047);
xor U48466 (N_48466,N_47765,N_46311);
xor U48467 (N_48467,N_47989,N_47073);
nand U48468 (N_48468,N_46865,N_46387);
nand U48469 (N_48469,N_47286,N_46660);
nor U48470 (N_48470,N_46048,N_47869);
xor U48471 (N_48471,N_47899,N_46834);
or U48472 (N_48472,N_46902,N_47620);
and U48473 (N_48473,N_47100,N_47937);
xor U48474 (N_48474,N_47991,N_46963);
xnor U48475 (N_48475,N_47586,N_47313);
nand U48476 (N_48476,N_46170,N_47188);
or U48477 (N_48477,N_47409,N_47829);
nand U48478 (N_48478,N_47413,N_47591);
nor U48479 (N_48479,N_47934,N_47433);
or U48480 (N_48480,N_46674,N_47543);
or U48481 (N_48481,N_47532,N_47035);
nand U48482 (N_48482,N_47383,N_47518);
xor U48483 (N_48483,N_46051,N_46763);
or U48484 (N_48484,N_46940,N_46733);
nand U48485 (N_48485,N_47071,N_47481);
xnor U48486 (N_48486,N_46987,N_46256);
xor U48487 (N_48487,N_47630,N_46475);
nor U48488 (N_48488,N_47847,N_46041);
and U48489 (N_48489,N_46197,N_46898);
xor U48490 (N_48490,N_46385,N_46194);
nor U48491 (N_48491,N_46031,N_47417);
xnor U48492 (N_48492,N_46884,N_47243);
and U48493 (N_48493,N_47885,N_46264);
nor U48494 (N_48494,N_46040,N_46091);
xnor U48495 (N_48495,N_46747,N_47361);
or U48496 (N_48496,N_47217,N_47036);
xnor U48497 (N_48497,N_46033,N_46805);
or U48498 (N_48498,N_47257,N_47517);
nand U48499 (N_48499,N_47782,N_47272);
nor U48500 (N_48500,N_47032,N_47054);
xnor U48501 (N_48501,N_46445,N_47491);
or U48502 (N_48502,N_46462,N_46476);
nor U48503 (N_48503,N_46598,N_47418);
xnor U48504 (N_48504,N_46959,N_46929);
or U48505 (N_48505,N_46113,N_46263);
xnor U48506 (N_48506,N_47357,N_47058);
nand U48507 (N_48507,N_46212,N_47303);
nor U48508 (N_48508,N_46949,N_47174);
nor U48509 (N_48509,N_46134,N_47162);
or U48510 (N_48510,N_46253,N_47145);
and U48511 (N_48511,N_47789,N_47823);
nor U48512 (N_48512,N_46685,N_47826);
and U48513 (N_48513,N_46890,N_46099);
nor U48514 (N_48514,N_47911,N_46493);
or U48515 (N_48515,N_46321,N_46218);
nand U48516 (N_48516,N_47008,N_46002);
nor U48517 (N_48517,N_47795,N_47940);
or U48518 (N_48518,N_47098,N_46405);
nand U48519 (N_48519,N_46716,N_47218);
and U48520 (N_48520,N_46124,N_46267);
xnor U48521 (N_48521,N_46162,N_46178);
and U48522 (N_48522,N_46027,N_46255);
nor U48523 (N_48523,N_47176,N_47390);
and U48524 (N_48524,N_47097,N_46123);
xor U48525 (N_48525,N_47828,N_47483);
or U48526 (N_48526,N_47126,N_47298);
nor U48527 (N_48527,N_46180,N_46231);
nor U48528 (N_48528,N_47300,N_47771);
and U48529 (N_48529,N_47752,N_47469);
nor U48530 (N_48530,N_46687,N_46055);
or U48531 (N_48531,N_46053,N_47559);
nor U48532 (N_48532,N_46880,N_47608);
or U48533 (N_48533,N_47434,N_47149);
nor U48534 (N_48534,N_47918,N_47856);
or U48535 (N_48535,N_46793,N_46809);
xnor U48536 (N_48536,N_46454,N_46913);
nor U48537 (N_48537,N_46904,N_46444);
or U48538 (N_48538,N_46914,N_46525);
and U48539 (N_48539,N_47995,N_46785);
nor U48540 (N_48540,N_47192,N_47025);
nor U48541 (N_48541,N_46671,N_46447);
nand U48542 (N_48542,N_47295,N_47193);
nor U48543 (N_48543,N_47191,N_46107);
nand U48544 (N_48544,N_47380,N_47614);
nor U48545 (N_48545,N_46276,N_47610);
xor U48546 (N_48546,N_46404,N_47157);
nor U48547 (N_48547,N_46470,N_47247);
xor U48548 (N_48548,N_47727,N_46819);
xor U48549 (N_48549,N_47411,N_47737);
and U48550 (N_48550,N_46599,N_46543);
nor U48551 (N_48551,N_47397,N_47626);
or U48552 (N_48552,N_46181,N_46069);
and U48553 (N_48553,N_46150,N_46101);
nor U48554 (N_48554,N_47304,N_46727);
xnor U48555 (N_48555,N_47400,N_46161);
and U48556 (N_48556,N_46997,N_46066);
and U48557 (N_48557,N_46110,N_47121);
and U48558 (N_48558,N_47055,N_46955);
xor U48559 (N_48559,N_46990,N_46905);
nand U48560 (N_48560,N_47521,N_47059);
nand U48561 (N_48561,N_46569,N_47336);
xnor U48562 (N_48562,N_47450,N_47691);
and U48563 (N_48563,N_47274,N_46103);
nor U48564 (N_48564,N_47171,N_47010);
nor U48565 (N_48565,N_47951,N_46974);
nor U48566 (N_48566,N_46752,N_47080);
nand U48567 (N_48567,N_46127,N_46855);
nand U48568 (N_48568,N_46641,N_47797);
or U48569 (N_48569,N_46652,N_46157);
xnor U48570 (N_48570,N_47180,N_47209);
or U48571 (N_48571,N_46252,N_46779);
xor U48572 (N_48572,N_47811,N_46750);
or U48573 (N_48573,N_47028,N_46678);
or U48574 (N_48574,N_47287,N_47189);
xnor U48575 (N_48575,N_47589,N_47526);
xnor U48576 (N_48576,N_47101,N_46937);
nand U48577 (N_48577,N_46818,N_47522);
nor U48578 (N_48578,N_46563,N_46688);
nor U48579 (N_48579,N_46562,N_47183);
xor U48580 (N_48580,N_47117,N_47916);
xor U48581 (N_48581,N_46232,N_46953);
nand U48582 (N_48582,N_46958,N_47780);
nand U48583 (N_48583,N_46351,N_46070);
xor U48584 (N_48584,N_46883,N_46783);
or U48585 (N_48585,N_47422,N_46381);
nand U48586 (N_48586,N_47698,N_47343);
xor U48587 (N_48587,N_47027,N_46488);
xor U48588 (N_48588,N_46025,N_47766);
and U48589 (N_48589,N_47742,N_46596);
or U48590 (N_48590,N_47211,N_46319);
and U48591 (N_48591,N_46244,N_47625);
and U48592 (N_48592,N_47593,N_46786);
or U48593 (N_48593,N_47084,N_47686);
and U48594 (N_48594,N_46886,N_47536);
and U48595 (N_48595,N_46128,N_46238);
or U48596 (N_48596,N_46487,N_47227);
nand U48597 (N_48597,N_47309,N_47987);
and U48598 (N_48598,N_46831,N_47166);
or U48599 (N_48599,N_47229,N_46221);
or U48600 (N_48600,N_47880,N_46473);
nand U48601 (N_48601,N_47800,N_46006);
nor U48602 (N_48602,N_46922,N_46211);
or U48603 (N_48603,N_47642,N_46700);
xor U48604 (N_48604,N_46522,N_46464);
or U48605 (N_48605,N_46655,N_46358);
nor U48606 (N_48606,N_46414,N_46847);
xor U48607 (N_48607,N_47746,N_47932);
or U48608 (N_48608,N_46035,N_46258);
nand U48609 (N_48609,N_46948,N_46459);
xnor U48610 (N_48610,N_46976,N_46313);
or U48611 (N_48611,N_46821,N_47753);
or U48612 (N_48612,N_47231,N_46437);
xor U48613 (N_48613,N_46133,N_46147);
or U48614 (N_48614,N_46962,N_47550);
xnor U48615 (N_48615,N_47386,N_47276);
nand U48616 (N_48616,N_46054,N_47096);
nand U48617 (N_48617,N_46036,N_46290);
nand U48618 (N_48618,N_46177,N_46323);
or U48619 (N_48619,N_47339,N_47327);
or U48620 (N_48620,N_46185,N_46111);
and U48621 (N_48621,N_46292,N_46012);
nor U48622 (N_48622,N_46076,N_46875);
or U48623 (N_48623,N_46973,N_46395);
xor U48624 (N_48624,N_46882,N_46341);
and U48625 (N_48625,N_47074,N_47618);
nor U48626 (N_48626,N_46664,N_46528);
nor U48627 (N_48627,N_47460,N_47950);
xor U48628 (N_48628,N_46679,N_46353);
nor U48629 (N_48629,N_47389,N_46117);
and U48630 (N_48630,N_47366,N_47429);
xor U48631 (N_48631,N_46838,N_46732);
nand U48632 (N_48632,N_46028,N_46260);
and U48633 (N_48633,N_46329,N_46706);
and U48634 (N_48634,N_47699,N_47236);
nand U48635 (N_48635,N_47924,N_47702);
nand U48636 (N_48636,N_46961,N_47949);
xor U48637 (N_48637,N_46864,N_47616);
xor U48638 (N_48638,N_47037,N_47955);
nand U48639 (N_48639,N_47640,N_46060);
or U48640 (N_48640,N_47775,N_46201);
and U48641 (N_48641,N_46608,N_46626);
or U48642 (N_48642,N_46823,N_47170);
or U48643 (N_48643,N_47472,N_46171);
or U48644 (N_48644,N_46981,N_47957);
nand U48645 (N_48645,N_46398,N_47245);
nand U48646 (N_48646,N_46455,N_46383);
xor U48647 (N_48647,N_46484,N_47553);
or U48648 (N_48648,N_47615,N_47228);
or U48649 (N_48649,N_46738,N_46533);
xnor U48650 (N_48650,N_46615,N_47696);
nand U48651 (N_48651,N_46559,N_47496);
and U48652 (N_48652,N_46388,N_47046);
and U48653 (N_48653,N_47596,N_47285);
nand U48654 (N_48654,N_47793,N_46550);
xor U48655 (N_48655,N_46270,N_47783);
nand U48656 (N_48656,N_46034,N_47634);
nand U48657 (N_48657,N_46680,N_47919);
nor U48658 (N_48658,N_47468,N_46192);
nand U48659 (N_48659,N_47613,N_46651);
nor U48660 (N_48660,N_47896,N_47774);
or U48661 (N_48661,N_47929,N_46494);
nand U48662 (N_48662,N_47572,N_46479);
nand U48663 (N_48663,N_47541,N_46357);
nor U48664 (N_48664,N_46382,N_47086);
or U48665 (N_48665,N_46396,N_47540);
xnor U48666 (N_48666,N_46234,N_47421);
and U48667 (N_48667,N_47049,N_46524);
or U48668 (N_48668,N_47952,N_46888);
or U48669 (N_48669,N_46184,N_46593);
xor U48670 (N_48670,N_46531,N_46777);
nand U48671 (N_48671,N_47441,N_47943);
xnor U48672 (N_48672,N_47069,N_46731);
xnor U48673 (N_48673,N_46240,N_46828);
and U48674 (N_48674,N_47875,N_46196);
nand U48675 (N_48675,N_47412,N_46941);
nor U48676 (N_48676,N_46944,N_47944);
xnor U48677 (N_48677,N_47122,N_46376);
and U48678 (N_48678,N_46984,N_47060);
nor U48679 (N_48679,N_46453,N_46523);
nor U48680 (N_48680,N_46757,N_47544);
nor U48681 (N_48681,N_46708,N_46280);
xor U48682 (N_48682,N_47142,N_46924);
nand U48683 (N_48683,N_46046,N_46268);
nand U48684 (N_48684,N_47398,N_46266);
and U48685 (N_48685,N_47063,N_46574);
and U48686 (N_48686,N_47824,N_47023);
and U48687 (N_48687,N_46555,N_47085);
nor U48688 (N_48688,N_46335,N_47725);
xor U48689 (N_48689,N_46621,N_47976);
or U48690 (N_48690,N_47498,N_47244);
nor U48691 (N_48691,N_46970,N_47649);
nand U48692 (N_48692,N_46000,N_46765);
or U48693 (N_48693,N_46568,N_46966);
xnor U48694 (N_48694,N_47301,N_47476);
xor U48695 (N_48695,N_46443,N_46945);
nand U48696 (N_48696,N_46005,N_46998);
nor U48697 (N_48697,N_46637,N_46799);
nand U48698 (N_48698,N_46659,N_47679);
xnor U48699 (N_48699,N_46814,N_47146);
or U48700 (N_48700,N_46098,N_46530);
nand U48701 (N_48701,N_47395,N_46456);
nor U48702 (N_48702,N_46952,N_47133);
and U48703 (N_48703,N_47956,N_47904);
nand U48704 (N_48704,N_46803,N_46190);
or U48705 (N_48705,N_47370,N_47464);
nor U48706 (N_48706,N_46427,N_46217);
or U48707 (N_48707,N_47206,N_46878);
nand U48708 (N_48708,N_47109,N_47486);
nor U48709 (N_48709,N_47402,N_46210);
xnor U48710 (N_48710,N_46631,N_47718);
nand U48711 (N_48711,N_47358,N_47256);
nand U48712 (N_48712,N_46686,N_47399);
and U48713 (N_48713,N_46705,N_47076);
or U48714 (N_48714,N_47454,N_47852);
and U48715 (N_48715,N_46153,N_47892);
xnor U48716 (N_48716,N_47764,N_46458);
and U48717 (N_48717,N_46297,N_46215);
nor U48718 (N_48718,N_47248,N_46377);
or U48719 (N_48719,N_47479,N_47053);
or U48720 (N_48720,N_46118,N_46918);
and U48721 (N_48721,N_46469,N_47404);
and U48722 (N_48722,N_46724,N_46390);
or U48723 (N_48723,N_47401,N_47512);
or U48724 (N_48724,N_46595,N_46594);
and U48725 (N_48725,N_46843,N_47198);
nor U48726 (N_48726,N_46155,N_46219);
nor U48727 (N_48727,N_47693,N_47426);
xor U48728 (N_48728,N_47638,N_47646);
xor U48729 (N_48729,N_46534,N_46737);
nand U48730 (N_48730,N_46769,N_47222);
or U48731 (N_48731,N_46166,N_47360);
nor U48732 (N_48732,N_47251,N_47794);
xnor U48733 (N_48733,N_47898,N_47138);
nor U48734 (N_48734,N_47213,N_46225);
nand U48735 (N_48735,N_46030,N_46557);
xnor U48736 (N_48736,N_46149,N_47571);
nor U48737 (N_48737,N_46135,N_46160);
and U48738 (N_48738,N_47169,N_47238);
nor U48739 (N_48739,N_46993,N_47051);
and U48740 (N_48740,N_47431,N_47451);
nand U48741 (N_48741,N_46985,N_46143);
or U48742 (N_48742,N_46285,N_47585);
nand U48743 (N_48743,N_47455,N_46947);
xor U48744 (N_48744,N_47437,N_47818);
nor U48745 (N_48745,N_47478,N_47552);
xnor U48746 (N_48746,N_46300,N_47760);
nor U48747 (N_48747,N_46359,N_46753);
nor U48748 (N_48748,N_47645,N_46343);
nand U48749 (N_48749,N_46536,N_47321);
nand U48750 (N_48750,N_46366,N_47196);
and U48751 (N_48751,N_46934,N_47813);
or U48752 (N_48752,N_47435,N_47866);
xnor U48753 (N_48753,N_46842,N_46172);
xor U48754 (N_48754,N_47834,N_46806);
xor U48755 (N_48755,N_46333,N_47583);
or U48756 (N_48756,N_47504,N_46202);
and U48757 (N_48757,N_46369,N_47500);
xor U48758 (N_48758,N_47510,N_47678);
or U48759 (N_48759,N_46839,N_47977);
and U48760 (N_48760,N_47759,N_46725);
nand U48761 (N_48761,N_46449,N_46896);
or U48762 (N_48762,N_47153,N_47855);
and U48763 (N_48763,N_47447,N_47607);
nor U48764 (N_48764,N_47299,N_47558);
nor U48765 (N_48765,N_46920,N_47210);
or U48766 (N_48766,N_46662,N_47779);
nor U48767 (N_48767,N_46322,N_46573);
or U48768 (N_48768,N_46526,N_47485);
nor U48769 (N_48769,N_47598,N_46817);
nand U48770 (N_48770,N_46283,N_47966);
xnor U48771 (N_48771,N_47601,N_47072);
nor U48772 (N_48772,N_47788,N_47009);
or U48773 (N_48773,N_47007,N_47790);
or U48774 (N_48774,N_46417,N_47420);
and U48775 (N_48775,N_46500,N_47308);
nand U48776 (N_48776,N_46243,N_47688);
nand U48777 (N_48777,N_46485,N_47722);
nand U48778 (N_48778,N_47661,N_47650);
and U48779 (N_48779,N_47017,N_47195);
nand U48780 (N_48780,N_46146,N_46174);
nor U48781 (N_48781,N_47241,N_46951);
nor U48782 (N_48782,N_46246,N_47938);
and U48783 (N_48783,N_47713,N_47150);
xor U48784 (N_48784,N_46348,N_47594);
nand U48785 (N_48785,N_47621,N_46661);
nand U48786 (N_48786,N_46397,N_46815);
nor U48787 (N_48787,N_46537,N_47920);
xor U48788 (N_48788,N_46848,N_46228);
nand U48789 (N_48789,N_46954,N_47612);
or U48790 (N_48790,N_46121,N_47288);
or U48791 (N_48791,N_47861,N_47897);
nor U48792 (N_48792,N_46696,N_46646);
and U48793 (N_48793,N_46164,N_46721);
or U48794 (N_48794,N_46386,N_47816);
nor U48795 (N_48795,N_47158,N_47240);
nand U48796 (N_48796,N_47482,N_46213);
or U48797 (N_48797,N_46131,N_47075);
and U48798 (N_48798,N_46613,N_46541);
or U48799 (N_48799,N_46804,N_47769);
nand U48800 (N_48800,N_46910,N_47936);
nand U48801 (N_48801,N_47224,N_47982);
and U48802 (N_48802,N_46032,N_47501);
or U48803 (N_48803,N_47662,N_46798);
nand U48804 (N_48804,N_47253,N_46115);
nor U48805 (N_48805,N_47160,N_47127);
or U48806 (N_48806,N_46227,N_47432);
nand U48807 (N_48807,N_47461,N_46558);
and U48808 (N_48808,N_46513,N_46770);
and U48809 (N_48809,N_47958,N_46001);
xnor U48810 (N_48810,N_46109,N_47668);
xnor U48811 (N_48811,N_46647,N_47307);
nand U48812 (N_48812,N_46116,N_46364);
nand U48813 (N_48813,N_46093,N_46617);
nand U48814 (N_48814,N_47837,N_46375);
xnor U48815 (N_48815,N_47291,N_47871);
xor U48816 (N_48816,N_47151,N_47629);
nand U48817 (N_48817,N_46433,N_47136);
and U48818 (N_48818,N_47930,N_46551);
and U48819 (N_48819,N_47045,N_47664);
or U48820 (N_48820,N_46269,N_46399);
or U48821 (N_48821,N_47168,N_46105);
and U48822 (N_48822,N_47564,N_47034);
xnor U48823 (N_48823,N_46840,N_47720);
or U48824 (N_48824,N_47026,N_46072);
xor U48825 (N_48825,N_46468,N_47996);
and U48826 (N_48826,N_46787,N_47250);
nand U48827 (N_48827,N_47804,N_47953);
nand U48828 (N_48828,N_46436,N_47267);
and U48829 (N_48829,N_47148,N_46619);
nand U48830 (N_48830,N_47474,N_46251);
nor U48831 (N_48831,N_47721,N_46331);
nand U48832 (N_48832,N_47566,N_46906);
nor U48833 (N_48833,N_46782,N_47962);
and U48834 (N_48834,N_47744,N_47677);
nor U48835 (N_48835,N_47990,N_46589);
xor U48836 (N_48836,N_46438,N_47527);
or U48837 (N_48837,N_46760,N_47470);
xor U48838 (N_48838,N_47378,N_47423);
or U48839 (N_48839,N_47147,N_46179);
or U48840 (N_48840,N_47843,N_47425);
nor U48841 (N_48841,N_46575,N_47511);
xnor U48842 (N_48842,N_46020,N_46418);
nor U48843 (N_48843,N_46684,N_47660);
or U48844 (N_48844,N_47873,N_46709);
or U48845 (N_48845,N_47306,N_46083);
and U48846 (N_48846,N_46374,N_46935);
or U48847 (N_48847,N_47266,N_47581);
nor U48848 (N_48848,N_46606,N_47708);
xor U48849 (N_48849,N_46857,N_47014);
xor U48850 (N_48850,N_46023,N_47863);
or U48851 (N_48851,N_47709,N_46490);
nand U48852 (N_48852,N_46874,N_47001);
nor U48853 (N_48853,N_46204,N_47969);
or U48854 (N_48854,N_47705,N_46503);
xnor U48855 (N_48855,N_47967,N_46912);
xor U48856 (N_48856,N_47015,N_46605);
or U48857 (N_48857,N_46029,N_47931);
xor U48858 (N_48858,N_47965,N_47330);
nor U48859 (N_48859,N_47641,N_46499);
xnor U48860 (N_48860,N_47465,N_46189);
or U48861 (N_48861,N_47214,N_47459);
xor U48862 (N_48862,N_46774,N_46790);
nand U48863 (N_48863,N_47547,N_47563);
xor U48864 (N_48864,N_47340,N_46451);
and U48865 (N_48865,N_46609,N_46730);
xnor U48866 (N_48866,N_46701,N_46501);
and U48867 (N_48867,N_46778,N_46653);
xnor U48868 (N_48868,N_47851,N_46584);
nand U48869 (N_48869,N_47644,N_47876);
and U48870 (N_48870,N_47263,N_47405);
and U48871 (N_48871,N_47860,N_47156);
or U48872 (N_48872,N_46933,N_46756);
and U48873 (N_48873,N_46719,N_46694);
or U48874 (N_48874,N_47216,N_47821);
xor U48875 (N_48875,N_47311,N_47376);
xor U48876 (N_48876,N_47595,N_47888);
nor U48877 (N_48877,N_46075,N_47315);
nor U48878 (N_48878,N_47373,N_47839);
nand U48879 (N_48879,N_47685,N_47385);
or U48880 (N_48880,N_46287,N_46999);
nand U48881 (N_48881,N_47554,N_47044);
xnor U48882 (N_48882,N_47002,N_46570);
nand U48883 (N_48883,N_47318,N_47687);
nand U48884 (N_48884,N_46325,N_46186);
nand U48885 (N_48885,N_47602,N_47065);
nor U48886 (N_48886,N_46712,N_47326);
and U48887 (N_48887,N_46707,N_46867);
xnor U48888 (N_48888,N_46038,N_47271);
xor U48889 (N_48889,N_47933,N_47908);
xnor U48890 (N_48890,N_47865,N_47773);
or U48891 (N_48891,N_46539,N_46675);
or U48892 (N_48892,N_46327,N_46198);
or U48893 (N_48893,N_47587,N_47600);
nor U48894 (N_48894,N_46826,N_47269);
nor U48895 (N_48895,N_46911,N_47040);
nor U48896 (N_48896,N_47745,N_46423);
nand U48897 (N_48897,N_47473,N_46590);
nand U48898 (N_48898,N_46429,N_47803);
and U48899 (N_48899,N_46677,N_46837);
nand U48900 (N_48900,N_46901,N_46665);
nor U48901 (N_48901,N_46975,N_46891);
nor U48902 (N_48902,N_47341,N_46063);
nand U48903 (N_48903,N_47038,N_47576);
nor U48904 (N_48904,N_46784,N_47255);
and U48905 (N_48905,N_47161,N_46895);
or U48906 (N_48906,N_46199,N_46480);
and U48907 (N_48907,N_46704,N_47103);
nand U48908 (N_48908,N_47830,N_47449);
nand U48909 (N_48909,N_46078,N_47808);
xor U48910 (N_48910,N_46188,N_46833);
or U48911 (N_48911,N_46394,N_47611);
nor U48912 (N_48912,N_47909,N_47706);
nor U48913 (N_48913,N_47365,N_47740);
and U48914 (N_48914,N_47556,N_46305);
xnor U48915 (N_48915,N_46371,N_47106);
xor U48916 (N_48916,N_47119,N_47577);
and U48917 (N_48917,N_47355,N_47533);
nand U48918 (N_48918,N_47246,N_46812);
xnor U48919 (N_48919,N_46510,N_47814);
xor U48920 (N_48920,N_46432,N_47728);
nand U48921 (N_48921,N_46623,N_46862);
nor U48922 (N_48922,N_46863,N_46794);
or U48923 (N_48923,N_47208,N_47749);
xor U48924 (N_48924,N_46547,N_47726);
or U48925 (N_48925,N_46759,N_46356);
nor U48926 (N_48926,N_46690,N_46045);
xor U48927 (N_48927,N_46257,N_46336);
xnor U48928 (N_48928,N_47163,N_47858);
nor U48929 (N_48929,N_47806,N_46994);
nor U48930 (N_48930,N_46676,N_46279);
nand U48931 (N_48931,N_46577,N_47155);
and U48932 (N_48932,N_46791,N_47013);
nand U48933 (N_48933,N_47374,N_46634);
nand U48934 (N_48934,N_46361,N_46463);
or U48935 (N_48935,N_46019,N_46373);
xor U48936 (N_48936,N_46294,N_46214);
and U48937 (N_48937,N_46749,N_46205);
and U48938 (N_48938,N_46648,N_47181);
and U48939 (N_48939,N_47194,N_47719);
and U48940 (N_48940,N_47948,N_46535);
nor U48941 (N_48941,N_47910,N_46163);
nand U48942 (N_48942,N_47796,N_47857);
or U48943 (N_48943,N_46632,N_46491);
nor U48944 (N_48944,N_46699,N_47738);
nand U48945 (N_48945,N_47867,N_46504);
or U48946 (N_48946,N_47333,N_47921);
xnor U48947 (N_48947,N_46538,N_47215);
nand U48948 (N_48948,N_47353,N_46393);
or U48949 (N_48949,N_46037,N_47000);
and U48950 (N_48950,N_46220,N_46165);
nor U48951 (N_48951,N_46844,N_47781);
xnor U48952 (N_48952,N_46141,N_46142);
or U48953 (N_48953,N_46964,N_46474);
or U48954 (N_48954,N_46349,N_46209);
nor U48955 (N_48955,N_47763,N_47173);
xnor U48956 (N_48956,N_46080,N_47347);
nand U48957 (N_48957,N_46520,N_46620);
nand U48958 (N_48958,N_46097,N_47408);
nand U48959 (N_48959,N_47971,N_47672);
or U48960 (N_48960,N_46100,N_47831);
xor U48961 (N_48961,N_46306,N_47877);
nor U48962 (N_48962,N_47495,N_47643);
nor U48963 (N_48963,N_46928,N_47139);
nor U48964 (N_48964,N_46086,N_47016);
nand U48965 (N_48965,N_47316,N_47551);
or U48966 (N_48966,N_47239,N_46050);
nand U48967 (N_48967,N_47886,N_46576);
nor U48968 (N_48968,N_46275,N_47406);
or U48969 (N_48969,N_46729,N_47599);
and U48970 (N_48970,N_46639,N_46579);
xor U48971 (N_48971,N_47633,N_46084);
nand U48972 (N_48972,N_46096,N_47264);
or U48973 (N_48973,N_47778,N_46936);
xor U48974 (N_48974,N_46391,N_46136);
nand U48975 (N_48975,N_46603,N_47375);
and U48976 (N_48976,N_46193,N_46683);
xor U48977 (N_48977,N_47052,N_47665);
nor U48978 (N_48978,N_47810,N_46191);
xnor U48979 (N_48979,N_47108,N_46742);
or U48980 (N_48980,N_46448,N_47890);
nand U48981 (N_48981,N_47212,N_47941);
and U48982 (N_48982,N_47582,N_46094);
nor U48983 (N_48983,N_47505,N_46461);
nand U48984 (N_48984,N_47822,N_47490);
xor U48985 (N_48985,N_47835,N_46206);
nor U48986 (N_48986,N_46872,N_46334);
nand U48987 (N_48987,N_46991,N_46850);
nor U48988 (N_48988,N_46893,N_47177);
or U48989 (N_48989,N_47033,N_47862);
xor U48990 (N_48990,N_46483,N_47317);
nand U48991 (N_48991,N_46073,N_46362);
or U48992 (N_48992,N_47832,N_46428);
xor U48993 (N_48993,N_46380,N_46011);
or U48994 (N_48994,N_47515,N_46441);
or U48995 (N_48995,N_47203,N_46168);
nand U48996 (N_48996,N_46529,N_46067);
or U48997 (N_48997,N_46758,N_47531);
nor U48998 (N_48998,N_47731,N_47292);
and U48999 (N_48999,N_46728,N_46726);
and U49000 (N_49000,N_46458,N_46833);
nor U49001 (N_49001,N_46348,N_46391);
or U49002 (N_49002,N_47102,N_46500);
nand U49003 (N_49003,N_46311,N_47337);
nor U49004 (N_49004,N_46986,N_46675);
xnor U49005 (N_49005,N_46001,N_47180);
nand U49006 (N_49006,N_46120,N_46081);
nand U49007 (N_49007,N_46357,N_47782);
nand U49008 (N_49008,N_46541,N_46579);
nor U49009 (N_49009,N_46942,N_47106);
nor U49010 (N_49010,N_47717,N_46384);
and U49011 (N_49011,N_47435,N_46715);
nor U49012 (N_49012,N_47525,N_47762);
nand U49013 (N_49013,N_46382,N_46217);
and U49014 (N_49014,N_46979,N_47183);
or U49015 (N_49015,N_46300,N_47758);
nor U49016 (N_49016,N_47897,N_47938);
or U49017 (N_49017,N_47302,N_46108);
xnor U49018 (N_49018,N_47583,N_47429);
and U49019 (N_49019,N_47937,N_47170);
xnor U49020 (N_49020,N_46522,N_46684);
nand U49021 (N_49021,N_47794,N_47090);
nand U49022 (N_49022,N_47373,N_46414);
or U49023 (N_49023,N_47508,N_47290);
nor U49024 (N_49024,N_46458,N_47670);
and U49025 (N_49025,N_46462,N_47336);
or U49026 (N_49026,N_47827,N_46993);
nor U49027 (N_49027,N_47094,N_47893);
nand U49028 (N_49028,N_47780,N_46300);
or U49029 (N_49029,N_46332,N_47354);
and U49030 (N_49030,N_46826,N_46423);
and U49031 (N_49031,N_46405,N_46967);
nor U49032 (N_49032,N_47886,N_46914);
nor U49033 (N_49033,N_46089,N_46884);
nand U49034 (N_49034,N_47307,N_47885);
and U49035 (N_49035,N_46691,N_47906);
nor U49036 (N_49036,N_46543,N_47945);
or U49037 (N_49037,N_47646,N_47460);
and U49038 (N_49038,N_47335,N_46801);
or U49039 (N_49039,N_46397,N_47266);
or U49040 (N_49040,N_47350,N_46214);
and U49041 (N_49041,N_47043,N_47541);
xnor U49042 (N_49042,N_46483,N_47641);
nor U49043 (N_49043,N_47778,N_46227);
xnor U49044 (N_49044,N_47971,N_46911);
or U49045 (N_49045,N_46893,N_46827);
nor U49046 (N_49046,N_46168,N_47489);
nand U49047 (N_49047,N_47229,N_47359);
xnor U49048 (N_49048,N_47506,N_47761);
nand U49049 (N_49049,N_47240,N_46323);
xor U49050 (N_49050,N_46527,N_46235);
xnor U49051 (N_49051,N_47471,N_46993);
nand U49052 (N_49052,N_47354,N_47170);
or U49053 (N_49053,N_47121,N_47929);
and U49054 (N_49054,N_47725,N_46115);
or U49055 (N_49055,N_46078,N_47046);
nand U49056 (N_49056,N_46135,N_46189);
nand U49057 (N_49057,N_47047,N_46724);
and U49058 (N_49058,N_46064,N_47707);
xnor U49059 (N_49059,N_46797,N_46035);
xnor U49060 (N_49060,N_46111,N_47283);
or U49061 (N_49061,N_46170,N_47962);
xor U49062 (N_49062,N_46091,N_46934);
or U49063 (N_49063,N_46702,N_46295);
nand U49064 (N_49064,N_47495,N_47634);
or U49065 (N_49065,N_47978,N_46552);
nand U49066 (N_49066,N_46112,N_46365);
nand U49067 (N_49067,N_46247,N_47792);
or U49068 (N_49068,N_47804,N_47553);
and U49069 (N_49069,N_47919,N_46606);
xor U49070 (N_49070,N_46697,N_46666);
and U49071 (N_49071,N_47455,N_47240);
xor U49072 (N_49072,N_47781,N_47319);
nor U49073 (N_49073,N_47918,N_46505);
nor U49074 (N_49074,N_47510,N_46872);
nor U49075 (N_49075,N_46008,N_46402);
and U49076 (N_49076,N_47659,N_47541);
or U49077 (N_49077,N_47616,N_46970);
or U49078 (N_49078,N_46854,N_46323);
nand U49079 (N_49079,N_46815,N_47719);
nor U49080 (N_49080,N_46779,N_47792);
nor U49081 (N_49081,N_46965,N_46731);
nor U49082 (N_49082,N_46791,N_47205);
or U49083 (N_49083,N_46760,N_46539);
nor U49084 (N_49084,N_47945,N_47841);
or U49085 (N_49085,N_47109,N_46059);
nand U49086 (N_49086,N_47631,N_46674);
nand U49087 (N_49087,N_46990,N_46105);
xor U49088 (N_49088,N_46069,N_47802);
nor U49089 (N_49089,N_46167,N_47012);
nand U49090 (N_49090,N_47939,N_47967);
xnor U49091 (N_49091,N_47569,N_47858);
or U49092 (N_49092,N_47110,N_47895);
xnor U49093 (N_49093,N_47516,N_47181);
nor U49094 (N_49094,N_47811,N_46989);
and U49095 (N_49095,N_46965,N_47903);
xor U49096 (N_49096,N_46697,N_47149);
or U49097 (N_49097,N_47554,N_46641);
or U49098 (N_49098,N_46277,N_46247);
or U49099 (N_49099,N_46396,N_47463);
nor U49100 (N_49100,N_46804,N_47482);
nor U49101 (N_49101,N_46197,N_46969);
and U49102 (N_49102,N_46528,N_46069);
nand U49103 (N_49103,N_47584,N_47331);
nor U49104 (N_49104,N_46001,N_46782);
nor U49105 (N_49105,N_47197,N_46267);
nor U49106 (N_49106,N_46836,N_46292);
xnor U49107 (N_49107,N_47634,N_46063);
and U49108 (N_49108,N_47316,N_46665);
or U49109 (N_49109,N_46405,N_47226);
nor U49110 (N_49110,N_46066,N_46224);
xor U49111 (N_49111,N_47524,N_47777);
nor U49112 (N_49112,N_47504,N_47920);
or U49113 (N_49113,N_46384,N_47088);
and U49114 (N_49114,N_46351,N_46164);
nand U49115 (N_49115,N_47499,N_47378);
or U49116 (N_49116,N_46297,N_46781);
xor U49117 (N_49117,N_46205,N_46840);
and U49118 (N_49118,N_46110,N_46888);
and U49119 (N_49119,N_47276,N_47909);
xnor U49120 (N_49120,N_47232,N_47881);
and U49121 (N_49121,N_47585,N_47913);
and U49122 (N_49122,N_47787,N_47900);
nand U49123 (N_49123,N_46249,N_46316);
xor U49124 (N_49124,N_47281,N_46854);
nor U49125 (N_49125,N_46126,N_47060);
xor U49126 (N_49126,N_47056,N_46499);
or U49127 (N_49127,N_47929,N_47644);
and U49128 (N_49128,N_47276,N_47116);
nand U49129 (N_49129,N_46367,N_47316);
and U49130 (N_49130,N_46718,N_46754);
or U49131 (N_49131,N_46487,N_47631);
or U49132 (N_49132,N_46923,N_47370);
and U49133 (N_49133,N_46616,N_47659);
xnor U49134 (N_49134,N_46944,N_46458);
and U49135 (N_49135,N_47808,N_46790);
nor U49136 (N_49136,N_47479,N_46766);
and U49137 (N_49137,N_47840,N_46271);
or U49138 (N_49138,N_46363,N_46881);
or U49139 (N_49139,N_46256,N_46145);
nand U49140 (N_49140,N_47439,N_46777);
nor U49141 (N_49141,N_47272,N_47721);
nor U49142 (N_49142,N_46218,N_47450);
nand U49143 (N_49143,N_46304,N_47518);
nor U49144 (N_49144,N_47120,N_47835);
nor U49145 (N_49145,N_47828,N_47808);
xnor U49146 (N_49146,N_47379,N_47553);
nor U49147 (N_49147,N_47106,N_47497);
or U49148 (N_49148,N_47177,N_47213);
or U49149 (N_49149,N_47523,N_47245);
nand U49150 (N_49150,N_47187,N_47779);
nor U49151 (N_49151,N_46218,N_47763);
xor U49152 (N_49152,N_46080,N_47480);
nor U49153 (N_49153,N_47108,N_46149);
nand U49154 (N_49154,N_47699,N_47061);
xnor U49155 (N_49155,N_47924,N_47352);
or U49156 (N_49156,N_47112,N_47924);
or U49157 (N_49157,N_47894,N_46418);
and U49158 (N_49158,N_46963,N_47194);
or U49159 (N_49159,N_46547,N_47927);
nand U49160 (N_49160,N_46556,N_47179);
nor U49161 (N_49161,N_46665,N_47529);
and U49162 (N_49162,N_47941,N_46527);
nor U49163 (N_49163,N_47381,N_46285);
nor U49164 (N_49164,N_46161,N_46110);
nor U49165 (N_49165,N_46500,N_47824);
and U49166 (N_49166,N_47723,N_46439);
nand U49167 (N_49167,N_47112,N_46990);
or U49168 (N_49168,N_46255,N_46810);
nand U49169 (N_49169,N_46914,N_47202);
xnor U49170 (N_49170,N_46778,N_47667);
nor U49171 (N_49171,N_47849,N_46489);
nor U49172 (N_49172,N_46703,N_46856);
nor U49173 (N_49173,N_46815,N_46179);
xnor U49174 (N_49174,N_46677,N_47407);
and U49175 (N_49175,N_46891,N_46426);
nor U49176 (N_49176,N_47677,N_46385);
nor U49177 (N_49177,N_47059,N_47464);
xnor U49178 (N_49178,N_47940,N_46589);
nand U49179 (N_49179,N_47434,N_46784);
and U49180 (N_49180,N_46128,N_47108);
and U49181 (N_49181,N_47962,N_46460);
or U49182 (N_49182,N_47318,N_46518);
nand U49183 (N_49183,N_46119,N_46854);
or U49184 (N_49184,N_46907,N_47034);
nand U49185 (N_49185,N_46856,N_47477);
xor U49186 (N_49186,N_47571,N_47297);
and U49187 (N_49187,N_47202,N_47018);
xor U49188 (N_49188,N_46660,N_46118);
and U49189 (N_49189,N_47114,N_47678);
nor U49190 (N_49190,N_47957,N_47976);
and U49191 (N_49191,N_46723,N_47574);
nor U49192 (N_49192,N_46815,N_47832);
nand U49193 (N_49193,N_47858,N_47414);
nand U49194 (N_49194,N_46317,N_47134);
xnor U49195 (N_49195,N_47229,N_46988);
nor U49196 (N_49196,N_46054,N_46048);
and U49197 (N_49197,N_46077,N_47968);
and U49198 (N_49198,N_47239,N_47725);
nor U49199 (N_49199,N_47717,N_47158);
and U49200 (N_49200,N_46286,N_46595);
xnor U49201 (N_49201,N_46005,N_46535);
nand U49202 (N_49202,N_47799,N_46016);
and U49203 (N_49203,N_46199,N_46793);
xnor U49204 (N_49204,N_47843,N_47587);
xor U49205 (N_49205,N_46903,N_47792);
or U49206 (N_49206,N_47863,N_46210);
xnor U49207 (N_49207,N_47127,N_47191);
or U49208 (N_49208,N_46458,N_47345);
or U49209 (N_49209,N_47763,N_46511);
and U49210 (N_49210,N_47198,N_46336);
or U49211 (N_49211,N_47727,N_46182);
and U49212 (N_49212,N_46639,N_47213);
nand U49213 (N_49213,N_46664,N_47297);
and U49214 (N_49214,N_47049,N_46293);
or U49215 (N_49215,N_47782,N_47672);
nand U49216 (N_49216,N_46050,N_46974);
and U49217 (N_49217,N_46939,N_47310);
nand U49218 (N_49218,N_46913,N_47021);
nand U49219 (N_49219,N_47605,N_46148);
nand U49220 (N_49220,N_46635,N_46676);
xor U49221 (N_49221,N_46252,N_46668);
nand U49222 (N_49222,N_47997,N_46341);
nor U49223 (N_49223,N_46158,N_47022);
and U49224 (N_49224,N_46842,N_46665);
nand U49225 (N_49225,N_47915,N_46958);
nor U49226 (N_49226,N_47619,N_46405);
or U49227 (N_49227,N_46986,N_46947);
nor U49228 (N_49228,N_47067,N_46038);
xor U49229 (N_49229,N_47490,N_46281);
nand U49230 (N_49230,N_46572,N_46149);
or U49231 (N_49231,N_47717,N_46071);
or U49232 (N_49232,N_46714,N_46564);
nand U49233 (N_49233,N_47066,N_46021);
nor U49234 (N_49234,N_47016,N_47590);
and U49235 (N_49235,N_47340,N_47062);
xor U49236 (N_49236,N_47762,N_46724);
nand U49237 (N_49237,N_47519,N_47736);
and U49238 (N_49238,N_47035,N_46952);
xor U49239 (N_49239,N_46121,N_46860);
nor U49240 (N_49240,N_47350,N_46371);
xor U49241 (N_49241,N_46722,N_46147);
and U49242 (N_49242,N_46827,N_47212);
or U49243 (N_49243,N_47684,N_46748);
xnor U49244 (N_49244,N_47869,N_47203);
nor U49245 (N_49245,N_46673,N_47634);
nor U49246 (N_49246,N_47478,N_47420);
and U49247 (N_49247,N_47799,N_47005);
and U49248 (N_49248,N_46788,N_47867);
nor U49249 (N_49249,N_46169,N_46749);
and U49250 (N_49250,N_46913,N_46831);
xnor U49251 (N_49251,N_46967,N_46240);
nor U49252 (N_49252,N_47897,N_46739);
or U49253 (N_49253,N_46042,N_47206);
xor U49254 (N_49254,N_47763,N_46737);
and U49255 (N_49255,N_46022,N_46929);
nor U49256 (N_49256,N_47049,N_47371);
and U49257 (N_49257,N_47519,N_47211);
nand U49258 (N_49258,N_47619,N_46515);
or U49259 (N_49259,N_46807,N_47346);
or U49260 (N_49260,N_47011,N_46043);
nor U49261 (N_49261,N_47273,N_47332);
and U49262 (N_49262,N_47372,N_47228);
nand U49263 (N_49263,N_46443,N_47221);
or U49264 (N_49264,N_46848,N_47931);
nand U49265 (N_49265,N_47343,N_47327);
and U49266 (N_49266,N_46016,N_46188);
nand U49267 (N_49267,N_47385,N_47564);
or U49268 (N_49268,N_46581,N_47957);
xor U49269 (N_49269,N_46794,N_47947);
xor U49270 (N_49270,N_47703,N_46110);
xnor U49271 (N_49271,N_46867,N_47567);
or U49272 (N_49272,N_46140,N_46459);
nor U49273 (N_49273,N_47264,N_46346);
or U49274 (N_49274,N_46860,N_47940);
or U49275 (N_49275,N_47059,N_47862);
xor U49276 (N_49276,N_47294,N_47231);
and U49277 (N_49277,N_47306,N_47533);
nand U49278 (N_49278,N_47242,N_46206);
nand U49279 (N_49279,N_46906,N_46793);
and U49280 (N_49280,N_47452,N_47072);
nand U49281 (N_49281,N_46594,N_47705);
nor U49282 (N_49282,N_47249,N_46112);
and U49283 (N_49283,N_46158,N_47348);
and U49284 (N_49284,N_46729,N_47489);
and U49285 (N_49285,N_46842,N_47070);
or U49286 (N_49286,N_47431,N_47610);
nand U49287 (N_49287,N_46368,N_47281);
and U49288 (N_49288,N_47344,N_46916);
nor U49289 (N_49289,N_46540,N_46180);
and U49290 (N_49290,N_46574,N_46744);
nor U49291 (N_49291,N_47781,N_47302);
nor U49292 (N_49292,N_47096,N_46217);
nand U49293 (N_49293,N_46788,N_46483);
or U49294 (N_49294,N_47539,N_47935);
xor U49295 (N_49295,N_47949,N_46454);
nand U49296 (N_49296,N_47330,N_47961);
nor U49297 (N_49297,N_46979,N_46940);
nor U49298 (N_49298,N_46870,N_47517);
xor U49299 (N_49299,N_46604,N_47311);
or U49300 (N_49300,N_46523,N_46987);
xor U49301 (N_49301,N_46829,N_47011);
and U49302 (N_49302,N_47424,N_47796);
nor U49303 (N_49303,N_46570,N_47212);
nor U49304 (N_49304,N_46626,N_46360);
nor U49305 (N_49305,N_47469,N_46866);
or U49306 (N_49306,N_46964,N_47811);
or U49307 (N_49307,N_46863,N_47744);
or U49308 (N_49308,N_46731,N_46743);
nor U49309 (N_49309,N_46074,N_47089);
xor U49310 (N_49310,N_46634,N_47028);
nor U49311 (N_49311,N_47841,N_47551);
nor U49312 (N_49312,N_47390,N_47430);
or U49313 (N_49313,N_47350,N_46454);
nand U49314 (N_49314,N_46406,N_46215);
or U49315 (N_49315,N_46423,N_46769);
or U49316 (N_49316,N_46082,N_46939);
nor U49317 (N_49317,N_47218,N_46629);
xnor U49318 (N_49318,N_46748,N_46514);
xnor U49319 (N_49319,N_47947,N_46602);
nand U49320 (N_49320,N_47390,N_47050);
nor U49321 (N_49321,N_47890,N_46704);
and U49322 (N_49322,N_47825,N_46380);
or U49323 (N_49323,N_47738,N_46986);
or U49324 (N_49324,N_47885,N_46095);
or U49325 (N_49325,N_47225,N_47945);
and U49326 (N_49326,N_46895,N_47866);
nand U49327 (N_49327,N_47299,N_47830);
or U49328 (N_49328,N_46182,N_46213);
and U49329 (N_49329,N_46962,N_46664);
nor U49330 (N_49330,N_46786,N_47025);
xnor U49331 (N_49331,N_47262,N_47232);
or U49332 (N_49332,N_46444,N_47899);
or U49333 (N_49333,N_46736,N_46303);
or U49334 (N_49334,N_47482,N_47413);
or U49335 (N_49335,N_46594,N_46572);
nand U49336 (N_49336,N_47291,N_46977);
xnor U49337 (N_49337,N_47442,N_46487);
xor U49338 (N_49338,N_46628,N_46857);
and U49339 (N_49339,N_47900,N_46763);
or U49340 (N_49340,N_46993,N_47449);
nand U49341 (N_49341,N_46231,N_46864);
xnor U49342 (N_49342,N_46685,N_47507);
nor U49343 (N_49343,N_46742,N_47437);
nand U49344 (N_49344,N_47950,N_47014);
nor U49345 (N_49345,N_46477,N_47221);
xor U49346 (N_49346,N_47481,N_47596);
xnor U49347 (N_49347,N_47340,N_47613);
xor U49348 (N_49348,N_47255,N_46349);
nand U49349 (N_49349,N_47594,N_46071);
nor U49350 (N_49350,N_46231,N_47646);
nand U49351 (N_49351,N_46679,N_46231);
and U49352 (N_49352,N_47216,N_47282);
and U49353 (N_49353,N_47520,N_46776);
nand U49354 (N_49354,N_46371,N_46582);
and U49355 (N_49355,N_47486,N_46266);
xnor U49356 (N_49356,N_47800,N_46968);
and U49357 (N_49357,N_47965,N_47456);
nor U49358 (N_49358,N_46019,N_46508);
xnor U49359 (N_49359,N_47046,N_47771);
nand U49360 (N_49360,N_47110,N_47260);
nand U49361 (N_49361,N_47603,N_46735);
xor U49362 (N_49362,N_47520,N_47825);
and U49363 (N_49363,N_47088,N_47207);
and U49364 (N_49364,N_47388,N_47831);
nor U49365 (N_49365,N_47845,N_47645);
nor U49366 (N_49366,N_47322,N_46241);
nand U49367 (N_49367,N_47106,N_46358);
xor U49368 (N_49368,N_46963,N_46694);
xnor U49369 (N_49369,N_46831,N_46025);
nor U49370 (N_49370,N_47121,N_46541);
nor U49371 (N_49371,N_47312,N_47006);
or U49372 (N_49372,N_46503,N_47873);
and U49373 (N_49373,N_47724,N_46217);
or U49374 (N_49374,N_47147,N_46326);
nor U49375 (N_49375,N_47670,N_47509);
or U49376 (N_49376,N_47909,N_46631);
nor U49377 (N_49377,N_46642,N_46539);
xnor U49378 (N_49378,N_46403,N_46065);
nor U49379 (N_49379,N_46060,N_47033);
or U49380 (N_49380,N_47801,N_47142);
nand U49381 (N_49381,N_46990,N_46297);
and U49382 (N_49382,N_46972,N_46733);
and U49383 (N_49383,N_47325,N_47817);
or U49384 (N_49384,N_46546,N_47147);
or U49385 (N_49385,N_47850,N_46842);
nand U49386 (N_49386,N_46624,N_47046);
nor U49387 (N_49387,N_46911,N_47184);
and U49388 (N_49388,N_46399,N_46160);
nand U49389 (N_49389,N_46033,N_46841);
nor U49390 (N_49390,N_47582,N_47895);
xnor U49391 (N_49391,N_47293,N_47828);
nor U49392 (N_49392,N_47563,N_47449);
or U49393 (N_49393,N_46914,N_46795);
and U49394 (N_49394,N_46585,N_46835);
and U49395 (N_49395,N_46233,N_46968);
nand U49396 (N_49396,N_46240,N_46946);
nor U49397 (N_49397,N_47818,N_46933);
nor U49398 (N_49398,N_46014,N_46731);
and U49399 (N_49399,N_46745,N_47559);
xnor U49400 (N_49400,N_47590,N_47326);
nor U49401 (N_49401,N_47986,N_47422);
or U49402 (N_49402,N_46828,N_46531);
xnor U49403 (N_49403,N_46984,N_46028);
and U49404 (N_49404,N_47361,N_46092);
xnor U49405 (N_49405,N_46082,N_47647);
nand U49406 (N_49406,N_47489,N_46276);
xor U49407 (N_49407,N_47073,N_47567);
and U49408 (N_49408,N_47393,N_47730);
nor U49409 (N_49409,N_47462,N_46695);
nand U49410 (N_49410,N_47500,N_47092);
xor U49411 (N_49411,N_46527,N_46289);
and U49412 (N_49412,N_47020,N_47828);
xnor U49413 (N_49413,N_47250,N_47791);
and U49414 (N_49414,N_46040,N_47722);
and U49415 (N_49415,N_47240,N_46957);
xor U49416 (N_49416,N_46768,N_47996);
xnor U49417 (N_49417,N_47592,N_46619);
nand U49418 (N_49418,N_47447,N_46852);
nand U49419 (N_49419,N_47758,N_47248);
nor U49420 (N_49420,N_46679,N_46278);
and U49421 (N_49421,N_47997,N_46597);
nor U49422 (N_49422,N_47352,N_47737);
and U49423 (N_49423,N_46536,N_46056);
nor U49424 (N_49424,N_46555,N_47098);
nand U49425 (N_49425,N_46725,N_47265);
nand U49426 (N_49426,N_47970,N_47425);
and U49427 (N_49427,N_46065,N_47463);
or U49428 (N_49428,N_46264,N_46150);
nand U49429 (N_49429,N_46195,N_46775);
nor U49430 (N_49430,N_47172,N_46576);
xor U49431 (N_49431,N_47754,N_46295);
xnor U49432 (N_49432,N_47955,N_47615);
xor U49433 (N_49433,N_47851,N_47271);
or U49434 (N_49434,N_46124,N_47634);
or U49435 (N_49435,N_46253,N_46185);
nand U49436 (N_49436,N_46857,N_46094);
nand U49437 (N_49437,N_46538,N_47670);
and U49438 (N_49438,N_46060,N_47145);
or U49439 (N_49439,N_46890,N_47893);
nor U49440 (N_49440,N_47464,N_46051);
nor U49441 (N_49441,N_46373,N_47110);
or U49442 (N_49442,N_47372,N_46412);
nor U49443 (N_49443,N_47381,N_47689);
xor U49444 (N_49444,N_46061,N_47395);
or U49445 (N_49445,N_47870,N_46128);
nand U49446 (N_49446,N_46380,N_47967);
nand U49447 (N_49447,N_46193,N_46855);
nand U49448 (N_49448,N_46783,N_47836);
nand U49449 (N_49449,N_47774,N_47282);
nand U49450 (N_49450,N_46254,N_47330);
xor U49451 (N_49451,N_46107,N_47281);
and U49452 (N_49452,N_46083,N_47760);
xnor U49453 (N_49453,N_46005,N_47018);
and U49454 (N_49454,N_46958,N_47548);
and U49455 (N_49455,N_47524,N_47364);
xnor U49456 (N_49456,N_47603,N_46105);
or U49457 (N_49457,N_46873,N_46346);
and U49458 (N_49458,N_47643,N_46284);
nor U49459 (N_49459,N_46155,N_47698);
nor U49460 (N_49460,N_47821,N_46402);
nand U49461 (N_49461,N_47361,N_47449);
and U49462 (N_49462,N_47048,N_46300);
nor U49463 (N_49463,N_47140,N_47903);
or U49464 (N_49464,N_47500,N_47321);
nor U49465 (N_49465,N_47823,N_47259);
nand U49466 (N_49466,N_46189,N_47851);
nand U49467 (N_49467,N_47232,N_46993);
nor U49468 (N_49468,N_47266,N_47530);
xor U49469 (N_49469,N_47967,N_47303);
nor U49470 (N_49470,N_46488,N_47793);
and U49471 (N_49471,N_46413,N_47057);
and U49472 (N_49472,N_46348,N_46104);
xor U49473 (N_49473,N_47768,N_46718);
xnor U49474 (N_49474,N_47051,N_46709);
or U49475 (N_49475,N_46558,N_46552);
xor U49476 (N_49476,N_47159,N_47936);
and U49477 (N_49477,N_46358,N_47383);
and U49478 (N_49478,N_47849,N_47422);
and U49479 (N_49479,N_47873,N_46385);
and U49480 (N_49480,N_46436,N_46289);
or U49481 (N_49481,N_46481,N_47087);
or U49482 (N_49482,N_46314,N_47069);
and U49483 (N_49483,N_46714,N_47398);
nand U49484 (N_49484,N_47810,N_47858);
xnor U49485 (N_49485,N_46580,N_46004);
nor U49486 (N_49486,N_46139,N_47816);
or U49487 (N_49487,N_47350,N_46101);
xor U49488 (N_49488,N_46892,N_47110);
nor U49489 (N_49489,N_46243,N_47712);
nor U49490 (N_49490,N_46056,N_47634);
or U49491 (N_49491,N_46434,N_47608);
and U49492 (N_49492,N_47935,N_46020);
nor U49493 (N_49493,N_47133,N_47536);
nand U49494 (N_49494,N_46035,N_46735);
xor U49495 (N_49495,N_46358,N_47572);
and U49496 (N_49496,N_47602,N_47801);
and U49497 (N_49497,N_46989,N_47895);
xor U49498 (N_49498,N_46689,N_46579);
nor U49499 (N_49499,N_46260,N_47039);
and U49500 (N_49500,N_47634,N_46624);
or U49501 (N_49501,N_46877,N_46370);
or U49502 (N_49502,N_47546,N_46379);
nor U49503 (N_49503,N_46489,N_47002);
nand U49504 (N_49504,N_46458,N_46449);
or U49505 (N_49505,N_47437,N_46390);
nor U49506 (N_49506,N_46609,N_47517);
nor U49507 (N_49507,N_47719,N_46205);
and U49508 (N_49508,N_47231,N_47430);
xnor U49509 (N_49509,N_46701,N_47259);
nand U49510 (N_49510,N_47665,N_46399);
nand U49511 (N_49511,N_46182,N_46014);
nor U49512 (N_49512,N_47090,N_47311);
xor U49513 (N_49513,N_47742,N_47833);
and U49514 (N_49514,N_47486,N_46455);
or U49515 (N_49515,N_46693,N_46723);
xor U49516 (N_49516,N_47849,N_46404);
and U49517 (N_49517,N_47441,N_47199);
nor U49518 (N_49518,N_46549,N_46971);
and U49519 (N_49519,N_46582,N_47726);
and U49520 (N_49520,N_46065,N_46709);
or U49521 (N_49521,N_47904,N_47679);
xor U49522 (N_49522,N_47203,N_46632);
nand U49523 (N_49523,N_47026,N_46276);
or U49524 (N_49524,N_47569,N_47506);
and U49525 (N_49525,N_46793,N_46061);
nor U49526 (N_49526,N_47723,N_46966);
xnor U49527 (N_49527,N_47548,N_47721);
nand U49528 (N_49528,N_47103,N_47639);
and U49529 (N_49529,N_47711,N_47405);
and U49530 (N_49530,N_47777,N_47133);
or U49531 (N_49531,N_47180,N_47694);
nor U49532 (N_49532,N_46378,N_46970);
or U49533 (N_49533,N_47153,N_46239);
and U49534 (N_49534,N_47552,N_47830);
and U49535 (N_49535,N_46671,N_46345);
or U49536 (N_49536,N_46377,N_47496);
nor U49537 (N_49537,N_47205,N_46061);
nor U49538 (N_49538,N_46243,N_46809);
and U49539 (N_49539,N_46987,N_47760);
xnor U49540 (N_49540,N_46152,N_47319);
nor U49541 (N_49541,N_47915,N_47752);
or U49542 (N_49542,N_46026,N_46237);
or U49543 (N_49543,N_47874,N_47127);
or U49544 (N_49544,N_46294,N_47904);
nor U49545 (N_49545,N_47589,N_46223);
or U49546 (N_49546,N_47278,N_46815);
or U49547 (N_49547,N_46627,N_46763);
nand U49548 (N_49548,N_46822,N_47763);
nand U49549 (N_49549,N_46283,N_47261);
or U49550 (N_49550,N_46724,N_47568);
or U49551 (N_49551,N_47806,N_46359);
nand U49552 (N_49552,N_47746,N_46459);
nand U49553 (N_49553,N_47306,N_47251);
and U49554 (N_49554,N_46587,N_46263);
nand U49555 (N_49555,N_47895,N_46518);
or U49556 (N_49556,N_47738,N_47019);
and U49557 (N_49557,N_46730,N_46080);
nor U49558 (N_49558,N_47891,N_47240);
nor U49559 (N_49559,N_46027,N_46169);
or U49560 (N_49560,N_46940,N_46901);
nor U49561 (N_49561,N_46075,N_46386);
nand U49562 (N_49562,N_47694,N_46424);
or U49563 (N_49563,N_46060,N_46089);
or U49564 (N_49564,N_47741,N_47499);
and U49565 (N_49565,N_47825,N_47015);
nor U49566 (N_49566,N_47408,N_46559);
xnor U49567 (N_49567,N_47503,N_46414);
nand U49568 (N_49568,N_47525,N_47897);
or U49569 (N_49569,N_46699,N_47655);
nor U49570 (N_49570,N_46743,N_46149);
xnor U49571 (N_49571,N_47588,N_47277);
nand U49572 (N_49572,N_47285,N_46866);
and U49573 (N_49573,N_46531,N_46917);
or U49574 (N_49574,N_46722,N_47043);
or U49575 (N_49575,N_47092,N_46530);
xnor U49576 (N_49576,N_46721,N_47254);
xnor U49577 (N_49577,N_46936,N_46314);
nor U49578 (N_49578,N_47046,N_46076);
and U49579 (N_49579,N_47554,N_47155);
xnor U49580 (N_49580,N_47084,N_47282);
xnor U49581 (N_49581,N_46240,N_46979);
or U49582 (N_49582,N_46927,N_46982);
xor U49583 (N_49583,N_47297,N_47187);
xnor U49584 (N_49584,N_46604,N_47370);
xor U49585 (N_49585,N_47594,N_46568);
xor U49586 (N_49586,N_46331,N_47953);
xnor U49587 (N_49587,N_47502,N_46687);
nand U49588 (N_49588,N_47530,N_47295);
xor U49589 (N_49589,N_47606,N_46803);
nand U49590 (N_49590,N_46589,N_46750);
nor U49591 (N_49591,N_47603,N_47645);
and U49592 (N_49592,N_47399,N_47058);
and U49593 (N_49593,N_47203,N_47646);
nand U49594 (N_49594,N_46070,N_46483);
and U49595 (N_49595,N_47322,N_46781);
or U49596 (N_49596,N_47896,N_46054);
nor U49597 (N_49597,N_47499,N_46159);
nand U49598 (N_49598,N_47925,N_47061);
nand U49599 (N_49599,N_47488,N_46366);
nor U49600 (N_49600,N_47904,N_46040);
nor U49601 (N_49601,N_46414,N_46416);
xor U49602 (N_49602,N_47240,N_46574);
or U49603 (N_49603,N_46438,N_46516);
nor U49604 (N_49604,N_47449,N_46735);
xnor U49605 (N_49605,N_47139,N_46816);
nor U49606 (N_49606,N_46959,N_47277);
or U49607 (N_49607,N_46003,N_47761);
nor U49608 (N_49608,N_46162,N_47407);
xnor U49609 (N_49609,N_47597,N_47687);
xnor U49610 (N_49610,N_46685,N_47486);
and U49611 (N_49611,N_46136,N_47567);
nor U49612 (N_49612,N_46010,N_46766);
xnor U49613 (N_49613,N_47327,N_46392);
nor U49614 (N_49614,N_47230,N_47085);
nor U49615 (N_49615,N_46925,N_47620);
nor U49616 (N_49616,N_46979,N_47595);
or U49617 (N_49617,N_46402,N_46013);
nand U49618 (N_49618,N_47793,N_46130);
nand U49619 (N_49619,N_47254,N_46323);
and U49620 (N_49620,N_46855,N_47856);
xnor U49621 (N_49621,N_47225,N_46621);
nand U49622 (N_49622,N_46630,N_47655);
and U49623 (N_49623,N_46921,N_47298);
nor U49624 (N_49624,N_47730,N_47376);
xor U49625 (N_49625,N_47489,N_46404);
xnor U49626 (N_49626,N_46273,N_46298);
xnor U49627 (N_49627,N_47926,N_46384);
or U49628 (N_49628,N_46111,N_47370);
xor U49629 (N_49629,N_46705,N_46868);
or U49630 (N_49630,N_47826,N_46677);
nor U49631 (N_49631,N_47887,N_47888);
xnor U49632 (N_49632,N_46385,N_46721);
nor U49633 (N_49633,N_46327,N_47105);
xnor U49634 (N_49634,N_46271,N_46607);
or U49635 (N_49635,N_46221,N_46876);
or U49636 (N_49636,N_46797,N_46890);
and U49637 (N_49637,N_47671,N_47806);
nand U49638 (N_49638,N_47451,N_46833);
or U49639 (N_49639,N_47077,N_47080);
or U49640 (N_49640,N_46663,N_46780);
xnor U49641 (N_49641,N_47094,N_47240);
xor U49642 (N_49642,N_46679,N_46319);
nand U49643 (N_49643,N_47736,N_47657);
or U49644 (N_49644,N_47297,N_46102);
and U49645 (N_49645,N_47866,N_47404);
nand U49646 (N_49646,N_47345,N_46489);
nand U49647 (N_49647,N_46300,N_47729);
nand U49648 (N_49648,N_46853,N_47754);
nand U49649 (N_49649,N_46621,N_46576);
nor U49650 (N_49650,N_46925,N_47097);
nor U49651 (N_49651,N_46761,N_47237);
and U49652 (N_49652,N_47911,N_46267);
and U49653 (N_49653,N_46043,N_47716);
nor U49654 (N_49654,N_47728,N_47429);
xnor U49655 (N_49655,N_47840,N_46225);
nor U49656 (N_49656,N_46009,N_47265);
nand U49657 (N_49657,N_46004,N_47570);
xor U49658 (N_49658,N_46715,N_46177);
or U49659 (N_49659,N_46883,N_46099);
xnor U49660 (N_49660,N_47414,N_46984);
xnor U49661 (N_49661,N_46770,N_46692);
or U49662 (N_49662,N_46479,N_47301);
xnor U49663 (N_49663,N_46733,N_47237);
or U49664 (N_49664,N_46309,N_46152);
nor U49665 (N_49665,N_46577,N_46047);
xnor U49666 (N_49666,N_47101,N_47759);
nand U49667 (N_49667,N_46160,N_47067);
nor U49668 (N_49668,N_47891,N_47777);
nor U49669 (N_49669,N_47382,N_47146);
and U49670 (N_49670,N_46153,N_46410);
nand U49671 (N_49671,N_46870,N_46344);
nor U49672 (N_49672,N_46690,N_46856);
or U49673 (N_49673,N_46252,N_47181);
and U49674 (N_49674,N_46407,N_46425);
nor U49675 (N_49675,N_46252,N_47012);
xnor U49676 (N_49676,N_46465,N_46050);
or U49677 (N_49677,N_47019,N_46593);
or U49678 (N_49678,N_47053,N_46294);
or U49679 (N_49679,N_46699,N_47392);
nor U49680 (N_49680,N_46841,N_46745);
nand U49681 (N_49681,N_46584,N_46918);
nand U49682 (N_49682,N_47413,N_47724);
or U49683 (N_49683,N_46288,N_47006);
or U49684 (N_49684,N_46969,N_47098);
nor U49685 (N_49685,N_46247,N_47407);
and U49686 (N_49686,N_47444,N_46801);
nor U49687 (N_49687,N_47820,N_46563);
and U49688 (N_49688,N_46686,N_46961);
or U49689 (N_49689,N_47848,N_47787);
or U49690 (N_49690,N_46211,N_46680);
or U49691 (N_49691,N_47059,N_46797);
nand U49692 (N_49692,N_46090,N_47032);
and U49693 (N_49693,N_47832,N_46663);
and U49694 (N_49694,N_46227,N_46634);
nor U49695 (N_49695,N_47346,N_47690);
nor U49696 (N_49696,N_47957,N_46533);
nor U49697 (N_49697,N_46748,N_46700);
or U49698 (N_49698,N_47222,N_46024);
and U49699 (N_49699,N_46627,N_47274);
xor U49700 (N_49700,N_46098,N_47184);
xor U49701 (N_49701,N_47424,N_47586);
nor U49702 (N_49702,N_46692,N_47129);
nor U49703 (N_49703,N_47004,N_46009);
nor U49704 (N_49704,N_47905,N_47769);
and U49705 (N_49705,N_47014,N_46825);
nand U49706 (N_49706,N_47955,N_47870);
nand U49707 (N_49707,N_46230,N_47447);
xor U49708 (N_49708,N_47320,N_46397);
or U49709 (N_49709,N_46489,N_47366);
and U49710 (N_49710,N_46999,N_46923);
nand U49711 (N_49711,N_47692,N_47156);
nand U49712 (N_49712,N_46329,N_47143);
nor U49713 (N_49713,N_46550,N_47309);
nor U49714 (N_49714,N_46850,N_46264);
nor U49715 (N_49715,N_47016,N_46446);
and U49716 (N_49716,N_46055,N_47598);
or U49717 (N_49717,N_46735,N_47443);
nand U49718 (N_49718,N_47777,N_46382);
and U49719 (N_49719,N_47201,N_47177);
nand U49720 (N_49720,N_46657,N_46142);
nand U49721 (N_49721,N_46823,N_46500);
and U49722 (N_49722,N_47467,N_46866);
or U49723 (N_49723,N_46782,N_47747);
nand U49724 (N_49724,N_47232,N_46452);
xnor U49725 (N_49725,N_47690,N_47809);
nor U49726 (N_49726,N_46411,N_46988);
nor U49727 (N_49727,N_46416,N_47662);
and U49728 (N_49728,N_46305,N_47546);
nand U49729 (N_49729,N_46521,N_46831);
and U49730 (N_49730,N_46769,N_47947);
nor U49731 (N_49731,N_46671,N_47594);
and U49732 (N_49732,N_47319,N_47633);
xor U49733 (N_49733,N_47249,N_47466);
or U49734 (N_49734,N_47389,N_46598);
and U49735 (N_49735,N_46696,N_47966);
nand U49736 (N_49736,N_47744,N_47189);
and U49737 (N_49737,N_47305,N_46985);
nand U49738 (N_49738,N_47682,N_46537);
nor U49739 (N_49739,N_46490,N_46764);
or U49740 (N_49740,N_46940,N_47017);
and U49741 (N_49741,N_46991,N_46772);
and U49742 (N_49742,N_47615,N_46588);
nor U49743 (N_49743,N_46600,N_46481);
xnor U49744 (N_49744,N_47347,N_46115);
and U49745 (N_49745,N_47204,N_46569);
and U49746 (N_49746,N_47965,N_47274);
nand U49747 (N_49747,N_46593,N_47462);
and U49748 (N_49748,N_47529,N_47231);
or U49749 (N_49749,N_47827,N_47429);
nor U49750 (N_49750,N_47955,N_46515);
xor U49751 (N_49751,N_47161,N_46912);
nor U49752 (N_49752,N_46436,N_47039);
and U49753 (N_49753,N_47938,N_46295);
xnor U49754 (N_49754,N_46502,N_46485);
nor U49755 (N_49755,N_47317,N_46270);
and U49756 (N_49756,N_46401,N_46327);
nand U49757 (N_49757,N_46868,N_47082);
or U49758 (N_49758,N_46818,N_46796);
and U49759 (N_49759,N_46227,N_46623);
nor U49760 (N_49760,N_46821,N_47477);
and U49761 (N_49761,N_46926,N_46519);
or U49762 (N_49762,N_47439,N_47018);
nand U49763 (N_49763,N_46294,N_47980);
and U49764 (N_49764,N_46822,N_46091);
and U49765 (N_49765,N_47515,N_47333);
nand U49766 (N_49766,N_47422,N_46428);
nor U49767 (N_49767,N_47800,N_47207);
and U49768 (N_49768,N_47824,N_46153);
and U49769 (N_49769,N_47343,N_47456);
and U49770 (N_49770,N_46833,N_46302);
or U49771 (N_49771,N_47756,N_46474);
or U49772 (N_49772,N_46431,N_46787);
and U49773 (N_49773,N_47005,N_46048);
nand U49774 (N_49774,N_47915,N_47042);
and U49775 (N_49775,N_46219,N_46774);
and U49776 (N_49776,N_46477,N_46533);
or U49777 (N_49777,N_47572,N_46990);
nor U49778 (N_49778,N_47305,N_47156);
nor U49779 (N_49779,N_46369,N_47886);
xor U49780 (N_49780,N_46337,N_46112);
xor U49781 (N_49781,N_46221,N_46071);
and U49782 (N_49782,N_47795,N_46164);
xor U49783 (N_49783,N_46743,N_46046);
nor U49784 (N_49784,N_46189,N_46930);
and U49785 (N_49785,N_47010,N_47599);
and U49786 (N_49786,N_47847,N_46415);
and U49787 (N_49787,N_47170,N_47482);
nand U49788 (N_49788,N_47317,N_46185);
xnor U49789 (N_49789,N_47387,N_46373);
or U49790 (N_49790,N_46246,N_47943);
and U49791 (N_49791,N_47883,N_46154);
or U49792 (N_49792,N_46852,N_46120);
nor U49793 (N_49793,N_46762,N_47513);
xor U49794 (N_49794,N_47030,N_46748);
xnor U49795 (N_49795,N_46000,N_47076);
xnor U49796 (N_49796,N_46581,N_47303);
or U49797 (N_49797,N_46503,N_47058);
nor U49798 (N_49798,N_46176,N_46184);
or U49799 (N_49799,N_47758,N_46223);
xnor U49800 (N_49800,N_47783,N_47835);
xnor U49801 (N_49801,N_46052,N_46807);
xnor U49802 (N_49802,N_46517,N_46152);
xnor U49803 (N_49803,N_47863,N_46574);
xor U49804 (N_49804,N_46554,N_47022);
xor U49805 (N_49805,N_47397,N_46664);
xor U49806 (N_49806,N_46951,N_46283);
nand U49807 (N_49807,N_46604,N_46910);
and U49808 (N_49808,N_47764,N_46787);
xnor U49809 (N_49809,N_46535,N_47841);
nand U49810 (N_49810,N_46461,N_46830);
and U49811 (N_49811,N_46849,N_47111);
nand U49812 (N_49812,N_46785,N_47980);
nor U49813 (N_49813,N_46496,N_46692);
nor U49814 (N_49814,N_46264,N_47231);
and U49815 (N_49815,N_46663,N_47823);
nor U49816 (N_49816,N_46316,N_47469);
nor U49817 (N_49817,N_46239,N_47910);
or U49818 (N_49818,N_47510,N_46136);
xor U49819 (N_49819,N_47332,N_47454);
nor U49820 (N_49820,N_47260,N_46009);
nand U49821 (N_49821,N_47596,N_46374);
nor U49822 (N_49822,N_47803,N_47691);
nand U49823 (N_49823,N_47792,N_47924);
and U49824 (N_49824,N_47571,N_47695);
nor U49825 (N_49825,N_47190,N_46036);
nand U49826 (N_49826,N_46025,N_47323);
nand U49827 (N_49827,N_46298,N_47261);
nand U49828 (N_49828,N_46632,N_46934);
xnor U49829 (N_49829,N_47441,N_46962);
nand U49830 (N_49830,N_46060,N_47975);
or U49831 (N_49831,N_47960,N_46838);
xor U49832 (N_49832,N_47841,N_46907);
and U49833 (N_49833,N_47805,N_47281);
nand U49834 (N_49834,N_46103,N_46063);
or U49835 (N_49835,N_47210,N_47610);
xor U49836 (N_49836,N_46675,N_46326);
xnor U49837 (N_49837,N_46682,N_46630);
and U49838 (N_49838,N_47555,N_46106);
or U49839 (N_49839,N_46852,N_46518);
or U49840 (N_49840,N_47693,N_46269);
and U49841 (N_49841,N_47136,N_46972);
and U49842 (N_49842,N_46886,N_47314);
nor U49843 (N_49843,N_46984,N_46762);
or U49844 (N_49844,N_46570,N_47820);
xnor U49845 (N_49845,N_47649,N_47086);
nor U49846 (N_49846,N_46663,N_47966);
nand U49847 (N_49847,N_47002,N_46850);
and U49848 (N_49848,N_46124,N_47652);
xnor U49849 (N_49849,N_47441,N_47189);
nor U49850 (N_49850,N_46574,N_46734);
or U49851 (N_49851,N_47640,N_46023);
nand U49852 (N_49852,N_46241,N_46869);
nor U49853 (N_49853,N_46578,N_46242);
nand U49854 (N_49854,N_47850,N_46462);
and U49855 (N_49855,N_47784,N_47685);
and U49856 (N_49856,N_47562,N_47658);
xor U49857 (N_49857,N_47121,N_47646);
and U49858 (N_49858,N_47526,N_46676);
and U49859 (N_49859,N_47108,N_47760);
or U49860 (N_49860,N_46638,N_46380);
xor U49861 (N_49861,N_46851,N_46800);
and U49862 (N_49862,N_47610,N_46378);
nand U49863 (N_49863,N_46120,N_47976);
nor U49864 (N_49864,N_46954,N_47275);
nor U49865 (N_49865,N_47856,N_47810);
nand U49866 (N_49866,N_46281,N_46579);
nand U49867 (N_49867,N_46525,N_47460);
or U49868 (N_49868,N_47780,N_47451);
nor U49869 (N_49869,N_47063,N_46153);
or U49870 (N_49870,N_46615,N_47887);
nor U49871 (N_49871,N_46905,N_46256);
or U49872 (N_49872,N_47696,N_47918);
xor U49873 (N_49873,N_47673,N_47111);
and U49874 (N_49874,N_46589,N_46201);
or U49875 (N_49875,N_47204,N_47677);
nor U49876 (N_49876,N_46293,N_47719);
xnor U49877 (N_49877,N_46767,N_46556);
or U49878 (N_49878,N_47275,N_47709);
nor U49879 (N_49879,N_47104,N_47810);
xnor U49880 (N_49880,N_47352,N_46163);
xor U49881 (N_49881,N_47293,N_47377);
nor U49882 (N_49882,N_47469,N_46181);
nor U49883 (N_49883,N_46616,N_47389);
nand U49884 (N_49884,N_46921,N_46086);
or U49885 (N_49885,N_46337,N_46099);
xor U49886 (N_49886,N_47662,N_47114);
xnor U49887 (N_49887,N_46722,N_47311);
and U49888 (N_49888,N_46084,N_47724);
nand U49889 (N_49889,N_46991,N_46268);
nor U49890 (N_49890,N_47719,N_47751);
xor U49891 (N_49891,N_47368,N_47525);
nor U49892 (N_49892,N_46072,N_47663);
or U49893 (N_49893,N_47374,N_47331);
or U49894 (N_49894,N_46308,N_46610);
or U49895 (N_49895,N_47494,N_47663);
nand U49896 (N_49896,N_47497,N_47147);
xor U49897 (N_49897,N_47226,N_46938);
or U49898 (N_49898,N_47430,N_46300);
and U49899 (N_49899,N_46017,N_46668);
xor U49900 (N_49900,N_46228,N_47557);
nand U49901 (N_49901,N_46534,N_47933);
xnor U49902 (N_49902,N_47067,N_46288);
xor U49903 (N_49903,N_47789,N_46422);
and U49904 (N_49904,N_47632,N_46793);
and U49905 (N_49905,N_47214,N_47810);
or U49906 (N_49906,N_47795,N_46417);
nand U49907 (N_49907,N_46973,N_46990);
xnor U49908 (N_49908,N_46751,N_47792);
nor U49909 (N_49909,N_46438,N_46224);
and U49910 (N_49910,N_47344,N_46950);
xnor U49911 (N_49911,N_47346,N_47504);
and U49912 (N_49912,N_47240,N_46908);
and U49913 (N_49913,N_46622,N_47166);
nand U49914 (N_49914,N_47306,N_47949);
nand U49915 (N_49915,N_46483,N_47470);
xnor U49916 (N_49916,N_47940,N_47746);
nor U49917 (N_49917,N_47212,N_46733);
or U49918 (N_49918,N_46576,N_46966);
nor U49919 (N_49919,N_47765,N_47927);
and U49920 (N_49920,N_47840,N_47058);
nor U49921 (N_49921,N_47603,N_47435);
xnor U49922 (N_49922,N_46868,N_47392);
or U49923 (N_49923,N_47759,N_46495);
and U49924 (N_49924,N_47842,N_47430);
xnor U49925 (N_49925,N_46543,N_47499);
nor U49926 (N_49926,N_46757,N_47682);
or U49927 (N_49927,N_46343,N_46775);
nor U49928 (N_49928,N_46138,N_47500);
nand U49929 (N_49929,N_47305,N_46459);
xnor U49930 (N_49930,N_47618,N_46540);
or U49931 (N_49931,N_46813,N_47913);
xnor U49932 (N_49932,N_47287,N_47474);
xnor U49933 (N_49933,N_46284,N_47541);
or U49934 (N_49934,N_47895,N_47840);
xor U49935 (N_49935,N_47269,N_46687);
nor U49936 (N_49936,N_47556,N_46537);
xor U49937 (N_49937,N_47266,N_47302);
and U49938 (N_49938,N_47707,N_47876);
and U49939 (N_49939,N_46576,N_46173);
nor U49940 (N_49940,N_46290,N_46507);
nor U49941 (N_49941,N_46864,N_47677);
or U49942 (N_49942,N_46560,N_47595);
or U49943 (N_49943,N_47211,N_47077);
nor U49944 (N_49944,N_47491,N_47639);
nor U49945 (N_49945,N_47170,N_46054);
nand U49946 (N_49946,N_46383,N_47468);
and U49947 (N_49947,N_47874,N_47380);
nor U49948 (N_49948,N_47874,N_47991);
xor U49949 (N_49949,N_47535,N_47222);
xor U49950 (N_49950,N_46779,N_47876);
xor U49951 (N_49951,N_47353,N_46744);
or U49952 (N_49952,N_46473,N_47717);
nor U49953 (N_49953,N_47658,N_46078);
or U49954 (N_49954,N_46657,N_47740);
or U49955 (N_49955,N_46083,N_47340);
xor U49956 (N_49956,N_47486,N_46299);
or U49957 (N_49957,N_46199,N_46207);
nand U49958 (N_49958,N_46202,N_47425);
nor U49959 (N_49959,N_46399,N_46517);
and U49960 (N_49960,N_46828,N_46700);
nand U49961 (N_49961,N_46429,N_46810);
nand U49962 (N_49962,N_47076,N_46147);
or U49963 (N_49963,N_46816,N_46987);
xor U49964 (N_49964,N_46057,N_47309);
nand U49965 (N_49965,N_47468,N_46024);
nand U49966 (N_49966,N_47799,N_47760);
xnor U49967 (N_49967,N_46232,N_47913);
nor U49968 (N_49968,N_47430,N_47137);
nand U49969 (N_49969,N_46036,N_46795);
and U49970 (N_49970,N_47786,N_46643);
or U49971 (N_49971,N_46690,N_47446);
and U49972 (N_49972,N_46333,N_46261);
nand U49973 (N_49973,N_47266,N_47084);
nor U49974 (N_49974,N_46947,N_47155);
and U49975 (N_49975,N_47815,N_47657);
xor U49976 (N_49976,N_46470,N_47785);
nor U49977 (N_49977,N_46579,N_47322);
xor U49978 (N_49978,N_46245,N_47949);
xnor U49979 (N_49979,N_47568,N_46471);
or U49980 (N_49980,N_47822,N_47205);
and U49981 (N_49981,N_47832,N_46013);
and U49982 (N_49982,N_46316,N_47427);
xor U49983 (N_49983,N_47904,N_47381);
or U49984 (N_49984,N_46854,N_46530);
nand U49985 (N_49985,N_46385,N_46236);
nand U49986 (N_49986,N_47374,N_46267);
nand U49987 (N_49987,N_46809,N_46972);
nor U49988 (N_49988,N_47901,N_46288);
and U49989 (N_49989,N_46890,N_46606);
and U49990 (N_49990,N_47339,N_46461);
xnor U49991 (N_49991,N_47998,N_47828);
nand U49992 (N_49992,N_46920,N_47139);
or U49993 (N_49993,N_47878,N_47870);
nand U49994 (N_49994,N_47889,N_46396);
or U49995 (N_49995,N_47160,N_46802);
nand U49996 (N_49996,N_47115,N_46667);
nor U49997 (N_49997,N_47532,N_46780);
nand U49998 (N_49998,N_46947,N_46542);
nand U49999 (N_49999,N_47120,N_47728);
and UO_0 (O_0,N_49114,N_49408);
and UO_1 (O_1,N_48612,N_48619);
or UO_2 (O_2,N_48815,N_48172);
nor UO_3 (O_3,N_48715,N_49106);
nand UO_4 (O_4,N_49868,N_48035);
nand UO_5 (O_5,N_49774,N_48994);
or UO_6 (O_6,N_49025,N_48290);
nand UO_7 (O_7,N_48644,N_48728);
and UO_8 (O_8,N_48890,N_49222);
or UO_9 (O_9,N_48697,N_48127);
and UO_10 (O_10,N_48719,N_48207);
nor UO_11 (O_11,N_49759,N_49919);
nand UO_12 (O_12,N_48914,N_48529);
or UO_13 (O_13,N_49179,N_49290);
and UO_14 (O_14,N_49543,N_49460);
nand UO_15 (O_15,N_49150,N_48282);
xnor UO_16 (O_16,N_48390,N_49932);
xnor UO_17 (O_17,N_48523,N_49535);
nor UO_18 (O_18,N_49062,N_48811);
nand UO_19 (O_19,N_48018,N_49484);
nor UO_20 (O_20,N_48797,N_49021);
nor UO_21 (O_21,N_48701,N_49322);
nor UO_22 (O_22,N_49555,N_48064);
xnor UO_23 (O_23,N_49233,N_49928);
nor UO_24 (O_24,N_49826,N_48957);
nor UO_25 (O_25,N_48541,N_48025);
nand UO_26 (O_26,N_49684,N_49040);
xor UO_27 (O_27,N_49955,N_49782);
xor UO_28 (O_28,N_48253,N_48120);
or UO_29 (O_29,N_49553,N_48497);
or UO_30 (O_30,N_48907,N_49175);
and UO_31 (O_31,N_48543,N_49466);
nand UO_32 (O_32,N_48109,N_48921);
nor UO_33 (O_33,N_48001,N_48533);
nor UO_34 (O_34,N_48349,N_49344);
nor UO_35 (O_35,N_49001,N_49378);
xor UO_36 (O_36,N_48175,N_48696);
xnor UO_37 (O_37,N_49951,N_48802);
or UO_38 (O_38,N_48501,N_48704);
nand UO_39 (O_39,N_48481,N_49956);
nor UO_40 (O_40,N_48969,N_48502);
or UO_41 (O_41,N_49144,N_49482);
and UO_42 (O_42,N_49686,N_48558);
or UO_43 (O_43,N_49756,N_48103);
nor UO_44 (O_44,N_49780,N_49889);
and UO_45 (O_45,N_49295,N_49767);
xnor UO_46 (O_46,N_49895,N_49638);
nor UO_47 (O_47,N_48688,N_48990);
or UO_48 (O_48,N_49178,N_49528);
and UO_49 (O_49,N_49827,N_49435);
and UO_50 (O_50,N_48414,N_49655);
or UO_51 (O_51,N_49550,N_49986);
nand UO_52 (O_52,N_49271,N_49239);
or UO_53 (O_53,N_48430,N_49861);
and UO_54 (O_54,N_49781,N_49352);
nor UO_55 (O_55,N_48032,N_49132);
xor UO_56 (O_56,N_49042,N_49002);
nor UO_57 (O_57,N_49672,N_48877);
nor UO_58 (O_58,N_48788,N_49419);
or UO_59 (O_59,N_49749,N_48183);
or UO_60 (O_60,N_48074,N_49665);
xor UO_61 (O_61,N_49515,N_49738);
and UO_62 (O_62,N_49149,N_49676);
nand UO_63 (O_63,N_48029,N_48416);
nor UO_64 (O_64,N_49246,N_49970);
or UO_65 (O_65,N_48265,N_48861);
or UO_66 (O_66,N_49280,N_49966);
and UO_67 (O_67,N_49923,N_49424);
nor UO_68 (O_68,N_48427,N_48708);
nand UO_69 (O_69,N_49799,N_48762);
xor UO_70 (O_70,N_48066,N_48984);
and UO_71 (O_71,N_49348,N_49567);
nand UO_72 (O_72,N_49566,N_48795);
and UO_73 (O_73,N_49965,N_48749);
or UO_74 (O_74,N_49719,N_48357);
and UO_75 (O_75,N_49772,N_48174);
xnor UO_76 (O_76,N_49403,N_48751);
or UO_77 (O_77,N_48522,N_48130);
nor UO_78 (O_78,N_49586,N_49085);
and UO_79 (O_79,N_49382,N_48593);
or UO_80 (O_80,N_48709,N_48671);
xnor UO_81 (O_81,N_49793,N_49924);
and UO_82 (O_82,N_49192,N_48091);
and UO_83 (O_83,N_49317,N_49547);
nor UO_84 (O_84,N_48810,N_49946);
xnor UO_85 (O_85,N_49584,N_48974);
nor UO_86 (O_86,N_48736,N_48968);
and UO_87 (O_87,N_48916,N_49691);
nand UO_88 (O_88,N_49366,N_48735);
or UO_89 (O_89,N_48942,N_49575);
and UO_90 (O_90,N_48006,N_48148);
or UO_91 (O_91,N_48666,N_48185);
and UO_92 (O_92,N_48125,N_48903);
or UO_93 (O_93,N_48426,N_49620);
nor UO_94 (O_94,N_48937,N_49959);
or UO_95 (O_95,N_49259,N_49390);
xnor UO_96 (O_96,N_48020,N_49639);
nand UO_97 (O_97,N_48888,N_48417);
and UO_98 (O_98,N_48197,N_48402);
xor UO_99 (O_99,N_48138,N_49707);
xnor UO_100 (O_100,N_49155,N_49860);
nor UO_101 (O_101,N_48613,N_48821);
and UO_102 (O_102,N_48875,N_48892);
xnor UO_103 (O_103,N_49830,N_49650);
nand UO_104 (O_104,N_49355,N_48482);
nand UO_105 (O_105,N_48269,N_48364);
or UO_106 (O_106,N_48019,N_49434);
nand UO_107 (O_107,N_48104,N_49729);
and UO_108 (O_108,N_49448,N_48013);
nor UO_109 (O_109,N_49506,N_49766);
nor UO_110 (O_110,N_48727,N_49548);
nand UO_111 (O_111,N_48947,N_48242);
and UO_112 (O_112,N_48980,N_48331);
nand UO_113 (O_113,N_49777,N_48279);
and UO_114 (O_114,N_49326,N_49358);
nand UO_115 (O_115,N_49972,N_49992);
or UO_116 (O_116,N_49661,N_48859);
or UO_117 (O_117,N_48303,N_48310);
or UO_118 (O_118,N_48599,N_49055);
nand UO_119 (O_119,N_48446,N_48561);
nand UO_120 (O_120,N_48324,N_49765);
nor UO_121 (O_121,N_49395,N_49373);
xor UO_122 (O_122,N_49779,N_49472);
and UO_123 (O_123,N_49188,N_49845);
xnor UO_124 (O_124,N_49809,N_48158);
nand UO_125 (O_125,N_49292,N_48531);
nor UO_126 (O_126,N_48461,N_48358);
xnor UO_127 (O_127,N_48484,N_49513);
nand UO_128 (O_128,N_49823,N_49595);
nor UO_129 (O_129,N_49388,N_49978);
or UO_130 (O_130,N_49272,N_48503);
or UO_131 (O_131,N_49576,N_48166);
nand UO_132 (O_132,N_48397,N_49337);
and UO_133 (O_133,N_49113,N_49585);
and UO_134 (O_134,N_49309,N_49467);
xor UO_135 (O_135,N_49255,N_48607);
or UO_136 (O_136,N_48705,N_48255);
nor UO_137 (O_137,N_49427,N_48630);
nand UO_138 (O_138,N_48500,N_49364);
xnor UO_139 (O_139,N_49379,N_48759);
xnor UO_140 (O_140,N_48748,N_49370);
xnor UO_141 (O_141,N_49079,N_49629);
and UO_142 (O_142,N_49439,N_49999);
or UO_143 (O_143,N_49457,N_49048);
nor UO_144 (O_144,N_49289,N_48377);
nand UO_145 (O_145,N_48210,N_49169);
nand UO_146 (O_146,N_49306,N_48520);
nand UO_147 (O_147,N_49402,N_49432);
or UO_148 (O_148,N_49561,N_49721);
xor UO_149 (O_149,N_49268,N_48793);
nor UO_150 (O_150,N_48784,N_49252);
nand UO_151 (O_151,N_48573,N_49194);
or UO_152 (O_152,N_49695,N_49708);
and UO_153 (O_153,N_49105,N_48830);
xor UO_154 (O_154,N_49596,N_49213);
nor UO_155 (O_155,N_49139,N_49703);
or UO_156 (O_156,N_49209,N_49750);
xnor UO_157 (O_157,N_48149,N_48118);
or UO_158 (O_158,N_49670,N_48171);
or UO_159 (O_159,N_49886,N_48654);
xnor UO_160 (O_160,N_48044,N_49478);
or UO_161 (O_161,N_48211,N_49559);
xnor UO_162 (O_162,N_48322,N_48660);
nor UO_163 (O_163,N_49897,N_49357);
nand UO_164 (O_164,N_48798,N_48702);
or UO_165 (O_165,N_49033,N_49597);
nand UO_166 (O_166,N_49912,N_49265);
nor UO_167 (O_167,N_49529,N_49303);
xnor UO_168 (O_168,N_49362,N_48931);
and UO_169 (O_169,N_48581,N_49302);
nand UO_170 (O_170,N_48356,N_49137);
and UO_171 (O_171,N_48090,N_49170);
nand UO_172 (O_172,N_49853,N_48447);
nor UO_173 (O_173,N_49146,N_48297);
xnor UO_174 (O_174,N_48274,N_49318);
xor UO_175 (O_175,N_48509,N_48477);
nor UO_176 (O_176,N_49680,N_48897);
and UO_177 (O_177,N_48733,N_49718);
and UO_178 (O_178,N_49801,N_48721);
nand UO_179 (O_179,N_49275,N_49702);
or UO_180 (O_180,N_49167,N_48929);
xnor UO_181 (O_181,N_49952,N_49143);
or UO_182 (O_182,N_49104,N_49570);
and UO_183 (O_183,N_48124,N_49125);
and UO_184 (O_184,N_48889,N_48764);
nand UO_185 (O_185,N_49443,N_49894);
or UO_186 (O_186,N_48480,N_49723);
or UO_187 (O_187,N_48079,N_48156);
nor UO_188 (O_188,N_49200,N_48161);
nor UO_189 (O_189,N_48268,N_48476);
xor UO_190 (O_190,N_48726,N_48567);
nor UO_191 (O_191,N_48063,N_48003);
and UO_192 (O_192,N_48273,N_49308);
nor UO_193 (O_193,N_48292,N_48456);
xor UO_194 (O_194,N_49995,N_48223);
and UO_195 (O_195,N_48308,N_49926);
xor UO_196 (O_196,N_49740,N_49900);
nor UO_197 (O_197,N_49623,N_49741);
and UO_198 (O_198,N_48505,N_48270);
or UO_199 (O_199,N_48881,N_49936);
xnor UO_200 (O_200,N_49345,N_49849);
nand UO_201 (O_201,N_48515,N_48344);
nor UO_202 (O_202,N_49206,N_49768);
nand UO_203 (O_203,N_49636,N_48668);
nand UO_204 (O_204,N_49097,N_49736);
nand UO_205 (O_205,N_48234,N_49735);
or UO_206 (O_206,N_48371,N_49260);
or UO_207 (O_207,N_48252,N_49128);
and UO_208 (O_208,N_48062,N_48394);
nand UO_209 (O_209,N_48664,N_48944);
nor UO_210 (O_210,N_48251,N_49591);
or UO_211 (O_211,N_49525,N_48530);
or UO_212 (O_212,N_48198,N_48452);
nand UO_213 (O_213,N_48878,N_48342);
or UO_214 (O_214,N_48047,N_48649);
xnor UO_215 (O_215,N_48934,N_48030);
nand UO_216 (O_216,N_49982,N_49825);
and UO_217 (O_217,N_48844,N_49404);
xnor UO_218 (O_218,N_49800,N_48400);
or UO_219 (O_219,N_49334,N_49834);
or UO_220 (O_220,N_49593,N_49744);
or UO_221 (O_221,N_48572,N_49993);
nor UO_222 (O_222,N_48408,N_48985);
nand UO_223 (O_223,N_48512,N_48084);
nor UO_224 (O_224,N_49305,N_48439);
and UO_225 (O_225,N_49314,N_49022);
or UO_226 (O_226,N_49376,N_49180);
or UO_227 (O_227,N_48862,N_49142);
xnor UO_228 (O_228,N_49354,N_48004);
nor UO_229 (O_229,N_49375,N_48898);
nand UO_230 (O_230,N_49577,N_48488);
or UO_231 (O_231,N_48469,N_49123);
xnor UO_232 (O_232,N_48335,N_49546);
and UO_233 (O_233,N_49507,N_48239);
or UO_234 (O_234,N_49006,N_49681);
and UO_235 (O_235,N_48110,N_48640);
nor UO_236 (O_236,N_49815,N_49207);
nor UO_237 (O_237,N_48662,N_49835);
nor UO_238 (O_238,N_48583,N_49653);
nand UO_239 (O_239,N_48359,N_48899);
nand UO_240 (O_240,N_48328,N_48620);
and UO_241 (O_241,N_48987,N_48221);
and UO_242 (O_242,N_49425,N_48673);
or UO_243 (O_243,N_48046,N_49925);
and UO_244 (O_244,N_49803,N_48904);
nor UO_245 (O_245,N_49950,N_49274);
nand UO_246 (O_246,N_48874,N_48803);
xor UO_247 (O_247,N_48615,N_48562);
xnor UO_248 (O_248,N_48055,N_48475);
xnor UO_249 (O_249,N_49581,N_49539);
or UO_250 (O_250,N_49784,N_48822);
nand UO_251 (O_251,N_48490,N_49698);
or UO_252 (O_252,N_49863,N_48078);
or UO_253 (O_253,N_48757,N_49399);
nor UO_254 (O_254,N_48636,N_49247);
nand UO_255 (O_255,N_48299,N_48319);
and UO_256 (O_256,N_49152,N_49266);
nor UO_257 (O_257,N_48566,N_49509);
or UO_258 (O_258,N_48168,N_48794);
or UO_259 (O_259,N_48824,N_48352);
or UO_260 (O_260,N_48232,N_49606);
and UO_261 (O_261,N_48679,N_49485);
nor UO_262 (O_262,N_49941,N_48329);
nor UO_263 (O_263,N_49182,N_48981);
nor UO_264 (O_264,N_48832,N_48425);
xor UO_265 (O_265,N_49565,N_49617);
or UO_266 (O_266,N_49521,N_49039);
nor UO_267 (O_267,N_49804,N_49571);
nand UO_268 (O_268,N_48286,N_49116);
and UO_269 (O_269,N_49898,N_48173);
nand UO_270 (O_270,N_48423,N_48909);
and UO_271 (O_271,N_49607,N_49762);
nand UO_272 (O_272,N_49444,N_49420);
nor UO_273 (O_273,N_48542,N_49287);
xnor UO_274 (O_274,N_48924,N_48521);
nand UO_275 (O_275,N_49563,N_48302);
or UO_276 (O_276,N_49628,N_49270);
nor UO_277 (O_277,N_48946,N_49938);
or UO_278 (O_278,N_49298,N_49331);
and UO_279 (O_279,N_49277,N_48864);
xnor UO_280 (O_280,N_49041,N_48202);
xor UO_281 (O_281,N_49341,N_48350);
nor UO_282 (O_282,N_48938,N_48433);
and UO_283 (O_283,N_48466,N_48353);
and UO_284 (O_284,N_48315,N_49284);
and UO_285 (O_285,N_49300,N_49961);
xnor UO_286 (O_286,N_48238,N_49028);
xnor UO_287 (O_287,N_48372,N_48415);
nand UO_288 (O_288,N_49962,N_49612);
nor UO_289 (O_289,N_48094,N_49102);
xor UO_290 (O_290,N_49872,N_48912);
nand UO_291 (O_291,N_48053,N_48841);
or UO_292 (O_292,N_49544,N_49909);
nand UO_293 (O_293,N_49820,N_49010);
xnor UO_294 (O_294,N_49592,N_48655);
and UO_295 (O_295,N_48203,N_48925);
nor UO_296 (O_296,N_49631,N_49742);
xnor UO_297 (O_297,N_49621,N_48687);
xor UO_298 (O_298,N_49229,N_49294);
or UO_299 (O_299,N_49086,N_48146);
or UO_300 (O_300,N_48072,N_49456);
xnor UO_301 (O_301,N_48266,N_49056);
and UO_302 (O_302,N_48754,N_49118);
nand UO_303 (O_303,N_48123,N_49013);
nor UO_304 (O_304,N_49664,N_48317);
xnor UO_305 (O_305,N_49881,N_49043);
and UO_306 (O_306,N_48605,N_49080);
nor UO_307 (O_307,N_48760,N_48559);
nand UO_308 (O_308,N_48193,N_48939);
nand UO_309 (O_309,N_48287,N_48164);
or UO_310 (O_310,N_48182,N_49453);
or UO_311 (O_311,N_49573,N_49396);
xnor UO_312 (O_312,N_48177,N_48386);
nor UO_313 (O_313,N_48196,N_48073);
or UO_314 (O_314,N_49542,N_49844);
xor UO_315 (O_315,N_48410,N_48839);
xor UO_316 (O_316,N_48403,N_48819);
nor UO_317 (O_317,N_49365,N_48406);
or UO_318 (O_318,N_48187,N_48382);
or UO_319 (O_319,N_49258,N_48431);
or UO_320 (O_320,N_49051,N_48000);
nand UO_321 (O_321,N_49988,N_49496);
nand UO_322 (O_322,N_48464,N_48846);
or UO_323 (O_323,N_49637,N_49915);
nand UO_324 (O_324,N_49154,N_49973);
and UO_325 (O_325,N_48143,N_49921);
xor UO_326 (O_326,N_48113,N_48453);
nand UO_327 (O_327,N_48855,N_48271);
and UO_328 (O_328,N_49746,N_48419);
nand UO_329 (O_329,N_48879,N_48711);
or UO_330 (O_330,N_49293,N_49700);
or UO_331 (O_331,N_49032,N_48033);
nor UO_332 (O_332,N_48420,N_49866);
xor UO_333 (O_333,N_48387,N_49004);
xor UO_334 (O_334,N_48858,N_48871);
and UO_335 (O_335,N_48970,N_49805);
or UO_336 (O_336,N_49890,N_48144);
or UO_337 (O_337,N_48102,N_48448);
nor UO_338 (O_338,N_49441,N_49216);
nor UO_339 (O_339,N_48507,N_48478);
nand UO_340 (O_340,N_49816,N_49089);
nand UO_341 (O_341,N_48463,N_48691);
nor UO_342 (O_342,N_48421,N_48071);
nor UO_343 (O_343,N_49286,N_48989);
xnor UO_344 (O_344,N_48021,N_48126);
or UO_345 (O_345,N_49416,N_48191);
xnor UO_346 (O_346,N_49888,N_49244);
or UO_347 (O_347,N_49046,N_49832);
and UO_348 (O_348,N_48472,N_48807);
or UO_349 (O_349,N_48634,N_49262);
and UO_350 (O_350,N_48495,N_49556);
nor UO_351 (O_351,N_49451,N_48093);
nor UO_352 (O_352,N_49217,N_48134);
nand UO_353 (O_353,N_48782,N_49405);
nand UO_354 (O_354,N_49121,N_48557);
nand UO_355 (O_355,N_48157,N_49241);
xnor UO_356 (O_356,N_49953,N_49459);
and UO_357 (O_357,N_49090,N_49944);
or UO_358 (O_358,N_48893,N_48996);
and UO_359 (O_359,N_49989,N_48219);
nor UO_360 (O_360,N_49622,N_48971);
nor UO_361 (O_361,N_48860,N_48216);
xnor UO_362 (O_362,N_48460,N_48958);
nand UO_363 (O_363,N_49099,N_48825);
or UO_364 (O_364,N_49437,N_48948);
and UO_365 (O_365,N_49191,N_48418);
and UO_366 (O_366,N_48789,N_49401);
and UO_367 (O_367,N_49417,N_49706);
and UO_368 (O_368,N_48444,N_49273);
xnor UO_369 (O_369,N_48313,N_48590);
nor UO_370 (O_370,N_49795,N_49634);
nor UO_371 (O_371,N_48532,N_48524);
nor UO_372 (O_372,N_48908,N_48220);
nor UO_373 (O_373,N_49733,N_48876);
or UO_374 (O_374,N_48236,N_48829);
or UO_375 (O_375,N_49157,N_49481);
nor UO_376 (O_376,N_48584,N_48121);
and UO_377 (O_377,N_49162,N_48443);
xnor UO_378 (O_378,N_49745,N_48621);
and UO_379 (O_379,N_49603,N_48539);
nor UO_380 (O_380,N_48873,N_48028);
nor UO_381 (O_381,N_48441,N_49892);
nand UO_382 (O_382,N_48128,N_49283);
nand UO_383 (O_383,N_48677,N_48301);
or UO_384 (O_384,N_48544,N_48375);
xnor UO_385 (O_385,N_48368,N_48678);
nor UO_386 (O_386,N_48289,N_49533);
and UO_387 (O_387,N_48224,N_48896);
and UO_388 (O_388,N_48913,N_49050);
xor UO_389 (O_389,N_48201,N_48905);
xnor UO_390 (O_390,N_49498,N_49383);
xor UO_391 (O_391,N_48645,N_49474);
xnor UO_392 (O_392,N_49541,N_48396);
or UO_393 (O_393,N_49771,N_49224);
nand UO_394 (O_394,N_49257,N_48627);
and UO_395 (O_395,N_49884,N_49579);
nand UO_396 (O_396,N_48643,N_48842);
xnor UO_397 (O_397,N_49748,N_49231);
or UO_398 (O_398,N_49465,N_49429);
nor UO_399 (O_399,N_49393,N_48546);
xnor UO_400 (O_400,N_48720,N_49847);
xor UO_401 (O_401,N_49426,N_49193);
and UO_402 (O_402,N_49014,N_49658);
xnor UO_403 (O_403,N_49878,N_49153);
nor UO_404 (O_404,N_49361,N_49490);
or UO_405 (O_405,N_49640,N_49101);
and UO_406 (O_406,N_49583,N_49831);
nor UO_407 (O_407,N_48730,N_48742);
and UO_408 (O_408,N_49856,N_48550);
and UO_409 (O_409,N_48525,N_48451);
nand UO_410 (O_410,N_48215,N_49811);
nor UO_411 (O_411,N_49410,N_48129);
nand UO_412 (O_412,N_48192,N_49939);
and UO_413 (O_413,N_48212,N_49107);
nor UO_414 (O_414,N_48283,N_49659);
xor UO_415 (O_415,N_48326,N_49726);
nand UO_416 (O_416,N_48384,N_49633);
nand UO_417 (O_417,N_49792,N_48717);
and UO_418 (O_418,N_48068,N_48095);
nor UO_419 (O_419,N_48056,N_49753);
xnor UO_420 (O_420,N_49971,N_49715);
or UO_421 (O_421,N_48150,N_48926);
xor UO_422 (O_422,N_48991,N_49391);
nand UO_423 (O_423,N_49369,N_48051);
nor UO_424 (O_424,N_49455,N_49501);
nand UO_425 (O_425,N_48295,N_49791);
nor UO_426 (O_426,N_49092,N_49787);
nand UO_427 (O_427,N_48670,N_48254);
nor UO_428 (O_428,N_48208,N_48307);
and UO_429 (O_429,N_48586,N_48962);
and UO_430 (O_430,N_48988,N_49321);
xnor UO_431 (O_431,N_49669,N_48052);
nor UO_432 (O_432,N_49312,N_48585);
nand UO_433 (O_433,N_49296,N_48769);
nor UO_434 (O_434,N_48776,N_49855);
nand UO_435 (O_435,N_48300,N_49491);
and UO_436 (O_436,N_48169,N_48152);
xor UO_437 (O_437,N_48600,N_49502);
nand UO_438 (O_438,N_48024,N_49632);
or UO_439 (O_439,N_49821,N_49047);
xor UO_440 (O_440,N_48465,N_49763);
xnor UO_441 (O_441,N_48411,N_48098);
xor UO_442 (O_442,N_49654,N_48015);
xnor UO_443 (O_443,N_49220,N_48949);
nand UO_444 (O_444,N_48724,N_48294);
or UO_445 (O_445,N_48930,N_48026);
nand UO_446 (O_446,N_48179,N_48647);
nor UO_447 (O_447,N_48247,N_48851);
nor UO_448 (O_448,N_48923,N_48682);
and UO_449 (O_449,N_48886,N_48494);
or UO_450 (O_450,N_48413,N_48200);
nor UO_451 (O_451,N_49689,N_48088);
nor UO_452 (O_452,N_48953,N_48955);
and UO_453 (O_453,N_48298,N_49016);
xnor UO_454 (O_454,N_49394,N_48389);
or UO_455 (O_455,N_49730,N_48610);
xor UO_456 (O_456,N_49987,N_49587);
xor UO_457 (O_457,N_48653,N_48993);
xnor UO_458 (O_458,N_48499,N_49788);
or UO_459 (O_459,N_48438,N_49885);
and UO_460 (O_460,N_49758,N_49673);
nand UO_461 (O_461,N_48333,N_49957);
nand UO_462 (O_462,N_49985,N_49574);
nand UO_463 (O_463,N_48434,N_49243);
and UO_464 (O_464,N_49119,N_48097);
xor UO_465 (O_465,N_48617,N_49072);
or UO_466 (O_466,N_48468,N_49031);
xor UO_467 (O_467,N_49688,N_49531);
or UO_468 (O_468,N_49757,N_49044);
xor UO_469 (O_469,N_48059,N_49342);
xor UO_470 (O_470,N_49183,N_49552);
xor UO_471 (O_471,N_49057,N_48493);
xnor UO_472 (O_472,N_48147,N_49026);
xor UO_473 (O_473,N_49796,N_48139);
nor UO_474 (O_474,N_48609,N_49906);
nand UO_475 (O_475,N_48901,N_48917);
or UO_476 (O_476,N_49947,N_49727);
xor UO_477 (O_477,N_49311,N_48260);
nor UO_478 (O_478,N_49147,N_49760);
or UO_479 (O_479,N_49610,N_48755);
or UO_480 (O_480,N_48932,N_48246);
xor UO_481 (O_481,N_48745,N_48054);
nand UO_482 (O_482,N_49601,N_49841);
or UO_483 (O_483,N_48263,N_49604);
nor UO_484 (O_484,N_48436,N_48880);
nor UO_485 (O_485,N_48278,N_49651);
nor UO_486 (O_486,N_49397,N_48399);
and UO_487 (O_487,N_49551,N_49174);
and UO_488 (O_488,N_48449,N_49902);
xor UO_489 (O_489,N_48616,N_48159);
nand UO_490 (O_490,N_49761,N_49232);
nor UO_491 (O_491,N_48111,N_48698);
or UO_492 (O_492,N_48831,N_49851);
nand UO_493 (O_493,N_49084,N_49045);
and UO_494 (O_494,N_49500,N_48746);
nor UO_495 (O_495,N_49339,N_49588);
nand UO_496 (O_496,N_49933,N_49127);
nand UO_497 (O_497,N_48462,N_49722);
nand UO_498 (O_498,N_49605,N_49646);
and UO_499 (O_499,N_49690,N_48758);
or UO_500 (O_500,N_48965,N_48982);
xor UO_501 (O_501,N_49415,N_49725);
nand UO_502 (O_502,N_48058,N_48906);
xor UO_503 (O_503,N_48706,N_49624);
nor UO_504 (O_504,N_48117,N_49857);
xnor UO_505 (O_505,N_48773,N_49005);
or UO_506 (O_506,N_49285,N_48943);
and UO_507 (O_507,N_49400,N_49469);
and UO_508 (O_508,N_48070,N_49446);
xor UO_509 (O_509,N_48304,N_48646);
nand UO_510 (O_510,N_48370,N_48309);
and UO_511 (O_511,N_48049,N_48281);
and UO_512 (O_512,N_49476,N_48045);
nand UO_513 (O_513,N_48911,N_48429);
and UO_514 (O_514,N_48205,N_49064);
or UO_515 (O_515,N_49649,N_49920);
and UO_516 (O_516,N_49368,N_49980);
nand UO_517 (O_517,N_49493,N_49353);
nor UO_518 (O_518,N_48092,N_48065);
xnor UO_519 (O_519,N_48935,N_49963);
xor UO_520 (O_520,N_48770,N_49203);
or UO_521 (O_521,N_49937,N_49008);
or UO_522 (O_522,N_48633,N_49590);
or UO_523 (O_523,N_49218,N_48763);
or UO_524 (O_524,N_49810,N_49903);
and UO_525 (O_525,N_48632,N_49411);
nor UO_526 (O_526,N_48217,N_48440);
and UO_527 (O_527,N_49196,N_49454);
nand UO_528 (O_528,N_48067,N_48801);
xor UO_529 (O_529,N_49163,N_48142);
nand UO_530 (O_530,N_49699,N_49330);
and UO_531 (O_531,N_48318,N_48738);
nor UO_532 (O_532,N_48817,N_49059);
nor UO_533 (O_533,N_49346,N_48628);
and UO_534 (O_534,N_48009,N_48321);
xor UO_535 (O_535,N_49728,N_48504);
nor UO_536 (O_536,N_49647,N_49824);
nor UO_537 (O_537,N_48392,N_49329);
xor UO_538 (O_538,N_48857,N_49098);
nand UO_539 (O_539,N_48703,N_49020);
and UO_540 (O_540,N_48737,N_49461);
nor UO_541 (O_541,N_49662,N_49307);
xnor UO_542 (O_542,N_48041,N_48178);
or UO_543 (O_543,N_48626,N_49609);
or UO_544 (O_544,N_48595,N_49789);
and UO_545 (O_545,N_48927,N_48783);
nor UO_546 (O_546,N_48554,N_48578);
nand UO_547 (O_547,N_48790,N_49024);
or UO_548 (O_548,N_48656,N_48369);
nor UO_549 (O_549,N_48272,N_48518);
or UO_550 (O_550,N_49807,N_48089);
nor UO_551 (O_551,N_49225,N_49108);
or UO_552 (O_552,N_49445,N_48775);
xor UO_553 (O_553,N_49027,N_49069);
nand UO_554 (O_554,N_48910,N_48340);
nor UO_555 (O_555,N_49948,N_48243);
xor UO_556 (O_556,N_49398,N_48099);
and UO_557 (O_557,N_48226,N_48087);
and UO_558 (O_558,N_48536,N_49517);
and UO_559 (O_559,N_48676,N_48107);
or UO_560 (O_560,N_49829,N_48141);
and UO_561 (O_561,N_48976,N_49301);
nor UO_562 (O_562,N_49679,N_49806);
xnor UO_563 (O_563,N_48293,N_49908);
nor UO_564 (O_564,N_48106,N_49077);
or UO_565 (O_565,N_49462,N_49199);
nor UO_566 (O_566,N_48186,N_49288);
or UO_567 (O_567,N_49211,N_48577);
nor UO_568 (O_568,N_48061,N_48547);
xnor UO_569 (O_569,N_48823,N_48597);
or UO_570 (O_570,N_48777,N_48638);
nand UO_571 (O_571,N_49785,N_49882);
and UO_572 (O_572,N_48005,N_49618);
or UO_573 (O_573,N_49136,N_49166);
xor UO_574 (O_574,N_48778,N_48674);
or UO_575 (O_575,N_49198,N_49421);
or UO_576 (O_576,N_48360,N_49245);
or UO_577 (O_577,N_48454,N_48552);
nor UO_578 (O_578,N_48498,N_48786);
or UO_579 (O_579,N_49983,N_49103);
or UO_580 (O_580,N_49641,N_48787);
or UO_581 (O_581,N_48850,N_48347);
or UO_582 (O_582,N_48952,N_49643);
nand UO_583 (O_583,N_49678,N_48661);
nand UO_584 (O_584,N_49371,N_48637);
nand UO_585 (O_585,N_49694,N_49635);
or UO_586 (O_586,N_48667,N_49433);
or UO_587 (O_587,N_49240,N_49109);
nor UO_588 (O_588,N_48866,N_49668);
nor UO_589 (O_589,N_49034,N_48527);
xor UO_590 (O_590,N_49126,N_49228);
xnor UO_591 (O_591,N_49325,N_49692);
or UO_592 (O_592,N_49023,N_48849);
nor UO_593 (O_593,N_49594,N_48296);
nor UO_594 (O_594,N_48514,N_48380);
xor UO_595 (O_595,N_48043,N_48816);
xor UO_596 (O_596,N_48050,N_48391);
nand UO_597 (O_597,N_48564,N_48218);
nor UO_598 (O_598,N_48940,N_49018);
xor UO_599 (O_599,N_48635,N_49599);
or UO_600 (O_600,N_48826,N_49991);
nand UO_601 (O_601,N_49859,N_49904);
nor UO_602 (O_602,N_48479,N_48933);
and UO_603 (O_603,N_49115,N_49819);
or UO_604 (O_604,N_48603,N_49929);
nor UO_605 (O_605,N_48027,N_48284);
nor UO_606 (O_606,N_49168,N_49112);
xor UO_607 (O_607,N_48534,N_48407);
nand UO_608 (O_608,N_48657,N_49797);
and UO_609 (O_609,N_48992,N_48834);
nand UO_610 (O_610,N_49627,N_48435);
or UO_611 (O_611,N_48034,N_48741);
nor UO_612 (O_612,N_49711,N_48508);
or UO_613 (O_613,N_48853,N_48474);
xor UO_614 (O_614,N_49786,N_49385);
nor UO_615 (O_615,N_48184,N_49843);
or UO_616 (O_616,N_48471,N_49159);
and UO_617 (O_617,N_48483,N_49248);
xor UO_618 (O_618,N_48569,N_48785);
or UO_619 (O_619,N_48383,N_48568);
nand UO_620 (O_620,N_49176,N_48155);
or UO_621 (O_621,N_48332,N_49710);
nand UO_622 (O_622,N_49614,N_49773);
xnor UO_623 (O_623,N_48154,N_48902);
and UO_624 (O_624,N_49360,N_48170);
nor UO_625 (O_625,N_48153,N_48663);
and UO_626 (O_626,N_49158,N_49495);
nand UO_627 (O_627,N_48404,N_49310);
nor UO_628 (O_628,N_49755,N_48076);
xnor UO_629 (O_629,N_49716,N_49648);
or UO_630 (O_630,N_48845,N_49464);
xnor UO_631 (O_631,N_48553,N_49842);
and UO_632 (O_632,N_48928,N_49138);
nor UO_633 (O_633,N_49095,N_48345);
nor UO_634 (O_634,N_49324,N_49914);
nand UO_635 (O_635,N_48596,N_49580);
and UO_636 (O_636,N_49712,N_49075);
nor UO_637 (O_637,N_48428,N_48048);
xnor UO_638 (O_638,N_49751,N_48791);
or UO_639 (O_639,N_49510,N_49049);
and UO_640 (O_640,N_48999,N_49177);
nand UO_641 (O_641,N_49221,N_49076);
xnor UO_642 (O_642,N_48843,N_49124);
or UO_643 (O_643,N_49009,N_48555);
and UO_644 (O_644,N_49778,N_48686);
and UO_645 (O_645,N_48422,N_49440);
nor UO_646 (O_646,N_49931,N_48629);
and UO_647 (O_647,N_48771,N_49899);
or UO_648 (O_648,N_48812,N_48496);
nand UO_649 (O_649,N_49351,N_49486);
nand UO_650 (O_650,N_49675,N_48548);
or UO_651 (O_651,N_48037,N_48779);
nand UO_652 (O_652,N_49141,N_49905);
and UO_653 (O_653,N_49494,N_49333);
or UO_654 (O_654,N_49017,N_48057);
nand UO_655 (O_655,N_49367,N_48767);
nor UO_656 (O_656,N_49747,N_49873);
xor UO_657 (O_657,N_48229,N_48075);
nor UO_658 (O_658,N_49078,N_49671);
nand UO_659 (O_659,N_48725,N_48576);
nor UO_660 (O_660,N_48133,N_49223);
and UO_661 (O_661,N_49564,N_49261);
or UO_662 (O_662,N_48225,N_49572);
or UO_663 (O_663,N_49477,N_49392);
or UO_664 (O_664,N_49852,N_49549);
nor UO_665 (O_665,N_49458,N_49865);
and UO_666 (O_666,N_48806,N_49949);
or UO_667 (O_667,N_49447,N_49219);
or UO_668 (O_668,N_49015,N_48545);
or UO_669 (O_669,N_48244,N_48108);
xnor UO_670 (O_670,N_48180,N_49463);
nand UO_671 (O_671,N_48181,N_49374);
nor UO_672 (O_672,N_49409,N_48036);
or UO_673 (O_673,N_49091,N_48689);
or UO_674 (O_674,N_48966,N_49422);
xor UO_675 (O_675,N_48800,N_49279);
xnor UO_676 (O_676,N_49930,N_49315);
or UO_677 (O_677,N_49297,N_48038);
xnor UO_678 (O_678,N_48516,N_48250);
nand UO_679 (O_679,N_49423,N_49066);
xor UO_680 (O_680,N_49065,N_48565);
and UO_681 (O_681,N_49067,N_49867);
nand UO_682 (O_682,N_48848,N_49656);
xnor UO_683 (O_683,N_48723,N_48665);
xnor UO_684 (O_684,N_49299,N_49164);
xor UO_685 (O_685,N_48022,N_49615);
xor UO_686 (O_686,N_48276,N_48997);
or UO_687 (O_687,N_49475,N_48401);
and UO_688 (O_688,N_48373,N_49195);
or UO_689 (O_689,N_49524,N_48618);
or UO_690 (O_690,N_49942,N_49226);
xnor UO_691 (O_691,N_49783,N_48865);
and UO_692 (O_692,N_49214,N_49320);
nor UO_693 (O_693,N_49269,N_48228);
nand UO_694 (O_694,N_48393,N_48395);
or UO_695 (O_695,N_48838,N_48870);
nor UO_696 (O_696,N_49387,N_49645);
or UO_697 (O_697,N_49007,N_49251);
xor UO_698 (O_698,N_49468,N_49887);
nand UO_699 (O_699,N_49488,N_48894);
nor UO_700 (O_700,N_49717,N_48941);
xor UO_701 (O_701,N_49503,N_49316);
or UO_702 (O_702,N_48895,N_49840);
or UO_703 (O_703,N_49743,N_48338);
or UO_704 (O_704,N_48114,N_49532);
or UO_705 (O_705,N_49452,N_49724);
and UO_706 (O_706,N_49850,N_48115);
nor UO_707 (O_707,N_48625,N_48374);
nand UO_708 (O_708,N_49350,N_48828);
and UO_709 (O_709,N_49630,N_49087);
xor UO_710 (O_710,N_49910,N_48750);
and UO_711 (O_711,N_49349,N_49505);
xor UO_712 (O_712,N_48799,N_49483);
nor UO_713 (O_713,N_48227,N_49470);
nor UO_714 (O_714,N_49871,N_49701);
nand UO_715 (O_715,N_49642,N_49869);
or UO_716 (O_716,N_48261,N_49975);
nor UO_717 (O_717,N_49133,N_48487);
or UO_718 (O_718,N_48964,N_48563);
nor UO_719 (O_719,N_49436,N_49083);
xnor UO_720 (O_720,N_48233,N_49111);
and UO_721 (O_721,N_48796,N_48096);
nor UO_722 (O_722,N_48206,N_48012);
or UO_723 (O_723,N_49332,N_48351);
nand UO_724 (O_724,N_48262,N_48920);
or UO_725 (O_725,N_48808,N_48014);
nor UO_726 (O_726,N_48222,N_49663);
nor UO_727 (O_727,N_49858,N_48589);
and UO_728 (O_728,N_48343,N_49833);
xnor UO_729 (O_729,N_49714,N_48641);
nor UO_730 (O_730,N_48489,N_48492);
xnor UO_731 (O_731,N_49407,N_48780);
xnor UO_732 (O_732,N_48766,N_49560);
nor UO_733 (O_733,N_49818,N_48348);
or UO_734 (O_734,N_49967,N_48140);
xnor UO_735 (O_735,N_48336,N_48060);
nor UO_736 (O_736,N_49492,N_49117);
and UO_737 (O_737,N_49839,N_49974);
xnor UO_738 (O_738,N_48887,N_49602);
and UO_739 (O_739,N_48450,N_49173);
and UO_740 (O_740,N_48379,N_49406);
nor UO_741 (O_741,N_49666,N_49854);
or UO_742 (O_742,N_49883,N_48537);
nor UO_743 (O_743,N_49359,N_48235);
or UO_744 (O_744,N_48388,N_49934);
or UO_745 (O_745,N_48311,N_48575);
and UO_746 (O_746,N_48713,N_48077);
and UO_747 (O_747,N_48639,N_48362);
nand UO_748 (O_748,N_49917,N_48986);
nor UO_749 (O_749,N_49110,N_49278);
xnor UO_750 (O_750,N_49927,N_48258);
or UO_751 (O_751,N_48007,N_49916);
nand UO_752 (O_752,N_48836,N_48611);
nand UO_753 (O_753,N_49874,N_49540);
nand UO_754 (O_754,N_49511,N_48891);
and UO_755 (O_755,N_48341,N_48069);
or UO_756 (O_756,N_48683,N_48031);
or UO_757 (O_757,N_49135,N_48852);
xor UO_758 (O_758,N_49731,N_48945);
nand UO_759 (O_759,N_49471,N_49250);
nor UO_760 (O_760,N_49693,N_48606);
nand UO_761 (O_761,N_49626,N_49201);
nand UO_762 (O_762,N_49338,N_48761);
or UO_763 (O_763,N_49236,N_48972);
xnor UO_764 (O_764,N_48085,N_49657);
nor UO_765 (O_765,N_48650,N_49754);
or UO_766 (O_766,N_49430,N_49998);
and UO_767 (O_767,N_49181,N_49732);
nand UO_768 (O_768,N_48259,N_49386);
nand UO_769 (O_769,N_49019,N_48473);
or UO_770 (O_770,N_49235,N_48695);
xnor UO_771 (O_771,N_48813,N_48040);
or UO_772 (O_772,N_48840,N_48556);
xnor UO_773 (O_773,N_48339,N_48039);
nor UO_774 (O_774,N_49922,N_48672);
nand UO_775 (O_775,N_48209,N_48961);
and UO_776 (O_776,N_49372,N_49068);
and UO_777 (O_777,N_49990,N_48511);
nor UO_778 (O_778,N_49896,N_48692);
nand UO_779 (O_779,N_48919,N_49012);
and UO_780 (O_780,N_48820,N_48734);
nand UO_781 (O_781,N_48485,N_48361);
nand UO_782 (O_782,N_49082,N_49568);
nor UO_783 (O_783,N_49313,N_48774);
or UO_784 (O_784,N_48681,N_48591);
or UO_785 (O_785,N_48743,N_49504);
nor UO_786 (O_786,N_49412,N_49093);
nand UO_787 (O_787,N_49389,N_49363);
nand UO_788 (O_788,N_49071,N_49449);
or UO_789 (O_789,N_49512,N_48847);
or UO_790 (O_790,N_48432,N_49130);
and UO_791 (O_791,N_49264,N_48105);
and UO_792 (O_792,N_49227,N_49134);
nand UO_793 (O_793,N_48756,N_48685);
and UO_794 (O_794,N_48867,N_49611);
and UO_795 (O_795,N_48241,N_48747);
or UO_796 (O_796,N_48275,N_48967);
nand UO_797 (O_797,N_49720,N_48437);
nand UO_798 (O_798,N_49608,N_48470);
nor UO_799 (O_799,N_49145,N_48963);
nand UO_800 (O_800,N_48540,N_49242);
xnor UO_801 (O_801,N_48792,N_48598);
nand UO_802 (O_802,N_48412,N_48245);
nor UO_803 (O_803,N_48739,N_49148);
xor UO_804 (O_804,N_49557,N_49081);
nor UO_805 (O_805,N_48082,N_48190);
and UO_806 (O_806,N_49598,N_49848);
xor UO_807 (O_807,N_48648,N_48249);
and UO_808 (O_808,N_48714,N_48579);
and UO_809 (O_809,N_48995,N_49822);
nor UO_810 (O_810,N_49518,N_48884);
nand UO_811 (O_811,N_48256,N_48549);
or UO_812 (O_812,N_48135,N_48587);
nor UO_813 (O_813,N_49035,N_48312);
nor UO_814 (O_814,N_49737,N_49003);
and UO_815 (O_815,N_48856,N_48264);
and UO_816 (O_816,N_49323,N_49891);
xnor UO_817 (O_817,N_49940,N_48002);
nand UO_818 (O_818,N_48160,N_49558);
nand UO_819 (O_819,N_48868,N_48869);
or UO_820 (O_820,N_49281,N_49613);
nand UO_821 (O_821,N_49901,N_48833);
and UO_822 (O_822,N_49380,N_49094);
xnor UO_823 (O_823,N_48684,N_48837);
nand UO_824 (O_824,N_49499,N_49739);
nor UO_825 (O_825,N_49249,N_49073);
and UO_826 (O_826,N_49487,N_49384);
or UO_827 (O_827,N_49197,N_49011);
xor UO_828 (O_828,N_49096,N_49674);
nor UO_829 (O_829,N_49202,N_49347);
and UO_830 (O_830,N_49131,N_48960);
xnor UO_831 (O_831,N_48119,N_48983);
xnor UO_832 (O_832,N_48277,N_49263);
or UO_833 (O_833,N_48213,N_49770);
and UO_834 (O_834,N_48240,N_48280);
xor UO_835 (O_835,N_49589,N_49438);
or UO_836 (O_836,N_48863,N_49600);
and UO_837 (O_837,N_48017,N_48330);
xor UO_838 (O_838,N_49291,N_49625);
xnor UO_839 (O_839,N_48631,N_49828);
nor UO_840 (O_840,N_49545,N_49667);
or UO_841 (O_841,N_49215,N_48080);
xor UO_842 (O_842,N_48956,N_48722);
xor UO_843 (O_843,N_48112,N_48768);
or UO_844 (O_844,N_48355,N_49519);
nor UO_845 (O_845,N_49208,N_49997);
xor UO_846 (O_846,N_48291,N_48136);
nor UO_847 (O_847,N_49074,N_48574);
or UO_848 (O_848,N_49230,N_49813);
xor UO_849 (O_849,N_49038,N_49238);
nand UO_850 (O_850,N_48580,N_49336);
nor UO_851 (O_851,N_48642,N_49812);
and UO_852 (O_852,N_49253,N_48950);
nor UO_853 (O_853,N_48918,N_48320);
and UO_854 (O_854,N_49151,N_49660);
nand UO_855 (O_855,N_48405,N_49969);
nor UO_856 (O_856,N_48376,N_49254);
xor UO_857 (O_857,N_48690,N_49709);
xnor UO_858 (O_858,N_48710,N_49480);
or UO_859 (O_859,N_49414,N_49582);
nor UO_860 (O_860,N_48486,N_48975);
nor UO_861 (O_861,N_48506,N_48188);
nand UO_862 (O_862,N_49327,N_49713);
and UO_863 (O_863,N_49473,N_49237);
nor UO_864 (O_864,N_48716,N_49619);
or UO_865 (O_865,N_49977,N_49205);
nor UO_866 (O_866,N_49060,N_48316);
nor UO_867 (O_867,N_49156,N_49794);
xnor UO_868 (O_868,N_49893,N_49817);
nor UO_869 (O_869,N_48409,N_49798);
xor UO_870 (O_870,N_48010,N_48614);
or UO_871 (O_871,N_48455,N_49562);
nand UO_872 (O_872,N_48979,N_49996);
nor UO_873 (O_873,N_48189,N_49960);
xnor UO_874 (O_874,N_48081,N_48346);
or UO_875 (O_875,N_49734,N_48571);
and UO_876 (O_876,N_48592,N_49569);
nand UO_877 (O_877,N_49554,N_48922);
xor UO_878 (O_878,N_48457,N_49161);
xor UO_879 (O_879,N_49976,N_49527);
or UO_880 (O_880,N_49814,N_49431);
or UO_881 (O_881,N_48398,N_48519);
xnor UO_882 (O_882,N_48623,N_48885);
nor UO_883 (O_883,N_48132,N_48378);
nor UO_884 (O_884,N_48366,N_48385);
nor UO_885 (O_885,N_49377,N_49413);
xor UO_886 (O_886,N_49000,N_49687);
and UO_887 (O_887,N_49063,N_48602);
or UO_888 (O_888,N_48936,N_48588);
and UO_889 (O_889,N_48805,N_48753);
nor UO_890 (O_890,N_49876,N_49335);
nor UO_891 (O_891,N_48538,N_48528);
nand UO_892 (O_892,N_48608,N_48257);
xnor UO_893 (O_893,N_49058,N_48381);
or UO_894 (O_894,N_49340,N_49256);
nand UO_895 (O_895,N_48288,N_49036);
and UO_896 (O_896,N_49522,N_49945);
and UO_897 (O_897,N_49862,N_48237);
xor UO_898 (O_898,N_49875,N_48601);
nor UO_899 (O_899,N_48337,N_49186);
nor UO_900 (O_900,N_49276,N_48582);
or UO_901 (O_901,N_49578,N_48551);
or UO_902 (O_902,N_48367,N_49802);
nand UO_903 (O_903,N_48365,N_49979);
nor UO_904 (O_904,N_48740,N_48363);
nand UO_905 (O_905,N_48248,N_48145);
and UO_906 (O_906,N_49204,N_48176);
nand UO_907 (O_907,N_48978,N_48163);
nor UO_908 (O_908,N_49489,N_48306);
or UO_909 (O_909,N_48459,N_49968);
and UO_910 (O_910,N_48951,N_49526);
nand UO_911 (O_911,N_49029,N_48323);
xnor UO_912 (O_912,N_49165,N_48827);
nand UO_913 (O_913,N_49129,N_48804);
or UO_914 (O_914,N_49682,N_49536);
or UO_915 (O_915,N_48732,N_48267);
nor UO_916 (O_916,N_49054,N_49907);
nand UO_917 (O_917,N_48882,N_49172);
and UO_918 (O_918,N_49836,N_48424);
xnor UO_919 (O_919,N_48973,N_48131);
and UO_920 (O_920,N_48285,N_48214);
or UO_921 (O_921,N_48652,N_48083);
nand UO_922 (O_922,N_48814,N_48458);
or UO_923 (O_923,N_48526,N_48604);
nor UO_924 (O_924,N_49696,N_49356);
or UO_925 (O_925,N_48535,N_49190);
and UO_926 (O_926,N_49683,N_48809);
and UO_927 (O_927,N_48835,N_48101);
nand UO_928 (O_928,N_49508,N_49520);
nor UO_929 (O_929,N_49497,N_48954);
nor UO_930 (O_930,N_48086,N_48959);
and UO_931 (O_931,N_49879,N_49776);
xor UO_932 (O_932,N_49685,N_48872);
nand UO_933 (O_933,N_48570,N_48731);
and UO_934 (O_934,N_48122,N_49808);
or UO_935 (O_935,N_48204,N_49184);
nor UO_936 (O_936,N_48675,N_48016);
and UO_937 (O_937,N_49030,N_49870);
and UO_938 (O_938,N_48167,N_48137);
and UO_939 (O_939,N_48594,N_49752);
xnor UO_940 (O_940,N_49122,N_48354);
nand UO_941 (O_941,N_49140,N_49994);
nor UO_942 (O_942,N_48314,N_49644);
or UO_943 (O_943,N_49282,N_48305);
or UO_944 (O_944,N_49418,N_48772);
nand UO_945 (O_945,N_48729,N_48334);
and UO_946 (O_946,N_48744,N_49877);
xnor UO_947 (O_947,N_49775,N_49790);
nand UO_948 (O_948,N_48854,N_49864);
and UO_949 (O_949,N_49185,N_49984);
nor UO_950 (O_950,N_49837,N_49120);
or UO_951 (O_951,N_48818,N_49537);
or UO_952 (O_952,N_48325,N_48517);
or UO_953 (O_953,N_49037,N_48915);
nand UO_954 (O_954,N_48622,N_48694);
nand UO_955 (O_955,N_49769,N_49704);
nor UO_956 (O_956,N_49764,N_49534);
nand UO_957 (O_957,N_49943,N_49616);
and UO_958 (O_958,N_49652,N_48707);
or UO_959 (O_959,N_49428,N_48151);
nor UO_960 (O_960,N_48165,N_48042);
or UO_961 (O_961,N_48442,N_49981);
and UO_962 (O_962,N_49913,N_48680);
or UO_963 (O_963,N_48669,N_48195);
or UO_964 (O_964,N_49523,N_48327);
or UO_965 (O_965,N_49304,N_48718);
or UO_966 (O_966,N_49880,N_49838);
nor UO_967 (O_967,N_49212,N_49052);
or UO_968 (O_968,N_49538,N_48765);
nand UO_969 (O_969,N_48513,N_49343);
and UO_970 (O_970,N_49187,N_48752);
nor UO_971 (O_971,N_49697,N_48693);
nor UO_972 (O_972,N_49171,N_48651);
nor UO_973 (O_973,N_49189,N_48023);
nand UO_974 (O_974,N_49450,N_49160);
nand UO_975 (O_975,N_49479,N_48008);
nor UO_976 (O_976,N_49088,N_49677);
or UO_977 (O_977,N_48699,N_49442);
xnor UO_978 (O_978,N_49958,N_48230);
or UO_979 (O_979,N_48658,N_48194);
nor UO_980 (O_980,N_49053,N_48510);
nand UO_981 (O_981,N_49319,N_49964);
or UO_982 (O_982,N_49061,N_49267);
nor UO_983 (O_983,N_48199,N_48491);
nor UO_984 (O_984,N_49210,N_48883);
and UO_985 (O_985,N_48116,N_49328);
and UO_986 (O_986,N_48445,N_48700);
nor UO_987 (O_987,N_49516,N_48560);
nand UO_988 (O_988,N_48624,N_49911);
and UO_989 (O_989,N_49070,N_48712);
xnor UO_990 (O_990,N_49514,N_48100);
or UO_991 (O_991,N_48781,N_49846);
nand UO_992 (O_992,N_49234,N_48998);
and UO_993 (O_993,N_48977,N_49918);
nand UO_994 (O_994,N_49954,N_49935);
or UO_995 (O_995,N_48011,N_49100);
nor UO_996 (O_996,N_49381,N_49705);
and UO_997 (O_997,N_48231,N_48900);
xnor UO_998 (O_998,N_48162,N_49530);
and UO_999 (O_999,N_48467,N_48659);
and UO_1000 (O_1000,N_48353,N_48415);
nor UO_1001 (O_1001,N_48529,N_48065);
and UO_1002 (O_1002,N_48349,N_49170);
xnor UO_1003 (O_1003,N_48993,N_49956);
nand UO_1004 (O_1004,N_49848,N_49851);
nand UO_1005 (O_1005,N_49148,N_49415);
nor UO_1006 (O_1006,N_49630,N_49669);
or UO_1007 (O_1007,N_48390,N_49611);
nor UO_1008 (O_1008,N_49122,N_48635);
xnor UO_1009 (O_1009,N_48618,N_49556);
nand UO_1010 (O_1010,N_49773,N_48490);
nor UO_1011 (O_1011,N_48580,N_48596);
and UO_1012 (O_1012,N_49969,N_49329);
xor UO_1013 (O_1013,N_49868,N_49036);
xor UO_1014 (O_1014,N_49579,N_49299);
and UO_1015 (O_1015,N_49911,N_48611);
xnor UO_1016 (O_1016,N_48509,N_48087);
and UO_1017 (O_1017,N_49312,N_48316);
or UO_1018 (O_1018,N_49916,N_49345);
xnor UO_1019 (O_1019,N_48781,N_49637);
or UO_1020 (O_1020,N_48197,N_48270);
or UO_1021 (O_1021,N_49193,N_48326);
and UO_1022 (O_1022,N_48471,N_49882);
nand UO_1023 (O_1023,N_49274,N_48213);
or UO_1024 (O_1024,N_49957,N_49885);
or UO_1025 (O_1025,N_48486,N_49939);
nor UO_1026 (O_1026,N_49387,N_49403);
or UO_1027 (O_1027,N_49201,N_49643);
xnor UO_1028 (O_1028,N_49010,N_48216);
and UO_1029 (O_1029,N_48433,N_49957);
xor UO_1030 (O_1030,N_49560,N_49343);
or UO_1031 (O_1031,N_48712,N_48270);
nor UO_1032 (O_1032,N_48841,N_49452);
xnor UO_1033 (O_1033,N_48244,N_48019);
nor UO_1034 (O_1034,N_48219,N_49923);
xnor UO_1035 (O_1035,N_48046,N_48758);
or UO_1036 (O_1036,N_49510,N_48509);
or UO_1037 (O_1037,N_48222,N_48974);
and UO_1038 (O_1038,N_48295,N_48547);
nand UO_1039 (O_1039,N_48353,N_49950);
nand UO_1040 (O_1040,N_48177,N_48467);
xor UO_1041 (O_1041,N_48703,N_49901);
xor UO_1042 (O_1042,N_48225,N_49853);
nand UO_1043 (O_1043,N_49770,N_49231);
and UO_1044 (O_1044,N_48063,N_48337);
nand UO_1045 (O_1045,N_49876,N_48155);
nor UO_1046 (O_1046,N_48347,N_49697);
or UO_1047 (O_1047,N_48165,N_49012);
nand UO_1048 (O_1048,N_49601,N_49416);
or UO_1049 (O_1049,N_49424,N_48581);
nand UO_1050 (O_1050,N_49520,N_49036);
nor UO_1051 (O_1051,N_49749,N_48497);
nor UO_1052 (O_1052,N_48765,N_49015);
and UO_1053 (O_1053,N_49913,N_48508);
nor UO_1054 (O_1054,N_49646,N_48652);
xor UO_1055 (O_1055,N_49037,N_49082);
xor UO_1056 (O_1056,N_48210,N_49517);
nand UO_1057 (O_1057,N_49802,N_48421);
nor UO_1058 (O_1058,N_48223,N_49502);
nor UO_1059 (O_1059,N_48793,N_49287);
nand UO_1060 (O_1060,N_49101,N_49144);
xor UO_1061 (O_1061,N_49882,N_49226);
nor UO_1062 (O_1062,N_49321,N_48613);
and UO_1063 (O_1063,N_48896,N_48486);
and UO_1064 (O_1064,N_49616,N_48376);
or UO_1065 (O_1065,N_48049,N_49458);
or UO_1066 (O_1066,N_49722,N_48082);
nand UO_1067 (O_1067,N_49445,N_49540);
or UO_1068 (O_1068,N_49594,N_49397);
and UO_1069 (O_1069,N_48174,N_49420);
xor UO_1070 (O_1070,N_49827,N_48055);
and UO_1071 (O_1071,N_48238,N_48752);
nand UO_1072 (O_1072,N_48239,N_48594);
nor UO_1073 (O_1073,N_49730,N_48579);
or UO_1074 (O_1074,N_49091,N_49780);
nand UO_1075 (O_1075,N_49724,N_49579);
xor UO_1076 (O_1076,N_49047,N_49050);
nor UO_1077 (O_1077,N_48629,N_49999);
nor UO_1078 (O_1078,N_49441,N_48319);
nor UO_1079 (O_1079,N_49183,N_49860);
nor UO_1080 (O_1080,N_48789,N_49906);
nor UO_1081 (O_1081,N_48592,N_48420);
and UO_1082 (O_1082,N_49165,N_49213);
nand UO_1083 (O_1083,N_49386,N_48203);
and UO_1084 (O_1084,N_49068,N_49665);
or UO_1085 (O_1085,N_48142,N_49001);
nand UO_1086 (O_1086,N_49089,N_49905);
and UO_1087 (O_1087,N_48579,N_49500);
nor UO_1088 (O_1088,N_48637,N_48674);
nor UO_1089 (O_1089,N_49090,N_49106);
or UO_1090 (O_1090,N_48349,N_49149);
xnor UO_1091 (O_1091,N_48695,N_48550);
nand UO_1092 (O_1092,N_48237,N_49321);
xnor UO_1093 (O_1093,N_48874,N_49537);
and UO_1094 (O_1094,N_48833,N_49804);
and UO_1095 (O_1095,N_48864,N_49314);
nor UO_1096 (O_1096,N_48665,N_49275);
or UO_1097 (O_1097,N_49712,N_48452);
nand UO_1098 (O_1098,N_49570,N_49703);
or UO_1099 (O_1099,N_48800,N_49872);
nand UO_1100 (O_1100,N_48392,N_49752);
or UO_1101 (O_1101,N_48557,N_48797);
nor UO_1102 (O_1102,N_48486,N_48446);
xor UO_1103 (O_1103,N_49649,N_49373);
nor UO_1104 (O_1104,N_49601,N_49357);
nor UO_1105 (O_1105,N_49993,N_48500);
xor UO_1106 (O_1106,N_48182,N_48565);
nand UO_1107 (O_1107,N_49053,N_48616);
and UO_1108 (O_1108,N_49799,N_48779);
or UO_1109 (O_1109,N_48921,N_48298);
nor UO_1110 (O_1110,N_48099,N_48088);
nand UO_1111 (O_1111,N_48485,N_49510);
and UO_1112 (O_1112,N_49494,N_49293);
or UO_1113 (O_1113,N_49653,N_48210);
xor UO_1114 (O_1114,N_48790,N_49338);
and UO_1115 (O_1115,N_49606,N_49373);
and UO_1116 (O_1116,N_49923,N_49245);
or UO_1117 (O_1117,N_49292,N_49363);
nor UO_1118 (O_1118,N_48957,N_49370);
nor UO_1119 (O_1119,N_49428,N_48216);
nor UO_1120 (O_1120,N_49892,N_49594);
nor UO_1121 (O_1121,N_48205,N_48008);
nand UO_1122 (O_1122,N_48614,N_48324);
nor UO_1123 (O_1123,N_48901,N_49818);
or UO_1124 (O_1124,N_48459,N_49542);
or UO_1125 (O_1125,N_48678,N_48032);
and UO_1126 (O_1126,N_48913,N_49400);
nand UO_1127 (O_1127,N_48843,N_49749);
nand UO_1128 (O_1128,N_49567,N_49883);
nor UO_1129 (O_1129,N_48805,N_49303);
xnor UO_1130 (O_1130,N_49503,N_48593);
nor UO_1131 (O_1131,N_49456,N_49556);
and UO_1132 (O_1132,N_49216,N_49418);
or UO_1133 (O_1133,N_48434,N_49840);
or UO_1134 (O_1134,N_48462,N_49707);
nand UO_1135 (O_1135,N_49254,N_48618);
and UO_1136 (O_1136,N_49338,N_49743);
and UO_1137 (O_1137,N_49201,N_49001);
nor UO_1138 (O_1138,N_49843,N_49210);
and UO_1139 (O_1139,N_49422,N_48416);
or UO_1140 (O_1140,N_48673,N_48493);
nor UO_1141 (O_1141,N_49103,N_49850);
nand UO_1142 (O_1142,N_48243,N_48312);
or UO_1143 (O_1143,N_48530,N_49734);
and UO_1144 (O_1144,N_48561,N_48978);
and UO_1145 (O_1145,N_48170,N_49801);
or UO_1146 (O_1146,N_48606,N_49848);
nor UO_1147 (O_1147,N_49724,N_49881);
xor UO_1148 (O_1148,N_48526,N_49996);
or UO_1149 (O_1149,N_48359,N_48875);
nor UO_1150 (O_1150,N_48663,N_49250);
or UO_1151 (O_1151,N_48813,N_48802);
and UO_1152 (O_1152,N_49807,N_48199);
nand UO_1153 (O_1153,N_48447,N_49750);
xnor UO_1154 (O_1154,N_48258,N_49408);
or UO_1155 (O_1155,N_49235,N_49869);
nor UO_1156 (O_1156,N_49382,N_48101);
xor UO_1157 (O_1157,N_48477,N_48407);
xor UO_1158 (O_1158,N_49150,N_49605);
nor UO_1159 (O_1159,N_49231,N_49827);
and UO_1160 (O_1160,N_49579,N_49387);
or UO_1161 (O_1161,N_48335,N_48348);
or UO_1162 (O_1162,N_49014,N_49475);
nand UO_1163 (O_1163,N_49064,N_49553);
or UO_1164 (O_1164,N_48395,N_48953);
xnor UO_1165 (O_1165,N_48121,N_48380);
nor UO_1166 (O_1166,N_48293,N_48762);
or UO_1167 (O_1167,N_48196,N_48095);
nor UO_1168 (O_1168,N_49088,N_48858);
nor UO_1169 (O_1169,N_49183,N_48162);
or UO_1170 (O_1170,N_49956,N_48550);
nand UO_1171 (O_1171,N_49350,N_49789);
nand UO_1172 (O_1172,N_48505,N_49295);
xor UO_1173 (O_1173,N_48444,N_49491);
and UO_1174 (O_1174,N_48024,N_48207);
and UO_1175 (O_1175,N_49041,N_49724);
xnor UO_1176 (O_1176,N_48967,N_48931);
nor UO_1177 (O_1177,N_48299,N_49968);
nor UO_1178 (O_1178,N_49152,N_48303);
nand UO_1179 (O_1179,N_48127,N_48001);
nor UO_1180 (O_1180,N_48203,N_49942);
nor UO_1181 (O_1181,N_48085,N_48040);
xnor UO_1182 (O_1182,N_49974,N_48066);
and UO_1183 (O_1183,N_49908,N_48927);
nand UO_1184 (O_1184,N_48088,N_48571);
xnor UO_1185 (O_1185,N_48218,N_49885);
xnor UO_1186 (O_1186,N_48456,N_49235);
nor UO_1187 (O_1187,N_49884,N_49720);
and UO_1188 (O_1188,N_48654,N_49416);
nand UO_1189 (O_1189,N_49709,N_48250);
and UO_1190 (O_1190,N_49295,N_49495);
nor UO_1191 (O_1191,N_49932,N_48176);
and UO_1192 (O_1192,N_49378,N_48389);
and UO_1193 (O_1193,N_49916,N_49828);
nand UO_1194 (O_1194,N_48797,N_49250);
nand UO_1195 (O_1195,N_48390,N_49621);
nand UO_1196 (O_1196,N_48299,N_48204);
nand UO_1197 (O_1197,N_49376,N_48710);
nor UO_1198 (O_1198,N_49880,N_48425);
or UO_1199 (O_1199,N_48489,N_48282);
nand UO_1200 (O_1200,N_48334,N_49464);
or UO_1201 (O_1201,N_48307,N_48967);
nand UO_1202 (O_1202,N_48984,N_48271);
and UO_1203 (O_1203,N_49098,N_49811);
or UO_1204 (O_1204,N_49479,N_49769);
or UO_1205 (O_1205,N_49763,N_48960);
nand UO_1206 (O_1206,N_48908,N_49153);
and UO_1207 (O_1207,N_49141,N_49038);
nor UO_1208 (O_1208,N_49793,N_48083);
nor UO_1209 (O_1209,N_49297,N_49277);
nand UO_1210 (O_1210,N_49434,N_48570);
and UO_1211 (O_1211,N_48746,N_48318);
or UO_1212 (O_1212,N_48931,N_48583);
nand UO_1213 (O_1213,N_48330,N_48900);
or UO_1214 (O_1214,N_48550,N_49010);
nand UO_1215 (O_1215,N_49944,N_49484);
and UO_1216 (O_1216,N_49255,N_49276);
and UO_1217 (O_1217,N_49550,N_48425);
xnor UO_1218 (O_1218,N_48659,N_48641);
or UO_1219 (O_1219,N_48440,N_49535);
nand UO_1220 (O_1220,N_48062,N_48448);
nand UO_1221 (O_1221,N_49035,N_49474);
and UO_1222 (O_1222,N_48029,N_49261);
or UO_1223 (O_1223,N_48073,N_49315);
nand UO_1224 (O_1224,N_48852,N_49592);
or UO_1225 (O_1225,N_48138,N_49476);
xnor UO_1226 (O_1226,N_49329,N_48205);
nand UO_1227 (O_1227,N_49669,N_49892);
nand UO_1228 (O_1228,N_49211,N_49841);
and UO_1229 (O_1229,N_48670,N_49807);
nor UO_1230 (O_1230,N_49731,N_48134);
xor UO_1231 (O_1231,N_48273,N_49774);
or UO_1232 (O_1232,N_48276,N_48490);
and UO_1233 (O_1233,N_48866,N_49304);
nand UO_1234 (O_1234,N_49257,N_48077);
xor UO_1235 (O_1235,N_48027,N_48884);
and UO_1236 (O_1236,N_48278,N_49269);
xnor UO_1237 (O_1237,N_48421,N_48767);
nand UO_1238 (O_1238,N_48941,N_49702);
nor UO_1239 (O_1239,N_49962,N_48932);
nand UO_1240 (O_1240,N_48873,N_49479);
and UO_1241 (O_1241,N_49507,N_49362);
or UO_1242 (O_1242,N_49244,N_48250);
nor UO_1243 (O_1243,N_49821,N_48954);
and UO_1244 (O_1244,N_48036,N_48701);
xor UO_1245 (O_1245,N_48607,N_49210);
and UO_1246 (O_1246,N_48208,N_48435);
xor UO_1247 (O_1247,N_48772,N_49482);
xnor UO_1248 (O_1248,N_49930,N_48100);
xnor UO_1249 (O_1249,N_49157,N_48164);
nor UO_1250 (O_1250,N_48617,N_48616);
xnor UO_1251 (O_1251,N_48485,N_48043);
nor UO_1252 (O_1252,N_49249,N_49813);
nand UO_1253 (O_1253,N_49314,N_48624);
or UO_1254 (O_1254,N_49699,N_49462);
or UO_1255 (O_1255,N_49304,N_49928);
nand UO_1256 (O_1256,N_48916,N_48910);
xor UO_1257 (O_1257,N_49151,N_48492);
or UO_1258 (O_1258,N_48713,N_48907);
xnor UO_1259 (O_1259,N_49848,N_49168);
and UO_1260 (O_1260,N_48984,N_48507);
and UO_1261 (O_1261,N_49591,N_48777);
and UO_1262 (O_1262,N_48067,N_49562);
nand UO_1263 (O_1263,N_49141,N_49396);
nor UO_1264 (O_1264,N_49570,N_49921);
nand UO_1265 (O_1265,N_48849,N_48265);
nor UO_1266 (O_1266,N_49406,N_49495);
nor UO_1267 (O_1267,N_48108,N_48509);
xor UO_1268 (O_1268,N_48262,N_48953);
xnor UO_1269 (O_1269,N_48058,N_49014);
or UO_1270 (O_1270,N_48751,N_48320);
and UO_1271 (O_1271,N_48279,N_48431);
and UO_1272 (O_1272,N_49756,N_49015);
or UO_1273 (O_1273,N_48500,N_48685);
and UO_1274 (O_1274,N_48732,N_48990);
nand UO_1275 (O_1275,N_49615,N_49553);
or UO_1276 (O_1276,N_48944,N_48010);
or UO_1277 (O_1277,N_48424,N_49293);
nor UO_1278 (O_1278,N_49532,N_49651);
nor UO_1279 (O_1279,N_49673,N_48406);
nor UO_1280 (O_1280,N_48802,N_48585);
or UO_1281 (O_1281,N_49297,N_49629);
and UO_1282 (O_1282,N_49650,N_48027);
xnor UO_1283 (O_1283,N_49229,N_49039);
xor UO_1284 (O_1284,N_48571,N_49864);
nand UO_1285 (O_1285,N_48525,N_49221);
nand UO_1286 (O_1286,N_48790,N_49396);
nor UO_1287 (O_1287,N_48433,N_49376);
xnor UO_1288 (O_1288,N_48564,N_49353);
and UO_1289 (O_1289,N_49921,N_48665);
or UO_1290 (O_1290,N_48596,N_48338);
or UO_1291 (O_1291,N_48658,N_49342);
and UO_1292 (O_1292,N_49535,N_48543);
or UO_1293 (O_1293,N_48078,N_48370);
and UO_1294 (O_1294,N_48157,N_48839);
nor UO_1295 (O_1295,N_49269,N_49057);
xor UO_1296 (O_1296,N_49570,N_49102);
or UO_1297 (O_1297,N_49279,N_49052);
or UO_1298 (O_1298,N_49381,N_49004);
nor UO_1299 (O_1299,N_49381,N_49772);
and UO_1300 (O_1300,N_49131,N_48565);
and UO_1301 (O_1301,N_49109,N_48395);
xnor UO_1302 (O_1302,N_49751,N_49975);
nor UO_1303 (O_1303,N_49923,N_49227);
nand UO_1304 (O_1304,N_49794,N_48886);
and UO_1305 (O_1305,N_49306,N_49254);
xnor UO_1306 (O_1306,N_49585,N_48042);
xnor UO_1307 (O_1307,N_49772,N_49708);
nand UO_1308 (O_1308,N_48841,N_48725);
xor UO_1309 (O_1309,N_48213,N_49976);
nor UO_1310 (O_1310,N_48744,N_48799);
and UO_1311 (O_1311,N_48824,N_48021);
nand UO_1312 (O_1312,N_49605,N_49702);
nand UO_1313 (O_1313,N_48117,N_49443);
nor UO_1314 (O_1314,N_48516,N_48727);
nand UO_1315 (O_1315,N_48100,N_49702);
and UO_1316 (O_1316,N_48270,N_48624);
or UO_1317 (O_1317,N_48081,N_48301);
and UO_1318 (O_1318,N_48247,N_49931);
or UO_1319 (O_1319,N_48413,N_49422);
nor UO_1320 (O_1320,N_48371,N_49720);
nand UO_1321 (O_1321,N_49530,N_49774);
nor UO_1322 (O_1322,N_49912,N_49016);
xnor UO_1323 (O_1323,N_49972,N_49844);
xnor UO_1324 (O_1324,N_49252,N_49139);
and UO_1325 (O_1325,N_48058,N_48798);
xor UO_1326 (O_1326,N_48521,N_48082);
nor UO_1327 (O_1327,N_48105,N_49979);
nand UO_1328 (O_1328,N_49773,N_48527);
nand UO_1329 (O_1329,N_49057,N_48987);
xnor UO_1330 (O_1330,N_49661,N_48951);
or UO_1331 (O_1331,N_49723,N_48844);
nand UO_1332 (O_1332,N_49774,N_48922);
xor UO_1333 (O_1333,N_48767,N_48365);
nor UO_1334 (O_1334,N_49910,N_49711);
and UO_1335 (O_1335,N_49934,N_48591);
or UO_1336 (O_1336,N_48124,N_49600);
nor UO_1337 (O_1337,N_48282,N_48449);
and UO_1338 (O_1338,N_48655,N_49859);
nor UO_1339 (O_1339,N_49839,N_49109);
xor UO_1340 (O_1340,N_49001,N_49134);
and UO_1341 (O_1341,N_48069,N_48370);
xnor UO_1342 (O_1342,N_48894,N_49452);
xnor UO_1343 (O_1343,N_49140,N_48066);
and UO_1344 (O_1344,N_49463,N_48255);
xnor UO_1345 (O_1345,N_49709,N_48836);
and UO_1346 (O_1346,N_49856,N_49836);
or UO_1347 (O_1347,N_48813,N_49653);
or UO_1348 (O_1348,N_48435,N_48685);
xor UO_1349 (O_1349,N_48741,N_48814);
and UO_1350 (O_1350,N_49616,N_49828);
and UO_1351 (O_1351,N_49985,N_48748);
and UO_1352 (O_1352,N_48810,N_49521);
and UO_1353 (O_1353,N_49744,N_48680);
nor UO_1354 (O_1354,N_48803,N_48258);
xnor UO_1355 (O_1355,N_49910,N_49068);
or UO_1356 (O_1356,N_49774,N_48583);
nand UO_1357 (O_1357,N_48958,N_48785);
or UO_1358 (O_1358,N_48062,N_49315);
nor UO_1359 (O_1359,N_48429,N_48583);
nand UO_1360 (O_1360,N_48151,N_49532);
or UO_1361 (O_1361,N_49221,N_48851);
and UO_1362 (O_1362,N_48968,N_48729);
and UO_1363 (O_1363,N_49489,N_48891);
or UO_1364 (O_1364,N_48325,N_48710);
nand UO_1365 (O_1365,N_48099,N_48262);
or UO_1366 (O_1366,N_49727,N_49887);
and UO_1367 (O_1367,N_49304,N_49014);
xnor UO_1368 (O_1368,N_49397,N_48122);
and UO_1369 (O_1369,N_48499,N_48323);
or UO_1370 (O_1370,N_48592,N_48960);
xnor UO_1371 (O_1371,N_48183,N_49114);
nand UO_1372 (O_1372,N_48850,N_49409);
or UO_1373 (O_1373,N_49627,N_49725);
nand UO_1374 (O_1374,N_48363,N_48581);
or UO_1375 (O_1375,N_49694,N_48977);
and UO_1376 (O_1376,N_49055,N_48241);
nor UO_1377 (O_1377,N_49628,N_49203);
or UO_1378 (O_1378,N_48050,N_49231);
xnor UO_1379 (O_1379,N_48465,N_48719);
nand UO_1380 (O_1380,N_48168,N_49104);
or UO_1381 (O_1381,N_49404,N_49796);
xnor UO_1382 (O_1382,N_48446,N_49332);
xnor UO_1383 (O_1383,N_48857,N_48409);
xnor UO_1384 (O_1384,N_48362,N_49136);
and UO_1385 (O_1385,N_48564,N_48111);
and UO_1386 (O_1386,N_49299,N_49984);
nor UO_1387 (O_1387,N_49153,N_49536);
or UO_1388 (O_1388,N_49949,N_49833);
nor UO_1389 (O_1389,N_48683,N_48725);
nor UO_1390 (O_1390,N_48178,N_48909);
nand UO_1391 (O_1391,N_48086,N_49615);
xor UO_1392 (O_1392,N_49132,N_49366);
xor UO_1393 (O_1393,N_48504,N_48260);
nand UO_1394 (O_1394,N_48952,N_48425);
and UO_1395 (O_1395,N_49052,N_49456);
nand UO_1396 (O_1396,N_48316,N_48592);
or UO_1397 (O_1397,N_48494,N_49813);
nor UO_1398 (O_1398,N_49415,N_49814);
or UO_1399 (O_1399,N_49874,N_48204);
nor UO_1400 (O_1400,N_48482,N_49368);
nand UO_1401 (O_1401,N_49974,N_49377);
and UO_1402 (O_1402,N_49854,N_48977);
xnor UO_1403 (O_1403,N_48849,N_48349);
nor UO_1404 (O_1404,N_49174,N_48761);
nand UO_1405 (O_1405,N_49210,N_49865);
or UO_1406 (O_1406,N_48423,N_49657);
nor UO_1407 (O_1407,N_48922,N_49727);
xor UO_1408 (O_1408,N_49436,N_49025);
xor UO_1409 (O_1409,N_48118,N_48939);
or UO_1410 (O_1410,N_48826,N_48013);
xor UO_1411 (O_1411,N_48731,N_49886);
and UO_1412 (O_1412,N_49512,N_49414);
nand UO_1413 (O_1413,N_49256,N_48372);
xnor UO_1414 (O_1414,N_49943,N_48496);
or UO_1415 (O_1415,N_48642,N_49636);
or UO_1416 (O_1416,N_48388,N_49371);
nand UO_1417 (O_1417,N_48642,N_48293);
nand UO_1418 (O_1418,N_48239,N_49948);
nor UO_1419 (O_1419,N_49627,N_48535);
and UO_1420 (O_1420,N_49199,N_49001);
or UO_1421 (O_1421,N_48045,N_49168);
and UO_1422 (O_1422,N_49198,N_49534);
xor UO_1423 (O_1423,N_49139,N_49285);
and UO_1424 (O_1424,N_48620,N_49327);
nor UO_1425 (O_1425,N_48884,N_49491);
or UO_1426 (O_1426,N_48843,N_48198);
nand UO_1427 (O_1427,N_48625,N_49352);
nor UO_1428 (O_1428,N_48442,N_49603);
and UO_1429 (O_1429,N_48889,N_49944);
nor UO_1430 (O_1430,N_48593,N_48104);
xor UO_1431 (O_1431,N_48127,N_49526);
nor UO_1432 (O_1432,N_49401,N_49775);
nor UO_1433 (O_1433,N_49077,N_48241);
or UO_1434 (O_1434,N_48579,N_48619);
xor UO_1435 (O_1435,N_48424,N_49254);
nand UO_1436 (O_1436,N_48571,N_48926);
nand UO_1437 (O_1437,N_49604,N_49799);
nor UO_1438 (O_1438,N_49137,N_49092);
xnor UO_1439 (O_1439,N_48625,N_48613);
or UO_1440 (O_1440,N_48664,N_48650);
and UO_1441 (O_1441,N_48262,N_48197);
xnor UO_1442 (O_1442,N_49623,N_48738);
nor UO_1443 (O_1443,N_48543,N_48054);
xor UO_1444 (O_1444,N_48216,N_48198);
xor UO_1445 (O_1445,N_48414,N_49361);
nor UO_1446 (O_1446,N_49708,N_48055);
xor UO_1447 (O_1447,N_49297,N_49945);
nor UO_1448 (O_1448,N_49982,N_49166);
and UO_1449 (O_1449,N_48978,N_48071);
xnor UO_1450 (O_1450,N_48578,N_48085);
nand UO_1451 (O_1451,N_49329,N_48059);
nand UO_1452 (O_1452,N_49616,N_49296);
nand UO_1453 (O_1453,N_48538,N_48745);
xor UO_1454 (O_1454,N_48235,N_49271);
nor UO_1455 (O_1455,N_48580,N_48563);
and UO_1456 (O_1456,N_49384,N_49983);
and UO_1457 (O_1457,N_48403,N_48712);
xor UO_1458 (O_1458,N_48132,N_48691);
nand UO_1459 (O_1459,N_49295,N_49210);
xor UO_1460 (O_1460,N_48097,N_49786);
nand UO_1461 (O_1461,N_49424,N_49920);
nor UO_1462 (O_1462,N_48698,N_48320);
and UO_1463 (O_1463,N_49727,N_48946);
xnor UO_1464 (O_1464,N_48642,N_49564);
nor UO_1465 (O_1465,N_49385,N_48799);
and UO_1466 (O_1466,N_49642,N_49572);
xor UO_1467 (O_1467,N_48138,N_49016);
xor UO_1468 (O_1468,N_48757,N_49181);
xor UO_1469 (O_1469,N_49878,N_48378);
nor UO_1470 (O_1470,N_49538,N_49984);
and UO_1471 (O_1471,N_49641,N_49672);
nand UO_1472 (O_1472,N_49869,N_48855);
nand UO_1473 (O_1473,N_49233,N_48483);
xnor UO_1474 (O_1474,N_49488,N_49875);
nand UO_1475 (O_1475,N_48851,N_48383);
or UO_1476 (O_1476,N_48657,N_48894);
or UO_1477 (O_1477,N_49697,N_49883);
nor UO_1478 (O_1478,N_49394,N_49476);
nand UO_1479 (O_1479,N_48246,N_49348);
xor UO_1480 (O_1480,N_49766,N_48419);
or UO_1481 (O_1481,N_48217,N_49192);
or UO_1482 (O_1482,N_49752,N_49757);
or UO_1483 (O_1483,N_48111,N_48923);
nand UO_1484 (O_1484,N_48361,N_48270);
xnor UO_1485 (O_1485,N_49078,N_48246);
nand UO_1486 (O_1486,N_48148,N_49322);
nand UO_1487 (O_1487,N_49443,N_49033);
xnor UO_1488 (O_1488,N_48288,N_49882);
or UO_1489 (O_1489,N_49945,N_48243);
nand UO_1490 (O_1490,N_48407,N_49808);
or UO_1491 (O_1491,N_48480,N_48605);
and UO_1492 (O_1492,N_48893,N_49869);
and UO_1493 (O_1493,N_48320,N_49634);
nand UO_1494 (O_1494,N_48936,N_49247);
nor UO_1495 (O_1495,N_48470,N_48479);
and UO_1496 (O_1496,N_48201,N_48098);
or UO_1497 (O_1497,N_48790,N_48557);
nor UO_1498 (O_1498,N_49781,N_49526);
xnor UO_1499 (O_1499,N_48646,N_48198);
nand UO_1500 (O_1500,N_48103,N_49952);
nand UO_1501 (O_1501,N_49163,N_49249);
xor UO_1502 (O_1502,N_48561,N_48165);
nor UO_1503 (O_1503,N_48330,N_49038);
nor UO_1504 (O_1504,N_49764,N_49105);
nor UO_1505 (O_1505,N_49377,N_49267);
nand UO_1506 (O_1506,N_49252,N_49576);
xnor UO_1507 (O_1507,N_48522,N_49617);
xor UO_1508 (O_1508,N_48650,N_49547);
nand UO_1509 (O_1509,N_49485,N_49169);
and UO_1510 (O_1510,N_48779,N_48003);
xnor UO_1511 (O_1511,N_49817,N_49530);
xnor UO_1512 (O_1512,N_48423,N_48411);
nand UO_1513 (O_1513,N_49515,N_49916);
nor UO_1514 (O_1514,N_48598,N_49041);
nor UO_1515 (O_1515,N_48978,N_49482);
and UO_1516 (O_1516,N_48423,N_49816);
nor UO_1517 (O_1517,N_49097,N_49491);
and UO_1518 (O_1518,N_48721,N_48290);
xor UO_1519 (O_1519,N_49255,N_48127);
and UO_1520 (O_1520,N_49058,N_49647);
nor UO_1521 (O_1521,N_49345,N_49258);
or UO_1522 (O_1522,N_48356,N_49142);
and UO_1523 (O_1523,N_49210,N_49664);
nand UO_1524 (O_1524,N_49753,N_49667);
and UO_1525 (O_1525,N_48886,N_48476);
nor UO_1526 (O_1526,N_48954,N_48889);
and UO_1527 (O_1527,N_48643,N_49998);
nand UO_1528 (O_1528,N_49508,N_49957);
nor UO_1529 (O_1529,N_48687,N_48502);
or UO_1530 (O_1530,N_48133,N_48294);
nor UO_1531 (O_1531,N_48683,N_48760);
or UO_1532 (O_1532,N_49192,N_49401);
xnor UO_1533 (O_1533,N_48195,N_48559);
nor UO_1534 (O_1534,N_49066,N_49945);
nand UO_1535 (O_1535,N_49406,N_49137);
or UO_1536 (O_1536,N_49931,N_49244);
or UO_1537 (O_1537,N_49168,N_48991);
nor UO_1538 (O_1538,N_49645,N_49711);
and UO_1539 (O_1539,N_49145,N_48103);
nand UO_1540 (O_1540,N_49480,N_48876);
xnor UO_1541 (O_1541,N_48841,N_49612);
xnor UO_1542 (O_1542,N_49824,N_49268);
nand UO_1543 (O_1543,N_48659,N_49952);
nor UO_1544 (O_1544,N_48316,N_49233);
or UO_1545 (O_1545,N_48140,N_49627);
and UO_1546 (O_1546,N_49243,N_48819);
or UO_1547 (O_1547,N_49522,N_49657);
and UO_1548 (O_1548,N_49523,N_49568);
nand UO_1549 (O_1549,N_49657,N_49025);
nand UO_1550 (O_1550,N_49151,N_49835);
or UO_1551 (O_1551,N_48573,N_49362);
nor UO_1552 (O_1552,N_49486,N_49880);
xor UO_1553 (O_1553,N_48698,N_49993);
or UO_1554 (O_1554,N_49363,N_49260);
or UO_1555 (O_1555,N_49839,N_49193);
and UO_1556 (O_1556,N_48832,N_49375);
xnor UO_1557 (O_1557,N_48485,N_48674);
and UO_1558 (O_1558,N_49883,N_49560);
and UO_1559 (O_1559,N_48910,N_49539);
and UO_1560 (O_1560,N_49479,N_49889);
nand UO_1561 (O_1561,N_48441,N_48382);
and UO_1562 (O_1562,N_49636,N_49695);
nand UO_1563 (O_1563,N_48578,N_48433);
nand UO_1564 (O_1564,N_49864,N_49326);
nor UO_1565 (O_1565,N_49818,N_49436);
xor UO_1566 (O_1566,N_49277,N_49513);
nor UO_1567 (O_1567,N_49386,N_48755);
nor UO_1568 (O_1568,N_48196,N_48953);
and UO_1569 (O_1569,N_49369,N_49259);
nor UO_1570 (O_1570,N_48594,N_49389);
xnor UO_1571 (O_1571,N_49399,N_49952);
xnor UO_1572 (O_1572,N_48927,N_48288);
or UO_1573 (O_1573,N_49738,N_48746);
and UO_1574 (O_1574,N_49861,N_49099);
nand UO_1575 (O_1575,N_49959,N_48452);
xnor UO_1576 (O_1576,N_48549,N_48962);
and UO_1577 (O_1577,N_48016,N_49955);
nand UO_1578 (O_1578,N_48074,N_48162);
nor UO_1579 (O_1579,N_49571,N_49801);
or UO_1580 (O_1580,N_49292,N_48721);
xor UO_1581 (O_1581,N_48569,N_49531);
or UO_1582 (O_1582,N_49383,N_48559);
or UO_1583 (O_1583,N_48213,N_48550);
or UO_1584 (O_1584,N_49647,N_49110);
or UO_1585 (O_1585,N_49656,N_49870);
or UO_1586 (O_1586,N_48449,N_49388);
nor UO_1587 (O_1587,N_49159,N_49500);
nor UO_1588 (O_1588,N_48463,N_48512);
xnor UO_1589 (O_1589,N_48752,N_48646);
or UO_1590 (O_1590,N_48927,N_49309);
nand UO_1591 (O_1591,N_48459,N_49947);
xor UO_1592 (O_1592,N_49381,N_49120);
nor UO_1593 (O_1593,N_48983,N_48504);
xor UO_1594 (O_1594,N_49806,N_49396);
and UO_1595 (O_1595,N_49933,N_49226);
nor UO_1596 (O_1596,N_49453,N_48077);
or UO_1597 (O_1597,N_48013,N_49600);
xnor UO_1598 (O_1598,N_48591,N_48557);
or UO_1599 (O_1599,N_48712,N_48677);
or UO_1600 (O_1600,N_48446,N_48442);
and UO_1601 (O_1601,N_49726,N_49254);
xnor UO_1602 (O_1602,N_48127,N_48355);
nand UO_1603 (O_1603,N_48128,N_48614);
nor UO_1604 (O_1604,N_48579,N_48736);
nor UO_1605 (O_1605,N_49144,N_49715);
nand UO_1606 (O_1606,N_48550,N_49403);
xor UO_1607 (O_1607,N_49394,N_49583);
nand UO_1608 (O_1608,N_48832,N_48253);
nand UO_1609 (O_1609,N_48159,N_48479);
nor UO_1610 (O_1610,N_48339,N_48442);
nor UO_1611 (O_1611,N_49370,N_49962);
or UO_1612 (O_1612,N_49033,N_49746);
and UO_1613 (O_1613,N_48911,N_49808);
nor UO_1614 (O_1614,N_48943,N_49621);
xnor UO_1615 (O_1615,N_49274,N_48059);
nand UO_1616 (O_1616,N_49209,N_49002);
and UO_1617 (O_1617,N_49611,N_49069);
nor UO_1618 (O_1618,N_49827,N_49046);
or UO_1619 (O_1619,N_48442,N_48589);
nor UO_1620 (O_1620,N_49402,N_49270);
or UO_1621 (O_1621,N_49377,N_48499);
nand UO_1622 (O_1622,N_48926,N_49465);
or UO_1623 (O_1623,N_49400,N_49364);
xor UO_1624 (O_1624,N_49047,N_48766);
and UO_1625 (O_1625,N_49300,N_48810);
xor UO_1626 (O_1626,N_48427,N_49652);
nor UO_1627 (O_1627,N_48860,N_49705);
nand UO_1628 (O_1628,N_48975,N_49931);
and UO_1629 (O_1629,N_48842,N_48812);
nand UO_1630 (O_1630,N_49966,N_49248);
or UO_1631 (O_1631,N_49812,N_48709);
xor UO_1632 (O_1632,N_49667,N_48582);
nor UO_1633 (O_1633,N_48960,N_48585);
xnor UO_1634 (O_1634,N_48406,N_49812);
and UO_1635 (O_1635,N_49385,N_49439);
nand UO_1636 (O_1636,N_49410,N_49622);
xor UO_1637 (O_1637,N_48694,N_48112);
or UO_1638 (O_1638,N_48786,N_48771);
nand UO_1639 (O_1639,N_49038,N_48305);
nor UO_1640 (O_1640,N_49378,N_49944);
and UO_1641 (O_1641,N_48712,N_48042);
xor UO_1642 (O_1642,N_49651,N_48013);
nand UO_1643 (O_1643,N_48558,N_49790);
or UO_1644 (O_1644,N_49085,N_48329);
xor UO_1645 (O_1645,N_48171,N_48343);
nand UO_1646 (O_1646,N_48433,N_48894);
nand UO_1647 (O_1647,N_49909,N_49351);
and UO_1648 (O_1648,N_49555,N_48080);
or UO_1649 (O_1649,N_48751,N_49035);
xor UO_1650 (O_1650,N_48290,N_49988);
or UO_1651 (O_1651,N_48779,N_48916);
or UO_1652 (O_1652,N_48839,N_49909);
nor UO_1653 (O_1653,N_48665,N_48954);
and UO_1654 (O_1654,N_48000,N_49272);
nor UO_1655 (O_1655,N_48058,N_48105);
nor UO_1656 (O_1656,N_48792,N_49103);
nand UO_1657 (O_1657,N_49654,N_48295);
nor UO_1658 (O_1658,N_49439,N_49332);
or UO_1659 (O_1659,N_49899,N_49060);
xnor UO_1660 (O_1660,N_48717,N_48147);
and UO_1661 (O_1661,N_49506,N_49058);
or UO_1662 (O_1662,N_48689,N_49787);
nand UO_1663 (O_1663,N_48007,N_49328);
and UO_1664 (O_1664,N_49887,N_49886);
xnor UO_1665 (O_1665,N_48120,N_49835);
nand UO_1666 (O_1666,N_49539,N_49748);
nand UO_1667 (O_1667,N_49999,N_49443);
or UO_1668 (O_1668,N_49511,N_49950);
and UO_1669 (O_1669,N_48309,N_49314);
xor UO_1670 (O_1670,N_49148,N_48354);
nand UO_1671 (O_1671,N_48205,N_49218);
or UO_1672 (O_1672,N_48396,N_48837);
nor UO_1673 (O_1673,N_49541,N_48392);
and UO_1674 (O_1674,N_49377,N_49427);
xor UO_1675 (O_1675,N_49017,N_48547);
and UO_1676 (O_1676,N_48601,N_49321);
xor UO_1677 (O_1677,N_48566,N_48692);
nor UO_1678 (O_1678,N_48979,N_48364);
xnor UO_1679 (O_1679,N_48477,N_49361);
nor UO_1680 (O_1680,N_49235,N_48802);
nor UO_1681 (O_1681,N_49956,N_49139);
and UO_1682 (O_1682,N_48865,N_48608);
nand UO_1683 (O_1683,N_48920,N_48403);
nand UO_1684 (O_1684,N_49182,N_48723);
or UO_1685 (O_1685,N_48151,N_48766);
nand UO_1686 (O_1686,N_49352,N_48077);
xor UO_1687 (O_1687,N_48820,N_49850);
and UO_1688 (O_1688,N_49847,N_49918);
nand UO_1689 (O_1689,N_49579,N_48976);
and UO_1690 (O_1690,N_48578,N_48189);
or UO_1691 (O_1691,N_49332,N_49546);
xnor UO_1692 (O_1692,N_48897,N_48190);
xor UO_1693 (O_1693,N_49792,N_49944);
nand UO_1694 (O_1694,N_48078,N_49000);
nor UO_1695 (O_1695,N_48719,N_48349);
nor UO_1696 (O_1696,N_49252,N_49962);
xnor UO_1697 (O_1697,N_48595,N_49909);
or UO_1698 (O_1698,N_49492,N_49005);
nand UO_1699 (O_1699,N_48297,N_49374);
or UO_1700 (O_1700,N_48489,N_48519);
and UO_1701 (O_1701,N_48501,N_49199);
nand UO_1702 (O_1702,N_48885,N_48953);
nor UO_1703 (O_1703,N_48733,N_49185);
nor UO_1704 (O_1704,N_48793,N_48451);
nor UO_1705 (O_1705,N_48799,N_48841);
nor UO_1706 (O_1706,N_48983,N_49582);
or UO_1707 (O_1707,N_48710,N_48242);
nand UO_1708 (O_1708,N_48945,N_48537);
nand UO_1709 (O_1709,N_48126,N_48628);
and UO_1710 (O_1710,N_49085,N_49663);
xnor UO_1711 (O_1711,N_49134,N_49007);
xnor UO_1712 (O_1712,N_49566,N_48106);
nor UO_1713 (O_1713,N_49434,N_49859);
nand UO_1714 (O_1714,N_48651,N_49695);
nor UO_1715 (O_1715,N_48265,N_48391);
and UO_1716 (O_1716,N_48377,N_48456);
and UO_1717 (O_1717,N_49557,N_49816);
nand UO_1718 (O_1718,N_49268,N_48127);
and UO_1719 (O_1719,N_48571,N_48895);
xnor UO_1720 (O_1720,N_48326,N_48718);
nand UO_1721 (O_1721,N_48374,N_48144);
or UO_1722 (O_1722,N_48023,N_48643);
nand UO_1723 (O_1723,N_48206,N_49122);
nand UO_1724 (O_1724,N_49911,N_48448);
nand UO_1725 (O_1725,N_48239,N_49385);
nand UO_1726 (O_1726,N_49964,N_48714);
nor UO_1727 (O_1727,N_48334,N_49861);
nor UO_1728 (O_1728,N_49904,N_49280);
and UO_1729 (O_1729,N_48178,N_48792);
nor UO_1730 (O_1730,N_48242,N_49823);
and UO_1731 (O_1731,N_48114,N_49181);
xor UO_1732 (O_1732,N_49596,N_48695);
or UO_1733 (O_1733,N_49149,N_48736);
nand UO_1734 (O_1734,N_48843,N_48458);
nand UO_1735 (O_1735,N_49262,N_49988);
and UO_1736 (O_1736,N_49085,N_48360);
nor UO_1737 (O_1737,N_48542,N_49443);
xor UO_1738 (O_1738,N_49651,N_49211);
xor UO_1739 (O_1739,N_49336,N_48670);
and UO_1740 (O_1740,N_48983,N_49666);
or UO_1741 (O_1741,N_49637,N_48543);
or UO_1742 (O_1742,N_49326,N_49417);
xor UO_1743 (O_1743,N_48805,N_48586);
nor UO_1744 (O_1744,N_48793,N_49909);
and UO_1745 (O_1745,N_48835,N_49811);
nand UO_1746 (O_1746,N_48429,N_48398);
xor UO_1747 (O_1747,N_48222,N_49398);
or UO_1748 (O_1748,N_49719,N_48455);
xor UO_1749 (O_1749,N_48823,N_48211);
nand UO_1750 (O_1750,N_49773,N_49050);
nand UO_1751 (O_1751,N_49050,N_48998);
and UO_1752 (O_1752,N_49356,N_49134);
nand UO_1753 (O_1753,N_49032,N_49647);
xnor UO_1754 (O_1754,N_49540,N_49897);
nand UO_1755 (O_1755,N_48518,N_49907);
and UO_1756 (O_1756,N_49542,N_49638);
nand UO_1757 (O_1757,N_48376,N_49247);
nand UO_1758 (O_1758,N_49181,N_49373);
or UO_1759 (O_1759,N_48925,N_48635);
nor UO_1760 (O_1760,N_49843,N_48544);
xor UO_1761 (O_1761,N_49469,N_49468);
nand UO_1762 (O_1762,N_49892,N_49990);
or UO_1763 (O_1763,N_48697,N_49759);
nor UO_1764 (O_1764,N_49650,N_49781);
nand UO_1765 (O_1765,N_49268,N_49600);
and UO_1766 (O_1766,N_49453,N_49548);
xor UO_1767 (O_1767,N_49492,N_49403);
nand UO_1768 (O_1768,N_48903,N_48907);
or UO_1769 (O_1769,N_48792,N_49773);
nand UO_1770 (O_1770,N_48999,N_48833);
or UO_1771 (O_1771,N_48855,N_48191);
xnor UO_1772 (O_1772,N_49337,N_48631);
nand UO_1773 (O_1773,N_48938,N_48844);
nor UO_1774 (O_1774,N_49055,N_49083);
nand UO_1775 (O_1775,N_48118,N_48297);
nor UO_1776 (O_1776,N_48884,N_48303);
or UO_1777 (O_1777,N_48208,N_48834);
nand UO_1778 (O_1778,N_48311,N_48038);
and UO_1779 (O_1779,N_49719,N_49579);
nor UO_1780 (O_1780,N_49228,N_49619);
xor UO_1781 (O_1781,N_48397,N_49193);
xnor UO_1782 (O_1782,N_48589,N_49812);
xnor UO_1783 (O_1783,N_48672,N_49889);
xnor UO_1784 (O_1784,N_49694,N_49865);
xor UO_1785 (O_1785,N_48603,N_49015);
xnor UO_1786 (O_1786,N_49254,N_49672);
xor UO_1787 (O_1787,N_48259,N_49264);
xnor UO_1788 (O_1788,N_48538,N_48277);
nor UO_1789 (O_1789,N_49361,N_49724);
or UO_1790 (O_1790,N_49120,N_48341);
nand UO_1791 (O_1791,N_49916,N_48558);
nor UO_1792 (O_1792,N_49954,N_48304);
and UO_1793 (O_1793,N_48040,N_48927);
xnor UO_1794 (O_1794,N_48400,N_48719);
xor UO_1795 (O_1795,N_48253,N_49266);
and UO_1796 (O_1796,N_49769,N_49532);
and UO_1797 (O_1797,N_48111,N_49617);
nor UO_1798 (O_1798,N_49642,N_48572);
nand UO_1799 (O_1799,N_48985,N_49680);
nor UO_1800 (O_1800,N_48105,N_49188);
or UO_1801 (O_1801,N_48554,N_49162);
nand UO_1802 (O_1802,N_49567,N_49258);
and UO_1803 (O_1803,N_48283,N_48687);
and UO_1804 (O_1804,N_48385,N_49132);
xor UO_1805 (O_1805,N_49954,N_49421);
or UO_1806 (O_1806,N_49321,N_49496);
nand UO_1807 (O_1807,N_49982,N_48805);
nor UO_1808 (O_1808,N_49048,N_49181);
xnor UO_1809 (O_1809,N_48585,N_49838);
xnor UO_1810 (O_1810,N_48845,N_48450);
or UO_1811 (O_1811,N_48272,N_49314);
or UO_1812 (O_1812,N_48343,N_49588);
nor UO_1813 (O_1813,N_49040,N_49425);
and UO_1814 (O_1814,N_49563,N_48663);
xnor UO_1815 (O_1815,N_49452,N_48793);
xnor UO_1816 (O_1816,N_49691,N_48541);
or UO_1817 (O_1817,N_49355,N_48794);
nand UO_1818 (O_1818,N_49536,N_49004);
nor UO_1819 (O_1819,N_48114,N_49879);
xnor UO_1820 (O_1820,N_48225,N_48665);
and UO_1821 (O_1821,N_49170,N_49157);
nand UO_1822 (O_1822,N_49638,N_49710);
and UO_1823 (O_1823,N_48773,N_49136);
nor UO_1824 (O_1824,N_49782,N_48263);
xnor UO_1825 (O_1825,N_49389,N_48444);
or UO_1826 (O_1826,N_49644,N_49498);
or UO_1827 (O_1827,N_48668,N_49293);
or UO_1828 (O_1828,N_49979,N_49260);
xnor UO_1829 (O_1829,N_48834,N_48154);
nand UO_1830 (O_1830,N_49156,N_49522);
xnor UO_1831 (O_1831,N_48974,N_49104);
and UO_1832 (O_1832,N_48683,N_49680);
nand UO_1833 (O_1833,N_48809,N_48388);
and UO_1834 (O_1834,N_48912,N_48210);
xor UO_1835 (O_1835,N_48932,N_49657);
and UO_1836 (O_1836,N_48618,N_49406);
and UO_1837 (O_1837,N_49023,N_48580);
nor UO_1838 (O_1838,N_49420,N_49307);
xor UO_1839 (O_1839,N_48697,N_49420);
and UO_1840 (O_1840,N_49150,N_49383);
nor UO_1841 (O_1841,N_48302,N_49849);
and UO_1842 (O_1842,N_48135,N_48398);
or UO_1843 (O_1843,N_49958,N_49429);
xor UO_1844 (O_1844,N_49549,N_48879);
and UO_1845 (O_1845,N_48343,N_49338);
nand UO_1846 (O_1846,N_49900,N_49796);
or UO_1847 (O_1847,N_49164,N_48790);
or UO_1848 (O_1848,N_48713,N_48900);
and UO_1849 (O_1849,N_48040,N_48511);
xor UO_1850 (O_1850,N_49240,N_49613);
xor UO_1851 (O_1851,N_49498,N_49589);
or UO_1852 (O_1852,N_49060,N_49399);
and UO_1853 (O_1853,N_48969,N_49771);
xor UO_1854 (O_1854,N_49333,N_49992);
nand UO_1855 (O_1855,N_49250,N_48409);
nor UO_1856 (O_1856,N_49312,N_48735);
and UO_1857 (O_1857,N_48293,N_49658);
nor UO_1858 (O_1858,N_48865,N_48837);
nor UO_1859 (O_1859,N_49965,N_48217);
xor UO_1860 (O_1860,N_49326,N_48718);
and UO_1861 (O_1861,N_48872,N_48234);
or UO_1862 (O_1862,N_49828,N_48809);
nand UO_1863 (O_1863,N_49685,N_48248);
and UO_1864 (O_1864,N_48642,N_48583);
nor UO_1865 (O_1865,N_49076,N_49595);
or UO_1866 (O_1866,N_49061,N_48074);
or UO_1867 (O_1867,N_49306,N_49998);
nand UO_1868 (O_1868,N_48573,N_49414);
nor UO_1869 (O_1869,N_48111,N_48250);
or UO_1870 (O_1870,N_48074,N_49077);
or UO_1871 (O_1871,N_48239,N_48684);
and UO_1872 (O_1872,N_48881,N_49985);
xor UO_1873 (O_1873,N_49214,N_49020);
nor UO_1874 (O_1874,N_48450,N_49140);
or UO_1875 (O_1875,N_49066,N_49781);
and UO_1876 (O_1876,N_49331,N_49236);
or UO_1877 (O_1877,N_49373,N_49705);
and UO_1878 (O_1878,N_48002,N_49410);
nor UO_1879 (O_1879,N_48519,N_48323);
nor UO_1880 (O_1880,N_48853,N_48046);
or UO_1881 (O_1881,N_48303,N_49556);
nor UO_1882 (O_1882,N_49276,N_49189);
nand UO_1883 (O_1883,N_49230,N_48746);
xor UO_1884 (O_1884,N_49140,N_49318);
or UO_1885 (O_1885,N_49944,N_48183);
xnor UO_1886 (O_1886,N_49544,N_49530);
xor UO_1887 (O_1887,N_48993,N_48251);
and UO_1888 (O_1888,N_49488,N_48136);
xor UO_1889 (O_1889,N_48623,N_49473);
nand UO_1890 (O_1890,N_48060,N_48463);
nand UO_1891 (O_1891,N_49760,N_49808);
or UO_1892 (O_1892,N_48402,N_49249);
nor UO_1893 (O_1893,N_49553,N_49111);
nor UO_1894 (O_1894,N_48570,N_48253);
nand UO_1895 (O_1895,N_49369,N_49171);
nand UO_1896 (O_1896,N_48036,N_48732);
xor UO_1897 (O_1897,N_49503,N_48424);
or UO_1898 (O_1898,N_49940,N_49879);
nor UO_1899 (O_1899,N_48436,N_48460);
or UO_1900 (O_1900,N_49285,N_48255);
and UO_1901 (O_1901,N_49095,N_48560);
and UO_1902 (O_1902,N_49972,N_48531);
nand UO_1903 (O_1903,N_49947,N_48470);
or UO_1904 (O_1904,N_48651,N_49074);
xnor UO_1905 (O_1905,N_49221,N_48777);
xnor UO_1906 (O_1906,N_48739,N_48486);
or UO_1907 (O_1907,N_49062,N_48241);
nand UO_1908 (O_1908,N_48041,N_48254);
or UO_1909 (O_1909,N_48328,N_49531);
nand UO_1910 (O_1910,N_48625,N_49648);
xnor UO_1911 (O_1911,N_48718,N_48325);
xnor UO_1912 (O_1912,N_48459,N_48427);
and UO_1913 (O_1913,N_48923,N_49587);
or UO_1914 (O_1914,N_48380,N_49823);
nand UO_1915 (O_1915,N_48240,N_48846);
or UO_1916 (O_1916,N_49247,N_48983);
and UO_1917 (O_1917,N_48664,N_48559);
nor UO_1918 (O_1918,N_49251,N_48031);
nor UO_1919 (O_1919,N_48070,N_48233);
or UO_1920 (O_1920,N_48164,N_48239);
nor UO_1921 (O_1921,N_48123,N_49239);
nor UO_1922 (O_1922,N_48924,N_49839);
or UO_1923 (O_1923,N_49668,N_49681);
xnor UO_1924 (O_1924,N_49385,N_49226);
or UO_1925 (O_1925,N_48691,N_48797);
xor UO_1926 (O_1926,N_49247,N_48103);
xnor UO_1927 (O_1927,N_48054,N_49824);
or UO_1928 (O_1928,N_49103,N_48706);
nand UO_1929 (O_1929,N_49857,N_48062);
nand UO_1930 (O_1930,N_48512,N_49771);
and UO_1931 (O_1931,N_48205,N_48375);
or UO_1932 (O_1932,N_49407,N_48713);
xnor UO_1933 (O_1933,N_48655,N_48915);
or UO_1934 (O_1934,N_49405,N_48674);
nor UO_1935 (O_1935,N_49722,N_49787);
or UO_1936 (O_1936,N_48645,N_48824);
xor UO_1937 (O_1937,N_49275,N_48355);
and UO_1938 (O_1938,N_49299,N_49001);
or UO_1939 (O_1939,N_49773,N_48305);
or UO_1940 (O_1940,N_49255,N_48475);
and UO_1941 (O_1941,N_48930,N_48340);
or UO_1942 (O_1942,N_48764,N_48878);
nand UO_1943 (O_1943,N_48443,N_48217);
nand UO_1944 (O_1944,N_48554,N_49051);
nand UO_1945 (O_1945,N_49101,N_49540);
and UO_1946 (O_1946,N_49297,N_48545);
xnor UO_1947 (O_1947,N_48636,N_49192);
nor UO_1948 (O_1948,N_48777,N_48660);
nor UO_1949 (O_1949,N_48306,N_49211);
nand UO_1950 (O_1950,N_49610,N_48249);
nand UO_1951 (O_1951,N_48238,N_49019);
or UO_1952 (O_1952,N_49083,N_48474);
and UO_1953 (O_1953,N_48724,N_49662);
or UO_1954 (O_1954,N_49728,N_49979);
xor UO_1955 (O_1955,N_49969,N_49809);
and UO_1956 (O_1956,N_48167,N_49319);
and UO_1957 (O_1957,N_49603,N_48421);
nand UO_1958 (O_1958,N_49300,N_49928);
nor UO_1959 (O_1959,N_48670,N_49128);
xor UO_1960 (O_1960,N_48921,N_49251);
and UO_1961 (O_1961,N_49169,N_48005);
xnor UO_1962 (O_1962,N_49978,N_48469);
xor UO_1963 (O_1963,N_49053,N_49041);
and UO_1964 (O_1964,N_48555,N_49000);
xor UO_1965 (O_1965,N_49053,N_49134);
xor UO_1966 (O_1966,N_49182,N_49037);
and UO_1967 (O_1967,N_49503,N_49420);
nand UO_1968 (O_1968,N_49272,N_49717);
nand UO_1969 (O_1969,N_49795,N_48108);
and UO_1970 (O_1970,N_48955,N_49553);
nor UO_1971 (O_1971,N_49013,N_48901);
and UO_1972 (O_1972,N_48159,N_48266);
or UO_1973 (O_1973,N_48441,N_49919);
and UO_1974 (O_1974,N_48446,N_49952);
nor UO_1975 (O_1975,N_49443,N_48658);
nor UO_1976 (O_1976,N_48649,N_49876);
or UO_1977 (O_1977,N_48218,N_49982);
or UO_1978 (O_1978,N_49288,N_49503);
nor UO_1979 (O_1979,N_48088,N_48409);
or UO_1980 (O_1980,N_48932,N_49522);
xnor UO_1981 (O_1981,N_49106,N_48059);
nor UO_1982 (O_1982,N_48793,N_48993);
xor UO_1983 (O_1983,N_49977,N_49608);
xor UO_1984 (O_1984,N_48189,N_48337);
nand UO_1985 (O_1985,N_48495,N_49898);
and UO_1986 (O_1986,N_49865,N_49556);
nand UO_1987 (O_1987,N_49804,N_49629);
nor UO_1988 (O_1988,N_49967,N_48002);
or UO_1989 (O_1989,N_49268,N_49538);
or UO_1990 (O_1990,N_49245,N_49005);
or UO_1991 (O_1991,N_48400,N_48464);
and UO_1992 (O_1992,N_48617,N_48933);
or UO_1993 (O_1993,N_49653,N_49758);
or UO_1994 (O_1994,N_49983,N_49636);
and UO_1995 (O_1995,N_49705,N_49064);
and UO_1996 (O_1996,N_48959,N_48619);
xnor UO_1997 (O_1997,N_49597,N_49058);
and UO_1998 (O_1998,N_49863,N_48508);
xor UO_1999 (O_1999,N_49506,N_49148);
nand UO_2000 (O_2000,N_49403,N_48227);
nor UO_2001 (O_2001,N_49347,N_49843);
nor UO_2002 (O_2002,N_48775,N_49341);
nor UO_2003 (O_2003,N_49709,N_49505);
or UO_2004 (O_2004,N_49217,N_49707);
xnor UO_2005 (O_2005,N_49110,N_48831);
and UO_2006 (O_2006,N_49207,N_48806);
and UO_2007 (O_2007,N_49209,N_48284);
nor UO_2008 (O_2008,N_48890,N_49638);
xor UO_2009 (O_2009,N_48546,N_49254);
nor UO_2010 (O_2010,N_48382,N_48749);
xor UO_2011 (O_2011,N_49184,N_48712);
nor UO_2012 (O_2012,N_49988,N_48633);
xor UO_2013 (O_2013,N_49739,N_48815);
and UO_2014 (O_2014,N_48280,N_49311);
and UO_2015 (O_2015,N_48880,N_49912);
nand UO_2016 (O_2016,N_49539,N_48879);
or UO_2017 (O_2017,N_48489,N_48708);
and UO_2018 (O_2018,N_49629,N_48456);
nand UO_2019 (O_2019,N_49396,N_49888);
nand UO_2020 (O_2020,N_49615,N_48557);
xor UO_2021 (O_2021,N_48272,N_48752);
xor UO_2022 (O_2022,N_48649,N_48984);
and UO_2023 (O_2023,N_49625,N_49283);
nand UO_2024 (O_2024,N_48891,N_48396);
and UO_2025 (O_2025,N_48339,N_48592);
xor UO_2026 (O_2026,N_48622,N_49539);
or UO_2027 (O_2027,N_48834,N_48062);
xnor UO_2028 (O_2028,N_48958,N_48708);
nor UO_2029 (O_2029,N_49943,N_48265);
or UO_2030 (O_2030,N_48223,N_49708);
xnor UO_2031 (O_2031,N_48848,N_49037);
nand UO_2032 (O_2032,N_48477,N_48112);
nand UO_2033 (O_2033,N_49801,N_49019);
xor UO_2034 (O_2034,N_49494,N_49215);
and UO_2035 (O_2035,N_48471,N_48776);
nor UO_2036 (O_2036,N_49036,N_48395);
nor UO_2037 (O_2037,N_49678,N_48831);
nor UO_2038 (O_2038,N_49646,N_48575);
or UO_2039 (O_2039,N_48168,N_49015);
nor UO_2040 (O_2040,N_49820,N_48044);
nor UO_2041 (O_2041,N_49931,N_49188);
or UO_2042 (O_2042,N_49417,N_48966);
nand UO_2043 (O_2043,N_48945,N_48991);
or UO_2044 (O_2044,N_48037,N_49629);
or UO_2045 (O_2045,N_49140,N_48222);
nor UO_2046 (O_2046,N_49350,N_49120);
xor UO_2047 (O_2047,N_49159,N_49673);
nand UO_2048 (O_2048,N_48369,N_49678);
nand UO_2049 (O_2049,N_49032,N_48934);
xor UO_2050 (O_2050,N_48711,N_48272);
and UO_2051 (O_2051,N_48450,N_49365);
nand UO_2052 (O_2052,N_48888,N_49604);
nor UO_2053 (O_2053,N_49642,N_48915);
nand UO_2054 (O_2054,N_48056,N_49558);
xor UO_2055 (O_2055,N_49245,N_48568);
or UO_2056 (O_2056,N_48573,N_48569);
nor UO_2057 (O_2057,N_48056,N_49932);
and UO_2058 (O_2058,N_49352,N_48663);
or UO_2059 (O_2059,N_48904,N_48295);
nand UO_2060 (O_2060,N_49978,N_49602);
or UO_2061 (O_2061,N_49570,N_49055);
and UO_2062 (O_2062,N_49097,N_49041);
xor UO_2063 (O_2063,N_49891,N_49975);
xnor UO_2064 (O_2064,N_49328,N_48965);
xnor UO_2065 (O_2065,N_49885,N_49117);
xor UO_2066 (O_2066,N_48468,N_48962);
nand UO_2067 (O_2067,N_48246,N_48689);
nand UO_2068 (O_2068,N_48338,N_49875);
and UO_2069 (O_2069,N_48457,N_49691);
nor UO_2070 (O_2070,N_48223,N_49047);
nor UO_2071 (O_2071,N_49888,N_48364);
xnor UO_2072 (O_2072,N_48575,N_48770);
or UO_2073 (O_2073,N_48815,N_48698);
or UO_2074 (O_2074,N_49225,N_48581);
or UO_2075 (O_2075,N_49608,N_49605);
and UO_2076 (O_2076,N_49625,N_48765);
nor UO_2077 (O_2077,N_49853,N_48895);
nand UO_2078 (O_2078,N_49394,N_48622);
xnor UO_2079 (O_2079,N_49001,N_49846);
xor UO_2080 (O_2080,N_48108,N_48941);
nor UO_2081 (O_2081,N_48738,N_48398);
or UO_2082 (O_2082,N_48157,N_49407);
xor UO_2083 (O_2083,N_49372,N_49374);
nand UO_2084 (O_2084,N_49708,N_48122);
and UO_2085 (O_2085,N_49690,N_49622);
nand UO_2086 (O_2086,N_48233,N_48412);
or UO_2087 (O_2087,N_49990,N_49924);
nand UO_2088 (O_2088,N_49478,N_48997);
nand UO_2089 (O_2089,N_48741,N_48768);
and UO_2090 (O_2090,N_48483,N_48754);
nand UO_2091 (O_2091,N_48105,N_48824);
nand UO_2092 (O_2092,N_48789,N_48558);
xnor UO_2093 (O_2093,N_49900,N_49245);
xor UO_2094 (O_2094,N_48155,N_49452);
or UO_2095 (O_2095,N_48378,N_49355);
or UO_2096 (O_2096,N_48414,N_49252);
xnor UO_2097 (O_2097,N_49063,N_49826);
nand UO_2098 (O_2098,N_48750,N_48821);
xnor UO_2099 (O_2099,N_48576,N_49322);
or UO_2100 (O_2100,N_48383,N_49166);
xnor UO_2101 (O_2101,N_48934,N_49056);
xor UO_2102 (O_2102,N_48757,N_49956);
xnor UO_2103 (O_2103,N_49063,N_49448);
and UO_2104 (O_2104,N_49444,N_49678);
xnor UO_2105 (O_2105,N_48225,N_49160);
and UO_2106 (O_2106,N_49322,N_48785);
and UO_2107 (O_2107,N_48858,N_48053);
xor UO_2108 (O_2108,N_48184,N_49483);
nand UO_2109 (O_2109,N_49625,N_48141);
nand UO_2110 (O_2110,N_49496,N_49182);
nand UO_2111 (O_2111,N_49122,N_49069);
nand UO_2112 (O_2112,N_49969,N_49633);
nand UO_2113 (O_2113,N_48924,N_48262);
nor UO_2114 (O_2114,N_49692,N_49182);
nand UO_2115 (O_2115,N_48534,N_48743);
or UO_2116 (O_2116,N_49289,N_49231);
and UO_2117 (O_2117,N_49428,N_49025);
or UO_2118 (O_2118,N_48616,N_49696);
nand UO_2119 (O_2119,N_49966,N_48579);
nand UO_2120 (O_2120,N_49139,N_48888);
and UO_2121 (O_2121,N_48799,N_48681);
nand UO_2122 (O_2122,N_49675,N_48809);
and UO_2123 (O_2123,N_48183,N_48276);
nand UO_2124 (O_2124,N_49136,N_49758);
nand UO_2125 (O_2125,N_48958,N_48860);
and UO_2126 (O_2126,N_49416,N_49619);
nor UO_2127 (O_2127,N_49088,N_49212);
nand UO_2128 (O_2128,N_49106,N_49425);
nor UO_2129 (O_2129,N_48317,N_48958);
or UO_2130 (O_2130,N_48282,N_49184);
nor UO_2131 (O_2131,N_48619,N_49476);
or UO_2132 (O_2132,N_49552,N_48260);
xnor UO_2133 (O_2133,N_49560,N_48696);
nor UO_2134 (O_2134,N_49587,N_49809);
nor UO_2135 (O_2135,N_48142,N_48444);
nand UO_2136 (O_2136,N_49069,N_49343);
and UO_2137 (O_2137,N_49670,N_49007);
nor UO_2138 (O_2138,N_48242,N_48748);
or UO_2139 (O_2139,N_49919,N_49926);
xnor UO_2140 (O_2140,N_48760,N_49212);
nand UO_2141 (O_2141,N_48882,N_48995);
or UO_2142 (O_2142,N_49142,N_49848);
nor UO_2143 (O_2143,N_49022,N_48699);
nand UO_2144 (O_2144,N_49655,N_49104);
xnor UO_2145 (O_2145,N_49181,N_48974);
or UO_2146 (O_2146,N_49896,N_49828);
nand UO_2147 (O_2147,N_48888,N_48491);
or UO_2148 (O_2148,N_48880,N_48738);
xnor UO_2149 (O_2149,N_49302,N_48024);
or UO_2150 (O_2150,N_49533,N_48527);
or UO_2151 (O_2151,N_49887,N_48291);
or UO_2152 (O_2152,N_49165,N_48897);
nor UO_2153 (O_2153,N_49262,N_48353);
xnor UO_2154 (O_2154,N_49545,N_48492);
nor UO_2155 (O_2155,N_49417,N_48896);
xor UO_2156 (O_2156,N_49978,N_48524);
nand UO_2157 (O_2157,N_48311,N_48613);
nand UO_2158 (O_2158,N_48818,N_49500);
or UO_2159 (O_2159,N_48275,N_48630);
nor UO_2160 (O_2160,N_49387,N_48188);
xor UO_2161 (O_2161,N_48918,N_49882);
nor UO_2162 (O_2162,N_49640,N_49228);
and UO_2163 (O_2163,N_49218,N_48039);
nand UO_2164 (O_2164,N_48543,N_49794);
or UO_2165 (O_2165,N_48673,N_49844);
nor UO_2166 (O_2166,N_49599,N_48540);
and UO_2167 (O_2167,N_49826,N_48493);
xor UO_2168 (O_2168,N_49140,N_48228);
and UO_2169 (O_2169,N_49054,N_49121);
xnor UO_2170 (O_2170,N_49081,N_48806);
or UO_2171 (O_2171,N_49629,N_48566);
nor UO_2172 (O_2172,N_48429,N_48394);
xor UO_2173 (O_2173,N_49518,N_49024);
nand UO_2174 (O_2174,N_48321,N_48512);
or UO_2175 (O_2175,N_49641,N_48150);
and UO_2176 (O_2176,N_48976,N_49457);
xnor UO_2177 (O_2177,N_49232,N_49916);
and UO_2178 (O_2178,N_48951,N_49044);
nand UO_2179 (O_2179,N_49811,N_49340);
xor UO_2180 (O_2180,N_48195,N_48688);
or UO_2181 (O_2181,N_48281,N_48091);
xor UO_2182 (O_2182,N_49530,N_48812);
and UO_2183 (O_2183,N_48395,N_49151);
nand UO_2184 (O_2184,N_49618,N_48342);
and UO_2185 (O_2185,N_49723,N_48143);
xnor UO_2186 (O_2186,N_48348,N_49096);
nand UO_2187 (O_2187,N_49096,N_49142);
and UO_2188 (O_2188,N_49654,N_48649);
nand UO_2189 (O_2189,N_48330,N_49452);
or UO_2190 (O_2190,N_49404,N_49963);
and UO_2191 (O_2191,N_49318,N_49545);
nor UO_2192 (O_2192,N_48033,N_49278);
xnor UO_2193 (O_2193,N_49978,N_48428);
or UO_2194 (O_2194,N_49749,N_48653);
and UO_2195 (O_2195,N_49216,N_49944);
and UO_2196 (O_2196,N_48010,N_49152);
or UO_2197 (O_2197,N_48657,N_48326);
nand UO_2198 (O_2198,N_49142,N_48197);
and UO_2199 (O_2199,N_49582,N_48797);
or UO_2200 (O_2200,N_49092,N_49493);
nand UO_2201 (O_2201,N_49749,N_48103);
or UO_2202 (O_2202,N_49172,N_48967);
or UO_2203 (O_2203,N_48264,N_48146);
xnor UO_2204 (O_2204,N_49896,N_49600);
nor UO_2205 (O_2205,N_48947,N_49814);
xnor UO_2206 (O_2206,N_48134,N_48346);
nor UO_2207 (O_2207,N_49354,N_49411);
and UO_2208 (O_2208,N_49444,N_49015);
and UO_2209 (O_2209,N_49031,N_48984);
nor UO_2210 (O_2210,N_49963,N_48827);
and UO_2211 (O_2211,N_49373,N_49295);
xor UO_2212 (O_2212,N_49640,N_48325);
and UO_2213 (O_2213,N_48997,N_48604);
and UO_2214 (O_2214,N_49878,N_49352);
xnor UO_2215 (O_2215,N_49529,N_48314);
nand UO_2216 (O_2216,N_48984,N_49842);
nor UO_2217 (O_2217,N_49102,N_48752);
nand UO_2218 (O_2218,N_49655,N_48796);
xnor UO_2219 (O_2219,N_49816,N_48829);
xor UO_2220 (O_2220,N_49872,N_48391);
nor UO_2221 (O_2221,N_49764,N_49173);
or UO_2222 (O_2222,N_48899,N_48618);
nand UO_2223 (O_2223,N_48718,N_49327);
nor UO_2224 (O_2224,N_48709,N_49940);
xor UO_2225 (O_2225,N_48489,N_48036);
xnor UO_2226 (O_2226,N_48913,N_49481);
xor UO_2227 (O_2227,N_49302,N_49221);
nor UO_2228 (O_2228,N_48571,N_49382);
and UO_2229 (O_2229,N_48640,N_49244);
or UO_2230 (O_2230,N_49530,N_48447);
nor UO_2231 (O_2231,N_48812,N_49233);
xnor UO_2232 (O_2232,N_49238,N_48347);
nand UO_2233 (O_2233,N_49173,N_49392);
and UO_2234 (O_2234,N_49668,N_48425);
xnor UO_2235 (O_2235,N_49235,N_49339);
nand UO_2236 (O_2236,N_49858,N_49602);
nor UO_2237 (O_2237,N_48430,N_48991);
nand UO_2238 (O_2238,N_48159,N_49387);
and UO_2239 (O_2239,N_49136,N_48267);
xnor UO_2240 (O_2240,N_49646,N_48404);
or UO_2241 (O_2241,N_49791,N_49596);
xor UO_2242 (O_2242,N_49049,N_49740);
nand UO_2243 (O_2243,N_48313,N_48806);
xnor UO_2244 (O_2244,N_49883,N_48054);
or UO_2245 (O_2245,N_49407,N_48304);
xor UO_2246 (O_2246,N_48259,N_48070);
xnor UO_2247 (O_2247,N_48663,N_48467);
xor UO_2248 (O_2248,N_48486,N_48668);
or UO_2249 (O_2249,N_48845,N_49306);
nand UO_2250 (O_2250,N_48716,N_48981);
and UO_2251 (O_2251,N_48851,N_48015);
xor UO_2252 (O_2252,N_49158,N_49871);
nand UO_2253 (O_2253,N_48550,N_48778);
nor UO_2254 (O_2254,N_48024,N_48929);
and UO_2255 (O_2255,N_48221,N_48050);
xor UO_2256 (O_2256,N_49796,N_48116);
or UO_2257 (O_2257,N_49034,N_48411);
nor UO_2258 (O_2258,N_48967,N_48679);
nand UO_2259 (O_2259,N_49661,N_48978);
xor UO_2260 (O_2260,N_49271,N_48014);
and UO_2261 (O_2261,N_48284,N_49303);
and UO_2262 (O_2262,N_49188,N_48830);
nor UO_2263 (O_2263,N_48745,N_49128);
nor UO_2264 (O_2264,N_49484,N_48880);
nor UO_2265 (O_2265,N_49459,N_49386);
and UO_2266 (O_2266,N_48907,N_48055);
nand UO_2267 (O_2267,N_48614,N_48726);
nor UO_2268 (O_2268,N_48646,N_49756);
or UO_2269 (O_2269,N_49678,N_48485);
xor UO_2270 (O_2270,N_48938,N_48965);
nor UO_2271 (O_2271,N_48994,N_48546);
nand UO_2272 (O_2272,N_49266,N_48162);
and UO_2273 (O_2273,N_49184,N_48210);
xnor UO_2274 (O_2274,N_49927,N_49126);
xor UO_2275 (O_2275,N_49298,N_49670);
or UO_2276 (O_2276,N_48496,N_48388);
xnor UO_2277 (O_2277,N_49935,N_49127);
or UO_2278 (O_2278,N_48737,N_48923);
nor UO_2279 (O_2279,N_48145,N_48737);
and UO_2280 (O_2280,N_48886,N_48984);
xor UO_2281 (O_2281,N_48150,N_49411);
xnor UO_2282 (O_2282,N_48649,N_49575);
and UO_2283 (O_2283,N_49852,N_48750);
nor UO_2284 (O_2284,N_49741,N_48591);
xor UO_2285 (O_2285,N_48869,N_49608);
or UO_2286 (O_2286,N_48845,N_49975);
nand UO_2287 (O_2287,N_49521,N_48884);
and UO_2288 (O_2288,N_49953,N_49230);
xnor UO_2289 (O_2289,N_49713,N_48593);
or UO_2290 (O_2290,N_48621,N_49094);
xnor UO_2291 (O_2291,N_49972,N_49202);
and UO_2292 (O_2292,N_48697,N_48609);
or UO_2293 (O_2293,N_49343,N_48093);
or UO_2294 (O_2294,N_49251,N_49824);
xor UO_2295 (O_2295,N_48406,N_48834);
xnor UO_2296 (O_2296,N_49583,N_49526);
nor UO_2297 (O_2297,N_48873,N_48272);
or UO_2298 (O_2298,N_48420,N_49147);
nand UO_2299 (O_2299,N_49892,N_49486);
or UO_2300 (O_2300,N_48955,N_49428);
nor UO_2301 (O_2301,N_49199,N_49128);
and UO_2302 (O_2302,N_48236,N_49742);
and UO_2303 (O_2303,N_48403,N_48025);
nor UO_2304 (O_2304,N_48270,N_48217);
and UO_2305 (O_2305,N_49968,N_48838);
and UO_2306 (O_2306,N_49724,N_48009);
xnor UO_2307 (O_2307,N_48053,N_49294);
or UO_2308 (O_2308,N_49854,N_48826);
and UO_2309 (O_2309,N_48427,N_49065);
nand UO_2310 (O_2310,N_49523,N_49607);
and UO_2311 (O_2311,N_49672,N_48662);
nand UO_2312 (O_2312,N_48971,N_48041);
nor UO_2313 (O_2313,N_48166,N_48223);
and UO_2314 (O_2314,N_48071,N_48798);
xor UO_2315 (O_2315,N_48070,N_49507);
nand UO_2316 (O_2316,N_49303,N_48762);
nor UO_2317 (O_2317,N_49410,N_49122);
nand UO_2318 (O_2318,N_48367,N_48724);
nand UO_2319 (O_2319,N_49273,N_48302);
or UO_2320 (O_2320,N_49628,N_48716);
nand UO_2321 (O_2321,N_48080,N_48345);
nand UO_2322 (O_2322,N_49441,N_49722);
nand UO_2323 (O_2323,N_49529,N_49449);
xor UO_2324 (O_2324,N_49023,N_49574);
and UO_2325 (O_2325,N_49828,N_49278);
or UO_2326 (O_2326,N_48119,N_48503);
and UO_2327 (O_2327,N_48075,N_49069);
xor UO_2328 (O_2328,N_48962,N_49886);
and UO_2329 (O_2329,N_48457,N_48720);
and UO_2330 (O_2330,N_48164,N_49392);
nand UO_2331 (O_2331,N_49861,N_49554);
or UO_2332 (O_2332,N_48561,N_48893);
nor UO_2333 (O_2333,N_48567,N_48233);
xnor UO_2334 (O_2334,N_48981,N_49187);
xnor UO_2335 (O_2335,N_49756,N_49244);
xnor UO_2336 (O_2336,N_49020,N_48894);
nand UO_2337 (O_2337,N_48424,N_48964);
or UO_2338 (O_2338,N_49433,N_49939);
and UO_2339 (O_2339,N_49354,N_49120);
and UO_2340 (O_2340,N_49012,N_49836);
and UO_2341 (O_2341,N_48510,N_49245);
nand UO_2342 (O_2342,N_48330,N_48469);
or UO_2343 (O_2343,N_49523,N_48715);
or UO_2344 (O_2344,N_49693,N_49259);
or UO_2345 (O_2345,N_48620,N_49320);
xnor UO_2346 (O_2346,N_48287,N_49294);
or UO_2347 (O_2347,N_48308,N_48899);
or UO_2348 (O_2348,N_49117,N_48587);
nand UO_2349 (O_2349,N_48485,N_49968);
xor UO_2350 (O_2350,N_49892,N_48484);
nand UO_2351 (O_2351,N_49132,N_49846);
nor UO_2352 (O_2352,N_48675,N_49660);
nand UO_2353 (O_2353,N_48526,N_49023);
and UO_2354 (O_2354,N_48875,N_48723);
nand UO_2355 (O_2355,N_48146,N_48426);
xor UO_2356 (O_2356,N_48568,N_49535);
and UO_2357 (O_2357,N_49655,N_48970);
or UO_2358 (O_2358,N_49615,N_48901);
or UO_2359 (O_2359,N_48500,N_48680);
xor UO_2360 (O_2360,N_49106,N_49706);
or UO_2361 (O_2361,N_48113,N_48937);
xor UO_2362 (O_2362,N_49170,N_49110);
or UO_2363 (O_2363,N_48991,N_49201);
nand UO_2364 (O_2364,N_48382,N_48485);
xnor UO_2365 (O_2365,N_48172,N_49298);
nand UO_2366 (O_2366,N_48772,N_48082);
or UO_2367 (O_2367,N_49018,N_49023);
xnor UO_2368 (O_2368,N_48816,N_49961);
nor UO_2369 (O_2369,N_48159,N_49237);
or UO_2370 (O_2370,N_48053,N_49794);
or UO_2371 (O_2371,N_49455,N_48475);
nor UO_2372 (O_2372,N_49321,N_48009);
nor UO_2373 (O_2373,N_49187,N_48305);
xnor UO_2374 (O_2374,N_49911,N_49936);
nand UO_2375 (O_2375,N_48832,N_49041);
nand UO_2376 (O_2376,N_49247,N_48841);
or UO_2377 (O_2377,N_48304,N_49955);
xor UO_2378 (O_2378,N_48198,N_48211);
or UO_2379 (O_2379,N_49648,N_49145);
nand UO_2380 (O_2380,N_49716,N_48088);
xnor UO_2381 (O_2381,N_49794,N_49724);
nand UO_2382 (O_2382,N_49772,N_48917);
or UO_2383 (O_2383,N_49188,N_49052);
nor UO_2384 (O_2384,N_49849,N_48427);
or UO_2385 (O_2385,N_48620,N_49809);
nand UO_2386 (O_2386,N_48620,N_49542);
nand UO_2387 (O_2387,N_48534,N_49809);
nand UO_2388 (O_2388,N_49502,N_48548);
nor UO_2389 (O_2389,N_49485,N_48839);
nand UO_2390 (O_2390,N_49111,N_49719);
nor UO_2391 (O_2391,N_49453,N_48289);
and UO_2392 (O_2392,N_48314,N_48493);
or UO_2393 (O_2393,N_49235,N_49086);
nand UO_2394 (O_2394,N_49197,N_48036);
and UO_2395 (O_2395,N_48242,N_49915);
and UO_2396 (O_2396,N_48213,N_48449);
nor UO_2397 (O_2397,N_48543,N_49487);
nor UO_2398 (O_2398,N_49967,N_49937);
nand UO_2399 (O_2399,N_49550,N_48137);
xnor UO_2400 (O_2400,N_48502,N_49908);
xor UO_2401 (O_2401,N_49411,N_49234);
or UO_2402 (O_2402,N_49889,N_49213);
nor UO_2403 (O_2403,N_49734,N_48871);
nor UO_2404 (O_2404,N_49063,N_49376);
nor UO_2405 (O_2405,N_49136,N_48153);
or UO_2406 (O_2406,N_49349,N_49613);
nand UO_2407 (O_2407,N_49977,N_48077);
nor UO_2408 (O_2408,N_49947,N_48228);
xnor UO_2409 (O_2409,N_48929,N_49946);
nor UO_2410 (O_2410,N_49560,N_49941);
or UO_2411 (O_2411,N_48063,N_49899);
nor UO_2412 (O_2412,N_49244,N_48131);
nor UO_2413 (O_2413,N_49034,N_49380);
and UO_2414 (O_2414,N_48368,N_48939);
and UO_2415 (O_2415,N_48886,N_48662);
or UO_2416 (O_2416,N_48457,N_48791);
nand UO_2417 (O_2417,N_49564,N_49273);
xor UO_2418 (O_2418,N_48099,N_48563);
and UO_2419 (O_2419,N_49165,N_49171);
or UO_2420 (O_2420,N_48071,N_48280);
and UO_2421 (O_2421,N_48680,N_48183);
and UO_2422 (O_2422,N_49039,N_49280);
or UO_2423 (O_2423,N_49679,N_49886);
xor UO_2424 (O_2424,N_49271,N_49249);
or UO_2425 (O_2425,N_49663,N_48195);
xnor UO_2426 (O_2426,N_49754,N_49976);
nor UO_2427 (O_2427,N_49229,N_48012);
or UO_2428 (O_2428,N_49581,N_48320);
xnor UO_2429 (O_2429,N_48043,N_49331);
xor UO_2430 (O_2430,N_48273,N_48277);
or UO_2431 (O_2431,N_49012,N_48373);
nor UO_2432 (O_2432,N_48722,N_49125);
or UO_2433 (O_2433,N_49273,N_49916);
nand UO_2434 (O_2434,N_48488,N_48238);
and UO_2435 (O_2435,N_49675,N_48357);
nor UO_2436 (O_2436,N_49575,N_49945);
nor UO_2437 (O_2437,N_48609,N_48845);
or UO_2438 (O_2438,N_49079,N_48898);
nand UO_2439 (O_2439,N_49105,N_49447);
nand UO_2440 (O_2440,N_49149,N_49968);
nand UO_2441 (O_2441,N_49430,N_49010);
xor UO_2442 (O_2442,N_48221,N_49798);
xnor UO_2443 (O_2443,N_49081,N_49858);
or UO_2444 (O_2444,N_49559,N_48253);
or UO_2445 (O_2445,N_48889,N_49045);
and UO_2446 (O_2446,N_49080,N_49698);
nor UO_2447 (O_2447,N_49802,N_49287);
and UO_2448 (O_2448,N_48498,N_49880);
xnor UO_2449 (O_2449,N_49138,N_49924);
xnor UO_2450 (O_2450,N_49936,N_48995);
nand UO_2451 (O_2451,N_49325,N_49096);
and UO_2452 (O_2452,N_48249,N_49744);
and UO_2453 (O_2453,N_48674,N_48793);
or UO_2454 (O_2454,N_49898,N_48116);
nand UO_2455 (O_2455,N_49361,N_48403);
nand UO_2456 (O_2456,N_49131,N_48992);
and UO_2457 (O_2457,N_48738,N_49741);
nor UO_2458 (O_2458,N_48143,N_48621);
nor UO_2459 (O_2459,N_48999,N_48278);
and UO_2460 (O_2460,N_48458,N_48175);
nor UO_2461 (O_2461,N_49499,N_48525);
or UO_2462 (O_2462,N_49689,N_48533);
nand UO_2463 (O_2463,N_48365,N_48857);
or UO_2464 (O_2464,N_49002,N_49062);
nand UO_2465 (O_2465,N_49996,N_48131);
nor UO_2466 (O_2466,N_49533,N_48664);
nand UO_2467 (O_2467,N_49619,N_49817);
xor UO_2468 (O_2468,N_48519,N_49357);
or UO_2469 (O_2469,N_48857,N_49751);
and UO_2470 (O_2470,N_49398,N_48158);
and UO_2471 (O_2471,N_49860,N_48624);
nor UO_2472 (O_2472,N_49860,N_49085);
xor UO_2473 (O_2473,N_49986,N_48982);
xnor UO_2474 (O_2474,N_48915,N_49257);
xnor UO_2475 (O_2475,N_48111,N_48383);
nor UO_2476 (O_2476,N_48578,N_48188);
xnor UO_2477 (O_2477,N_48634,N_49715);
nor UO_2478 (O_2478,N_49213,N_49091);
nor UO_2479 (O_2479,N_49797,N_48876);
nand UO_2480 (O_2480,N_49536,N_49064);
nand UO_2481 (O_2481,N_48760,N_49253);
and UO_2482 (O_2482,N_49143,N_49266);
nand UO_2483 (O_2483,N_49434,N_48816);
nand UO_2484 (O_2484,N_49986,N_48884);
nor UO_2485 (O_2485,N_49646,N_48052);
nand UO_2486 (O_2486,N_49472,N_49211);
nand UO_2487 (O_2487,N_49015,N_49404);
and UO_2488 (O_2488,N_49349,N_48980);
nor UO_2489 (O_2489,N_48292,N_48003);
nor UO_2490 (O_2490,N_48439,N_48546);
nor UO_2491 (O_2491,N_48832,N_48434);
and UO_2492 (O_2492,N_48376,N_48400);
xnor UO_2493 (O_2493,N_48989,N_49433);
nand UO_2494 (O_2494,N_49430,N_49368);
nor UO_2495 (O_2495,N_48128,N_48873);
nand UO_2496 (O_2496,N_49615,N_48340);
and UO_2497 (O_2497,N_49845,N_49662);
and UO_2498 (O_2498,N_49305,N_48752);
and UO_2499 (O_2499,N_49162,N_49428);
or UO_2500 (O_2500,N_49739,N_48975);
and UO_2501 (O_2501,N_49454,N_48398);
nor UO_2502 (O_2502,N_48667,N_49399);
nand UO_2503 (O_2503,N_48922,N_48156);
nand UO_2504 (O_2504,N_49416,N_48838);
xor UO_2505 (O_2505,N_48293,N_48648);
nand UO_2506 (O_2506,N_48107,N_49487);
nand UO_2507 (O_2507,N_49035,N_48398);
or UO_2508 (O_2508,N_49036,N_49613);
or UO_2509 (O_2509,N_49599,N_49951);
nand UO_2510 (O_2510,N_49003,N_49782);
nand UO_2511 (O_2511,N_48324,N_48787);
xor UO_2512 (O_2512,N_48529,N_48097);
or UO_2513 (O_2513,N_48354,N_49882);
nor UO_2514 (O_2514,N_48243,N_49311);
xor UO_2515 (O_2515,N_48503,N_49915);
or UO_2516 (O_2516,N_48629,N_49953);
and UO_2517 (O_2517,N_49065,N_49264);
or UO_2518 (O_2518,N_48884,N_48265);
nor UO_2519 (O_2519,N_48933,N_49839);
nand UO_2520 (O_2520,N_49860,N_49961);
nand UO_2521 (O_2521,N_48483,N_49312);
xor UO_2522 (O_2522,N_48478,N_49685);
nor UO_2523 (O_2523,N_49536,N_48234);
and UO_2524 (O_2524,N_49731,N_48194);
or UO_2525 (O_2525,N_48287,N_48700);
xnor UO_2526 (O_2526,N_49398,N_49296);
xor UO_2527 (O_2527,N_49305,N_49128);
xnor UO_2528 (O_2528,N_49820,N_49789);
nor UO_2529 (O_2529,N_48860,N_48668);
nand UO_2530 (O_2530,N_49380,N_49039);
and UO_2531 (O_2531,N_48096,N_49501);
xor UO_2532 (O_2532,N_48489,N_49604);
nand UO_2533 (O_2533,N_49017,N_49677);
and UO_2534 (O_2534,N_48874,N_49803);
xor UO_2535 (O_2535,N_48736,N_48883);
or UO_2536 (O_2536,N_48148,N_48411);
and UO_2537 (O_2537,N_48501,N_49406);
nand UO_2538 (O_2538,N_49505,N_49779);
nor UO_2539 (O_2539,N_49918,N_49012);
nand UO_2540 (O_2540,N_48607,N_48124);
nor UO_2541 (O_2541,N_49870,N_49078);
and UO_2542 (O_2542,N_48491,N_49258);
nor UO_2543 (O_2543,N_48523,N_48743);
nand UO_2544 (O_2544,N_48630,N_48039);
xor UO_2545 (O_2545,N_49462,N_48062);
and UO_2546 (O_2546,N_49758,N_48336);
nand UO_2547 (O_2547,N_49237,N_49872);
or UO_2548 (O_2548,N_49921,N_48019);
nor UO_2549 (O_2549,N_49091,N_49003);
nand UO_2550 (O_2550,N_49010,N_49149);
nand UO_2551 (O_2551,N_48453,N_48969);
xnor UO_2552 (O_2552,N_49269,N_49986);
or UO_2553 (O_2553,N_48127,N_48870);
nor UO_2554 (O_2554,N_49961,N_49534);
xnor UO_2555 (O_2555,N_48750,N_49599);
nand UO_2556 (O_2556,N_48473,N_48549);
xor UO_2557 (O_2557,N_49092,N_48265);
nand UO_2558 (O_2558,N_49214,N_49429);
and UO_2559 (O_2559,N_48576,N_49951);
or UO_2560 (O_2560,N_49972,N_48491);
nand UO_2561 (O_2561,N_49339,N_48069);
nand UO_2562 (O_2562,N_48933,N_49762);
nand UO_2563 (O_2563,N_48053,N_49714);
and UO_2564 (O_2564,N_48175,N_49224);
nor UO_2565 (O_2565,N_48854,N_49601);
nand UO_2566 (O_2566,N_49896,N_49964);
nor UO_2567 (O_2567,N_48317,N_49369);
xnor UO_2568 (O_2568,N_49673,N_48230);
and UO_2569 (O_2569,N_49848,N_49048);
or UO_2570 (O_2570,N_48265,N_49307);
nor UO_2571 (O_2571,N_48641,N_48586);
nor UO_2572 (O_2572,N_49075,N_48684);
nand UO_2573 (O_2573,N_49794,N_49676);
or UO_2574 (O_2574,N_49881,N_48246);
or UO_2575 (O_2575,N_48140,N_49605);
nor UO_2576 (O_2576,N_48571,N_49235);
or UO_2577 (O_2577,N_48317,N_48386);
nand UO_2578 (O_2578,N_48028,N_49812);
nor UO_2579 (O_2579,N_48035,N_49702);
nor UO_2580 (O_2580,N_48800,N_48915);
nand UO_2581 (O_2581,N_49161,N_49976);
nor UO_2582 (O_2582,N_48791,N_49204);
nor UO_2583 (O_2583,N_49033,N_48833);
nor UO_2584 (O_2584,N_48974,N_49737);
nand UO_2585 (O_2585,N_49318,N_49461);
nand UO_2586 (O_2586,N_48972,N_49609);
and UO_2587 (O_2587,N_49749,N_49917);
xnor UO_2588 (O_2588,N_48847,N_48703);
xor UO_2589 (O_2589,N_49880,N_49235);
nand UO_2590 (O_2590,N_48011,N_49105);
xor UO_2591 (O_2591,N_49088,N_49884);
and UO_2592 (O_2592,N_49823,N_48555);
or UO_2593 (O_2593,N_48232,N_48624);
or UO_2594 (O_2594,N_49810,N_49197);
and UO_2595 (O_2595,N_49847,N_48671);
and UO_2596 (O_2596,N_48723,N_48058);
and UO_2597 (O_2597,N_48610,N_49833);
xor UO_2598 (O_2598,N_49147,N_48378);
and UO_2599 (O_2599,N_49339,N_49174);
or UO_2600 (O_2600,N_48744,N_49274);
nand UO_2601 (O_2601,N_48027,N_48133);
or UO_2602 (O_2602,N_49229,N_49211);
xnor UO_2603 (O_2603,N_48236,N_48857);
nor UO_2604 (O_2604,N_48857,N_48018);
nor UO_2605 (O_2605,N_49484,N_49695);
and UO_2606 (O_2606,N_49840,N_49956);
and UO_2607 (O_2607,N_49355,N_48938);
nand UO_2608 (O_2608,N_49256,N_49849);
xnor UO_2609 (O_2609,N_48819,N_49784);
xnor UO_2610 (O_2610,N_48745,N_48530);
and UO_2611 (O_2611,N_48279,N_49237);
or UO_2612 (O_2612,N_48175,N_48725);
xnor UO_2613 (O_2613,N_49430,N_49316);
or UO_2614 (O_2614,N_49513,N_49598);
xnor UO_2615 (O_2615,N_48184,N_48109);
nor UO_2616 (O_2616,N_49110,N_49246);
and UO_2617 (O_2617,N_49117,N_48893);
nand UO_2618 (O_2618,N_48448,N_48523);
or UO_2619 (O_2619,N_48523,N_49911);
or UO_2620 (O_2620,N_48111,N_49741);
nor UO_2621 (O_2621,N_48618,N_48967);
nand UO_2622 (O_2622,N_48113,N_48360);
xnor UO_2623 (O_2623,N_48206,N_48616);
nand UO_2624 (O_2624,N_49025,N_49288);
and UO_2625 (O_2625,N_49460,N_48630);
and UO_2626 (O_2626,N_49988,N_49063);
and UO_2627 (O_2627,N_48813,N_48275);
nand UO_2628 (O_2628,N_49215,N_48046);
xnor UO_2629 (O_2629,N_49976,N_49009);
nor UO_2630 (O_2630,N_49648,N_49437);
xor UO_2631 (O_2631,N_48735,N_49581);
or UO_2632 (O_2632,N_49547,N_49289);
or UO_2633 (O_2633,N_49207,N_48053);
nand UO_2634 (O_2634,N_48199,N_48010);
nand UO_2635 (O_2635,N_49630,N_48041);
or UO_2636 (O_2636,N_48470,N_48150);
nand UO_2637 (O_2637,N_49606,N_48059);
xor UO_2638 (O_2638,N_49657,N_49915);
or UO_2639 (O_2639,N_48137,N_48023);
nor UO_2640 (O_2640,N_49040,N_48741);
and UO_2641 (O_2641,N_49412,N_48675);
nand UO_2642 (O_2642,N_49942,N_49195);
xnor UO_2643 (O_2643,N_49276,N_49143);
and UO_2644 (O_2644,N_49332,N_48552);
nand UO_2645 (O_2645,N_48233,N_48087);
xor UO_2646 (O_2646,N_48351,N_49633);
and UO_2647 (O_2647,N_48280,N_48424);
nand UO_2648 (O_2648,N_48818,N_48652);
and UO_2649 (O_2649,N_48122,N_49150);
xnor UO_2650 (O_2650,N_48648,N_48991);
and UO_2651 (O_2651,N_49947,N_49696);
nand UO_2652 (O_2652,N_48083,N_48469);
and UO_2653 (O_2653,N_49061,N_48114);
nand UO_2654 (O_2654,N_48885,N_48483);
nand UO_2655 (O_2655,N_49655,N_48306);
nor UO_2656 (O_2656,N_49019,N_48335);
nor UO_2657 (O_2657,N_48777,N_48501);
nor UO_2658 (O_2658,N_49394,N_48696);
and UO_2659 (O_2659,N_48572,N_49901);
nand UO_2660 (O_2660,N_49091,N_48544);
nor UO_2661 (O_2661,N_49806,N_49086);
and UO_2662 (O_2662,N_48339,N_48149);
and UO_2663 (O_2663,N_48915,N_49589);
xnor UO_2664 (O_2664,N_48508,N_48249);
nor UO_2665 (O_2665,N_49297,N_49092);
xor UO_2666 (O_2666,N_49849,N_49591);
and UO_2667 (O_2667,N_48018,N_48340);
nor UO_2668 (O_2668,N_49231,N_49048);
and UO_2669 (O_2669,N_49615,N_49297);
or UO_2670 (O_2670,N_48138,N_48957);
and UO_2671 (O_2671,N_48067,N_49447);
and UO_2672 (O_2672,N_48241,N_49845);
nor UO_2673 (O_2673,N_48103,N_48545);
nand UO_2674 (O_2674,N_49815,N_49168);
xnor UO_2675 (O_2675,N_48941,N_49913);
and UO_2676 (O_2676,N_49247,N_48515);
nand UO_2677 (O_2677,N_48638,N_49084);
and UO_2678 (O_2678,N_49612,N_49515);
and UO_2679 (O_2679,N_49763,N_49431);
xor UO_2680 (O_2680,N_49073,N_49384);
or UO_2681 (O_2681,N_49738,N_48059);
and UO_2682 (O_2682,N_48995,N_48862);
xor UO_2683 (O_2683,N_48850,N_49503);
or UO_2684 (O_2684,N_49237,N_49824);
or UO_2685 (O_2685,N_49046,N_49237);
nor UO_2686 (O_2686,N_49451,N_48562);
nor UO_2687 (O_2687,N_48993,N_49510);
or UO_2688 (O_2688,N_49674,N_49425);
xnor UO_2689 (O_2689,N_48010,N_48997);
or UO_2690 (O_2690,N_48204,N_48856);
and UO_2691 (O_2691,N_49199,N_49112);
xor UO_2692 (O_2692,N_48062,N_49379);
nor UO_2693 (O_2693,N_49547,N_48290);
nand UO_2694 (O_2694,N_48840,N_49870);
or UO_2695 (O_2695,N_48839,N_49130);
xnor UO_2696 (O_2696,N_48059,N_48463);
nor UO_2697 (O_2697,N_48691,N_48932);
nor UO_2698 (O_2698,N_49443,N_49279);
or UO_2699 (O_2699,N_49837,N_48560);
and UO_2700 (O_2700,N_48600,N_48061);
xnor UO_2701 (O_2701,N_49490,N_48338);
nor UO_2702 (O_2702,N_48226,N_49237);
xor UO_2703 (O_2703,N_49028,N_48790);
and UO_2704 (O_2704,N_48126,N_48091);
nand UO_2705 (O_2705,N_49165,N_49790);
and UO_2706 (O_2706,N_48349,N_48420);
or UO_2707 (O_2707,N_48180,N_49953);
xnor UO_2708 (O_2708,N_49333,N_48881);
or UO_2709 (O_2709,N_48514,N_49863);
nand UO_2710 (O_2710,N_48475,N_48884);
or UO_2711 (O_2711,N_49008,N_48746);
and UO_2712 (O_2712,N_48386,N_49759);
nor UO_2713 (O_2713,N_49438,N_48645);
nor UO_2714 (O_2714,N_48790,N_49694);
nand UO_2715 (O_2715,N_49495,N_48778);
and UO_2716 (O_2716,N_49408,N_49240);
and UO_2717 (O_2717,N_49043,N_48688);
or UO_2718 (O_2718,N_48724,N_48469);
nand UO_2719 (O_2719,N_49357,N_49632);
nor UO_2720 (O_2720,N_49186,N_48634);
nor UO_2721 (O_2721,N_49067,N_48799);
xor UO_2722 (O_2722,N_49208,N_49109);
nand UO_2723 (O_2723,N_49244,N_49976);
nand UO_2724 (O_2724,N_48858,N_49679);
and UO_2725 (O_2725,N_48555,N_48526);
nand UO_2726 (O_2726,N_49574,N_49033);
nand UO_2727 (O_2727,N_48619,N_48636);
nor UO_2728 (O_2728,N_48035,N_48325);
nor UO_2729 (O_2729,N_49014,N_49310);
xnor UO_2730 (O_2730,N_48085,N_49513);
and UO_2731 (O_2731,N_48544,N_48186);
xor UO_2732 (O_2732,N_48320,N_49736);
or UO_2733 (O_2733,N_49009,N_48269);
or UO_2734 (O_2734,N_48129,N_48206);
or UO_2735 (O_2735,N_48612,N_49417);
or UO_2736 (O_2736,N_48607,N_49462);
and UO_2737 (O_2737,N_48663,N_49682);
nand UO_2738 (O_2738,N_48666,N_49628);
nor UO_2739 (O_2739,N_49362,N_49159);
nand UO_2740 (O_2740,N_48023,N_49369);
xor UO_2741 (O_2741,N_48688,N_49724);
or UO_2742 (O_2742,N_49393,N_49082);
or UO_2743 (O_2743,N_48791,N_48467);
nor UO_2744 (O_2744,N_48406,N_49202);
nand UO_2745 (O_2745,N_49667,N_48009);
nand UO_2746 (O_2746,N_49727,N_48853);
xor UO_2747 (O_2747,N_49401,N_49810);
nor UO_2748 (O_2748,N_49033,N_49122);
xor UO_2749 (O_2749,N_49579,N_49726);
and UO_2750 (O_2750,N_48907,N_48177);
and UO_2751 (O_2751,N_49295,N_49159);
or UO_2752 (O_2752,N_49271,N_49733);
or UO_2753 (O_2753,N_48121,N_48830);
xnor UO_2754 (O_2754,N_49264,N_49851);
or UO_2755 (O_2755,N_49896,N_49444);
nor UO_2756 (O_2756,N_49139,N_49983);
or UO_2757 (O_2757,N_49593,N_49622);
nor UO_2758 (O_2758,N_49243,N_49339);
nor UO_2759 (O_2759,N_48095,N_48405);
nor UO_2760 (O_2760,N_49801,N_48124);
nand UO_2761 (O_2761,N_49770,N_49233);
nor UO_2762 (O_2762,N_48342,N_49551);
nand UO_2763 (O_2763,N_48884,N_48533);
nand UO_2764 (O_2764,N_49556,N_48930);
and UO_2765 (O_2765,N_49009,N_49470);
xor UO_2766 (O_2766,N_48155,N_49037);
and UO_2767 (O_2767,N_48651,N_49657);
or UO_2768 (O_2768,N_49608,N_49674);
and UO_2769 (O_2769,N_48139,N_48796);
or UO_2770 (O_2770,N_48750,N_48713);
nand UO_2771 (O_2771,N_48621,N_48776);
nor UO_2772 (O_2772,N_48385,N_49437);
and UO_2773 (O_2773,N_48692,N_48108);
xnor UO_2774 (O_2774,N_49192,N_48821);
or UO_2775 (O_2775,N_48550,N_49865);
nand UO_2776 (O_2776,N_48438,N_49495);
and UO_2777 (O_2777,N_49548,N_49313);
or UO_2778 (O_2778,N_49979,N_48965);
nand UO_2779 (O_2779,N_48912,N_48732);
xor UO_2780 (O_2780,N_48737,N_48395);
or UO_2781 (O_2781,N_49873,N_48987);
or UO_2782 (O_2782,N_49943,N_48171);
xor UO_2783 (O_2783,N_48194,N_48321);
nor UO_2784 (O_2784,N_49606,N_49256);
nand UO_2785 (O_2785,N_48439,N_49619);
xor UO_2786 (O_2786,N_49634,N_49236);
nand UO_2787 (O_2787,N_49664,N_49908);
nor UO_2788 (O_2788,N_48402,N_48097);
and UO_2789 (O_2789,N_49499,N_48863);
and UO_2790 (O_2790,N_49727,N_49438);
nor UO_2791 (O_2791,N_48928,N_49703);
or UO_2792 (O_2792,N_48222,N_49763);
or UO_2793 (O_2793,N_49839,N_48848);
and UO_2794 (O_2794,N_48166,N_49398);
and UO_2795 (O_2795,N_49997,N_48996);
and UO_2796 (O_2796,N_49255,N_48082);
and UO_2797 (O_2797,N_48100,N_49855);
nand UO_2798 (O_2798,N_48169,N_48305);
nor UO_2799 (O_2799,N_48241,N_49274);
xnor UO_2800 (O_2800,N_48817,N_48328);
and UO_2801 (O_2801,N_49661,N_48904);
or UO_2802 (O_2802,N_48624,N_49955);
or UO_2803 (O_2803,N_49594,N_49785);
nand UO_2804 (O_2804,N_49708,N_48733);
nand UO_2805 (O_2805,N_48284,N_49770);
xnor UO_2806 (O_2806,N_49382,N_48307);
nor UO_2807 (O_2807,N_49176,N_49668);
nand UO_2808 (O_2808,N_49575,N_48644);
nand UO_2809 (O_2809,N_49334,N_48645);
nand UO_2810 (O_2810,N_49591,N_48306);
nor UO_2811 (O_2811,N_48645,N_49999);
nor UO_2812 (O_2812,N_48408,N_49319);
nor UO_2813 (O_2813,N_49546,N_49824);
or UO_2814 (O_2814,N_49530,N_48473);
nor UO_2815 (O_2815,N_49957,N_48331);
nor UO_2816 (O_2816,N_48111,N_49702);
nand UO_2817 (O_2817,N_49577,N_49238);
and UO_2818 (O_2818,N_49577,N_49614);
xor UO_2819 (O_2819,N_48305,N_49929);
nand UO_2820 (O_2820,N_48743,N_49367);
and UO_2821 (O_2821,N_48277,N_49043);
nor UO_2822 (O_2822,N_48465,N_49885);
nor UO_2823 (O_2823,N_48691,N_48472);
and UO_2824 (O_2824,N_49133,N_48204);
and UO_2825 (O_2825,N_49136,N_48711);
nand UO_2826 (O_2826,N_48344,N_49907);
xor UO_2827 (O_2827,N_48682,N_48537);
nand UO_2828 (O_2828,N_48803,N_49422);
nand UO_2829 (O_2829,N_48583,N_49737);
or UO_2830 (O_2830,N_48484,N_48891);
xnor UO_2831 (O_2831,N_48313,N_49104);
xnor UO_2832 (O_2832,N_48945,N_49559);
or UO_2833 (O_2833,N_48093,N_49223);
xnor UO_2834 (O_2834,N_48305,N_49933);
or UO_2835 (O_2835,N_49606,N_48832);
nor UO_2836 (O_2836,N_49899,N_48811);
nor UO_2837 (O_2837,N_48491,N_48568);
nand UO_2838 (O_2838,N_49659,N_48647);
or UO_2839 (O_2839,N_48884,N_49075);
nand UO_2840 (O_2840,N_49426,N_49037);
nand UO_2841 (O_2841,N_49240,N_49907);
or UO_2842 (O_2842,N_49586,N_48900);
nor UO_2843 (O_2843,N_49225,N_48281);
xnor UO_2844 (O_2844,N_48311,N_48500);
xnor UO_2845 (O_2845,N_49721,N_48140);
or UO_2846 (O_2846,N_49655,N_49871);
or UO_2847 (O_2847,N_48630,N_49162);
nand UO_2848 (O_2848,N_48766,N_48553);
nor UO_2849 (O_2849,N_48487,N_48665);
or UO_2850 (O_2850,N_49250,N_49861);
or UO_2851 (O_2851,N_49213,N_49564);
or UO_2852 (O_2852,N_49051,N_49841);
nand UO_2853 (O_2853,N_49634,N_49635);
nor UO_2854 (O_2854,N_49923,N_48552);
xor UO_2855 (O_2855,N_48910,N_49427);
or UO_2856 (O_2856,N_48072,N_49885);
or UO_2857 (O_2857,N_49674,N_49927);
nor UO_2858 (O_2858,N_48865,N_48516);
nand UO_2859 (O_2859,N_48206,N_48585);
nand UO_2860 (O_2860,N_48097,N_49776);
nand UO_2861 (O_2861,N_48764,N_48158);
or UO_2862 (O_2862,N_49219,N_49396);
and UO_2863 (O_2863,N_49882,N_48559);
xor UO_2864 (O_2864,N_48702,N_48082);
xor UO_2865 (O_2865,N_48766,N_48228);
xor UO_2866 (O_2866,N_49650,N_48770);
xnor UO_2867 (O_2867,N_48580,N_48373);
nand UO_2868 (O_2868,N_49433,N_48144);
nand UO_2869 (O_2869,N_49819,N_49005);
xor UO_2870 (O_2870,N_48534,N_48212);
nand UO_2871 (O_2871,N_49818,N_49651);
xor UO_2872 (O_2872,N_48309,N_48007);
and UO_2873 (O_2873,N_49133,N_49708);
xor UO_2874 (O_2874,N_48776,N_48298);
and UO_2875 (O_2875,N_48823,N_49761);
nand UO_2876 (O_2876,N_49598,N_49053);
nor UO_2877 (O_2877,N_48500,N_48541);
or UO_2878 (O_2878,N_49795,N_49867);
nand UO_2879 (O_2879,N_48354,N_49108);
nor UO_2880 (O_2880,N_49790,N_49817);
nor UO_2881 (O_2881,N_49657,N_49000);
and UO_2882 (O_2882,N_48874,N_49007);
or UO_2883 (O_2883,N_48164,N_49993);
or UO_2884 (O_2884,N_48684,N_48386);
and UO_2885 (O_2885,N_48419,N_48981);
nand UO_2886 (O_2886,N_49873,N_49224);
nand UO_2887 (O_2887,N_48482,N_48051);
xnor UO_2888 (O_2888,N_48835,N_48727);
nand UO_2889 (O_2889,N_49869,N_48695);
nand UO_2890 (O_2890,N_49220,N_48496);
nand UO_2891 (O_2891,N_48539,N_48785);
or UO_2892 (O_2892,N_49028,N_48419);
nand UO_2893 (O_2893,N_49304,N_48005);
or UO_2894 (O_2894,N_48833,N_48534);
nor UO_2895 (O_2895,N_49855,N_48931);
and UO_2896 (O_2896,N_48936,N_49756);
and UO_2897 (O_2897,N_49442,N_48712);
nand UO_2898 (O_2898,N_49116,N_48357);
xnor UO_2899 (O_2899,N_48884,N_48905);
nand UO_2900 (O_2900,N_48543,N_49438);
xor UO_2901 (O_2901,N_48517,N_48675);
and UO_2902 (O_2902,N_49005,N_49666);
and UO_2903 (O_2903,N_49810,N_48778);
and UO_2904 (O_2904,N_49929,N_48344);
nand UO_2905 (O_2905,N_48048,N_48558);
and UO_2906 (O_2906,N_49294,N_49151);
or UO_2907 (O_2907,N_48705,N_49883);
xnor UO_2908 (O_2908,N_49692,N_49861);
xnor UO_2909 (O_2909,N_48780,N_48939);
and UO_2910 (O_2910,N_49590,N_49591);
xnor UO_2911 (O_2911,N_49337,N_49756);
nand UO_2912 (O_2912,N_48178,N_48239);
xnor UO_2913 (O_2913,N_49953,N_49143);
or UO_2914 (O_2914,N_48465,N_48797);
and UO_2915 (O_2915,N_48634,N_49672);
and UO_2916 (O_2916,N_48512,N_48296);
xnor UO_2917 (O_2917,N_48088,N_48779);
xnor UO_2918 (O_2918,N_49744,N_49228);
or UO_2919 (O_2919,N_49938,N_48426);
nand UO_2920 (O_2920,N_49222,N_49305);
xnor UO_2921 (O_2921,N_49497,N_49228);
and UO_2922 (O_2922,N_48395,N_49827);
xnor UO_2923 (O_2923,N_48368,N_49652);
nand UO_2924 (O_2924,N_48889,N_49284);
xor UO_2925 (O_2925,N_49998,N_48335);
and UO_2926 (O_2926,N_48499,N_49660);
xor UO_2927 (O_2927,N_49535,N_48209);
or UO_2928 (O_2928,N_49659,N_49893);
and UO_2929 (O_2929,N_49914,N_48212);
or UO_2930 (O_2930,N_49625,N_49162);
nand UO_2931 (O_2931,N_49250,N_48680);
xnor UO_2932 (O_2932,N_48622,N_48234);
nand UO_2933 (O_2933,N_49615,N_49550);
xor UO_2934 (O_2934,N_48648,N_49930);
and UO_2935 (O_2935,N_49276,N_48659);
nand UO_2936 (O_2936,N_49732,N_48412);
xnor UO_2937 (O_2937,N_49324,N_48561);
and UO_2938 (O_2938,N_49615,N_49468);
and UO_2939 (O_2939,N_48444,N_48310);
nor UO_2940 (O_2940,N_49949,N_49659);
or UO_2941 (O_2941,N_48387,N_48163);
or UO_2942 (O_2942,N_48948,N_48411);
xnor UO_2943 (O_2943,N_48791,N_49532);
xnor UO_2944 (O_2944,N_49828,N_49900);
or UO_2945 (O_2945,N_49637,N_49200);
nand UO_2946 (O_2946,N_49073,N_48092);
or UO_2947 (O_2947,N_49006,N_48150);
and UO_2948 (O_2948,N_49890,N_48064);
and UO_2949 (O_2949,N_48720,N_48544);
nor UO_2950 (O_2950,N_49599,N_49413);
xnor UO_2951 (O_2951,N_49791,N_49655);
or UO_2952 (O_2952,N_49433,N_49895);
nand UO_2953 (O_2953,N_49382,N_49261);
xor UO_2954 (O_2954,N_49520,N_49095);
nand UO_2955 (O_2955,N_48263,N_48593);
and UO_2956 (O_2956,N_48894,N_49505);
nand UO_2957 (O_2957,N_48953,N_48959);
nand UO_2958 (O_2958,N_49258,N_49923);
nor UO_2959 (O_2959,N_49913,N_48591);
or UO_2960 (O_2960,N_48115,N_49959);
nand UO_2961 (O_2961,N_48071,N_48136);
nor UO_2962 (O_2962,N_48733,N_49803);
and UO_2963 (O_2963,N_49614,N_49790);
or UO_2964 (O_2964,N_49863,N_48570);
xnor UO_2965 (O_2965,N_49970,N_49093);
and UO_2966 (O_2966,N_49524,N_48065);
xor UO_2967 (O_2967,N_48536,N_49766);
and UO_2968 (O_2968,N_48165,N_48285);
and UO_2969 (O_2969,N_49316,N_49724);
nor UO_2970 (O_2970,N_48313,N_49262);
and UO_2971 (O_2971,N_49662,N_49621);
xor UO_2972 (O_2972,N_49864,N_49552);
nor UO_2973 (O_2973,N_49753,N_49144);
or UO_2974 (O_2974,N_48192,N_48601);
xnor UO_2975 (O_2975,N_49883,N_48392);
or UO_2976 (O_2976,N_49754,N_48205);
nor UO_2977 (O_2977,N_48119,N_48872);
xor UO_2978 (O_2978,N_48271,N_48747);
and UO_2979 (O_2979,N_49101,N_49055);
nor UO_2980 (O_2980,N_49412,N_48791);
nor UO_2981 (O_2981,N_48793,N_48356);
and UO_2982 (O_2982,N_49862,N_49246);
xnor UO_2983 (O_2983,N_48783,N_49270);
and UO_2984 (O_2984,N_49591,N_49484);
nand UO_2985 (O_2985,N_49051,N_49178);
xnor UO_2986 (O_2986,N_48477,N_48569);
xnor UO_2987 (O_2987,N_49870,N_49061);
nor UO_2988 (O_2988,N_49466,N_48582);
nand UO_2989 (O_2989,N_48819,N_49230);
nand UO_2990 (O_2990,N_48435,N_48036);
nor UO_2991 (O_2991,N_48551,N_49357);
or UO_2992 (O_2992,N_49091,N_48208);
nand UO_2993 (O_2993,N_48881,N_48669);
nor UO_2994 (O_2994,N_49804,N_48038);
xnor UO_2995 (O_2995,N_49916,N_48582);
or UO_2996 (O_2996,N_49186,N_48127);
and UO_2997 (O_2997,N_48773,N_48920);
nand UO_2998 (O_2998,N_49952,N_49410);
or UO_2999 (O_2999,N_48622,N_49711);
and UO_3000 (O_3000,N_49056,N_49660);
nand UO_3001 (O_3001,N_49894,N_48256);
nor UO_3002 (O_3002,N_49400,N_49751);
nor UO_3003 (O_3003,N_49935,N_49260);
nand UO_3004 (O_3004,N_49249,N_48733);
and UO_3005 (O_3005,N_48840,N_48506);
nor UO_3006 (O_3006,N_48476,N_48995);
xnor UO_3007 (O_3007,N_49732,N_49935);
xnor UO_3008 (O_3008,N_49920,N_48606);
and UO_3009 (O_3009,N_49806,N_48535);
xnor UO_3010 (O_3010,N_48010,N_48312);
nor UO_3011 (O_3011,N_48676,N_48565);
nand UO_3012 (O_3012,N_49308,N_49345);
nand UO_3013 (O_3013,N_49443,N_48888);
or UO_3014 (O_3014,N_48882,N_48471);
nor UO_3015 (O_3015,N_48051,N_49964);
or UO_3016 (O_3016,N_49598,N_48318);
nor UO_3017 (O_3017,N_48161,N_48117);
nor UO_3018 (O_3018,N_48012,N_48873);
nand UO_3019 (O_3019,N_49815,N_48518);
xor UO_3020 (O_3020,N_48106,N_48259);
or UO_3021 (O_3021,N_48611,N_48350);
nand UO_3022 (O_3022,N_49309,N_48960);
or UO_3023 (O_3023,N_48792,N_49903);
or UO_3024 (O_3024,N_48751,N_49933);
or UO_3025 (O_3025,N_49874,N_48169);
or UO_3026 (O_3026,N_48349,N_48224);
nor UO_3027 (O_3027,N_49344,N_49294);
and UO_3028 (O_3028,N_49494,N_48255);
or UO_3029 (O_3029,N_48989,N_49013);
xnor UO_3030 (O_3030,N_49277,N_49404);
xor UO_3031 (O_3031,N_49891,N_49258);
or UO_3032 (O_3032,N_49615,N_49291);
and UO_3033 (O_3033,N_48516,N_48661);
and UO_3034 (O_3034,N_48212,N_49940);
or UO_3035 (O_3035,N_49804,N_48373);
or UO_3036 (O_3036,N_49126,N_49446);
xor UO_3037 (O_3037,N_48644,N_49845);
xor UO_3038 (O_3038,N_49624,N_48888);
nor UO_3039 (O_3039,N_48504,N_49711);
and UO_3040 (O_3040,N_49087,N_49669);
nand UO_3041 (O_3041,N_49336,N_48168);
or UO_3042 (O_3042,N_49821,N_49709);
nand UO_3043 (O_3043,N_49564,N_49038);
and UO_3044 (O_3044,N_49237,N_49276);
or UO_3045 (O_3045,N_48407,N_48526);
nor UO_3046 (O_3046,N_48663,N_48535);
xnor UO_3047 (O_3047,N_49816,N_48197);
or UO_3048 (O_3048,N_49733,N_49319);
xor UO_3049 (O_3049,N_48029,N_48219);
and UO_3050 (O_3050,N_48255,N_49325);
and UO_3051 (O_3051,N_48583,N_48360);
nor UO_3052 (O_3052,N_48371,N_48835);
xnor UO_3053 (O_3053,N_48624,N_49960);
xnor UO_3054 (O_3054,N_48877,N_48102);
and UO_3055 (O_3055,N_48930,N_49963);
nor UO_3056 (O_3056,N_49373,N_49355);
or UO_3057 (O_3057,N_48091,N_49223);
xor UO_3058 (O_3058,N_49565,N_49810);
nand UO_3059 (O_3059,N_48251,N_48370);
xor UO_3060 (O_3060,N_48121,N_49157);
nor UO_3061 (O_3061,N_49301,N_49614);
xnor UO_3062 (O_3062,N_49634,N_48890);
or UO_3063 (O_3063,N_49710,N_48961);
xnor UO_3064 (O_3064,N_49327,N_49295);
and UO_3065 (O_3065,N_48162,N_48429);
xor UO_3066 (O_3066,N_49068,N_49307);
xor UO_3067 (O_3067,N_48198,N_48038);
and UO_3068 (O_3068,N_48194,N_49263);
and UO_3069 (O_3069,N_48884,N_49493);
or UO_3070 (O_3070,N_49690,N_49026);
and UO_3071 (O_3071,N_48153,N_48473);
nor UO_3072 (O_3072,N_48933,N_49705);
nand UO_3073 (O_3073,N_49870,N_48727);
or UO_3074 (O_3074,N_48332,N_49054);
xnor UO_3075 (O_3075,N_48164,N_49418);
xor UO_3076 (O_3076,N_49447,N_49786);
nand UO_3077 (O_3077,N_49433,N_49876);
or UO_3078 (O_3078,N_49241,N_48911);
nor UO_3079 (O_3079,N_48987,N_48104);
and UO_3080 (O_3080,N_48428,N_48907);
xnor UO_3081 (O_3081,N_49337,N_49746);
and UO_3082 (O_3082,N_49702,N_49224);
xor UO_3083 (O_3083,N_48304,N_49383);
nand UO_3084 (O_3084,N_49129,N_48290);
and UO_3085 (O_3085,N_48109,N_48100);
nor UO_3086 (O_3086,N_48667,N_49943);
nand UO_3087 (O_3087,N_49071,N_49112);
xor UO_3088 (O_3088,N_48018,N_48740);
nand UO_3089 (O_3089,N_49753,N_49602);
nand UO_3090 (O_3090,N_48377,N_49823);
and UO_3091 (O_3091,N_49107,N_49389);
or UO_3092 (O_3092,N_49382,N_49596);
and UO_3093 (O_3093,N_48870,N_48718);
and UO_3094 (O_3094,N_48297,N_48794);
nand UO_3095 (O_3095,N_48908,N_48141);
nor UO_3096 (O_3096,N_49832,N_49000);
and UO_3097 (O_3097,N_49999,N_49913);
and UO_3098 (O_3098,N_49113,N_49474);
xor UO_3099 (O_3099,N_48986,N_49001);
nand UO_3100 (O_3100,N_48062,N_49835);
or UO_3101 (O_3101,N_49016,N_49699);
and UO_3102 (O_3102,N_49595,N_49494);
nor UO_3103 (O_3103,N_48400,N_49048);
nor UO_3104 (O_3104,N_48641,N_48233);
and UO_3105 (O_3105,N_48799,N_48066);
nand UO_3106 (O_3106,N_48566,N_48709);
or UO_3107 (O_3107,N_49139,N_48943);
and UO_3108 (O_3108,N_49376,N_48909);
xor UO_3109 (O_3109,N_49009,N_48480);
nand UO_3110 (O_3110,N_49415,N_48673);
nor UO_3111 (O_3111,N_49334,N_49403);
nand UO_3112 (O_3112,N_49386,N_49612);
nor UO_3113 (O_3113,N_49191,N_49970);
or UO_3114 (O_3114,N_49919,N_49646);
and UO_3115 (O_3115,N_48322,N_49292);
and UO_3116 (O_3116,N_48945,N_49852);
and UO_3117 (O_3117,N_49998,N_49343);
and UO_3118 (O_3118,N_48912,N_48039);
nand UO_3119 (O_3119,N_49860,N_48133);
nor UO_3120 (O_3120,N_48848,N_48901);
xnor UO_3121 (O_3121,N_49723,N_48464);
nand UO_3122 (O_3122,N_49380,N_48753);
xor UO_3123 (O_3123,N_49852,N_49521);
or UO_3124 (O_3124,N_48853,N_48003);
or UO_3125 (O_3125,N_49447,N_48940);
nor UO_3126 (O_3126,N_49502,N_49614);
xor UO_3127 (O_3127,N_49336,N_49801);
or UO_3128 (O_3128,N_49162,N_49708);
nor UO_3129 (O_3129,N_48569,N_48263);
or UO_3130 (O_3130,N_48675,N_48336);
nand UO_3131 (O_3131,N_49508,N_49609);
and UO_3132 (O_3132,N_48815,N_49406);
xnor UO_3133 (O_3133,N_48144,N_49610);
nor UO_3134 (O_3134,N_49596,N_49327);
nor UO_3135 (O_3135,N_49637,N_48528);
or UO_3136 (O_3136,N_49301,N_48183);
nor UO_3137 (O_3137,N_48502,N_48248);
nand UO_3138 (O_3138,N_48946,N_49070);
nand UO_3139 (O_3139,N_49753,N_49930);
or UO_3140 (O_3140,N_48069,N_49424);
or UO_3141 (O_3141,N_48878,N_49319);
nor UO_3142 (O_3142,N_49473,N_49201);
and UO_3143 (O_3143,N_49709,N_48540);
or UO_3144 (O_3144,N_48183,N_48476);
nor UO_3145 (O_3145,N_49773,N_48987);
nor UO_3146 (O_3146,N_49001,N_48919);
and UO_3147 (O_3147,N_49644,N_48117);
xor UO_3148 (O_3148,N_49841,N_48751);
nor UO_3149 (O_3149,N_48928,N_48871);
or UO_3150 (O_3150,N_48070,N_48739);
nand UO_3151 (O_3151,N_48978,N_48308);
nand UO_3152 (O_3152,N_48828,N_49867);
nand UO_3153 (O_3153,N_49587,N_48541);
and UO_3154 (O_3154,N_49686,N_49781);
and UO_3155 (O_3155,N_48161,N_48699);
nor UO_3156 (O_3156,N_49778,N_49270);
nand UO_3157 (O_3157,N_49315,N_48621);
nand UO_3158 (O_3158,N_49543,N_48891);
or UO_3159 (O_3159,N_48722,N_48416);
nand UO_3160 (O_3160,N_49874,N_48917);
xnor UO_3161 (O_3161,N_48174,N_48863);
xor UO_3162 (O_3162,N_48562,N_49053);
xnor UO_3163 (O_3163,N_49784,N_48180);
and UO_3164 (O_3164,N_48718,N_48202);
xor UO_3165 (O_3165,N_49612,N_49196);
nor UO_3166 (O_3166,N_48575,N_48225);
xnor UO_3167 (O_3167,N_48573,N_49821);
nor UO_3168 (O_3168,N_48898,N_48244);
nor UO_3169 (O_3169,N_48980,N_48447);
and UO_3170 (O_3170,N_49158,N_48258);
nand UO_3171 (O_3171,N_48168,N_49289);
or UO_3172 (O_3172,N_48856,N_48607);
or UO_3173 (O_3173,N_48265,N_49521);
nand UO_3174 (O_3174,N_48301,N_48421);
or UO_3175 (O_3175,N_49868,N_49069);
xor UO_3176 (O_3176,N_49653,N_49135);
or UO_3177 (O_3177,N_48067,N_49090);
nand UO_3178 (O_3178,N_48959,N_49417);
nand UO_3179 (O_3179,N_48672,N_49076);
nor UO_3180 (O_3180,N_48119,N_49517);
nor UO_3181 (O_3181,N_48044,N_49544);
and UO_3182 (O_3182,N_48665,N_49476);
and UO_3183 (O_3183,N_48159,N_48392);
nand UO_3184 (O_3184,N_48142,N_49628);
nor UO_3185 (O_3185,N_48867,N_48320);
or UO_3186 (O_3186,N_48356,N_48360);
or UO_3187 (O_3187,N_49407,N_48056);
nor UO_3188 (O_3188,N_49285,N_49506);
and UO_3189 (O_3189,N_48206,N_48622);
or UO_3190 (O_3190,N_48731,N_48838);
nand UO_3191 (O_3191,N_48278,N_48114);
nor UO_3192 (O_3192,N_48272,N_48040);
nand UO_3193 (O_3193,N_48871,N_49057);
nand UO_3194 (O_3194,N_48845,N_49955);
and UO_3195 (O_3195,N_49620,N_49682);
xor UO_3196 (O_3196,N_48620,N_49549);
nor UO_3197 (O_3197,N_49345,N_49132);
xnor UO_3198 (O_3198,N_49637,N_49107);
or UO_3199 (O_3199,N_49511,N_49520);
nor UO_3200 (O_3200,N_48405,N_49751);
and UO_3201 (O_3201,N_49862,N_48264);
nor UO_3202 (O_3202,N_48806,N_49257);
nand UO_3203 (O_3203,N_48051,N_49998);
nor UO_3204 (O_3204,N_48027,N_48051);
nand UO_3205 (O_3205,N_49123,N_48764);
nand UO_3206 (O_3206,N_48380,N_48495);
nor UO_3207 (O_3207,N_49540,N_48552);
or UO_3208 (O_3208,N_49662,N_49712);
nand UO_3209 (O_3209,N_49998,N_49811);
and UO_3210 (O_3210,N_49490,N_49141);
or UO_3211 (O_3211,N_48161,N_48181);
xnor UO_3212 (O_3212,N_48528,N_48887);
nor UO_3213 (O_3213,N_49851,N_49357);
or UO_3214 (O_3214,N_48329,N_48881);
xnor UO_3215 (O_3215,N_49719,N_48096);
nand UO_3216 (O_3216,N_49603,N_49955);
nor UO_3217 (O_3217,N_48929,N_49351);
nor UO_3218 (O_3218,N_49580,N_49972);
nor UO_3219 (O_3219,N_49472,N_48359);
nand UO_3220 (O_3220,N_49679,N_49602);
xor UO_3221 (O_3221,N_49041,N_48852);
or UO_3222 (O_3222,N_48788,N_48718);
or UO_3223 (O_3223,N_49569,N_48077);
and UO_3224 (O_3224,N_48434,N_49127);
or UO_3225 (O_3225,N_48009,N_48433);
and UO_3226 (O_3226,N_48071,N_48697);
nand UO_3227 (O_3227,N_49920,N_49705);
and UO_3228 (O_3228,N_49315,N_49929);
and UO_3229 (O_3229,N_49801,N_49401);
xnor UO_3230 (O_3230,N_49701,N_48781);
xnor UO_3231 (O_3231,N_49319,N_48077);
and UO_3232 (O_3232,N_49885,N_48386);
xor UO_3233 (O_3233,N_49147,N_48195);
and UO_3234 (O_3234,N_49020,N_49254);
or UO_3235 (O_3235,N_48671,N_49081);
nor UO_3236 (O_3236,N_49464,N_48549);
xnor UO_3237 (O_3237,N_48863,N_48965);
xor UO_3238 (O_3238,N_49763,N_49907);
xor UO_3239 (O_3239,N_49534,N_48538);
nor UO_3240 (O_3240,N_48426,N_49470);
nor UO_3241 (O_3241,N_49443,N_49475);
nand UO_3242 (O_3242,N_49027,N_48146);
or UO_3243 (O_3243,N_48918,N_48711);
xor UO_3244 (O_3244,N_49748,N_49944);
or UO_3245 (O_3245,N_48775,N_49644);
nand UO_3246 (O_3246,N_48739,N_48180);
nor UO_3247 (O_3247,N_48559,N_48011);
nand UO_3248 (O_3248,N_48409,N_48161);
xnor UO_3249 (O_3249,N_48618,N_48428);
nand UO_3250 (O_3250,N_48159,N_48025);
nand UO_3251 (O_3251,N_48021,N_48187);
nand UO_3252 (O_3252,N_48470,N_48314);
xor UO_3253 (O_3253,N_48244,N_49169);
xnor UO_3254 (O_3254,N_48336,N_48327);
and UO_3255 (O_3255,N_49751,N_48480);
nand UO_3256 (O_3256,N_48439,N_49270);
or UO_3257 (O_3257,N_48367,N_49886);
xnor UO_3258 (O_3258,N_49210,N_49627);
xnor UO_3259 (O_3259,N_48384,N_49601);
nor UO_3260 (O_3260,N_49867,N_48893);
xnor UO_3261 (O_3261,N_49703,N_48168);
nand UO_3262 (O_3262,N_48206,N_49654);
or UO_3263 (O_3263,N_48993,N_49547);
and UO_3264 (O_3264,N_49773,N_49958);
nor UO_3265 (O_3265,N_49281,N_49741);
nor UO_3266 (O_3266,N_49015,N_49500);
xor UO_3267 (O_3267,N_48384,N_48131);
or UO_3268 (O_3268,N_49289,N_49739);
xnor UO_3269 (O_3269,N_49710,N_49171);
nand UO_3270 (O_3270,N_48590,N_49451);
and UO_3271 (O_3271,N_48905,N_49420);
nor UO_3272 (O_3272,N_48923,N_48417);
xnor UO_3273 (O_3273,N_48030,N_48616);
or UO_3274 (O_3274,N_49892,N_48247);
and UO_3275 (O_3275,N_49385,N_48897);
nor UO_3276 (O_3276,N_49951,N_49608);
and UO_3277 (O_3277,N_48547,N_48491);
or UO_3278 (O_3278,N_48977,N_49896);
or UO_3279 (O_3279,N_49335,N_49763);
xor UO_3280 (O_3280,N_48132,N_49717);
nand UO_3281 (O_3281,N_48075,N_49818);
nor UO_3282 (O_3282,N_49011,N_49094);
nor UO_3283 (O_3283,N_48058,N_48337);
and UO_3284 (O_3284,N_48849,N_48710);
or UO_3285 (O_3285,N_49325,N_49679);
or UO_3286 (O_3286,N_48949,N_49691);
and UO_3287 (O_3287,N_49603,N_48487);
xnor UO_3288 (O_3288,N_48736,N_49950);
nand UO_3289 (O_3289,N_48073,N_49253);
or UO_3290 (O_3290,N_49982,N_49345);
nand UO_3291 (O_3291,N_49471,N_48320);
xnor UO_3292 (O_3292,N_48287,N_48930);
nor UO_3293 (O_3293,N_49635,N_49058);
nand UO_3294 (O_3294,N_48934,N_49277);
xor UO_3295 (O_3295,N_48836,N_49278);
nor UO_3296 (O_3296,N_48540,N_49444);
or UO_3297 (O_3297,N_48200,N_48545);
or UO_3298 (O_3298,N_49951,N_48206);
and UO_3299 (O_3299,N_49533,N_48562);
nand UO_3300 (O_3300,N_48566,N_48653);
nor UO_3301 (O_3301,N_49125,N_48533);
nor UO_3302 (O_3302,N_49558,N_49172);
nor UO_3303 (O_3303,N_49938,N_49792);
and UO_3304 (O_3304,N_49315,N_48769);
or UO_3305 (O_3305,N_48854,N_49815);
nand UO_3306 (O_3306,N_49533,N_48834);
nand UO_3307 (O_3307,N_48485,N_49070);
xnor UO_3308 (O_3308,N_49449,N_48942);
nor UO_3309 (O_3309,N_49189,N_48454);
nand UO_3310 (O_3310,N_49433,N_49096);
or UO_3311 (O_3311,N_49800,N_48590);
nor UO_3312 (O_3312,N_49390,N_49803);
nand UO_3313 (O_3313,N_49732,N_49363);
nand UO_3314 (O_3314,N_48360,N_48480);
nor UO_3315 (O_3315,N_49553,N_48055);
nor UO_3316 (O_3316,N_49448,N_49108);
xnor UO_3317 (O_3317,N_49941,N_48457);
or UO_3318 (O_3318,N_48587,N_48822);
xor UO_3319 (O_3319,N_49093,N_49546);
and UO_3320 (O_3320,N_49098,N_49621);
xnor UO_3321 (O_3321,N_48981,N_49192);
xnor UO_3322 (O_3322,N_48817,N_48469);
or UO_3323 (O_3323,N_49148,N_49938);
nand UO_3324 (O_3324,N_48320,N_48532);
nand UO_3325 (O_3325,N_48446,N_48198);
xor UO_3326 (O_3326,N_49146,N_49184);
xor UO_3327 (O_3327,N_48229,N_48555);
and UO_3328 (O_3328,N_48407,N_48977);
and UO_3329 (O_3329,N_49723,N_49076);
nand UO_3330 (O_3330,N_49955,N_48651);
xor UO_3331 (O_3331,N_49074,N_49133);
nor UO_3332 (O_3332,N_49507,N_49690);
nor UO_3333 (O_3333,N_49593,N_48910);
and UO_3334 (O_3334,N_48437,N_48302);
and UO_3335 (O_3335,N_49354,N_48797);
and UO_3336 (O_3336,N_48067,N_48051);
nor UO_3337 (O_3337,N_48823,N_49183);
nor UO_3338 (O_3338,N_48784,N_49484);
nor UO_3339 (O_3339,N_49679,N_48757);
nor UO_3340 (O_3340,N_48836,N_49028);
and UO_3341 (O_3341,N_48521,N_49861);
nand UO_3342 (O_3342,N_49516,N_48567);
nor UO_3343 (O_3343,N_48271,N_49949);
nor UO_3344 (O_3344,N_49582,N_48673);
xnor UO_3345 (O_3345,N_48777,N_49196);
or UO_3346 (O_3346,N_49200,N_49728);
xnor UO_3347 (O_3347,N_49688,N_48389);
nor UO_3348 (O_3348,N_48462,N_48602);
xnor UO_3349 (O_3349,N_48280,N_49666);
nor UO_3350 (O_3350,N_49427,N_48746);
or UO_3351 (O_3351,N_49961,N_49472);
nor UO_3352 (O_3352,N_48898,N_48962);
xnor UO_3353 (O_3353,N_48187,N_49453);
xnor UO_3354 (O_3354,N_48446,N_49548);
nand UO_3355 (O_3355,N_48907,N_48835);
and UO_3356 (O_3356,N_49155,N_49014);
xnor UO_3357 (O_3357,N_48105,N_49140);
and UO_3358 (O_3358,N_48629,N_49369);
or UO_3359 (O_3359,N_48327,N_49791);
and UO_3360 (O_3360,N_48980,N_49960);
nand UO_3361 (O_3361,N_48132,N_48736);
or UO_3362 (O_3362,N_48305,N_49232);
xor UO_3363 (O_3363,N_48758,N_49277);
nor UO_3364 (O_3364,N_48542,N_49315);
nor UO_3365 (O_3365,N_49120,N_48877);
nor UO_3366 (O_3366,N_48096,N_48211);
and UO_3367 (O_3367,N_49647,N_48132);
nand UO_3368 (O_3368,N_48494,N_48725);
nand UO_3369 (O_3369,N_49379,N_49158);
nand UO_3370 (O_3370,N_48480,N_48639);
nor UO_3371 (O_3371,N_48034,N_49254);
nor UO_3372 (O_3372,N_49756,N_49048);
and UO_3373 (O_3373,N_49497,N_48699);
nand UO_3374 (O_3374,N_49030,N_49363);
nand UO_3375 (O_3375,N_48936,N_48137);
xnor UO_3376 (O_3376,N_49429,N_48576);
nor UO_3377 (O_3377,N_48416,N_48428);
or UO_3378 (O_3378,N_49645,N_48523);
nor UO_3379 (O_3379,N_48610,N_49256);
and UO_3380 (O_3380,N_49534,N_49388);
nor UO_3381 (O_3381,N_48406,N_48165);
and UO_3382 (O_3382,N_48901,N_49568);
nor UO_3383 (O_3383,N_49867,N_48878);
nor UO_3384 (O_3384,N_48554,N_49411);
nand UO_3385 (O_3385,N_49694,N_48722);
nand UO_3386 (O_3386,N_49845,N_48554);
nor UO_3387 (O_3387,N_49980,N_49759);
nor UO_3388 (O_3388,N_49652,N_48668);
nor UO_3389 (O_3389,N_48085,N_49883);
or UO_3390 (O_3390,N_48012,N_49686);
nand UO_3391 (O_3391,N_49817,N_48624);
nand UO_3392 (O_3392,N_49048,N_49840);
nor UO_3393 (O_3393,N_48497,N_48764);
and UO_3394 (O_3394,N_48847,N_48269);
nand UO_3395 (O_3395,N_49573,N_49259);
or UO_3396 (O_3396,N_48076,N_49750);
and UO_3397 (O_3397,N_49717,N_49667);
nand UO_3398 (O_3398,N_48852,N_48203);
or UO_3399 (O_3399,N_48843,N_48613);
xor UO_3400 (O_3400,N_48011,N_49113);
nor UO_3401 (O_3401,N_49080,N_48692);
xnor UO_3402 (O_3402,N_49962,N_49598);
or UO_3403 (O_3403,N_48043,N_49316);
or UO_3404 (O_3404,N_49053,N_48546);
or UO_3405 (O_3405,N_49350,N_48808);
nor UO_3406 (O_3406,N_48606,N_49285);
nor UO_3407 (O_3407,N_49693,N_49442);
nor UO_3408 (O_3408,N_49588,N_49071);
nor UO_3409 (O_3409,N_49387,N_49553);
and UO_3410 (O_3410,N_49697,N_49640);
nor UO_3411 (O_3411,N_48144,N_48906);
and UO_3412 (O_3412,N_48210,N_49012);
and UO_3413 (O_3413,N_48446,N_48388);
or UO_3414 (O_3414,N_49947,N_48581);
or UO_3415 (O_3415,N_49739,N_49640);
or UO_3416 (O_3416,N_48374,N_48112);
nor UO_3417 (O_3417,N_48539,N_48514);
nor UO_3418 (O_3418,N_48039,N_48157);
xnor UO_3419 (O_3419,N_49279,N_48701);
nand UO_3420 (O_3420,N_48234,N_49105);
xnor UO_3421 (O_3421,N_48994,N_49246);
nor UO_3422 (O_3422,N_48871,N_49862);
and UO_3423 (O_3423,N_49626,N_48317);
nand UO_3424 (O_3424,N_49304,N_49973);
nand UO_3425 (O_3425,N_48903,N_49027);
xor UO_3426 (O_3426,N_48836,N_48005);
nand UO_3427 (O_3427,N_48308,N_48500);
or UO_3428 (O_3428,N_48390,N_48797);
xnor UO_3429 (O_3429,N_49348,N_48148);
xnor UO_3430 (O_3430,N_49614,N_49720);
or UO_3431 (O_3431,N_49965,N_48107);
and UO_3432 (O_3432,N_48225,N_48687);
and UO_3433 (O_3433,N_49889,N_48490);
or UO_3434 (O_3434,N_48046,N_48258);
and UO_3435 (O_3435,N_48030,N_49224);
and UO_3436 (O_3436,N_49586,N_48242);
and UO_3437 (O_3437,N_48197,N_49124);
and UO_3438 (O_3438,N_49533,N_49778);
nor UO_3439 (O_3439,N_48231,N_49745);
or UO_3440 (O_3440,N_48875,N_49429);
nor UO_3441 (O_3441,N_49810,N_49601);
or UO_3442 (O_3442,N_48903,N_48213);
nand UO_3443 (O_3443,N_48411,N_49865);
nor UO_3444 (O_3444,N_48188,N_48219);
or UO_3445 (O_3445,N_49631,N_49564);
nand UO_3446 (O_3446,N_48550,N_48607);
and UO_3447 (O_3447,N_48726,N_48299);
or UO_3448 (O_3448,N_49664,N_49294);
or UO_3449 (O_3449,N_49739,N_48178);
nor UO_3450 (O_3450,N_48213,N_48474);
or UO_3451 (O_3451,N_49277,N_49271);
or UO_3452 (O_3452,N_48583,N_49718);
or UO_3453 (O_3453,N_49082,N_48080);
nand UO_3454 (O_3454,N_49599,N_49237);
xor UO_3455 (O_3455,N_49576,N_48625);
xnor UO_3456 (O_3456,N_48261,N_48248);
xnor UO_3457 (O_3457,N_48214,N_48420);
nor UO_3458 (O_3458,N_48377,N_48506);
or UO_3459 (O_3459,N_49567,N_48542);
and UO_3460 (O_3460,N_48422,N_48940);
or UO_3461 (O_3461,N_48773,N_49930);
and UO_3462 (O_3462,N_48125,N_49198);
or UO_3463 (O_3463,N_49344,N_48822);
nand UO_3464 (O_3464,N_49803,N_48695);
and UO_3465 (O_3465,N_48171,N_49640);
and UO_3466 (O_3466,N_48504,N_49042);
xor UO_3467 (O_3467,N_49537,N_49928);
nor UO_3468 (O_3468,N_48898,N_48882);
or UO_3469 (O_3469,N_48152,N_48012);
and UO_3470 (O_3470,N_49834,N_48579);
and UO_3471 (O_3471,N_49613,N_49340);
nand UO_3472 (O_3472,N_49777,N_49351);
or UO_3473 (O_3473,N_49256,N_48144);
and UO_3474 (O_3474,N_48730,N_49904);
or UO_3475 (O_3475,N_48532,N_49224);
xnor UO_3476 (O_3476,N_49370,N_48801);
and UO_3477 (O_3477,N_49960,N_49188);
nand UO_3478 (O_3478,N_48894,N_49304);
xnor UO_3479 (O_3479,N_49974,N_49296);
or UO_3480 (O_3480,N_49813,N_48117);
nor UO_3481 (O_3481,N_49273,N_48306);
nand UO_3482 (O_3482,N_48504,N_49819);
or UO_3483 (O_3483,N_49821,N_48138);
or UO_3484 (O_3484,N_48320,N_49683);
or UO_3485 (O_3485,N_49050,N_48356);
or UO_3486 (O_3486,N_48726,N_48346);
or UO_3487 (O_3487,N_48833,N_49993);
nand UO_3488 (O_3488,N_49049,N_49173);
and UO_3489 (O_3489,N_48654,N_49413);
and UO_3490 (O_3490,N_49928,N_48926);
and UO_3491 (O_3491,N_49565,N_49834);
and UO_3492 (O_3492,N_48262,N_49329);
or UO_3493 (O_3493,N_48802,N_48551);
and UO_3494 (O_3494,N_48518,N_48827);
nor UO_3495 (O_3495,N_48486,N_49005);
or UO_3496 (O_3496,N_49662,N_49610);
nand UO_3497 (O_3497,N_49946,N_48661);
and UO_3498 (O_3498,N_48608,N_48043);
nor UO_3499 (O_3499,N_48371,N_49717);
nand UO_3500 (O_3500,N_48788,N_49182);
nor UO_3501 (O_3501,N_48961,N_48514);
or UO_3502 (O_3502,N_49564,N_48921);
or UO_3503 (O_3503,N_48111,N_49558);
nor UO_3504 (O_3504,N_49270,N_49169);
and UO_3505 (O_3505,N_49161,N_48232);
nor UO_3506 (O_3506,N_48821,N_49645);
nor UO_3507 (O_3507,N_48486,N_48109);
and UO_3508 (O_3508,N_48040,N_48195);
nand UO_3509 (O_3509,N_48411,N_48249);
nor UO_3510 (O_3510,N_48402,N_49348);
xnor UO_3511 (O_3511,N_48900,N_48464);
nor UO_3512 (O_3512,N_48218,N_48737);
or UO_3513 (O_3513,N_48525,N_49824);
and UO_3514 (O_3514,N_48720,N_48340);
nor UO_3515 (O_3515,N_49415,N_48249);
and UO_3516 (O_3516,N_49766,N_49493);
nand UO_3517 (O_3517,N_48413,N_48342);
xnor UO_3518 (O_3518,N_48804,N_48555);
nor UO_3519 (O_3519,N_49304,N_49969);
xnor UO_3520 (O_3520,N_49071,N_49852);
or UO_3521 (O_3521,N_48203,N_48951);
nand UO_3522 (O_3522,N_48465,N_48328);
nor UO_3523 (O_3523,N_48237,N_49012);
nor UO_3524 (O_3524,N_48875,N_49023);
xor UO_3525 (O_3525,N_49702,N_48554);
or UO_3526 (O_3526,N_48856,N_48842);
and UO_3527 (O_3527,N_48560,N_48348);
nand UO_3528 (O_3528,N_48089,N_48287);
nor UO_3529 (O_3529,N_49629,N_48609);
nand UO_3530 (O_3530,N_49240,N_49999);
xor UO_3531 (O_3531,N_48904,N_49763);
nand UO_3532 (O_3532,N_48246,N_49025);
and UO_3533 (O_3533,N_48707,N_48019);
or UO_3534 (O_3534,N_48554,N_49255);
xnor UO_3535 (O_3535,N_49730,N_48826);
nand UO_3536 (O_3536,N_48523,N_49336);
xnor UO_3537 (O_3537,N_49103,N_49916);
and UO_3538 (O_3538,N_49033,N_49706);
or UO_3539 (O_3539,N_49394,N_49594);
and UO_3540 (O_3540,N_48388,N_48871);
and UO_3541 (O_3541,N_49971,N_48263);
or UO_3542 (O_3542,N_48598,N_48725);
xor UO_3543 (O_3543,N_48239,N_48558);
xnor UO_3544 (O_3544,N_49670,N_49590);
nand UO_3545 (O_3545,N_48398,N_49969);
xnor UO_3546 (O_3546,N_48851,N_48050);
nand UO_3547 (O_3547,N_49423,N_49083);
and UO_3548 (O_3548,N_49091,N_49141);
xnor UO_3549 (O_3549,N_48041,N_48588);
and UO_3550 (O_3550,N_48359,N_48699);
and UO_3551 (O_3551,N_48581,N_48323);
and UO_3552 (O_3552,N_48506,N_49735);
nand UO_3553 (O_3553,N_48243,N_49480);
and UO_3554 (O_3554,N_48769,N_48833);
xnor UO_3555 (O_3555,N_49486,N_49053);
nand UO_3556 (O_3556,N_48594,N_48023);
xor UO_3557 (O_3557,N_49331,N_49374);
nand UO_3558 (O_3558,N_48287,N_49732);
xor UO_3559 (O_3559,N_48457,N_48528);
nand UO_3560 (O_3560,N_48623,N_48463);
and UO_3561 (O_3561,N_48018,N_48827);
nand UO_3562 (O_3562,N_49128,N_48837);
nand UO_3563 (O_3563,N_48332,N_48686);
or UO_3564 (O_3564,N_48248,N_49326);
or UO_3565 (O_3565,N_48105,N_49718);
and UO_3566 (O_3566,N_49045,N_49077);
nor UO_3567 (O_3567,N_48984,N_48849);
xor UO_3568 (O_3568,N_48322,N_49898);
xor UO_3569 (O_3569,N_48853,N_49365);
xnor UO_3570 (O_3570,N_49606,N_48456);
or UO_3571 (O_3571,N_48343,N_48119);
or UO_3572 (O_3572,N_49236,N_49812);
nor UO_3573 (O_3573,N_49516,N_49315);
nand UO_3574 (O_3574,N_48350,N_49466);
and UO_3575 (O_3575,N_48693,N_48688);
or UO_3576 (O_3576,N_48201,N_49967);
nand UO_3577 (O_3577,N_48654,N_48048);
xnor UO_3578 (O_3578,N_48709,N_48677);
nand UO_3579 (O_3579,N_48629,N_49371);
or UO_3580 (O_3580,N_48322,N_48282);
nor UO_3581 (O_3581,N_48411,N_48499);
nor UO_3582 (O_3582,N_48801,N_48604);
or UO_3583 (O_3583,N_49060,N_48232);
nand UO_3584 (O_3584,N_49279,N_48171);
and UO_3585 (O_3585,N_49865,N_48733);
or UO_3586 (O_3586,N_48125,N_49096);
and UO_3587 (O_3587,N_48897,N_48678);
nand UO_3588 (O_3588,N_48946,N_49404);
nand UO_3589 (O_3589,N_49117,N_48327);
or UO_3590 (O_3590,N_49510,N_48037);
xor UO_3591 (O_3591,N_48099,N_49136);
nand UO_3592 (O_3592,N_48575,N_49197);
nand UO_3593 (O_3593,N_49206,N_49825);
and UO_3594 (O_3594,N_48948,N_48647);
and UO_3595 (O_3595,N_48153,N_48398);
or UO_3596 (O_3596,N_49453,N_48165);
nand UO_3597 (O_3597,N_49620,N_49830);
nand UO_3598 (O_3598,N_49970,N_49782);
nor UO_3599 (O_3599,N_48429,N_49909);
or UO_3600 (O_3600,N_48733,N_48863);
nand UO_3601 (O_3601,N_48697,N_49665);
or UO_3602 (O_3602,N_48524,N_48835);
or UO_3603 (O_3603,N_49468,N_49338);
nand UO_3604 (O_3604,N_48415,N_49955);
and UO_3605 (O_3605,N_48586,N_49859);
and UO_3606 (O_3606,N_48787,N_49151);
or UO_3607 (O_3607,N_48178,N_49875);
or UO_3608 (O_3608,N_49025,N_49483);
or UO_3609 (O_3609,N_48737,N_49095);
nand UO_3610 (O_3610,N_48223,N_49967);
or UO_3611 (O_3611,N_48019,N_48067);
or UO_3612 (O_3612,N_48840,N_48011);
nor UO_3613 (O_3613,N_48677,N_49700);
xnor UO_3614 (O_3614,N_48630,N_49392);
nor UO_3615 (O_3615,N_48852,N_49063);
and UO_3616 (O_3616,N_48280,N_48911);
and UO_3617 (O_3617,N_48259,N_48430);
and UO_3618 (O_3618,N_48677,N_49596);
nor UO_3619 (O_3619,N_48023,N_49878);
nor UO_3620 (O_3620,N_48876,N_48209);
nand UO_3621 (O_3621,N_49988,N_48078);
nor UO_3622 (O_3622,N_49363,N_48686);
xnor UO_3623 (O_3623,N_48548,N_49020);
or UO_3624 (O_3624,N_49161,N_49611);
and UO_3625 (O_3625,N_49006,N_49790);
or UO_3626 (O_3626,N_48140,N_48541);
or UO_3627 (O_3627,N_49156,N_49198);
nand UO_3628 (O_3628,N_49445,N_49578);
nand UO_3629 (O_3629,N_48785,N_48276);
or UO_3630 (O_3630,N_49869,N_49337);
and UO_3631 (O_3631,N_49019,N_49159);
nand UO_3632 (O_3632,N_48565,N_49288);
or UO_3633 (O_3633,N_48002,N_49178);
or UO_3634 (O_3634,N_48506,N_49576);
nand UO_3635 (O_3635,N_49122,N_48424);
and UO_3636 (O_3636,N_48735,N_49141);
nand UO_3637 (O_3637,N_48113,N_49166);
nand UO_3638 (O_3638,N_49412,N_49167);
nand UO_3639 (O_3639,N_49050,N_48593);
xnor UO_3640 (O_3640,N_48873,N_48776);
and UO_3641 (O_3641,N_49296,N_48964);
nor UO_3642 (O_3642,N_48849,N_48892);
or UO_3643 (O_3643,N_49364,N_48794);
nor UO_3644 (O_3644,N_49312,N_49618);
xor UO_3645 (O_3645,N_48795,N_48970);
nand UO_3646 (O_3646,N_48633,N_48355);
nand UO_3647 (O_3647,N_48069,N_49430);
xor UO_3648 (O_3648,N_49899,N_49415);
nor UO_3649 (O_3649,N_49841,N_49039);
nand UO_3650 (O_3650,N_48297,N_49943);
nor UO_3651 (O_3651,N_49205,N_48696);
nand UO_3652 (O_3652,N_49440,N_49135);
xor UO_3653 (O_3653,N_49462,N_48049);
or UO_3654 (O_3654,N_49579,N_49284);
and UO_3655 (O_3655,N_49383,N_49304);
or UO_3656 (O_3656,N_49949,N_48046);
or UO_3657 (O_3657,N_48911,N_49997);
or UO_3658 (O_3658,N_48074,N_49393);
or UO_3659 (O_3659,N_48472,N_48830);
xnor UO_3660 (O_3660,N_48384,N_49783);
xor UO_3661 (O_3661,N_48584,N_48233);
nand UO_3662 (O_3662,N_49736,N_49842);
and UO_3663 (O_3663,N_48681,N_49531);
nand UO_3664 (O_3664,N_48577,N_48927);
nand UO_3665 (O_3665,N_48831,N_48434);
nand UO_3666 (O_3666,N_48104,N_49990);
nand UO_3667 (O_3667,N_49222,N_48207);
nand UO_3668 (O_3668,N_49518,N_48806);
and UO_3669 (O_3669,N_48057,N_49408);
and UO_3670 (O_3670,N_49031,N_48729);
nor UO_3671 (O_3671,N_49992,N_49759);
xnor UO_3672 (O_3672,N_48124,N_49809);
xor UO_3673 (O_3673,N_49561,N_48199);
xor UO_3674 (O_3674,N_49112,N_48661);
and UO_3675 (O_3675,N_49022,N_48708);
nor UO_3676 (O_3676,N_49420,N_49768);
xnor UO_3677 (O_3677,N_48164,N_49485);
xor UO_3678 (O_3678,N_49945,N_48421);
or UO_3679 (O_3679,N_48509,N_49427);
nor UO_3680 (O_3680,N_48896,N_49033);
nand UO_3681 (O_3681,N_48434,N_49350);
nor UO_3682 (O_3682,N_48004,N_48814);
nand UO_3683 (O_3683,N_49225,N_49292);
nor UO_3684 (O_3684,N_49158,N_48587);
nand UO_3685 (O_3685,N_48845,N_49444);
or UO_3686 (O_3686,N_49531,N_49163);
nand UO_3687 (O_3687,N_48947,N_48485);
or UO_3688 (O_3688,N_48575,N_48903);
xnor UO_3689 (O_3689,N_49301,N_49228);
or UO_3690 (O_3690,N_48494,N_48322);
nor UO_3691 (O_3691,N_49483,N_49833);
and UO_3692 (O_3692,N_48862,N_49057);
or UO_3693 (O_3693,N_48819,N_48361);
nand UO_3694 (O_3694,N_49810,N_49052);
or UO_3695 (O_3695,N_48357,N_48382);
or UO_3696 (O_3696,N_48767,N_49164);
xnor UO_3697 (O_3697,N_48115,N_48381);
and UO_3698 (O_3698,N_49334,N_49648);
nand UO_3699 (O_3699,N_49863,N_48733);
xor UO_3700 (O_3700,N_48686,N_48440);
nor UO_3701 (O_3701,N_49048,N_48895);
xor UO_3702 (O_3702,N_49045,N_49868);
and UO_3703 (O_3703,N_48010,N_48115);
and UO_3704 (O_3704,N_49694,N_48174);
or UO_3705 (O_3705,N_49883,N_49521);
nand UO_3706 (O_3706,N_48593,N_49017);
or UO_3707 (O_3707,N_49369,N_49759);
nor UO_3708 (O_3708,N_48321,N_49674);
xnor UO_3709 (O_3709,N_49135,N_48532);
xor UO_3710 (O_3710,N_48555,N_48206);
xor UO_3711 (O_3711,N_48837,N_49195);
or UO_3712 (O_3712,N_48533,N_49330);
and UO_3713 (O_3713,N_48846,N_49953);
or UO_3714 (O_3714,N_48832,N_48452);
nor UO_3715 (O_3715,N_48925,N_49576);
nor UO_3716 (O_3716,N_48293,N_48622);
xor UO_3717 (O_3717,N_49314,N_49205);
and UO_3718 (O_3718,N_48107,N_48088);
xnor UO_3719 (O_3719,N_49714,N_48241);
xor UO_3720 (O_3720,N_49637,N_48618);
and UO_3721 (O_3721,N_48436,N_48789);
nor UO_3722 (O_3722,N_49261,N_49872);
xnor UO_3723 (O_3723,N_48721,N_49876);
nor UO_3724 (O_3724,N_49558,N_49157);
and UO_3725 (O_3725,N_49015,N_49459);
or UO_3726 (O_3726,N_48241,N_48996);
or UO_3727 (O_3727,N_49863,N_48131);
xnor UO_3728 (O_3728,N_49512,N_48189);
xor UO_3729 (O_3729,N_48936,N_49430);
nand UO_3730 (O_3730,N_49640,N_48830);
nor UO_3731 (O_3731,N_48627,N_48202);
or UO_3732 (O_3732,N_48868,N_48741);
or UO_3733 (O_3733,N_49362,N_48284);
nand UO_3734 (O_3734,N_48865,N_48272);
nand UO_3735 (O_3735,N_48860,N_49961);
xor UO_3736 (O_3736,N_48118,N_49928);
and UO_3737 (O_3737,N_49993,N_49144);
xnor UO_3738 (O_3738,N_49703,N_48646);
and UO_3739 (O_3739,N_48204,N_49966);
nand UO_3740 (O_3740,N_49721,N_48513);
or UO_3741 (O_3741,N_48653,N_48850);
and UO_3742 (O_3742,N_48193,N_49600);
nor UO_3743 (O_3743,N_48705,N_49206);
nor UO_3744 (O_3744,N_49448,N_48217);
xor UO_3745 (O_3745,N_49850,N_49536);
nand UO_3746 (O_3746,N_48160,N_48344);
and UO_3747 (O_3747,N_49396,N_48630);
and UO_3748 (O_3748,N_49132,N_49826);
or UO_3749 (O_3749,N_48280,N_48348);
xnor UO_3750 (O_3750,N_49624,N_49363);
nand UO_3751 (O_3751,N_49149,N_49025);
nand UO_3752 (O_3752,N_48856,N_49568);
and UO_3753 (O_3753,N_49831,N_49248);
xnor UO_3754 (O_3754,N_48736,N_48403);
or UO_3755 (O_3755,N_48126,N_49168);
or UO_3756 (O_3756,N_49827,N_49288);
and UO_3757 (O_3757,N_48899,N_48432);
or UO_3758 (O_3758,N_49278,N_49700);
and UO_3759 (O_3759,N_48607,N_49401);
nand UO_3760 (O_3760,N_49032,N_49191);
and UO_3761 (O_3761,N_49656,N_48992);
and UO_3762 (O_3762,N_48518,N_49952);
or UO_3763 (O_3763,N_48376,N_49198);
nor UO_3764 (O_3764,N_49678,N_48560);
nor UO_3765 (O_3765,N_49590,N_48774);
nor UO_3766 (O_3766,N_48259,N_49924);
nand UO_3767 (O_3767,N_48640,N_48413);
xor UO_3768 (O_3768,N_49839,N_49228);
and UO_3769 (O_3769,N_49950,N_49333);
nand UO_3770 (O_3770,N_49937,N_49581);
or UO_3771 (O_3771,N_48198,N_48202);
nand UO_3772 (O_3772,N_48308,N_49101);
or UO_3773 (O_3773,N_49844,N_48612);
and UO_3774 (O_3774,N_48254,N_48705);
xor UO_3775 (O_3775,N_48700,N_49489);
and UO_3776 (O_3776,N_49295,N_48709);
and UO_3777 (O_3777,N_48876,N_49248);
nand UO_3778 (O_3778,N_49216,N_49059);
nand UO_3779 (O_3779,N_48699,N_49893);
and UO_3780 (O_3780,N_48286,N_48756);
nand UO_3781 (O_3781,N_48168,N_49266);
nor UO_3782 (O_3782,N_48177,N_48001);
nand UO_3783 (O_3783,N_49826,N_49422);
nor UO_3784 (O_3784,N_48656,N_49032);
or UO_3785 (O_3785,N_49905,N_48211);
and UO_3786 (O_3786,N_48553,N_49640);
xor UO_3787 (O_3787,N_48925,N_48093);
xor UO_3788 (O_3788,N_49116,N_49025);
and UO_3789 (O_3789,N_48328,N_48957);
nand UO_3790 (O_3790,N_48819,N_49943);
and UO_3791 (O_3791,N_49960,N_48689);
nor UO_3792 (O_3792,N_49908,N_48862);
or UO_3793 (O_3793,N_49015,N_48483);
nor UO_3794 (O_3794,N_48506,N_49310);
nor UO_3795 (O_3795,N_48869,N_48922);
nor UO_3796 (O_3796,N_49872,N_48698);
nor UO_3797 (O_3797,N_49255,N_49904);
nand UO_3798 (O_3798,N_49969,N_49854);
or UO_3799 (O_3799,N_48009,N_48312);
or UO_3800 (O_3800,N_48846,N_48929);
nand UO_3801 (O_3801,N_48008,N_48599);
nand UO_3802 (O_3802,N_48540,N_48948);
nor UO_3803 (O_3803,N_48915,N_48680);
xnor UO_3804 (O_3804,N_49821,N_48341);
nand UO_3805 (O_3805,N_49040,N_48017);
nand UO_3806 (O_3806,N_49573,N_49587);
nand UO_3807 (O_3807,N_49043,N_48260);
nor UO_3808 (O_3808,N_49709,N_49420);
and UO_3809 (O_3809,N_49907,N_49616);
or UO_3810 (O_3810,N_49048,N_48478);
or UO_3811 (O_3811,N_48131,N_49203);
nor UO_3812 (O_3812,N_48800,N_48329);
nor UO_3813 (O_3813,N_48401,N_48099);
xor UO_3814 (O_3814,N_48907,N_48929);
and UO_3815 (O_3815,N_49940,N_49907);
nand UO_3816 (O_3816,N_48083,N_48330);
and UO_3817 (O_3817,N_49396,N_49462);
nand UO_3818 (O_3818,N_48419,N_49911);
nor UO_3819 (O_3819,N_49153,N_48461);
xor UO_3820 (O_3820,N_48277,N_49101);
and UO_3821 (O_3821,N_49131,N_49983);
nor UO_3822 (O_3822,N_48761,N_49685);
and UO_3823 (O_3823,N_49558,N_49551);
nand UO_3824 (O_3824,N_48309,N_48859);
nor UO_3825 (O_3825,N_49972,N_48927);
and UO_3826 (O_3826,N_48833,N_49424);
nor UO_3827 (O_3827,N_48220,N_49815);
or UO_3828 (O_3828,N_49236,N_48475);
xnor UO_3829 (O_3829,N_48472,N_48750);
or UO_3830 (O_3830,N_49073,N_49635);
or UO_3831 (O_3831,N_48546,N_48599);
xnor UO_3832 (O_3832,N_48998,N_48477);
and UO_3833 (O_3833,N_49381,N_48364);
nor UO_3834 (O_3834,N_49543,N_48933);
or UO_3835 (O_3835,N_49930,N_49023);
xor UO_3836 (O_3836,N_49097,N_49534);
and UO_3837 (O_3837,N_49953,N_48157);
nor UO_3838 (O_3838,N_48538,N_49160);
and UO_3839 (O_3839,N_49074,N_49756);
xor UO_3840 (O_3840,N_48706,N_49401);
nand UO_3841 (O_3841,N_48620,N_48294);
nand UO_3842 (O_3842,N_49582,N_49120);
or UO_3843 (O_3843,N_48478,N_48766);
and UO_3844 (O_3844,N_49356,N_48521);
nand UO_3845 (O_3845,N_48265,N_49018);
and UO_3846 (O_3846,N_49129,N_48173);
or UO_3847 (O_3847,N_48931,N_49023);
xnor UO_3848 (O_3848,N_49250,N_48695);
and UO_3849 (O_3849,N_49133,N_48635);
nor UO_3850 (O_3850,N_48684,N_49051);
xnor UO_3851 (O_3851,N_48633,N_49979);
nor UO_3852 (O_3852,N_49051,N_48542);
nand UO_3853 (O_3853,N_48819,N_49674);
xnor UO_3854 (O_3854,N_48148,N_48014);
or UO_3855 (O_3855,N_49668,N_49978);
nand UO_3856 (O_3856,N_48857,N_49962);
or UO_3857 (O_3857,N_49517,N_49887);
or UO_3858 (O_3858,N_49147,N_49052);
or UO_3859 (O_3859,N_48785,N_49586);
nor UO_3860 (O_3860,N_49837,N_49205);
and UO_3861 (O_3861,N_49406,N_48359);
and UO_3862 (O_3862,N_49239,N_48683);
nand UO_3863 (O_3863,N_48045,N_49615);
nand UO_3864 (O_3864,N_49963,N_48864);
or UO_3865 (O_3865,N_49422,N_49360);
xor UO_3866 (O_3866,N_48160,N_48803);
nand UO_3867 (O_3867,N_49709,N_48455);
xnor UO_3868 (O_3868,N_49255,N_48456);
nor UO_3869 (O_3869,N_48894,N_49220);
or UO_3870 (O_3870,N_48637,N_48343);
nor UO_3871 (O_3871,N_49543,N_48606);
xnor UO_3872 (O_3872,N_49963,N_48322);
nand UO_3873 (O_3873,N_48683,N_49761);
or UO_3874 (O_3874,N_49360,N_48475);
xor UO_3875 (O_3875,N_48344,N_49024);
nand UO_3876 (O_3876,N_49134,N_48650);
or UO_3877 (O_3877,N_49304,N_49376);
xor UO_3878 (O_3878,N_49859,N_48206);
or UO_3879 (O_3879,N_49357,N_49820);
and UO_3880 (O_3880,N_49662,N_49413);
xnor UO_3881 (O_3881,N_48012,N_48378);
xnor UO_3882 (O_3882,N_49855,N_48339);
nor UO_3883 (O_3883,N_49539,N_49342);
and UO_3884 (O_3884,N_49902,N_49774);
nor UO_3885 (O_3885,N_49783,N_49815);
xor UO_3886 (O_3886,N_49189,N_48135);
nand UO_3887 (O_3887,N_48092,N_48060);
and UO_3888 (O_3888,N_49311,N_49660);
or UO_3889 (O_3889,N_48745,N_48566);
xnor UO_3890 (O_3890,N_49271,N_49612);
nand UO_3891 (O_3891,N_49855,N_49006);
and UO_3892 (O_3892,N_49587,N_49754);
xnor UO_3893 (O_3893,N_48458,N_49783);
nand UO_3894 (O_3894,N_49045,N_48266);
nand UO_3895 (O_3895,N_49462,N_48035);
and UO_3896 (O_3896,N_48506,N_48189);
nand UO_3897 (O_3897,N_48291,N_49611);
nor UO_3898 (O_3898,N_49708,N_48427);
and UO_3899 (O_3899,N_48464,N_48650);
nor UO_3900 (O_3900,N_48539,N_48322);
xor UO_3901 (O_3901,N_49402,N_48710);
or UO_3902 (O_3902,N_48727,N_49612);
or UO_3903 (O_3903,N_48207,N_49174);
or UO_3904 (O_3904,N_49209,N_48643);
nand UO_3905 (O_3905,N_49777,N_49409);
or UO_3906 (O_3906,N_49953,N_49729);
nor UO_3907 (O_3907,N_49465,N_49058);
nand UO_3908 (O_3908,N_48481,N_48498);
xnor UO_3909 (O_3909,N_48667,N_49051);
or UO_3910 (O_3910,N_49573,N_48724);
nand UO_3911 (O_3911,N_48369,N_48403);
xor UO_3912 (O_3912,N_49478,N_49344);
and UO_3913 (O_3913,N_49532,N_49017);
or UO_3914 (O_3914,N_48141,N_48829);
nand UO_3915 (O_3915,N_48514,N_49455);
and UO_3916 (O_3916,N_49499,N_49759);
xnor UO_3917 (O_3917,N_48453,N_49299);
nor UO_3918 (O_3918,N_48930,N_48073);
xnor UO_3919 (O_3919,N_49457,N_49373);
and UO_3920 (O_3920,N_49099,N_48138);
nand UO_3921 (O_3921,N_49587,N_48648);
nand UO_3922 (O_3922,N_49961,N_48915);
or UO_3923 (O_3923,N_48841,N_49096);
xor UO_3924 (O_3924,N_49964,N_49890);
nor UO_3925 (O_3925,N_49356,N_49375);
and UO_3926 (O_3926,N_49480,N_48761);
nor UO_3927 (O_3927,N_48424,N_48402);
and UO_3928 (O_3928,N_48161,N_48285);
xor UO_3929 (O_3929,N_48003,N_48119);
or UO_3930 (O_3930,N_48934,N_48513);
or UO_3931 (O_3931,N_48876,N_48011);
nand UO_3932 (O_3932,N_48903,N_49430);
or UO_3933 (O_3933,N_49930,N_48750);
or UO_3934 (O_3934,N_49098,N_49941);
xor UO_3935 (O_3935,N_49789,N_49275);
or UO_3936 (O_3936,N_48465,N_48347);
and UO_3937 (O_3937,N_49297,N_49075);
or UO_3938 (O_3938,N_49746,N_49327);
nor UO_3939 (O_3939,N_49981,N_49520);
nand UO_3940 (O_3940,N_48988,N_49859);
and UO_3941 (O_3941,N_49683,N_48666);
nand UO_3942 (O_3942,N_49801,N_49929);
or UO_3943 (O_3943,N_49540,N_48011);
and UO_3944 (O_3944,N_49099,N_49786);
xnor UO_3945 (O_3945,N_48796,N_49016);
nor UO_3946 (O_3946,N_48220,N_48095);
or UO_3947 (O_3947,N_49245,N_49640);
xnor UO_3948 (O_3948,N_49889,N_48743);
nand UO_3949 (O_3949,N_49801,N_48509);
and UO_3950 (O_3950,N_49181,N_49593);
xor UO_3951 (O_3951,N_49703,N_49135);
and UO_3952 (O_3952,N_48084,N_49412);
nand UO_3953 (O_3953,N_49751,N_48695);
nor UO_3954 (O_3954,N_48819,N_48801);
and UO_3955 (O_3955,N_48200,N_49933);
or UO_3956 (O_3956,N_49261,N_49926);
and UO_3957 (O_3957,N_49419,N_49215);
and UO_3958 (O_3958,N_48956,N_48026);
nand UO_3959 (O_3959,N_48045,N_49646);
and UO_3960 (O_3960,N_48210,N_48451);
xor UO_3961 (O_3961,N_48376,N_48895);
nor UO_3962 (O_3962,N_49786,N_48401);
nand UO_3963 (O_3963,N_49978,N_48423);
nor UO_3964 (O_3964,N_49037,N_48074);
and UO_3965 (O_3965,N_49335,N_48900);
and UO_3966 (O_3966,N_49526,N_49050);
or UO_3967 (O_3967,N_49855,N_48195);
xnor UO_3968 (O_3968,N_49625,N_49838);
and UO_3969 (O_3969,N_48168,N_49546);
or UO_3970 (O_3970,N_49161,N_49726);
xor UO_3971 (O_3971,N_49688,N_48690);
and UO_3972 (O_3972,N_48005,N_49316);
nand UO_3973 (O_3973,N_49663,N_49435);
nor UO_3974 (O_3974,N_48731,N_48686);
and UO_3975 (O_3975,N_48048,N_48116);
nor UO_3976 (O_3976,N_49501,N_48387);
nand UO_3977 (O_3977,N_48142,N_48507);
nor UO_3978 (O_3978,N_49491,N_49147);
or UO_3979 (O_3979,N_49900,N_49950);
and UO_3980 (O_3980,N_48464,N_49783);
or UO_3981 (O_3981,N_49567,N_49600);
nor UO_3982 (O_3982,N_48009,N_49044);
or UO_3983 (O_3983,N_48520,N_48906);
and UO_3984 (O_3984,N_48207,N_49252);
xnor UO_3985 (O_3985,N_49285,N_48827);
and UO_3986 (O_3986,N_49516,N_48578);
nor UO_3987 (O_3987,N_49531,N_49712);
or UO_3988 (O_3988,N_48799,N_48327);
or UO_3989 (O_3989,N_49738,N_49058);
and UO_3990 (O_3990,N_48651,N_48503);
xnor UO_3991 (O_3991,N_49507,N_48925);
and UO_3992 (O_3992,N_49743,N_48582);
nor UO_3993 (O_3993,N_49354,N_48887);
xnor UO_3994 (O_3994,N_48073,N_49505);
or UO_3995 (O_3995,N_49451,N_49374);
nand UO_3996 (O_3996,N_48034,N_49583);
nor UO_3997 (O_3997,N_49523,N_49459);
and UO_3998 (O_3998,N_48343,N_49943);
nor UO_3999 (O_3999,N_48185,N_49038);
and UO_4000 (O_4000,N_48639,N_49643);
and UO_4001 (O_4001,N_48964,N_48679);
nor UO_4002 (O_4002,N_49196,N_48499);
nor UO_4003 (O_4003,N_48420,N_49388);
and UO_4004 (O_4004,N_49915,N_49099);
xor UO_4005 (O_4005,N_48677,N_49355);
nor UO_4006 (O_4006,N_48046,N_49353);
or UO_4007 (O_4007,N_48375,N_49242);
and UO_4008 (O_4008,N_49555,N_49969);
and UO_4009 (O_4009,N_49710,N_48677);
nand UO_4010 (O_4010,N_49928,N_48748);
and UO_4011 (O_4011,N_48034,N_49879);
or UO_4012 (O_4012,N_48981,N_48512);
nor UO_4013 (O_4013,N_48137,N_49789);
nor UO_4014 (O_4014,N_48532,N_49018);
nand UO_4015 (O_4015,N_49243,N_49239);
and UO_4016 (O_4016,N_49516,N_49309);
nor UO_4017 (O_4017,N_48833,N_49359);
nor UO_4018 (O_4018,N_48776,N_48681);
or UO_4019 (O_4019,N_49640,N_49178);
nor UO_4020 (O_4020,N_48442,N_49321);
nor UO_4021 (O_4021,N_48585,N_49749);
xnor UO_4022 (O_4022,N_48386,N_49460);
and UO_4023 (O_4023,N_49929,N_48840);
xnor UO_4024 (O_4024,N_48474,N_49293);
nand UO_4025 (O_4025,N_48050,N_48107);
and UO_4026 (O_4026,N_49915,N_48303);
nor UO_4027 (O_4027,N_48919,N_49194);
nand UO_4028 (O_4028,N_48719,N_49013);
or UO_4029 (O_4029,N_49527,N_49806);
or UO_4030 (O_4030,N_48145,N_48424);
nand UO_4031 (O_4031,N_48586,N_49617);
nor UO_4032 (O_4032,N_49460,N_49648);
nor UO_4033 (O_4033,N_48060,N_48826);
xnor UO_4034 (O_4034,N_49150,N_48535);
or UO_4035 (O_4035,N_48685,N_49882);
or UO_4036 (O_4036,N_48934,N_49143);
xor UO_4037 (O_4037,N_49991,N_48890);
nand UO_4038 (O_4038,N_48964,N_49214);
nor UO_4039 (O_4039,N_49330,N_49082);
or UO_4040 (O_4040,N_48086,N_49573);
xor UO_4041 (O_4041,N_49890,N_49127);
or UO_4042 (O_4042,N_48652,N_49408);
nor UO_4043 (O_4043,N_48660,N_49953);
xor UO_4044 (O_4044,N_48955,N_49265);
xnor UO_4045 (O_4045,N_49353,N_48674);
or UO_4046 (O_4046,N_49490,N_48267);
and UO_4047 (O_4047,N_49424,N_49160);
nor UO_4048 (O_4048,N_49214,N_48395);
or UO_4049 (O_4049,N_49610,N_48217);
xnor UO_4050 (O_4050,N_48642,N_49132);
xor UO_4051 (O_4051,N_49821,N_49348);
or UO_4052 (O_4052,N_49991,N_49965);
nor UO_4053 (O_4053,N_48184,N_49940);
and UO_4054 (O_4054,N_48177,N_49799);
or UO_4055 (O_4055,N_49850,N_49619);
nand UO_4056 (O_4056,N_48499,N_48888);
or UO_4057 (O_4057,N_48514,N_48241);
nor UO_4058 (O_4058,N_48871,N_48993);
nor UO_4059 (O_4059,N_49256,N_49506);
nor UO_4060 (O_4060,N_48913,N_48126);
or UO_4061 (O_4061,N_49900,N_48329);
xnor UO_4062 (O_4062,N_49446,N_48620);
nand UO_4063 (O_4063,N_48508,N_49731);
nand UO_4064 (O_4064,N_48724,N_49313);
or UO_4065 (O_4065,N_49176,N_48661);
and UO_4066 (O_4066,N_49666,N_48449);
or UO_4067 (O_4067,N_49703,N_49946);
nor UO_4068 (O_4068,N_48423,N_48101);
xnor UO_4069 (O_4069,N_48291,N_48686);
and UO_4070 (O_4070,N_49119,N_48420);
or UO_4071 (O_4071,N_48376,N_49529);
nand UO_4072 (O_4072,N_49246,N_48267);
xnor UO_4073 (O_4073,N_49299,N_48131);
nand UO_4074 (O_4074,N_49021,N_49002);
and UO_4075 (O_4075,N_49710,N_48393);
xor UO_4076 (O_4076,N_48926,N_48708);
and UO_4077 (O_4077,N_48501,N_49542);
nor UO_4078 (O_4078,N_49828,N_48545);
or UO_4079 (O_4079,N_48268,N_49804);
nor UO_4080 (O_4080,N_48271,N_49719);
nand UO_4081 (O_4081,N_49609,N_49042);
and UO_4082 (O_4082,N_48136,N_49585);
xor UO_4083 (O_4083,N_48662,N_48986);
nand UO_4084 (O_4084,N_49642,N_49976);
nand UO_4085 (O_4085,N_48537,N_49429);
and UO_4086 (O_4086,N_48067,N_48666);
xor UO_4087 (O_4087,N_48700,N_49596);
xnor UO_4088 (O_4088,N_49624,N_49967);
xor UO_4089 (O_4089,N_49284,N_49675);
nand UO_4090 (O_4090,N_48363,N_48059);
nand UO_4091 (O_4091,N_49601,N_49344);
nor UO_4092 (O_4092,N_49170,N_48604);
xor UO_4093 (O_4093,N_48236,N_49210);
xor UO_4094 (O_4094,N_49425,N_49716);
xnor UO_4095 (O_4095,N_49267,N_49037);
or UO_4096 (O_4096,N_48894,N_48910);
xor UO_4097 (O_4097,N_49816,N_49360);
or UO_4098 (O_4098,N_49936,N_49269);
or UO_4099 (O_4099,N_49753,N_49220);
and UO_4100 (O_4100,N_49706,N_49166);
and UO_4101 (O_4101,N_49803,N_48351);
xor UO_4102 (O_4102,N_48216,N_49069);
nor UO_4103 (O_4103,N_49178,N_49406);
or UO_4104 (O_4104,N_48927,N_49817);
xor UO_4105 (O_4105,N_48098,N_49183);
and UO_4106 (O_4106,N_49477,N_48718);
nor UO_4107 (O_4107,N_48190,N_49270);
and UO_4108 (O_4108,N_49633,N_49152);
and UO_4109 (O_4109,N_49358,N_48099);
and UO_4110 (O_4110,N_48892,N_48667);
nand UO_4111 (O_4111,N_49973,N_49092);
and UO_4112 (O_4112,N_48255,N_49833);
nor UO_4113 (O_4113,N_49913,N_49989);
or UO_4114 (O_4114,N_48549,N_48508);
and UO_4115 (O_4115,N_49686,N_49469);
xor UO_4116 (O_4116,N_49692,N_48721);
nand UO_4117 (O_4117,N_48312,N_49617);
or UO_4118 (O_4118,N_49950,N_48621);
nand UO_4119 (O_4119,N_49903,N_48247);
nor UO_4120 (O_4120,N_48962,N_49674);
nand UO_4121 (O_4121,N_48940,N_49619);
nor UO_4122 (O_4122,N_49338,N_48949);
nand UO_4123 (O_4123,N_49542,N_49240);
and UO_4124 (O_4124,N_49525,N_49018);
xnor UO_4125 (O_4125,N_49001,N_48833);
and UO_4126 (O_4126,N_48720,N_48821);
nand UO_4127 (O_4127,N_48150,N_48459);
xor UO_4128 (O_4128,N_49509,N_48391);
nor UO_4129 (O_4129,N_49990,N_49772);
or UO_4130 (O_4130,N_49648,N_49920);
nand UO_4131 (O_4131,N_49226,N_49215);
or UO_4132 (O_4132,N_48449,N_49031);
xor UO_4133 (O_4133,N_49026,N_48273);
or UO_4134 (O_4134,N_48637,N_48012);
xor UO_4135 (O_4135,N_49491,N_48065);
nor UO_4136 (O_4136,N_49444,N_49808);
nor UO_4137 (O_4137,N_49366,N_48090);
and UO_4138 (O_4138,N_49357,N_48739);
and UO_4139 (O_4139,N_48927,N_49686);
or UO_4140 (O_4140,N_49380,N_48871);
nand UO_4141 (O_4141,N_49309,N_48995);
nor UO_4142 (O_4142,N_48510,N_48383);
or UO_4143 (O_4143,N_49953,N_48806);
nand UO_4144 (O_4144,N_49383,N_48969);
nand UO_4145 (O_4145,N_49107,N_48734);
xnor UO_4146 (O_4146,N_48414,N_49902);
nand UO_4147 (O_4147,N_49651,N_48568);
and UO_4148 (O_4148,N_49487,N_49500);
nor UO_4149 (O_4149,N_48378,N_48615);
or UO_4150 (O_4150,N_49164,N_48254);
xnor UO_4151 (O_4151,N_49134,N_49848);
nand UO_4152 (O_4152,N_49618,N_48399);
nand UO_4153 (O_4153,N_49684,N_48813);
nand UO_4154 (O_4154,N_48876,N_48621);
xnor UO_4155 (O_4155,N_49037,N_48248);
nand UO_4156 (O_4156,N_48112,N_48086);
nor UO_4157 (O_4157,N_49500,N_49499);
and UO_4158 (O_4158,N_49254,N_48828);
xor UO_4159 (O_4159,N_48196,N_48688);
xor UO_4160 (O_4160,N_49269,N_49341);
or UO_4161 (O_4161,N_48619,N_49320);
nand UO_4162 (O_4162,N_49212,N_49321);
or UO_4163 (O_4163,N_49628,N_48185);
xnor UO_4164 (O_4164,N_49470,N_48625);
or UO_4165 (O_4165,N_48446,N_49431);
nand UO_4166 (O_4166,N_49922,N_48518);
and UO_4167 (O_4167,N_48409,N_49838);
or UO_4168 (O_4168,N_48933,N_48016);
and UO_4169 (O_4169,N_49318,N_48788);
and UO_4170 (O_4170,N_49368,N_48794);
xnor UO_4171 (O_4171,N_49749,N_48525);
nand UO_4172 (O_4172,N_49388,N_49592);
and UO_4173 (O_4173,N_49604,N_49624);
or UO_4174 (O_4174,N_49678,N_49699);
or UO_4175 (O_4175,N_49366,N_49389);
xor UO_4176 (O_4176,N_48798,N_49891);
and UO_4177 (O_4177,N_48507,N_49218);
nor UO_4178 (O_4178,N_48726,N_48323);
nand UO_4179 (O_4179,N_49984,N_49176);
or UO_4180 (O_4180,N_48173,N_48449);
xnor UO_4181 (O_4181,N_48167,N_49060);
nand UO_4182 (O_4182,N_49879,N_49641);
or UO_4183 (O_4183,N_49770,N_48068);
nand UO_4184 (O_4184,N_49570,N_48208);
or UO_4185 (O_4185,N_49565,N_48359);
nor UO_4186 (O_4186,N_48566,N_48549);
nor UO_4187 (O_4187,N_48797,N_49969);
nor UO_4188 (O_4188,N_48655,N_49340);
or UO_4189 (O_4189,N_48364,N_48495);
nand UO_4190 (O_4190,N_49660,N_48294);
xor UO_4191 (O_4191,N_49066,N_49327);
nand UO_4192 (O_4192,N_49913,N_49025);
or UO_4193 (O_4193,N_49564,N_48090);
and UO_4194 (O_4194,N_49366,N_49688);
nor UO_4195 (O_4195,N_48726,N_48714);
nor UO_4196 (O_4196,N_48714,N_49360);
or UO_4197 (O_4197,N_48045,N_48624);
and UO_4198 (O_4198,N_48296,N_48990);
or UO_4199 (O_4199,N_48971,N_48178);
or UO_4200 (O_4200,N_49207,N_49046);
xnor UO_4201 (O_4201,N_48423,N_49820);
and UO_4202 (O_4202,N_48286,N_49884);
xnor UO_4203 (O_4203,N_48139,N_48979);
nor UO_4204 (O_4204,N_49459,N_49666);
or UO_4205 (O_4205,N_48659,N_49987);
and UO_4206 (O_4206,N_48665,N_49781);
or UO_4207 (O_4207,N_48335,N_48371);
nor UO_4208 (O_4208,N_49640,N_49788);
nor UO_4209 (O_4209,N_49210,N_48602);
or UO_4210 (O_4210,N_49335,N_48252);
nand UO_4211 (O_4211,N_48266,N_49993);
and UO_4212 (O_4212,N_49233,N_49833);
or UO_4213 (O_4213,N_49671,N_48235);
nand UO_4214 (O_4214,N_49126,N_48355);
or UO_4215 (O_4215,N_48505,N_49786);
or UO_4216 (O_4216,N_49559,N_48230);
and UO_4217 (O_4217,N_48418,N_48460);
and UO_4218 (O_4218,N_49878,N_49544);
nand UO_4219 (O_4219,N_49035,N_48634);
nor UO_4220 (O_4220,N_49126,N_48724);
or UO_4221 (O_4221,N_48089,N_48484);
nor UO_4222 (O_4222,N_49943,N_48367);
or UO_4223 (O_4223,N_48525,N_48757);
or UO_4224 (O_4224,N_48514,N_48247);
xor UO_4225 (O_4225,N_48907,N_48815);
and UO_4226 (O_4226,N_48109,N_49347);
nand UO_4227 (O_4227,N_49460,N_48940);
xor UO_4228 (O_4228,N_48561,N_48336);
xor UO_4229 (O_4229,N_48624,N_48790);
and UO_4230 (O_4230,N_48042,N_49293);
and UO_4231 (O_4231,N_49229,N_48653);
nand UO_4232 (O_4232,N_49834,N_48359);
nand UO_4233 (O_4233,N_49058,N_49153);
nand UO_4234 (O_4234,N_49414,N_49121);
or UO_4235 (O_4235,N_49940,N_49652);
nand UO_4236 (O_4236,N_48350,N_49092);
xnor UO_4237 (O_4237,N_49605,N_48657);
nand UO_4238 (O_4238,N_49195,N_48462);
nor UO_4239 (O_4239,N_49613,N_48651);
and UO_4240 (O_4240,N_49393,N_49716);
nand UO_4241 (O_4241,N_49946,N_48920);
nand UO_4242 (O_4242,N_48217,N_49621);
or UO_4243 (O_4243,N_48951,N_48735);
nand UO_4244 (O_4244,N_48262,N_49719);
nor UO_4245 (O_4245,N_48715,N_49798);
and UO_4246 (O_4246,N_48721,N_48365);
nor UO_4247 (O_4247,N_49050,N_49793);
nor UO_4248 (O_4248,N_48826,N_49735);
or UO_4249 (O_4249,N_48128,N_49277);
and UO_4250 (O_4250,N_48059,N_48163);
nand UO_4251 (O_4251,N_49030,N_49265);
xnor UO_4252 (O_4252,N_49596,N_49624);
and UO_4253 (O_4253,N_49866,N_48014);
xnor UO_4254 (O_4254,N_49290,N_48476);
xor UO_4255 (O_4255,N_49627,N_49114);
xnor UO_4256 (O_4256,N_48626,N_49137);
nand UO_4257 (O_4257,N_49308,N_49954);
and UO_4258 (O_4258,N_49485,N_48169);
or UO_4259 (O_4259,N_49821,N_48278);
nor UO_4260 (O_4260,N_49283,N_48767);
xor UO_4261 (O_4261,N_49090,N_48411);
nand UO_4262 (O_4262,N_48288,N_48740);
xor UO_4263 (O_4263,N_48070,N_49735);
xnor UO_4264 (O_4264,N_48088,N_48286);
and UO_4265 (O_4265,N_49515,N_49024);
nor UO_4266 (O_4266,N_49244,N_48153);
xnor UO_4267 (O_4267,N_48146,N_49921);
and UO_4268 (O_4268,N_49759,N_49670);
or UO_4269 (O_4269,N_49302,N_48730);
xnor UO_4270 (O_4270,N_48226,N_49296);
xnor UO_4271 (O_4271,N_49312,N_48673);
and UO_4272 (O_4272,N_49195,N_49886);
and UO_4273 (O_4273,N_49006,N_48991);
or UO_4274 (O_4274,N_48437,N_49859);
xor UO_4275 (O_4275,N_48409,N_49828);
nor UO_4276 (O_4276,N_48445,N_49226);
nor UO_4277 (O_4277,N_49728,N_49752);
and UO_4278 (O_4278,N_49696,N_49022);
xnor UO_4279 (O_4279,N_49918,N_49483);
or UO_4280 (O_4280,N_49152,N_49146);
or UO_4281 (O_4281,N_48381,N_49496);
or UO_4282 (O_4282,N_48607,N_48660);
or UO_4283 (O_4283,N_49985,N_49681);
xnor UO_4284 (O_4284,N_49327,N_49898);
and UO_4285 (O_4285,N_49472,N_48244);
xor UO_4286 (O_4286,N_48287,N_48673);
and UO_4287 (O_4287,N_49885,N_48067);
nor UO_4288 (O_4288,N_48623,N_48027);
nor UO_4289 (O_4289,N_49351,N_49180);
nand UO_4290 (O_4290,N_49658,N_48423);
nand UO_4291 (O_4291,N_48051,N_49901);
nor UO_4292 (O_4292,N_49986,N_48075);
and UO_4293 (O_4293,N_48843,N_49714);
or UO_4294 (O_4294,N_48669,N_49218);
nor UO_4295 (O_4295,N_49083,N_48405);
nand UO_4296 (O_4296,N_48605,N_49477);
xor UO_4297 (O_4297,N_48273,N_49191);
or UO_4298 (O_4298,N_48665,N_48749);
xor UO_4299 (O_4299,N_49765,N_49698);
nor UO_4300 (O_4300,N_49431,N_48394);
nand UO_4301 (O_4301,N_49494,N_49575);
and UO_4302 (O_4302,N_48338,N_48031);
xnor UO_4303 (O_4303,N_49680,N_49608);
nand UO_4304 (O_4304,N_48626,N_49701);
nor UO_4305 (O_4305,N_49884,N_49941);
xnor UO_4306 (O_4306,N_49358,N_48337);
nand UO_4307 (O_4307,N_48115,N_48260);
and UO_4308 (O_4308,N_48158,N_48450);
nand UO_4309 (O_4309,N_48983,N_48263);
xor UO_4310 (O_4310,N_49643,N_48807);
and UO_4311 (O_4311,N_49073,N_49995);
nand UO_4312 (O_4312,N_49113,N_48424);
nor UO_4313 (O_4313,N_49470,N_49371);
xor UO_4314 (O_4314,N_48450,N_49072);
and UO_4315 (O_4315,N_48320,N_49665);
xor UO_4316 (O_4316,N_49975,N_48685);
and UO_4317 (O_4317,N_48860,N_48830);
or UO_4318 (O_4318,N_49210,N_49926);
or UO_4319 (O_4319,N_49701,N_48848);
and UO_4320 (O_4320,N_48431,N_49064);
nor UO_4321 (O_4321,N_49848,N_48685);
or UO_4322 (O_4322,N_48584,N_49507);
xor UO_4323 (O_4323,N_48581,N_48408);
xor UO_4324 (O_4324,N_49123,N_49907);
and UO_4325 (O_4325,N_48992,N_49860);
and UO_4326 (O_4326,N_48333,N_49515);
or UO_4327 (O_4327,N_48624,N_48863);
nor UO_4328 (O_4328,N_49866,N_49082);
and UO_4329 (O_4329,N_48273,N_48211);
or UO_4330 (O_4330,N_49012,N_49070);
xnor UO_4331 (O_4331,N_49973,N_49665);
nand UO_4332 (O_4332,N_48816,N_48897);
nor UO_4333 (O_4333,N_49765,N_48895);
or UO_4334 (O_4334,N_48509,N_48851);
and UO_4335 (O_4335,N_49806,N_49152);
nand UO_4336 (O_4336,N_49305,N_48740);
xnor UO_4337 (O_4337,N_48114,N_49075);
xnor UO_4338 (O_4338,N_48777,N_48401);
or UO_4339 (O_4339,N_49560,N_49235);
nand UO_4340 (O_4340,N_48899,N_49770);
and UO_4341 (O_4341,N_49150,N_48297);
xnor UO_4342 (O_4342,N_49883,N_49578);
nand UO_4343 (O_4343,N_49272,N_48762);
nor UO_4344 (O_4344,N_49257,N_48860);
nand UO_4345 (O_4345,N_48012,N_48227);
nand UO_4346 (O_4346,N_49197,N_49587);
xor UO_4347 (O_4347,N_49531,N_48921);
or UO_4348 (O_4348,N_48480,N_49279);
or UO_4349 (O_4349,N_48814,N_48049);
xor UO_4350 (O_4350,N_49831,N_49008);
and UO_4351 (O_4351,N_49306,N_48878);
xnor UO_4352 (O_4352,N_48896,N_49022);
xor UO_4353 (O_4353,N_49048,N_48887);
xor UO_4354 (O_4354,N_48075,N_49627);
xor UO_4355 (O_4355,N_48786,N_49744);
or UO_4356 (O_4356,N_48896,N_49656);
nand UO_4357 (O_4357,N_48718,N_48332);
nand UO_4358 (O_4358,N_49514,N_48157);
and UO_4359 (O_4359,N_48952,N_49111);
and UO_4360 (O_4360,N_49894,N_49689);
or UO_4361 (O_4361,N_49638,N_49197);
or UO_4362 (O_4362,N_49088,N_49412);
nand UO_4363 (O_4363,N_49559,N_48222);
and UO_4364 (O_4364,N_49809,N_49428);
or UO_4365 (O_4365,N_49993,N_49592);
nor UO_4366 (O_4366,N_49727,N_48860);
nand UO_4367 (O_4367,N_48747,N_49932);
and UO_4368 (O_4368,N_48604,N_49719);
or UO_4369 (O_4369,N_48517,N_48042);
nand UO_4370 (O_4370,N_48392,N_49707);
nor UO_4371 (O_4371,N_49392,N_49487);
xor UO_4372 (O_4372,N_48563,N_49935);
xor UO_4373 (O_4373,N_49301,N_48697);
xnor UO_4374 (O_4374,N_48236,N_49117);
nor UO_4375 (O_4375,N_49556,N_49539);
xnor UO_4376 (O_4376,N_48701,N_49796);
or UO_4377 (O_4377,N_48171,N_49340);
nor UO_4378 (O_4378,N_48490,N_48784);
and UO_4379 (O_4379,N_49625,N_49117);
xnor UO_4380 (O_4380,N_49864,N_48908);
or UO_4381 (O_4381,N_49979,N_49737);
nor UO_4382 (O_4382,N_48838,N_49967);
xnor UO_4383 (O_4383,N_48879,N_49174);
nand UO_4384 (O_4384,N_48026,N_48585);
xor UO_4385 (O_4385,N_49140,N_49691);
nor UO_4386 (O_4386,N_49351,N_48306);
nor UO_4387 (O_4387,N_48771,N_48943);
or UO_4388 (O_4388,N_48019,N_48902);
and UO_4389 (O_4389,N_48321,N_48767);
xor UO_4390 (O_4390,N_48348,N_48854);
nor UO_4391 (O_4391,N_48639,N_48150);
xor UO_4392 (O_4392,N_49197,N_48857);
nor UO_4393 (O_4393,N_48855,N_48278);
and UO_4394 (O_4394,N_49012,N_48732);
and UO_4395 (O_4395,N_48035,N_48247);
or UO_4396 (O_4396,N_48309,N_49900);
or UO_4397 (O_4397,N_48991,N_49809);
nand UO_4398 (O_4398,N_49531,N_49140);
xor UO_4399 (O_4399,N_48650,N_48400);
and UO_4400 (O_4400,N_49777,N_48357);
or UO_4401 (O_4401,N_49753,N_49801);
xnor UO_4402 (O_4402,N_49693,N_48956);
nor UO_4403 (O_4403,N_49184,N_48700);
and UO_4404 (O_4404,N_48788,N_48577);
and UO_4405 (O_4405,N_49168,N_49433);
nor UO_4406 (O_4406,N_49985,N_48943);
xnor UO_4407 (O_4407,N_48536,N_48546);
nand UO_4408 (O_4408,N_48660,N_49858);
nand UO_4409 (O_4409,N_48089,N_48843);
xnor UO_4410 (O_4410,N_49339,N_48349);
or UO_4411 (O_4411,N_48680,N_48325);
nor UO_4412 (O_4412,N_48247,N_49206);
and UO_4413 (O_4413,N_48494,N_48816);
or UO_4414 (O_4414,N_49993,N_49023);
and UO_4415 (O_4415,N_49047,N_49380);
xnor UO_4416 (O_4416,N_49021,N_48387);
xnor UO_4417 (O_4417,N_49388,N_49530);
nor UO_4418 (O_4418,N_48091,N_49737);
nand UO_4419 (O_4419,N_48594,N_49451);
nand UO_4420 (O_4420,N_48755,N_49276);
or UO_4421 (O_4421,N_48515,N_48049);
xnor UO_4422 (O_4422,N_48212,N_49372);
xor UO_4423 (O_4423,N_48680,N_49649);
xnor UO_4424 (O_4424,N_49630,N_48381);
xor UO_4425 (O_4425,N_49470,N_48843);
and UO_4426 (O_4426,N_49223,N_49016);
nand UO_4427 (O_4427,N_48275,N_49263);
xnor UO_4428 (O_4428,N_48567,N_49502);
or UO_4429 (O_4429,N_49342,N_48490);
xnor UO_4430 (O_4430,N_48792,N_49456);
nor UO_4431 (O_4431,N_49574,N_49113);
nor UO_4432 (O_4432,N_48640,N_48538);
xnor UO_4433 (O_4433,N_49172,N_48442);
and UO_4434 (O_4434,N_48793,N_48040);
nor UO_4435 (O_4435,N_49524,N_48734);
and UO_4436 (O_4436,N_49870,N_48087);
or UO_4437 (O_4437,N_48043,N_48222);
or UO_4438 (O_4438,N_48623,N_49328);
xor UO_4439 (O_4439,N_48565,N_48976);
or UO_4440 (O_4440,N_49966,N_48713);
or UO_4441 (O_4441,N_49007,N_49504);
nand UO_4442 (O_4442,N_49031,N_48661);
or UO_4443 (O_4443,N_49279,N_49654);
nand UO_4444 (O_4444,N_48867,N_49274);
nor UO_4445 (O_4445,N_48189,N_48463);
xnor UO_4446 (O_4446,N_49721,N_49047);
and UO_4447 (O_4447,N_49783,N_49500);
or UO_4448 (O_4448,N_49282,N_48681);
nor UO_4449 (O_4449,N_48640,N_49041);
or UO_4450 (O_4450,N_49931,N_48912);
or UO_4451 (O_4451,N_48671,N_49234);
xnor UO_4452 (O_4452,N_48352,N_49536);
xnor UO_4453 (O_4453,N_48978,N_48693);
and UO_4454 (O_4454,N_49400,N_49094);
xnor UO_4455 (O_4455,N_48059,N_49976);
xnor UO_4456 (O_4456,N_49193,N_49748);
or UO_4457 (O_4457,N_48682,N_48695);
xor UO_4458 (O_4458,N_48530,N_49514);
nand UO_4459 (O_4459,N_49724,N_49552);
xnor UO_4460 (O_4460,N_48627,N_49744);
nand UO_4461 (O_4461,N_49857,N_49021);
and UO_4462 (O_4462,N_48183,N_48096);
nand UO_4463 (O_4463,N_48807,N_49084);
nor UO_4464 (O_4464,N_48584,N_48627);
and UO_4465 (O_4465,N_48540,N_48851);
and UO_4466 (O_4466,N_48149,N_49980);
and UO_4467 (O_4467,N_49998,N_49221);
and UO_4468 (O_4468,N_48513,N_48701);
nand UO_4469 (O_4469,N_49275,N_48616);
nand UO_4470 (O_4470,N_48511,N_49931);
or UO_4471 (O_4471,N_49071,N_49492);
xor UO_4472 (O_4472,N_48122,N_48462);
and UO_4473 (O_4473,N_48811,N_49583);
nor UO_4474 (O_4474,N_49244,N_48665);
xor UO_4475 (O_4475,N_48380,N_49910);
or UO_4476 (O_4476,N_49974,N_48297);
or UO_4477 (O_4477,N_48837,N_48080);
or UO_4478 (O_4478,N_49666,N_49860);
xor UO_4479 (O_4479,N_48883,N_49635);
or UO_4480 (O_4480,N_49543,N_49063);
xor UO_4481 (O_4481,N_49296,N_48183);
and UO_4482 (O_4482,N_48643,N_49777);
nand UO_4483 (O_4483,N_48220,N_49974);
and UO_4484 (O_4484,N_48205,N_48424);
and UO_4485 (O_4485,N_48848,N_48131);
nand UO_4486 (O_4486,N_49295,N_49010);
and UO_4487 (O_4487,N_49877,N_49281);
and UO_4488 (O_4488,N_48039,N_49633);
or UO_4489 (O_4489,N_49033,N_49765);
and UO_4490 (O_4490,N_49553,N_49350);
nor UO_4491 (O_4491,N_49088,N_48030);
nand UO_4492 (O_4492,N_48464,N_49629);
and UO_4493 (O_4493,N_48837,N_49429);
nand UO_4494 (O_4494,N_48006,N_49464);
and UO_4495 (O_4495,N_48121,N_48469);
and UO_4496 (O_4496,N_49077,N_48211);
nand UO_4497 (O_4497,N_49905,N_49428);
nor UO_4498 (O_4498,N_49218,N_49768);
nor UO_4499 (O_4499,N_49183,N_48384);
and UO_4500 (O_4500,N_48505,N_49711);
nor UO_4501 (O_4501,N_49895,N_48083);
and UO_4502 (O_4502,N_49509,N_49615);
nand UO_4503 (O_4503,N_48816,N_49490);
nor UO_4504 (O_4504,N_48983,N_48093);
xnor UO_4505 (O_4505,N_49990,N_48535);
and UO_4506 (O_4506,N_49594,N_49340);
nor UO_4507 (O_4507,N_49710,N_49467);
or UO_4508 (O_4508,N_49831,N_48545);
and UO_4509 (O_4509,N_48786,N_48845);
and UO_4510 (O_4510,N_48107,N_48372);
and UO_4511 (O_4511,N_48353,N_48922);
or UO_4512 (O_4512,N_49885,N_48204);
or UO_4513 (O_4513,N_49581,N_49366);
or UO_4514 (O_4514,N_49706,N_48914);
and UO_4515 (O_4515,N_48898,N_48637);
xor UO_4516 (O_4516,N_48461,N_48450);
and UO_4517 (O_4517,N_48664,N_49860);
nor UO_4518 (O_4518,N_49053,N_49385);
nor UO_4519 (O_4519,N_48974,N_48459);
nand UO_4520 (O_4520,N_49820,N_49334);
xor UO_4521 (O_4521,N_49258,N_48090);
and UO_4522 (O_4522,N_49096,N_48074);
or UO_4523 (O_4523,N_49370,N_49263);
and UO_4524 (O_4524,N_48725,N_49064);
nand UO_4525 (O_4525,N_48723,N_49658);
xor UO_4526 (O_4526,N_49861,N_49190);
and UO_4527 (O_4527,N_48731,N_49211);
nand UO_4528 (O_4528,N_48690,N_49821);
nor UO_4529 (O_4529,N_49138,N_48761);
xor UO_4530 (O_4530,N_49879,N_49871);
nor UO_4531 (O_4531,N_49554,N_48177);
or UO_4532 (O_4532,N_48088,N_48406);
nand UO_4533 (O_4533,N_49754,N_48509);
or UO_4534 (O_4534,N_48619,N_48534);
nor UO_4535 (O_4535,N_48419,N_49659);
or UO_4536 (O_4536,N_48204,N_48126);
xnor UO_4537 (O_4537,N_49025,N_49214);
xnor UO_4538 (O_4538,N_48452,N_49213);
nand UO_4539 (O_4539,N_49379,N_48549);
nand UO_4540 (O_4540,N_48839,N_48471);
xnor UO_4541 (O_4541,N_49135,N_48764);
and UO_4542 (O_4542,N_48704,N_49845);
or UO_4543 (O_4543,N_48531,N_48025);
nor UO_4544 (O_4544,N_49135,N_48725);
and UO_4545 (O_4545,N_49631,N_48234);
and UO_4546 (O_4546,N_49162,N_49821);
nand UO_4547 (O_4547,N_48913,N_49962);
or UO_4548 (O_4548,N_48154,N_49980);
xnor UO_4549 (O_4549,N_48947,N_49453);
and UO_4550 (O_4550,N_49216,N_48343);
and UO_4551 (O_4551,N_48028,N_48063);
nand UO_4552 (O_4552,N_48795,N_49928);
and UO_4553 (O_4553,N_49567,N_49293);
nand UO_4554 (O_4554,N_49984,N_48356);
or UO_4555 (O_4555,N_48953,N_49689);
nand UO_4556 (O_4556,N_49191,N_49683);
nand UO_4557 (O_4557,N_48771,N_49438);
nor UO_4558 (O_4558,N_48840,N_48278);
nand UO_4559 (O_4559,N_48814,N_48659);
nor UO_4560 (O_4560,N_48774,N_49304);
or UO_4561 (O_4561,N_48678,N_49706);
or UO_4562 (O_4562,N_49898,N_48796);
nor UO_4563 (O_4563,N_48963,N_49712);
or UO_4564 (O_4564,N_48908,N_48511);
xor UO_4565 (O_4565,N_49049,N_49101);
or UO_4566 (O_4566,N_48284,N_48694);
and UO_4567 (O_4567,N_48028,N_48166);
xnor UO_4568 (O_4568,N_48272,N_49937);
nand UO_4569 (O_4569,N_48447,N_48529);
xor UO_4570 (O_4570,N_48762,N_48003);
and UO_4571 (O_4571,N_49032,N_48758);
xor UO_4572 (O_4572,N_48521,N_49946);
xnor UO_4573 (O_4573,N_49323,N_49682);
nand UO_4574 (O_4574,N_49968,N_49564);
nor UO_4575 (O_4575,N_48970,N_49927);
nand UO_4576 (O_4576,N_49796,N_48425);
or UO_4577 (O_4577,N_48125,N_48084);
nor UO_4578 (O_4578,N_49011,N_49898);
or UO_4579 (O_4579,N_48830,N_48277);
nor UO_4580 (O_4580,N_49663,N_48948);
xnor UO_4581 (O_4581,N_49158,N_48626);
nand UO_4582 (O_4582,N_48203,N_48702);
xnor UO_4583 (O_4583,N_48412,N_49783);
nand UO_4584 (O_4584,N_48446,N_49485);
xnor UO_4585 (O_4585,N_48259,N_49854);
nor UO_4586 (O_4586,N_48218,N_49353);
or UO_4587 (O_4587,N_48877,N_48894);
xnor UO_4588 (O_4588,N_48312,N_48158);
or UO_4589 (O_4589,N_48342,N_49651);
xor UO_4590 (O_4590,N_49787,N_48530);
nor UO_4591 (O_4591,N_48152,N_48508);
and UO_4592 (O_4592,N_49447,N_48522);
nor UO_4593 (O_4593,N_48051,N_49460);
or UO_4594 (O_4594,N_49894,N_48311);
or UO_4595 (O_4595,N_49853,N_48155);
xnor UO_4596 (O_4596,N_49041,N_49433);
xor UO_4597 (O_4597,N_49602,N_48334);
and UO_4598 (O_4598,N_48567,N_49195);
nand UO_4599 (O_4599,N_49054,N_48333);
and UO_4600 (O_4600,N_48759,N_49860);
or UO_4601 (O_4601,N_48327,N_49617);
nor UO_4602 (O_4602,N_49779,N_49526);
nand UO_4603 (O_4603,N_49137,N_49454);
and UO_4604 (O_4604,N_48633,N_48184);
nand UO_4605 (O_4605,N_49360,N_48029);
and UO_4606 (O_4606,N_49898,N_48067);
nand UO_4607 (O_4607,N_49109,N_48749);
and UO_4608 (O_4608,N_49808,N_49147);
xnor UO_4609 (O_4609,N_48540,N_48754);
xnor UO_4610 (O_4610,N_49061,N_49461);
nor UO_4611 (O_4611,N_48520,N_48153);
or UO_4612 (O_4612,N_49414,N_48822);
and UO_4613 (O_4613,N_48145,N_49565);
nand UO_4614 (O_4614,N_49427,N_48955);
xnor UO_4615 (O_4615,N_48482,N_49996);
or UO_4616 (O_4616,N_48050,N_48462);
nor UO_4617 (O_4617,N_48092,N_48310);
xnor UO_4618 (O_4618,N_48753,N_49752);
and UO_4619 (O_4619,N_48292,N_49641);
xor UO_4620 (O_4620,N_48181,N_48638);
or UO_4621 (O_4621,N_49117,N_49479);
and UO_4622 (O_4622,N_49033,N_49112);
xor UO_4623 (O_4623,N_49845,N_49905);
or UO_4624 (O_4624,N_48201,N_48687);
and UO_4625 (O_4625,N_49226,N_49064);
nand UO_4626 (O_4626,N_48677,N_48863);
nand UO_4627 (O_4627,N_48040,N_48265);
xnor UO_4628 (O_4628,N_49340,N_48708);
nand UO_4629 (O_4629,N_49587,N_49019);
nand UO_4630 (O_4630,N_49001,N_49482);
or UO_4631 (O_4631,N_48946,N_49418);
or UO_4632 (O_4632,N_48556,N_49560);
and UO_4633 (O_4633,N_49114,N_48950);
nand UO_4634 (O_4634,N_49590,N_49073);
nand UO_4635 (O_4635,N_48500,N_48682);
nand UO_4636 (O_4636,N_48072,N_48194);
nand UO_4637 (O_4637,N_49031,N_48951);
xnor UO_4638 (O_4638,N_48767,N_48741);
or UO_4639 (O_4639,N_48498,N_49625);
xnor UO_4640 (O_4640,N_49378,N_48179);
and UO_4641 (O_4641,N_49077,N_49325);
nor UO_4642 (O_4642,N_49075,N_49177);
nand UO_4643 (O_4643,N_49577,N_49941);
xnor UO_4644 (O_4644,N_49345,N_49130);
xnor UO_4645 (O_4645,N_48773,N_48826);
xor UO_4646 (O_4646,N_49071,N_48707);
nand UO_4647 (O_4647,N_49650,N_48488);
and UO_4648 (O_4648,N_48942,N_49192);
nand UO_4649 (O_4649,N_48849,N_48284);
xnor UO_4650 (O_4650,N_49169,N_48143);
nand UO_4651 (O_4651,N_48536,N_48556);
nor UO_4652 (O_4652,N_49851,N_48390);
nor UO_4653 (O_4653,N_48045,N_49281);
nor UO_4654 (O_4654,N_49216,N_48952);
or UO_4655 (O_4655,N_48281,N_48715);
nor UO_4656 (O_4656,N_48580,N_49682);
xor UO_4657 (O_4657,N_49068,N_48013);
nand UO_4658 (O_4658,N_49309,N_48656);
and UO_4659 (O_4659,N_48855,N_49020);
nor UO_4660 (O_4660,N_49608,N_49403);
xnor UO_4661 (O_4661,N_48445,N_48835);
nand UO_4662 (O_4662,N_48551,N_48226);
nand UO_4663 (O_4663,N_49835,N_49807);
and UO_4664 (O_4664,N_48613,N_49490);
nor UO_4665 (O_4665,N_49012,N_49290);
xnor UO_4666 (O_4666,N_48529,N_48542);
xor UO_4667 (O_4667,N_48005,N_49753);
nor UO_4668 (O_4668,N_49889,N_49820);
nand UO_4669 (O_4669,N_49396,N_49245);
nor UO_4670 (O_4670,N_49208,N_49723);
and UO_4671 (O_4671,N_49020,N_48577);
nand UO_4672 (O_4672,N_48761,N_48014);
nand UO_4673 (O_4673,N_49007,N_49108);
nand UO_4674 (O_4674,N_48683,N_48051);
and UO_4675 (O_4675,N_49463,N_49381);
xnor UO_4676 (O_4676,N_48494,N_49121);
nand UO_4677 (O_4677,N_49516,N_48042);
or UO_4678 (O_4678,N_48558,N_49883);
nor UO_4679 (O_4679,N_48705,N_49616);
or UO_4680 (O_4680,N_48042,N_49223);
or UO_4681 (O_4681,N_49707,N_48251);
nand UO_4682 (O_4682,N_49881,N_48617);
and UO_4683 (O_4683,N_48073,N_49020);
nor UO_4684 (O_4684,N_49748,N_49945);
xor UO_4685 (O_4685,N_49531,N_48699);
or UO_4686 (O_4686,N_49544,N_48459);
nor UO_4687 (O_4687,N_49623,N_48680);
nor UO_4688 (O_4688,N_48602,N_49228);
nor UO_4689 (O_4689,N_49705,N_49770);
xor UO_4690 (O_4690,N_49493,N_49100);
nand UO_4691 (O_4691,N_48990,N_48816);
nand UO_4692 (O_4692,N_49535,N_49792);
or UO_4693 (O_4693,N_48054,N_49850);
nor UO_4694 (O_4694,N_48540,N_49574);
xor UO_4695 (O_4695,N_49186,N_48430);
nor UO_4696 (O_4696,N_48400,N_49079);
xnor UO_4697 (O_4697,N_48210,N_48942);
nor UO_4698 (O_4698,N_48685,N_48073);
or UO_4699 (O_4699,N_48786,N_49776);
nand UO_4700 (O_4700,N_48320,N_48274);
and UO_4701 (O_4701,N_48722,N_49900);
or UO_4702 (O_4702,N_48491,N_48085);
nand UO_4703 (O_4703,N_48762,N_49947);
xnor UO_4704 (O_4704,N_48261,N_49797);
or UO_4705 (O_4705,N_48557,N_48780);
xnor UO_4706 (O_4706,N_48689,N_49781);
nand UO_4707 (O_4707,N_48112,N_48110);
or UO_4708 (O_4708,N_49653,N_48510);
or UO_4709 (O_4709,N_49101,N_49250);
nor UO_4710 (O_4710,N_49228,N_49410);
xor UO_4711 (O_4711,N_48186,N_49059);
nand UO_4712 (O_4712,N_49774,N_48499);
and UO_4713 (O_4713,N_49364,N_48887);
nor UO_4714 (O_4714,N_49891,N_48954);
nor UO_4715 (O_4715,N_48381,N_49583);
or UO_4716 (O_4716,N_48199,N_49549);
xnor UO_4717 (O_4717,N_48366,N_48016);
nand UO_4718 (O_4718,N_49495,N_48392);
nor UO_4719 (O_4719,N_49729,N_49879);
nor UO_4720 (O_4720,N_49456,N_48393);
nor UO_4721 (O_4721,N_49080,N_48392);
xor UO_4722 (O_4722,N_48116,N_48932);
and UO_4723 (O_4723,N_49387,N_49582);
or UO_4724 (O_4724,N_48829,N_49427);
nand UO_4725 (O_4725,N_49307,N_49314);
xnor UO_4726 (O_4726,N_48476,N_48214);
nor UO_4727 (O_4727,N_49015,N_49552);
or UO_4728 (O_4728,N_49078,N_48366);
nor UO_4729 (O_4729,N_48526,N_48081);
or UO_4730 (O_4730,N_49498,N_48031);
nor UO_4731 (O_4731,N_49683,N_49607);
or UO_4732 (O_4732,N_49169,N_49349);
and UO_4733 (O_4733,N_49776,N_49471);
or UO_4734 (O_4734,N_48178,N_48647);
or UO_4735 (O_4735,N_48323,N_49114);
nand UO_4736 (O_4736,N_49872,N_49898);
and UO_4737 (O_4737,N_49623,N_48315);
and UO_4738 (O_4738,N_49411,N_48184);
xnor UO_4739 (O_4739,N_49067,N_48208);
nor UO_4740 (O_4740,N_48658,N_48696);
xor UO_4741 (O_4741,N_48173,N_48266);
or UO_4742 (O_4742,N_49980,N_49641);
and UO_4743 (O_4743,N_48354,N_49483);
nor UO_4744 (O_4744,N_49302,N_49501);
and UO_4745 (O_4745,N_48773,N_49071);
or UO_4746 (O_4746,N_48942,N_48321);
xor UO_4747 (O_4747,N_48442,N_48975);
and UO_4748 (O_4748,N_49856,N_49724);
nor UO_4749 (O_4749,N_48672,N_48748);
nand UO_4750 (O_4750,N_49567,N_48426);
and UO_4751 (O_4751,N_49959,N_48440);
xor UO_4752 (O_4752,N_49201,N_48225);
nand UO_4753 (O_4753,N_49474,N_48078);
or UO_4754 (O_4754,N_49147,N_48870);
nand UO_4755 (O_4755,N_48532,N_49694);
or UO_4756 (O_4756,N_48715,N_49903);
and UO_4757 (O_4757,N_49273,N_49340);
and UO_4758 (O_4758,N_48926,N_49678);
or UO_4759 (O_4759,N_49414,N_49011);
nand UO_4760 (O_4760,N_49925,N_48739);
nor UO_4761 (O_4761,N_49557,N_49420);
nand UO_4762 (O_4762,N_49921,N_48796);
xor UO_4763 (O_4763,N_48229,N_48774);
and UO_4764 (O_4764,N_49948,N_48048);
nand UO_4765 (O_4765,N_49725,N_49452);
nor UO_4766 (O_4766,N_48062,N_48345);
and UO_4767 (O_4767,N_48067,N_48451);
nand UO_4768 (O_4768,N_48863,N_49619);
or UO_4769 (O_4769,N_48512,N_48732);
nor UO_4770 (O_4770,N_48603,N_49177);
nor UO_4771 (O_4771,N_48386,N_48150);
xor UO_4772 (O_4772,N_49561,N_49776);
and UO_4773 (O_4773,N_49290,N_48079);
nor UO_4774 (O_4774,N_49429,N_49986);
xor UO_4775 (O_4775,N_48778,N_49425);
nand UO_4776 (O_4776,N_48184,N_48835);
nand UO_4777 (O_4777,N_48168,N_48176);
or UO_4778 (O_4778,N_49494,N_49535);
or UO_4779 (O_4779,N_48033,N_48939);
xnor UO_4780 (O_4780,N_48657,N_49405);
xnor UO_4781 (O_4781,N_49442,N_48380);
and UO_4782 (O_4782,N_48618,N_49599);
or UO_4783 (O_4783,N_49093,N_49584);
or UO_4784 (O_4784,N_48099,N_48859);
xnor UO_4785 (O_4785,N_48433,N_48251);
nand UO_4786 (O_4786,N_48748,N_49897);
or UO_4787 (O_4787,N_49013,N_49762);
or UO_4788 (O_4788,N_48555,N_49700);
and UO_4789 (O_4789,N_49601,N_48402);
nand UO_4790 (O_4790,N_48601,N_48426);
nand UO_4791 (O_4791,N_49391,N_49112);
nor UO_4792 (O_4792,N_48803,N_48784);
nor UO_4793 (O_4793,N_48072,N_48350);
and UO_4794 (O_4794,N_49441,N_48464);
and UO_4795 (O_4795,N_49484,N_48607);
nor UO_4796 (O_4796,N_48899,N_49249);
or UO_4797 (O_4797,N_49383,N_48606);
or UO_4798 (O_4798,N_49293,N_48662);
or UO_4799 (O_4799,N_49952,N_48145);
nand UO_4800 (O_4800,N_48331,N_48397);
and UO_4801 (O_4801,N_48089,N_49867);
nor UO_4802 (O_4802,N_48190,N_49333);
nand UO_4803 (O_4803,N_48611,N_49838);
nor UO_4804 (O_4804,N_48829,N_49681);
and UO_4805 (O_4805,N_48138,N_49725);
nor UO_4806 (O_4806,N_48059,N_48137);
xnor UO_4807 (O_4807,N_49142,N_48175);
xor UO_4808 (O_4808,N_49453,N_48473);
xor UO_4809 (O_4809,N_49417,N_48842);
or UO_4810 (O_4810,N_49154,N_49729);
nand UO_4811 (O_4811,N_48678,N_49154);
and UO_4812 (O_4812,N_49452,N_49436);
nor UO_4813 (O_4813,N_49847,N_49061);
nand UO_4814 (O_4814,N_48581,N_49298);
xor UO_4815 (O_4815,N_49043,N_49908);
nand UO_4816 (O_4816,N_49226,N_49456);
and UO_4817 (O_4817,N_49335,N_48392);
xnor UO_4818 (O_4818,N_49489,N_48701);
nor UO_4819 (O_4819,N_48850,N_48139);
and UO_4820 (O_4820,N_49822,N_48506);
nor UO_4821 (O_4821,N_49371,N_49146);
and UO_4822 (O_4822,N_48521,N_49626);
nand UO_4823 (O_4823,N_49870,N_48059);
nand UO_4824 (O_4824,N_49712,N_49390);
and UO_4825 (O_4825,N_48862,N_49410);
nor UO_4826 (O_4826,N_49907,N_49398);
and UO_4827 (O_4827,N_49073,N_49513);
and UO_4828 (O_4828,N_48701,N_48408);
xnor UO_4829 (O_4829,N_49878,N_48649);
or UO_4830 (O_4830,N_49250,N_48232);
nand UO_4831 (O_4831,N_49630,N_48511);
xnor UO_4832 (O_4832,N_48146,N_49078);
and UO_4833 (O_4833,N_48475,N_48638);
and UO_4834 (O_4834,N_48296,N_49304);
nor UO_4835 (O_4835,N_48496,N_49010);
or UO_4836 (O_4836,N_48805,N_49447);
nor UO_4837 (O_4837,N_49560,N_49642);
nor UO_4838 (O_4838,N_48858,N_49597);
nand UO_4839 (O_4839,N_48864,N_49536);
and UO_4840 (O_4840,N_49608,N_48100);
nor UO_4841 (O_4841,N_48212,N_48932);
or UO_4842 (O_4842,N_49142,N_49250);
or UO_4843 (O_4843,N_49403,N_49183);
nor UO_4844 (O_4844,N_49508,N_48473);
or UO_4845 (O_4845,N_49447,N_49611);
or UO_4846 (O_4846,N_48255,N_49547);
and UO_4847 (O_4847,N_49418,N_48109);
nor UO_4848 (O_4848,N_49058,N_48289);
xor UO_4849 (O_4849,N_48735,N_49191);
or UO_4850 (O_4850,N_49348,N_48682);
xor UO_4851 (O_4851,N_49703,N_49629);
or UO_4852 (O_4852,N_48971,N_49413);
and UO_4853 (O_4853,N_49465,N_49815);
or UO_4854 (O_4854,N_48735,N_49240);
nand UO_4855 (O_4855,N_49625,N_48166);
nand UO_4856 (O_4856,N_48137,N_49470);
xor UO_4857 (O_4857,N_49755,N_48430);
nand UO_4858 (O_4858,N_49398,N_49761);
xor UO_4859 (O_4859,N_49709,N_49813);
and UO_4860 (O_4860,N_48654,N_49620);
and UO_4861 (O_4861,N_49158,N_48778);
and UO_4862 (O_4862,N_49399,N_49113);
nor UO_4863 (O_4863,N_48148,N_49263);
or UO_4864 (O_4864,N_48438,N_48070);
xor UO_4865 (O_4865,N_49626,N_49418);
and UO_4866 (O_4866,N_48703,N_48030);
or UO_4867 (O_4867,N_49971,N_49162);
nor UO_4868 (O_4868,N_48055,N_48631);
xor UO_4869 (O_4869,N_49277,N_49799);
or UO_4870 (O_4870,N_49746,N_48144);
nand UO_4871 (O_4871,N_49350,N_49154);
nor UO_4872 (O_4872,N_48834,N_49989);
nand UO_4873 (O_4873,N_48369,N_48046);
xnor UO_4874 (O_4874,N_48875,N_49442);
xnor UO_4875 (O_4875,N_48104,N_49381);
and UO_4876 (O_4876,N_48451,N_49177);
or UO_4877 (O_4877,N_49330,N_48196);
nor UO_4878 (O_4878,N_48387,N_48860);
nand UO_4879 (O_4879,N_48312,N_49444);
xor UO_4880 (O_4880,N_49078,N_48447);
nand UO_4881 (O_4881,N_49418,N_49785);
nor UO_4882 (O_4882,N_48286,N_49795);
or UO_4883 (O_4883,N_48196,N_48381);
nor UO_4884 (O_4884,N_49401,N_49065);
or UO_4885 (O_4885,N_48294,N_48204);
nand UO_4886 (O_4886,N_48189,N_49206);
xor UO_4887 (O_4887,N_48843,N_48418);
nand UO_4888 (O_4888,N_49444,N_48985);
and UO_4889 (O_4889,N_49210,N_48496);
nor UO_4890 (O_4890,N_49028,N_48878);
and UO_4891 (O_4891,N_48473,N_48063);
or UO_4892 (O_4892,N_49233,N_49844);
or UO_4893 (O_4893,N_48253,N_48215);
or UO_4894 (O_4894,N_48072,N_49025);
nor UO_4895 (O_4895,N_49839,N_49721);
and UO_4896 (O_4896,N_48033,N_49292);
nor UO_4897 (O_4897,N_48432,N_48503);
nand UO_4898 (O_4898,N_48570,N_48934);
xor UO_4899 (O_4899,N_48952,N_49764);
xnor UO_4900 (O_4900,N_49168,N_49995);
or UO_4901 (O_4901,N_48097,N_49857);
nand UO_4902 (O_4902,N_48989,N_48275);
and UO_4903 (O_4903,N_48951,N_49131);
nand UO_4904 (O_4904,N_49315,N_49067);
and UO_4905 (O_4905,N_49942,N_48993);
nor UO_4906 (O_4906,N_48475,N_49412);
nand UO_4907 (O_4907,N_49372,N_49653);
and UO_4908 (O_4908,N_48907,N_49208);
xor UO_4909 (O_4909,N_49963,N_49400);
xor UO_4910 (O_4910,N_48850,N_49615);
xnor UO_4911 (O_4911,N_49316,N_48765);
and UO_4912 (O_4912,N_49371,N_49125);
and UO_4913 (O_4913,N_48756,N_49431);
and UO_4914 (O_4914,N_49808,N_48303);
and UO_4915 (O_4915,N_49380,N_48147);
or UO_4916 (O_4916,N_49202,N_49225);
and UO_4917 (O_4917,N_48787,N_48175);
and UO_4918 (O_4918,N_49643,N_48313);
nand UO_4919 (O_4919,N_49349,N_48900);
nand UO_4920 (O_4920,N_48279,N_49447);
or UO_4921 (O_4921,N_49666,N_48441);
nand UO_4922 (O_4922,N_48021,N_48169);
nand UO_4923 (O_4923,N_48052,N_49608);
nand UO_4924 (O_4924,N_48048,N_49096);
and UO_4925 (O_4925,N_48181,N_49394);
or UO_4926 (O_4926,N_49217,N_48380);
and UO_4927 (O_4927,N_49223,N_49621);
and UO_4928 (O_4928,N_48413,N_49250);
or UO_4929 (O_4929,N_49124,N_49713);
or UO_4930 (O_4930,N_48935,N_48552);
nor UO_4931 (O_4931,N_48925,N_48536);
or UO_4932 (O_4932,N_49617,N_49413);
nor UO_4933 (O_4933,N_48295,N_49400);
nand UO_4934 (O_4934,N_48839,N_49039);
or UO_4935 (O_4935,N_48912,N_48567);
nand UO_4936 (O_4936,N_48846,N_48063);
xnor UO_4937 (O_4937,N_48380,N_49199);
nand UO_4938 (O_4938,N_48007,N_48837);
and UO_4939 (O_4939,N_49936,N_48371);
and UO_4940 (O_4940,N_49998,N_48920);
nor UO_4941 (O_4941,N_49333,N_48737);
nand UO_4942 (O_4942,N_48144,N_49132);
or UO_4943 (O_4943,N_49271,N_49447);
nor UO_4944 (O_4944,N_48302,N_49790);
nand UO_4945 (O_4945,N_49774,N_48355);
and UO_4946 (O_4946,N_48511,N_48975);
nor UO_4947 (O_4947,N_48419,N_49544);
nand UO_4948 (O_4948,N_48357,N_49029);
and UO_4949 (O_4949,N_49954,N_49864);
xor UO_4950 (O_4950,N_49483,N_48409);
nor UO_4951 (O_4951,N_48732,N_49972);
nor UO_4952 (O_4952,N_49581,N_48104);
and UO_4953 (O_4953,N_48504,N_48046);
nand UO_4954 (O_4954,N_49861,N_49615);
nor UO_4955 (O_4955,N_49880,N_49241);
xor UO_4956 (O_4956,N_48048,N_48443);
xnor UO_4957 (O_4957,N_49319,N_49057);
and UO_4958 (O_4958,N_48613,N_48672);
and UO_4959 (O_4959,N_49475,N_49132);
nor UO_4960 (O_4960,N_49307,N_49087);
or UO_4961 (O_4961,N_49598,N_49677);
xnor UO_4962 (O_4962,N_49226,N_48801);
or UO_4963 (O_4963,N_49473,N_48427);
or UO_4964 (O_4964,N_48614,N_48874);
xnor UO_4965 (O_4965,N_49242,N_49471);
xnor UO_4966 (O_4966,N_48550,N_49546);
nor UO_4967 (O_4967,N_48693,N_49986);
xor UO_4968 (O_4968,N_48021,N_49180);
or UO_4969 (O_4969,N_49732,N_49981);
and UO_4970 (O_4970,N_49449,N_48340);
and UO_4971 (O_4971,N_48305,N_48129);
and UO_4972 (O_4972,N_48769,N_49374);
nand UO_4973 (O_4973,N_49229,N_48614);
or UO_4974 (O_4974,N_48067,N_48714);
or UO_4975 (O_4975,N_49482,N_48106);
nor UO_4976 (O_4976,N_48875,N_48866);
or UO_4977 (O_4977,N_48662,N_49685);
or UO_4978 (O_4978,N_49733,N_49099);
or UO_4979 (O_4979,N_49810,N_48161);
and UO_4980 (O_4980,N_49175,N_49084);
or UO_4981 (O_4981,N_48200,N_49241);
xor UO_4982 (O_4982,N_49722,N_48719);
or UO_4983 (O_4983,N_48271,N_49511);
nor UO_4984 (O_4984,N_48748,N_49579);
nand UO_4985 (O_4985,N_48161,N_48414);
nand UO_4986 (O_4986,N_48781,N_48104);
xnor UO_4987 (O_4987,N_48299,N_48209);
or UO_4988 (O_4988,N_48153,N_49040);
nand UO_4989 (O_4989,N_48705,N_49416);
and UO_4990 (O_4990,N_48770,N_48500);
nor UO_4991 (O_4991,N_49083,N_49856);
nand UO_4992 (O_4992,N_48115,N_49691);
or UO_4993 (O_4993,N_48441,N_48994);
xnor UO_4994 (O_4994,N_49336,N_49518);
and UO_4995 (O_4995,N_48109,N_48845);
xor UO_4996 (O_4996,N_49140,N_48155);
and UO_4997 (O_4997,N_49506,N_48193);
or UO_4998 (O_4998,N_49885,N_49139);
nand UO_4999 (O_4999,N_49071,N_48079);
endmodule