module basic_2000_20000_2500_80_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_139,In_1807);
xnor U1 (N_1,In_832,In_1536);
nor U2 (N_2,In_772,In_1234);
and U3 (N_3,In_1425,In_8);
and U4 (N_4,In_837,In_876);
or U5 (N_5,In_456,In_1135);
xor U6 (N_6,In_367,In_1081);
nand U7 (N_7,In_1576,In_778);
xnor U8 (N_8,In_416,In_157);
and U9 (N_9,In_723,In_1609);
nand U10 (N_10,In_1132,In_288);
nand U11 (N_11,In_119,In_1697);
nand U12 (N_12,In_1730,In_1461);
or U13 (N_13,In_373,In_314);
or U14 (N_14,In_1365,In_223);
and U15 (N_15,In_1404,In_1717);
or U16 (N_16,In_1284,In_1847);
or U17 (N_17,In_101,In_506);
nand U18 (N_18,In_1999,In_829);
xor U19 (N_19,In_1995,In_1192);
nand U20 (N_20,In_111,In_1848);
xnor U21 (N_21,In_1016,In_20);
xnor U22 (N_22,In_1194,In_1785);
nand U23 (N_23,In_682,In_516);
nor U24 (N_24,In_287,In_540);
or U25 (N_25,In_1544,In_1187);
and U26 (N_26,In_535,In_366);
and U27 (N_27,In_1923,In_356);
xnor U28 (N_28,In_992,In_951);
and U29 (N_29,In_197,In_53);
and U30 (N_30,In_991,In_1918);
and U31 (N_31,In_1587,In_418);
or U32 (N_32,In_1444,In_907);
nor U33 (N_33,In_1350,In_1331);
or U34 (N_34,In_938,In_150);
or U35 (N_35,In_250,In_461);
nor U36 (N_36,In_1631,In_521);
nand U37 (N_37,In_1176,In_1453);
nor U38 (N_38,In_1156,In_1966);
and U39 (N_39,In_795,In_33);
xor U40 (N_40,In_1754,In_1298);
and U41 (N_41,In_465,In_667);
xor U42 (N_42,In_980,In_495);
and U43 (N_43,In_1314,In_1560);
or U44 (N_44,In_445,In_713);
and U45 (N_45,In_1594,In_91);
and U46 (N_46,In_1709,In_1788);
or U47 (N_47,In_1446,In_344);
or U48 (N_48,In_638,In_700);
and U49 (N_49,In_42,In_1826);
nand U50 (N_50,In_689,In_626);
or U51 (N_51,In_136,In_843);
or U52 (N_52,In_1420,In_668);
nand U53 (N_53,In_811,In_95);
nand U54 (N_54,In_1993,In_72);
nand U55 (N_55,In_1075,In_470);
or U56 (N_56,In_1061,In_327);
nor U57 (N_57,In_168,In_1375);
and U58 (N_58,In_575,In_448);
nor U59 (N_59,In_458,In_1328);
nor U60 (N_60,In_1904,In_1539);
and U61 (N_61,In_972,In_1504);
and U62 (N_62,In_1191,In_192);
nor U63 (N_63,In_391,In_1128);
or U64 (N_64,In_1223,In_1636);
and U65 (N_65,In_1834,In_688);
nand U66 (N_66,In_186,In_1837);
xnor U67 (N_67,In_338,In_1556);
nor U68 (N_68,In_436,In_187);
and U69 (N_69,In_1033,In_612);
nand U70 (N_70,In_1347,In_633);
and U71 (N_71,In_800,In_785);
and U72 (N_72,In_1550,In_381);
nand U73 (N_73,In_1875,In_130);
and U74 (N_74,In_653,In_1805);
nand U75 (N_75,In_697,In_683);
xor U76 (N_76,In_299,In_1217);
or U77 (N_77,In_1242,In_153);
nor U78 (N_78,In_736,In_92);
nand U79 (N_79,In_350,In_580);
and U80 (N_80,In_774,In_1957);
xnor U81 (N_81,In_860,In_547);
and U82 (N_82,In_244,In_698);
nand U83 (N_83,In_218,In_686);
or U84 (N_84,In_452,In_1662);
nand U85 (N_85,In_1116,In_1778);
or U86 (N_86,In_1065,In_1094);
or U87 (N_87,In_372,In_1557);
and U88 (N_88,In_1817,In_3);
xnor U89 (N_89,In_519,In_83);
or U90 (N_90,In_1359,In_1044);
nand U91 (N_91,In_262,In_360);
or U92 (N_92,In_48,In_845);
and U93 (N_93,In_675,In_799);
xnor U94 (N_94,In_681,In_508);
and U95 (N_95,In_1086,In_1341);
xor U96 (N_96,In_896,In_396);
nand U97 (N_97,In_976,In_1253);
and U98 (N_98,In_1189,In_172);
nand U99 (N_99,In_507,In_1278);
xnor U100 (N_100,In_1247,In_1892);
and U101 (N_101,In_304,In_1100);
xor U102 (N_102,In_40,In_1394);
and U103 (N_103,In_1322,In_1275);
or U104 (N_104,In_1407,In_1241);
or U105 (N_105,In_79,In_1197);
nand U106 (N_106,In_1627,In_434);
or U107 (N_107,In_707,In_804);
or U108 (N_108,In_1392,In_1319);
xnor U109 (N_109,In_610,In_909);
nand U110 (N_110,In_430,In_1096);
xnor U111 (N_111,In_657,In_1795);
and U112 (N_112,In_929,In_443);
xor U113 (N_113,In_1027,In_243);
nand U114 (N_114,In_1545,In_676);
xor U115 (N_115,In_517,In_214);
and U116 (N_116,In_859,In_1206);
and U117 (N_117,In_1070,In_1887);
or U118 (N_118,In_1990,In_1614);
nand U119 (N_119,In_16,In_1690);
nand U120 (N_120,In_1751,In_558);
and U121 (N_121,In_1663,In_1437);
xor U122 (N_122,In_395,In_247);
and U123 (N_123,In_1244,In_428);
and U124 (N_124,In_987,In_1260);
or U125 (N_125,In_701,In_858);
nand U126 (N_126,In_363,In_228);
and U127 (N_127,In_1911,In_844);
and U128 (N_128,In_1939,In_1045);
xnor U129 (N_129,In_322,In_1502);
or U130 (N_130,In_1930,In_1926);
nor U131 (N_131,In_1787,In_1962);
xor U132 (N_132,In_311,In_303);
and U133 (N_133,In_892,In_450);
nand U134 (N_134,In_1546,In_114);
or U135 (N_135,In_1162,In_970);
or U136 (N_136,In_213,In_11);
nand U137 (N_137,In_1573,In_968);
or U138 (N_138,In_152,In_920);
xnor U139 (N_139,In_1415,In_1513);
or U140 (N_140,In_961,In_1441);
or U141 (N_141,In_605,In_1749);
nor U142 (N_142,In_971,In_673);
nor U143 (N_143,In_828,In_823);
or U144 (N_144,In_1389,In_273);
nor U145 (N_145,In_1616,In_487);
or U146 (N_146,In_394,In_1956);
nor U147 (N_147,In_1099,In_1903);
and U148 (N_148,In_446,In_725);
xnor U149 (N_149,In_543,In_1948);
and U150 (N_150,In_451,In_1548);
xnor U151 (N_151,In_50,In_1214);
or U152 (N_152,In_234,In_923);
nand U153 (N_153,In_814,In_1764);
and U154 (N_154,In_1882,In_132);
or U155 (N_155,In_1080,In_120);
nand U156 (N_156,In_1280,In_749);
or U157 (N_157,In_661,In_267);
xor U158 (N_158,In_1333,In_146);
or U159 (N_159,In_403,In_1184);
and U160 (N_160,In_998,In_985);
and U161 (N_161,In_1207,In_615);
xor U162 (N_162,In_1091,In_956);
nor U163 (N_163,In_75,In_1756);
or U164 (N_164,In_1257,In_177);
nor U165 (N_165,In_716,In_1179);
or U166 (N_166,In_239,In_622);
and U167 (N_167,In_1225,In_300);
xnor U168 (N_168,In_1929,In_385);
or U169 (N_169,In_1757,In_343);
nand U170 (N_170,In_1023,In_325);
nand U171 (N_171,In_307,In_1797);
nor U172 (N_172,In_313,In_522);
nor U173 (N_173,In_1680,In_1724);
nand U174 (N_174,In_245,In_687);
nor U175 (N_175,In_1079,In_1152);
and U176 (N_176,In_1725,In_1417);
or U177 (N_177,In_1024,In_1927);
nor U178 (N_178,In_1475,In_1133);
and U179 (N_179,In_1373,In_1038);
and U180 (N_180,In_1968,In_1581);
nor U181 (N_181,In_419,In_1564);
nor U182 (N_182,In_265,In_1501);
xor U183 (N_183,In_365,In_1281);
or U184 (N_184,In_1494,In_400);
xor U185 (N_185,In_1014,In_1316);
nor U186 (N_186,In_142,In_1237);
and U187 (N_187,In_1495,In_1409);
and U188 (N_188,In_36,In_207);
xnor U189 (N_189,In_726,In_431);
nor U190 (N_190,In_1822,In_1862);
and U191 (N_191,In_767,In_1050);
and U192 (N_192,In_1025,In_421);
nor U193 (N_193,In_497,In_754);
or U194 (N_194,In_126,In_1170);
or U195 (N_195,In_731,In_252);
nand U196 (N_196,In_379,In_398);
xnor U197 (N_197,In_1674,In_857);
xor U198 (N_198,In_729,In_1411);
or U199 (N_199,In_1367,In_1920);
xnor U200 (N_200,In_1734,In_1589);
nand U201 (N_201,In_1230,In_882);
or U202 (N_202,In_974,In_504);
nand U203 (N_203,In_1507,In_1881);
xnor U204 (N_204,In_108,In_442);
or U205 (N_205,In_1716,In_1036);
nor U206 (N_206,In_989,In_1992);
nor U207 (N_207,In_1173,In_1951);
nor U208 (N_208,In_1533,In_1579);
xor U209 (N_209,In_1028,In_1041);
nand U210 (N_210,In_1547,In_24);
nor U211 (N_211,In_935,In_948);
xnor U212 (N_212,In_251,In_276);
and U213 (N_213,In_1077,In_532);
xor U214 (N_214,In_576,In_341);
and U215 (N_215,In_203,In_335);
and U216 (N_216,In_526,In_55);
xnor U217 (N_217,In_997,In_70);
and U218 (N_218,In_831,In_925);
and U219 (N_219,In_1388,In_1824);
or U220 (N_220,In_1770,In_510);
nor U221 (N_221,In_1396,In_712);
or U222 (N_222,In_1376,In_1928);
xnor U223 (N_223,In_144,In_765);
nor U224 (N_224,In_1226,In_1511);
xor U225 (N_225,In_1888,In_427);
or U226 (N_226,In_1568,In_1413);
and U227 (N_227,In_1597,In_59);
nand U228 (N_228,In_710,In_1098);
nand U229 (N_229,In_1235,In_425);
nor U230 (N_230,In_1043,In_32);
xnor U231 (N_231,In_1739,In_1814);
and U232 (N_232,In_1503,In_815);
and U233 (N_233,In_1378,In_1783);
nand U234 (N_234,In_1048,In_1676);
xnor U235 (N_235,In_1924,In_1781);
nand U236 (N_236,In_794,In_389);
and U237 (N_237,In_460,In_1633);
and U238 (N_238,In_1729,In_1004);
and U239 (N_239,In_1171,In_1186);
and U240 (N_240,In_1440,In_1078);
xor U241 (N_241,In_35,In_1886);
or U242 (N_242,In_714,In_1645);
nand U243 (N_243,In_1895,In_1752);
xor U244 (N_244,In_560,In_1301);
or U245 (N_245,In_639,In_364);
xnor U246 (N_246,In_1285,In_520);
and U247 (N_247,In_1543,In_1800);
and U248 (N_248,In_1919,In_927);
nor U249 (N_249,In_1516,In_1017);
nand U250 (N_250,In_949,In_1753);
nor U251 (N_251,N_22,In_211);
xor U252 (N_252,In_1818,In_836);
nor U253 (N_253,In_1874,In_1653);
and U254 (N_254,In_1371,In_634);
and U255 (N_255,In_1965,In_212);
or U256 (N_256,In_435,In_354);
nand U257 (N_257,In_1514,In_1435);
nor U258 (N_258,In_1733,In_1528);
nand U259 (N_259,In_105,In_1141);
xnor U260 (N_260,In_679,In_1704);
nor U261 (N_261,In_1481,In_808);
nor U262 (N_262,N_175,In_1166);
xnor U263 (N_263,In_1529,In_256);
or U264 (N_264,N_13,In_69);
xnor U265 (N_265,In_337,In_586);
or U266 (N_266,In_1177,In_47);
xor U267 (N_267,In_208,In_1572);
xnor U268 (N_268,In_1908,In_1434);
or U269 (N_269,In_68,In_1710);
and U270 (N_270,In_1719,In_1356);
nor U271 (N_271,In_822,In_1037);
xnor U272 (N_272,In_1821,In_746);
nor U273 (N_273,In_34,In_43);
nand U274 (N_274,In_412,In_1866);
xor U275 (N_275,In_1427,In_724);
xnor U276 (N_276,In_750,In_492);
xnor U277 (N_277,In_1252,N_245);
nand U278 (N_278,N_222,In_764);
and U279 (N_279,In_509,N_28);
nand U280 (N_280,In_577,In_438);
nand U281 (N_281,In_1249,In_1873);
xnor U282 (N_282,In_711,N_238);
nor U283 (N_283,In_359,In_1483);
and U284 (N_284,In_1432,In_382);
or U285 (N_285,In_1088,N_166);
xor U286 (N_286,In_768,In_1212);
xnor U287 (N_287,N_68,In_915);
nand U288 (N_288,In_1022,In_1412);
nor U289 (N_289,In_913,In_810);
nor U290 (N_290,In_1921,In_1269);
xor U291 (N_291,In_637,In_399);
xnor U292 (N_292,In_1354,In_568);
and U293 (N_293,In_1360,In_1891);
xor U294 (N_294,In_1872,In_939);
nor U295 (N_295,In_1638,In_1496);
nand U296 (N_296,In_656,In_1700);
or U297 (N_297,In_1336,N_82);
or U298 (N_298,N_201,In_1932);
nor U299 (N_299,N_91,In_1019);
nand U300 (N_300,In_751,In_1679);
nand U301 (N_301,N_159,In_1711);
nand U302 (N_302,N_21,In_1215);
and U303 (N_303,In_1256,In_141);
or U304 (N_304,In_1468,In_14);
xor U305 (N_305,N_176,In_240);
xor U306 (N_306,In_1598,In_1876);
or U307 (N_307,In_328,In_620);
nor U308 (N_308,In_1899,In_1789);
nor U309 (N_309,In_1001,In_720);
nor U310 (N_310,N_180,In_1870);
nor U311 (N_311,In_690,In_1410);
nand U312 (N_312,In_894,In_1913);
nand U313 (N_313,N_114,N_167);
nor U314 (N_314,In_849,In_706);
nand U315 (N_315,In_691,In_1155);
and U316 (N_316,In_155,In_1900);
xnor U317 (N_317,In_246,In_1964);
and U318 (N_318,In_439,In_1339);
or U319 (N_319,In_1288,In_910);
and U320 (N_320,In_563,In_1276);
nand U321 (N_321,N_64,In_678);
and U322 (N_322,N_7,In_158);
and U323 (N_323,In_854,In_1148);
xnor U324 (N_324,In_1768,In_1279);
xor U325 (N_325,In_937,N_173);
and U326 (N_326,In_693,In_1071);
nand U327 (N_327,In_182,N_37);
nor U328 (N_328,In_1630,In_180);
xor U329 (N_329,In_1213,In_1657);
or U330 (N_330,In_1122,In_318);
nand U331 (N_331,In_73,In_618);
or U332 (N_332,N_67,N_188);
nand U333 (N_333,In_1224,In_23);
nand U334 (N_334,In_566,N_75);
nand U335 (N_335,In_296,In_1562);
or U336 (N_336,In_556,In_1157);
xor U337 (N_337,In_513,In_867);
xor U338 (N_338,In_151,In_1262);
xnor U339 (N_339,In_145,In_1765);
or U340 (N_340,In_1126,In_1426);
and U341 (N_341,In_1403,In_1815);
nand U342 (N_342,In_1448,N_0);
and U343 (N_343,In_826,In_1747);
nand U344 (N_344,In_1622,In_1291);
nor U345 (N_345,In_12,In_1537);
xor U346 (N_346,In_629,In_781);
and U347 (N_347,In_1705,In_596);
nor U348 (N_348,In_1334,In_1666);
and U349 (N_349,In_1541,In_1297);
or U350 (N_350,N_73,In_1332);
xor U351 (N_351,In_1641,In_787);
or U352 (N_352,In_740,In_1474);
and U353 (N_353,In_878,In_775);
nand U354 (N_354,In_1321,In_1853);
xnor U355 (N_355,In_171,In_1844);
and U356 (N_356,In_185,In_874);
xnor U357 (N_357,In_1055,In_1722);
nand U358 (N_358,In_1681,In_1574);
and U359 (N_359,In_1204,N_90);
xor U360 (N_360,In_312,In_94);
and U361 (N_361,In_1784,In_1062);
nor U362 (N_362,In_1060,In_1852);
and U363 (N_363,In_298,In_669);
and U364 (N_364,N_240,In_1151);
and U365 (N_365,In_630,In_226);
and U366 (N_366,In_604,In_699);
or U367 (N_367,N_66,N_204);
nor U368 (N_368,In_756,In_1200);
or U369 (N_369,In_942,In_1344);
nand U370 (N_370,In_643,In_84);
or U371 (N_371,In_198,N_210);
and U372 (N_372,N_70,In_550);
nor U373 (N_373,In_1101,In_1387);
nand U374 (N_374,In_1391,In_1012);
nand U375 (N_375,In_1105,In_1421);
or U376 (N_376,In_1490,In_926);
nand U377 (N_377,In_1652,In_293);
or U378 (N_378,N_41,In_1006);
nor U379 (N_379,In_533,In_1621);
or U380 (N_380,N_83,N_59);
or U381 (N_381,In_478,In_1009);
xnor U382 (N_382,In_202,In_309);
xnor U383 (N_383,N_103,In_283);
nor U384 (N_384,In_784,In_1205);
xnor U385 (N_385,In_397,In_717);
and U386 (N_386,In_319,In_1820);
and U387 (N_387,In_1402,In_1233);
xnor U388 (N_388,In_54,In_229);
nor U389 (N_389,In_762,In_1687);
nor U390 (N_390,N_226,In_217);
or U391 (N_391,In_830,In_1859);
nor U392 (N_392,In_1423,In_289);
nand U393 (N_393,In_1313,In_387);
and U394 (N_394,In_426,In_861);
nor U395 (N_395,In_952,In_869);
nand U396 (N_396,In_1454,In_1185);
xor U397 (N_397,In_993,N_27);
or U398 (N_398,In_1591,In_1610);
xnor U399 (N_399,In_315,In_1985);
nor U400 (N_400,In_565,In_640);
and U401 (N_401,In_17,In_1799);
nor U402 (N_402,N_115,In_1996);
or U403 (N_403,In_255,In_1465);
or U404 (N_404,In_872,In_1330);
and U405 (N_405,In_1248,In_902);
and U406 (N_406,In_1089,In_659);
nand U407 (N_407,In_805,N_77);
nor U408 (N_408,In_1084,In_1527);
and U409 (N_409,In_1129,N_214);
and U410 (N_410,In_1338,In_58);
nand U411 (N_411,In_392,In_413);
or U412 (N_412,In_747,In_1794);
xor U413 (N_413,In_1130,In_1046);
or U414 (N_414,In_248,N_4);
xnor U415 (N_415,In_1885,In_651);
nor U416 (N_416,In_1619,N_156);
xor U417 (N_417,In_1054,In_1819);
and U418 (N_418,In_1561,In_1406);
xor U419 (N_419,In_160,In_1586);
nand U420 (N_420,In_694,In_1526);
and U421 (N_421,In_818,In_1473);
xnor U422 (N_422,In_1210,In_1174);
nand U423 (N_423,In_30,In_9);
nand U424 (N_424,In_1369,In_1082);
nand U425 (N_425,N_6,In_1977);
xor U426 (N_426,In_601,In_1656);
nand U427 (N_427,In_388,In_21);
xnor U428 (N_428,In_931,In_677);
xnor U429 (N_429,In_965,In_1955);
xor U430 (N_430,In_483,In_269);
and U431 (N_431,N_26,N_95);
nor U432 (N_432,N_157,In_880);
nor U433 (N_433,N_126,In_1305);
xor U434 (N_434,In_1042,In_1689);
or U435 (N_435,In_644,In_1917);
nor U436 (N_436,In_227,In_1988);
xor U437 (N_437,In_621,N_242);
xor U438 (N_438,In_1097,In_1104);
nand U439 (N_439,In_1349,In_384);
or U440 (N_440,In_807,In_1505);
nand U441 (N_441,In_31,In_1726);
xnor U442 (N_442,In_25,In_1632);
nor U443 (N_443,In_147,In_1209);
and U444 (N_444,In_1251,In_542);
nor U445 (N_445,In_1601,N_236);
nor U446 (N_446,In_1310,In_888);
nor U447 (N_447,N_218,In_1779);
nor U448 (N_448,In_739,In_129);
nor U449 (N_449,In_1292,In_1792);
nor U450 (N_450,In_1457,In_149);
or U451 (N_451,N_18,In_1307);
nor U452 (N_452,In_1780,N_99);
or U453 (N_453,N_220,In_614);
or U454 (N_454,In_1802,N_160);
nand U455 (N_455,N_78,In_817);
xor U456 (N_456,In_128,In_1868);
and U457 (N_457,In_1487,N_230);
xnor U458 (N_458,In_635,N_224);
or U459 (N_459,In_140,N_174);
nand U460 (N_460,In_1090,In_233);
or U461 (N_461,In_904,In_195);
xor U462 (N_462,In_886,In_77);
xnor U463 (N_463,In_1958,In_1145);
xnor U464 (N_464,In_22,N_154);
or U465 (N_465,N_58,In_221);
xnor U466 (N_466,In_627,N_53);
or U467 (N_467,In_1949,In_969);
xnor U468 (N_468,In_1675,In_1769);
and U469 (N_469,In_986,N_50);
xor U470 (N_470,In_655,In_1637);
nand U471 (N_471,N_197,In_833);
xor U472 (N_472,In_589,In_1740);
and U473 (N_473,In_176,In_1353);
xor U474 (N_474,In_1467,In_231);
nor U475 (N_475,N_232,In_353);
xnor U476 (N_476,In_310,In_561);
xor U477 (N_477,In_1238,In_1981);
or U478 (N_478,In_1571,N_118);
xor U479 (N_479,N_164,In_1743);
nor U480 (N_480,In_1000,In_1879);
and U481 (N_481,In_333,N_190);
nor U482 (N_482,N_216,In_1201);
xnor U483 (N_483,N_212,In_625);
nor U484 (N_484,In_1243,In_1486);
nand U485 (N_485,In_1602,In_777);
and U486 (N_486,N_54,In_613);
or U487 (N_487,In_1290,In_1193);
nand U488 (N_488,In_523,N_110);
xnor U489 (N_489,In_1202,In_464);
nand U490 (N_490,In_743,In_463);
nor U491 (N_491,In_332,In_1345);
nand U492 (N_492,N_165,In_1745);
xor U493 (N_493,In_848,In_237);
nor U494 (N_494,N_87,In_1773);
nor U495 (N_495,In_1865,In_1265);
and U496 (N_496,In_409,In_1715);
nor U497 (N_497,In_454,In_1664);
xnor U498 (N_498,In_170,In_1003);
nor U499 (N_499,In_1693,In_1592);
and U500 (N_500,In_97,In_753);
xor U501 (N_501,In_1030,In_671);
nand U502 (N_502,N_333,N_462);
and U503 (N_503,In_1755,In_1352);
nand U504 (N_504,In_107,In_1500);
nand U505 (N_505,N_241,In_257);
nor U506 (N_506,In_475,In_1216);
xnor U507 (N_507,In_1748,In_1068);
nor U508 (N_508,N_374,In_1005);
nand U509 (N_509,In_903,N_61);
and U510 (N_510,In_124,N_38);
or U511 (N_511,In_1127,In_933);
xor U512 (N_512,In_734,In_1228);
and U513 (N_513,N_31,In_578);
nor U514 (N_514,In_1229,In_49);
xor U515 (N_515,N_52,In_1916);
xor U516 (N_516,In_928,In_444);
nand U517 (N_517,N_403,In_106);
nor U518 (N_518,In_1283,In_1617);
nand U519 (N_519,N_46,In_1855);
and U520 (N_520,In_518,In_1110);
nor U521 (N_521,In_559,In_471);
and U522 (N_522,In_199,In_966);
xnor U523 (N_523,N_217,N_463);
nor U524 (N_524,N_25,N_279);
xnor U525 (N_525,In_1741,In_1357);
or U526 (N_526,N_324,In_26);
xnor U527 (N_527,In_889,In_294);
or U528 (N_528,In_584,In_670);
nor U529 (N_529,In_87,N_171);
xnor U530 (N_530,In_264,In_1240);
nand U531 (N_531,N_256,In_1979);
or U532 (N_532,In_1946,In_1524);
and U533 (N_533,In_1810,In_870);
nand U534 (N_534,In_39,In_912);
xor U535 (N_535,In_1910,In_1976);
xor U536 (N_536,In_1335,In_7);
nand U537 (N_537,In_1830,In_1447);
nor U538 (N_538,In_1414,N_139);
and U539 (N_539,In_1258,In_1106);
and U540 (N_540,In_779,In_1158);
xor U541 (N_541,N_377,In_1020);
xnor U542 (N_542,N_437,In_1118);
or U543 (N_543,N_388,In_1945);
nor U544 (N_544,N_264,In_1239);
nor U545 (N_545,In_1970,In_551);
or U546 (N_546,In_875,In_1849);
or U547 (N_547,In_553,N_301);
nor U548 (N_548,In_840,N_142);
and U549 (N_549,N_475,N_124);
xor U550 (N_550,N_260,In_1850);
and U551 (N_551,In_1460,In_1998);
xor U552 (N_552,In_1940,In_847);
and U553 (N_553,In_1477,In_386);
xor U554 (N_554,In_1067,In_628);
or U555 (N_555,In_1960,In_1018);
or U556 (N_556,N_219,In_1472);
nor U557 (N_557,In_897,In_1076);
and U558 (N_558,N_393,In_1658);
nor U559 (N_559,N_111,In_405);
xor U560 (N_560,In_1655,N_223);
or U561 (N_561,In_63,In_1736);
and U562 (N_562,In_453,In_1218);
nor U563 (N_563,N_10,In_582);
or U564 (N_564,In_838,In_81);
or U565 (N_565,In_685,In_1161);
nand U566 (N_566,In_408,N_372);
xor U567 (N_567,N_102,In_769);
nand U568 (N_568,In_1989,In_719);
xor U569 (N_569,N_383,In_253);
or U570 (N_570,In_1530,N_370);
nor U571 (N_571,In_0,In_268);
or U572 (N_572,In_1914,In_164);
or U573 (N_573,N_398,In_737);
or U574 (N_574,In_631,In_954);
or U575 (N_575,N_72,In_241);
xor U576 (N_576,In_1294,N_117);
xor U577 (N_577,In_1509,In_324);
nor U578 (N_578,In_1603,In_945);
nor U579 (N_579,In_1738,In_1843);
or U580 (N_580,In_1115,In_118);
and U581 (N_581,In_1493,In_362);
or U582 (N_582,In_188,N_291);
xor U583 (N_583,In_1947,In_663);
nor U584 (N_584,In_447,In_205);
and U585 (N_585,N_93,In_1035);
xnor U586 (N_586,N_79,N_255);
and U587 (N_587,In_1801,N_357);
and U588 (N_588,In_215,In_1612);
and U589 (N_589,N_286,In_169);
nor U590 (N_590,In_469,In_1227);
nand U591 (N_591,N_395,N_433);
nor U592 (N_592,N_283,In_744);
or U593 (N_593,N_410,In_1685);
xnor U594 (N_594,N_263,In_1521);
xnor U595 (N_595,In_1140,In_1245);
or U596 (N_596,In_1678,In_1219);
and U597 (N_597,N_243,In_1125);
or U598 (N_598,In_1580,In_321);
nor U599 (N_599,In_85,In_1553);
nand U600 (N_600,In_156,In_133);
nor U601 (N_601,In_865,N_428);
or U602 (N_602,In_1445,In_856);
nor U603 (N_603,In_1464,N_427);
xnor U604 (N_604,N_289,In_567);
and U605 (N_605,In_1827,In_173);
and U606 (N_606,In_181,In_1578);
nor U607 (N_607,N_496,N_489);
nand U608 (N_608,N_490,N_495);
and U609 (N_609,In_664,In_1293);
xor U610 (N_610,N_341,N_48);
nor U611 (N_611,In_455,N_138);
xor U612 (N_612,In_964,In_86);
nor U613 (N_613,In_1400,N_376);
and U614 (N_614,N_334,N_181);
xor U615 (N_615,N_163,N_371);
xnor U616 (N_616,In_806,N_361);
or U617 (N_617,In_988,In_1300);
xnor U618 (N_618,In_930,In_1982);
and U619 (N_619,In_1950,In_1117);
or U620 (N_620,In_1969,In_165);
xnor U621 (N_621,In_1180,In_1484);
nand U622 (N_622,N_155,N_454);
and U623 (N_623,N_74,N_269);
xnor U624 (N_624,In_1701,In_38);
xor U625 (N_625,In_1750,N_69);
nor U626 (N_626,N_487,In_1327);
nor U627 (N_627,N_135,In_1302);
xnor U628 (N_628,In_457,In_1083);
or U629 (N_629,In_752,N_234);
nor U630 (N_630,In_1884,In_1804);
nand U631 (N_631,In_330,N_412);
nor U632 (N_632,In_466,In_718);
and U633 (N_633,N_132,In_329);
nor U634 (N_634,In_1577,In_123);
nand U635 (N_635,N_143,In_738);
nor U636 (N_636,N_396,In_757);
nor U637 (N_637,In_491,N_182);
xor U638 (N_638,N_119,In_1532);
and U639 (N_639,In_745,In_1199);
xor U640 (N_640,In_1361,In_1364);
and U641 (N_641,In_803,N_185);
nor U642 (N_642,N_3,N_258);
or U643 (N_643,In_1540,In_1549);
nand U644 (N_644,N_456,In_1342);
or U645 (N_645,In_357,In_1590);
nor U646 (N_646,In_1554,In_1871);
xnor U647 (N_647,In_1405,In_230);
or U648 (N_648,N_340,In_284);
nor U649 (N_649,In_121,In_674);
nand U650 (N_650,In_1845,N_296);
or U651 (N_651,N_319,In_1618);
nand U652 (N_652,In_1259,In_1190);
xnor U653 (N_653,N_105,N_172);
and U654 (N_654,In_1987,In_1395);
xor U655 (N_655,In_424,In_266);
xor U656 (N_656,In_963,In_429);
and U657 (N_657,N_473,In_786);
xnor U658 (N_658,In_1980,N_448);
and U659 (N_659,N_278,In_790);
or U660 (N_660,In_1836,In_109);
or U661 (N_661,N_71,In_1846);
nor U662 (N_662,In_71,In_474);
and U663 (N_663,In_238,In_573);
nor U664 (N_664,In_484,In_1829);
or U665 (N_665,N_42,In_13);
nor U666 (N_666,In_1123,In_1696);
nor U667 (N_667,In_984,N_129);
nor U668 (N_668,N_316,In_163);
or U669 (N_669,In_1380,N_452);
and U670 (N_670,In_1854,N_128);
nor U671 (N_671,N_295,In_1124);
and U672 (N_672,In_1640,N_418);
nand U673 (N_673,In_1471,In_1732);
or U674 (N_674,In_122,In_918);
and U675 (N_675,In_1142,In_1181);
or U676 (N_676,In_1673,In_1175);
xor U677 (N_677,In_1439,In_742);
nor U678 (N_678,In_1318,N_304);
or U679 (N_679,N_346,N_414);
xnor U680 (N_680,N_12,In_1051);
and U681 (N_681,N_362,In_1032);
nor U682 (N_682,N_310,In_1699);
and U683 (N_683,In_1498,In_1379);
and U684 (N_684,N_320,In_41);
xnor U685 (N_685,In_1299,N_113);
or U686 (N_686,In_479,In_728);
xor U687 (N_687,In_1144,In_1271);
nand U688 (N_688,In_1274,In_1975);
nand U689 (N_689,In_1760,N_24);
nand U690 (N_690,N_125,N_116);
xor U691 (N_691,In_189,In_1497);
and U692 (N_692,N_229,N_411);
and U693 (N_693,In_546,In_1518);
or U694 (N_694,N_49,In_1613);
xnor U695 (N_695,In_901,In_1902);
or U696 (N_696,N_480,In_1172);
nand U697 (N_697,In_1798,In_531);
and U698 (N_698,N_477,N_151);
or U699 (N_699,In_905,N_459);
and U700 (N_700,In_1268,In_704);
nand U701 (N_701,In_376,In_96);
or U702 (N_702,N_209,In_323);
nand U703 (N_703,In_665,In_1066);
and U704 (N_704,N_432,In_179);
and U705 (N_705,N_30,N_472);
or U706 (N_706,In_1761,In_1828);
or U707 (N_707,In_2,In_138);
or U708 (N_708,N_23,In_1644);
nor U709 (N_709,In_654,N_446);
xor U710 (N_710,In_602,In_1470);
xnor U711 (N_711,In_846,In_569);
nor U712 (N_712,N_259,In_1478);
xnor U713 (N_713,In_148,In_572);
xnor U714 (N_714,In_78,N_391);
xor U715 (N_715,N_2,N_43);
and U716 (N_716,In_1232,In_209);
or U717 (N_717,In_1056,In_1763);
nand U718 (N_718,In_459,In_1759);
and U719 (N_719,In_978,In_609);
xnor U720 (N_720,N_248,In_292);
and U721 (N_721,In_496,In_1111);
or U722 (N_722,In_709,In_871);
xor U723 (N_723,N_404,In_850);
or U724 (N_724,In_1838,In_536);
nand U725 (N_725,N_32,N_228);
and U726 (N_726,N_468,N_101);
xor U727 (N_727,In_598,In_358);
and U728 (N_728,In_1491,In_1273);
or U729 (N_729,In_1163,In_527);
and U730 (N_730,In_1665,In_1059);
nand U731 (N_731,In_117,In_1702);
nor U732 (N_732,N_302,N_408);
xor U733 (N_733,N_445,In_1776);
nand U734 (N_734,In_5,In_899);
nand U735 (N_735,In_539,In_1040);
xor U736 (N_736,N_29,N_330);
nor U737 (N_737,N_148,In_680);
nor U738 (N_738,In_1013,In_603);
and U739 (N_739,N_339,N_34);
or U740 (N_740,In_417,In_1137);
or U741 (N_741,In_1650,In_6);
nand U742 (N_742,In_1625,In_37);
nand U743 (N_743,N_327,In_1512);
xnor U744 (N_744,In_134,In_99);
nor U745 (N_745,In_1691,In_1462);
or U746 (N_746,In_619,In_1867);
xor U747 (N_747,N_499,N_356);
nand U748 (N_748,In_1069,In_748);
and U749 (N_749,N_127,In_295);
nor U750 (N_750,In_486,In_1994);
or U751 (N_751,N_566,N_666);
or U752 (N_752,N_97,In_1861);
xor U753 (N_753,In_1456,In_1164);
nor U754 (N_754,N_335,In_1523);
nand U755 (N_755,N_123,In_1306);
or U756 (N_756,In_1905,In_259);
and U757 (N_757,In_225,In_184);
xnor U758 (N_758,In_1723,In_616);
or U759 (N_759,N_554,In_873);
or U760 (N_760,In_1348,In_232);
nor U761 (N_761,In_741,In_1488);
xnor U762 (N_762,In_242,N_406);
or U763 (N_763,In_722,In_175);
and U764 (N_764,N_331,In_502);
nand U765 (N_765,In_1896,In_1346);
and U766 (N_766,In_793,N_63);
or U767 (N_767,In_798,In_236);
or U768 (N_768,N_676,In_1825);
nand U769 (N_769,N_434,In_193);
nand U770 (N_770,N_660,In_76);
and U771 (N_771,N_551,In_868);
and U772 (N_772,In_1295,In_1220);
or U773 (N_773,In_537,In_143);
nand U774 (N_774,In_796,In_1136);
and U775 (N_775,In_361,N_627);
xor U776 (N_776,N_634,In_1774);
or U777 (N_777,In_393,In_641);
nand U778 (N_778,In_1808,In_345);
or U779 (N_779,N_622,In_1329);
or U780 (N_780,In_10,In_316);
nor U781 (N_781,In_1160,N_718);
nand U782 (N_782,N_710,In_1858);
and U783 (N_783,In_773,In_611);
or U784 (N_784,In_1261,In_340);
and U785 (N_785,In_1029,In_646);
or U786 (N_786,N_276,In_1109);
or U787 (N_787,In_410,N_663);
xnor U788 (N_788,In_432,In_552);
nand U789 (N_789,In_587,In_1311);
or U790 (N_790,N_698,In_1131);
nand U791 (N_791,N_658,In_1558);
xnor U792 (N_792,In_1677,In_1583);
or U793 (N_793,N_161,In_308);
xnor U794 (N_794,N_250,In_990);
or U795 (N_795,In_1766,N_497);
nand U796 (N_796,N_645,In_921);
xor U797 (N_797,In_46,In_1355);
nor U798 (N_798,In_821,In_380);
and U799 (N_799,N_237,N_106);
nor U800 (N_800,In_1154,In_528);
and U801 (N_801,N_336,N_585);
nand U802 (N_802,In_1390,In_271);
or U803 (N_803,N_651,N_589);
and U804 (N_804,In_809,In_1431);
or U805 (N_805,In_1277,In_1519);
xnor U806 (N_806,N_614,In_285);
nand U807 (N_807,N_540,In_1011);
or U808 (N_808,In_632,N_415);
and U809 (N_809,In_498,N_17);
xnor U810 (N_810,In_599,N_729);
and U811 (N_811,N_630,In_159);
and U812 (N_812,In_1972,In_1195);
or U813 (N_813,N_380,In_1623);
and U814 (N_814,In_730,In_1198);
nor U815 (N_815,In_511,N_684);
nand U816 (N_816,In_1692,N_274);
nor U817 (N_817,N_519,In_1183);
nor U818 (N_818,In_973,In_1433);
or U819 (N_819,N_369,N_470);
nand U820 (N_820,In_695,In_1422);
xor U821 (N_821,In_881,N_652);
nor U822 (N_822,In_994,In_1264);
nor U823 (N_823,In_883,In_887);
nor U824 (N_824,In_1254,N_583);
and U825 (N_825,In_224,In_64);
nor U826 (N_826,In_1095,In_349);
or U827 (N_827,In_113,In_608);
or U828 (N_828,N_670,In_154);
nand U829 (N_829,N_623,N_130);
nand U830 (N_830,N_112,N_179);
nor U831 (N_831,In_326,N_579);
xnor U832 (N_832,In_249,In_884);
or U833 (N_833,In_623,N_713);
nor U834 (N_834,In_480,In_1007);
xnor U835 (N_835,In_1337,N_390);
nand U836 (N_836,In_346,In_1222);
nor U837 (N_837,In_423,In_1983);
nor U838 (N_838,N_703,N_604);
or U839 (N_839,In_28,N_550);
nand U840 (N_840,N_576,N_624);
nor U841 (N_841,In_895,N_533);
nand U842 (N_842,In_89,In_662);
and U843 (N_843,N_510,N_354);
and U844 (N_844,N_609,N_501);
or U845 (N_845,In_505,In_1894);
nand U846 (N_846,In_274,In_1897);
nor U847 (N_847,In_1525,N_625);
xor U848 (N_848,N_636,In_583);
nand U849 (N_849,In_819,N_607);
or U850 (N_850,In_650,N_695);
xor U851 (N_851,In_692,In_1901);
nand U852 (N_852,N_537,N_741);
nand U853 (N_853,N_261,In_1372);
or U854 (N_854,In_1877,In_222);
nand U855 (N_855,N_401,In_1718);
nand U856 (N_856,In_481,In_441);
and U857 (N_857,In_788,In_1270);
or U858 (N_858,N_581,N_169);
nand U859 (N_859,In_98,In_1864);
nor U860 (N_860,N_712,In_52);
and U861 (N_861,In_161,N_360);
and U862 (N_862,N_471,N_571);
xor U863 (N_863,In_1015,N_685);
nor U864 (N_864,N_665,In_1053);
nand U865 (N_865,N_578,In_1744);
xor U866 (N_866,N_555,In_272);
or U867 (N_867,In_776,N_641);
nor U868 (N_868,N_40,N_257);
or U869 (N_869,In_334,In_1713);
or U870 (N_870,In_1552,N_605);
and U871 (N_871,In_449,N_363);
or U872 (N_872,N_429,In_594);
and U873 (N_873,N_455,N_536);
nor U874 (N_874,N_737,In_62);
or U875 (N_875,In_1997,In_1401);
or U876 (N_876,N_638,N_387);
xnor U877 (N_877,In_863,N_534);
xnor U878 (N_878,N_491,In_1682);
or U879 (N_879,In_1139,In_1728);
xor U880 (N_880,In_1263,In_437);
nand U881 (N_881,In_4,In_1811);
and U882 (N_882,N_313,In_827);
nand U883 (N_883,N_514,N_275);
or U884 (N_884,In_1782,N_465);
and U885 (N_885,In_1660,N_667);
or U886 (N_886,N_426,In_936);
nor U887 (N_887,In_1515,In_1934);
nor U888 (N_888,In_331,In_1635);
nor U889 (N_889,In_879,In_1482);
nor U890 (N_890,N_701,N_120);
nor U891 (N_891,In_975,In_1479);
or U892 (N_892,In_1531,In_853);
nand U893 (N_893,In_88,N_134);
nor U894 (N_894,In_1906,In_1073);
or U895 (N_895,N_669,In_1424);
nand U896 (N_896,N_552,In_1374);
and U897 (N_897,N_569,N_318);
and U898 (N_898,In_297,N_205);
and U899 (N_899,N_521,In_780);
xnor U900 (N_900,In_1624,In_1085);
and U901 (N_901,In_1667,In_1842);
nor U902 (N_902,N_293,In_979);
and U903 (N_903,In_503,N_584);
and U904 (N_904,In_82,In_672);
xor U905 (N_905,In_1397,In_940);
xnor U906 (N_906,In_1510,In_1382);
nand U907 (N_907,N_724,N_62);
nor U908 (N_908,N_206,In_1074);
nand U909 (N_909,N_198,In_1803);
nor U910 (N_910,In_570,In_1121);
xnor U911 (N_911,In_103,In_167);
nand U912 (N_912,In_1708,N_734);
nor U913 (N_913,In_263,In_1315);
or U914 (N_914,In_1031,In_1551);
and U915 (N_915,In_390,N_677);
or U916 (N_916,N_482,In_67);
and U917 (N_917,N_717,In_494);
nor U918 (N_918,In_1694,N_203);
nand U919 (N_919,In_1476,In_1727);
or U920 (N_920,In_1878,N_305);
or U921 (N_921,N_358,N_326);
nor U922 (N_922,In_282,In_607);
and U923 (N_923,In_1775,In_914);
xnor U924 (N_924,In_1368,In_1890);
xnor U925 (N_925,In_590,N_606);
nor U926 (N_926,N_329,In_1064);
nand U927 (N_927,In_1767,N_121);
or U928 (N_928,In_1366,N_280);
nand U929 (N_929,In_1669,In_1385);
and U930 (N_930,N_5,N_251);
or U931 (N_931,In_1535,N_56);
or U932 (N_932,In_1506,In_885);
or U933 (N_933,In_1569,N_610);
or U934 (N_934,In_135,In_1737);
and U935 (N_935,In_1430,N_656);
and U936 (N_936,In_1542,In_65);
nor U937 (N_937,In_996,In_1942);
and U938 (N_938,N_731,N_342);
xnor U939 (N_939,In_1149,In_342);
and U940 (N_940,N_687,In_1272);
or U941 (N_941,N_270,In_983);
or U942 (N_942,N_322,N_478);
or U943 (N_943,In_490,N_588);
or U944 (N_944,In_721,N_266);
nor U945 (N_945,In_1058,N_443);
or U946 (N_946,N_133,N_285);
nor U947 (N_947,N_35,In_658);
or U948 (N_948,In_1841,In_339);
and U949 (N_949,In_1851,N_563);
and U950 (N_950,N_508,N_47);
nand U951 (N_951,In_934,In_708);
nor U952 (N_952,N_509,N_39);
and U953 (N_953,N_568,In_204);
nor U954 (N_954,N_267,N_621);
or U955 (N_955,In_732,N_122);
or U956 (N_956,In_1611,N_547);
nor U957 (N_957,N_744,N_690);
xor U958 (N_958,N_532,In_162);
and U959 (N_959,In_960,N_231);
nor U960 (N_960,N_743,In_562);
nand U961 (N_961,In_137,N_332);
xor U962 (N_962,In_110,In_355);
nor U963 (N_963,N_364,In_950);
nand U964 (N_964,In_1857,N_612);
nand U965 (N_965,In_1021,In_51);
xor U966 (N_966,N_386,N_141);
or U967 (N_967,In_1304,In_1686);
nand U968 (N_968,In_549,In_890);
nor U969 (N_969,In_1777,In_194);
or U970 (N_970,In_735,In_852);
or U971 (N_971,N_504,In_1672);
nand U972 (N_972,In_797,In_1706);
xor U973 (N_973,In_1714,In_1943);
xnor U974 (N_974,In_816,In_1236);
or U975 (N_975,N_338,In_201);
or U976 (N_976,In_1538,In_56);
xor U977 (N_977,N_586,In_834);
nor U978 (N_978,N_170,In_1047);
and U979 (N_979,In_1812,In_1026);
nand U980 (N_980,In_825,N_84);
nand U981 (N_981,In_1762,N_567);
nor U982 (N_982,In_1595,In_1605);
xor U983 (N_983,N_492,In_1296);
and U984 (N_984,N_299,N_647);
or U985 (N_985,N_19,N_506);
or U986 (N_986,In_1959,In_210);
or U987 (N_987,N_615,In_1);
nand U988 (N_988,N_535,N_348);
xnor U989 (N_989,N_575,N_655);
nand U990 (N_990,In_1358,In_1912);
xor U991 (N_991,N_644,In_922);
nor U992 (N_992,In_348,In_1898);
nor U993 (N_993,In_1869,N_45);
xor U994 (N_994,In_74,In_955);
xor U995 (N_995,N_233,In_1282);
or U996 (N_996,In_501,N_715);
xor U997 (N_997,In_1563,In_1167);
nand U998 (N_998,In_941,In_893);
and U999 (N_999,N_692,In_1646);
nand U1000 (N_1000,N_958,In_1114);
xor U1001 (N_1001,In_468,N_344);
and U1002 (N_1002,N_755,N_867);
nand U1003 (N_1003,N_150,In_281);
nand U1004 (N_1004,N_582,N_343);
and U1005 (N_1005,N_952,N_697);
nor U1006 (N_1006,In_727,N_976);
xnor U1007 (N_1007,In_1188,In_1384);
and U1008 (N_1008,N_846,N_539);
nor U1009 (N_1009,In_1991,N_144);
nand U1010 (N_1010,N_137,N_611);
nand U1011 (N_1011,In_1703,In_1585);
xnor U1012 (N_1012,In_1363,In_649);
or U1013 (N_1013,N_277,N_973);
or U1014 (N_1014,N_596,In_125);
or U1015 (N_1015,In_1596,N_460);
and U1016 (N_1016,N_405,In_1639);
and U1017 (N_1017,N_826,N_694);
nand U1018 (N_1018,N_735,N_350);
or U1019 (N_1019,In_383,In_541);
nor U1020 (N_1020,N_423,In_1954);
xor U1021 (N_1021,In_301,N_998);
nand U1022 (N_1022,N_700,In_1182);
or U1023 (N_1023,In_1370,In_112);
or U1024 (N_1024,N_392,N_787);
or U1025 (N_1025,In_302,N_668);
nand U1026 (N_1026,N_811,N_882);
or U1027 (N_1027,N_8,In_488);
xnor U1028 (N_1028,In_1570,N_187);
and U1029 (N_1029,N_881,N_805);
nand U1030 (N_1030,N_732,N_909);
xor U1031 (N_1031,N_966,N_828);
or U1032 (N_1032,In_1628,N_924);
nor U1033 (N_1033,N_708,N_913);
xor U1034 (N_1034,N_594,N_435);
nand U1035 (N_1035,In_1442,N_227);
nand U1036 (N_1036,N_920,N_809);
xor U1037 (N_1037,In_1039,N_945);
xnor U1038 (N_1038,N_671,In_1661);
xor U1039 (N_1039,N_347,N_840);
or U1040 (N_1040,N_733,N_199);
and U1041 (N_1041,N_152,N_851);
nand U1042 (N_1042,N_850,N_832);
or U1043 (N_1043,N_273,N_365);
or U1044 (N_1044,In_660,In_813);
and U1045 (N_1045,N_916,In_116);
xnor U1046 (N_1046,In_18,N_613);
nand U1047 (N_1047,N_253,N_893);
and U1048 (N_1048,N_980,N_936);
and U1049 (N_1049,In_1823,In_19);
nand U1050 (N_1050,N_702,N_545);
xnor U1051 (N_1051,In_1196,In_1103);
or U1052 (N_1052,N_937,In_336);
or U1053 (N_1053,In_898,N_494);
and U1054 (N_1054,In_485,N_894);
and U1055 (N_1055,In_1698,In_1647);
or U1056 (N_1056,N_483,N_810);
and U1057 (N_1057,N_60,N_928);
nand U1058 (N_1058,N_721,In_588);
nand U1059 (N_1059,N_951,In_1325);
nand U1060 (N_1060,N_730,N_899);
nand U1061 (N_1061,In_1648,N_917);
nor U1062 (N_1062,N_440,N_530);
xnor U1063 (N_1063,N_297,N_686);
nand U1064 (N_1064,In_866,N_792);
or U1065 (N_1065,N_89,N_748);
or U1066 (N_1066,N_511,In_1317);
or U1067 (N_1067,N_799,In_919);
and U1068 (N_1068,N_797,N_964);
xnor U1069 (N_1069,N_784,In_1793);
nor U1070 (N_1070,In_761,In_1634);
xnor U1071 (N_1071,In_482,N_654);
xor U1072 (N_1072,In_1984,N_523);
or U1073 (N_1073,In_60,In_924);
nor U1074 (N_1074,In_275,N_824);
nand U1075 (N_1075,N_961,N_562);
nor U1076 (N_1076,In_420,N_716);
xnor U1077 (N_1077,In_351,In_196);
xor U1078 (N_1078,In_414,In_1508);
xnor U1079 (N_1079,N_910,N_874);
xnor U1080 (N_1080,In_1377,N_960);
xnor U1081 (N_1081,N_680,N_312);
nor U1082 (N_1082,N_903,N_294);
nand U1083 (N_1083,N_726,In_770);
xor U1084 (N_1084,N_991,In_851);
and U1085 (N_1085,N_598,In_1499);
nand U1086 (N_1086,In_279,N_76);
nor U1087 (N_1087,In_206,In_1289);
nand U1088 (N_1088,In_953,N_949);
or U1089 (N_1089,In_1922,In_291);
or U1090 (N_1090,In_1416,In_906);
and U1091 (N_1091,N_884,N_308);
nand U1092 (N_1092,N_366,N_757);
and U1093 (N_1093,In_66,In_277);
and U1094 (N_1094,N_593,N_852);
xnor U1095 (N_1095,N_1,N_183);
nor U1096 (N_1096,N_760,N_9);
nand U1097 (N_1097,N_682,In_1399);
xor U1098 (N_1098,In_703,In_557);
nor U1099 (N_1099,In_835,N_430);
and U1100 (N_1100,N_531,N_451);
nand U1101 (N_1101,N_108,In_733);
xor U1102 (N_1102,In_1386,N_886);
or U1103 (N_1103,N_131,N_816);
nor U1104 (N_1104,N_927,In_1567);
or U1105 (N_1105,In_1450,In_591);
nand U1106 (N_1106,In_1323,N_848);
nand U1107 (N_1107,N_857,In_401);
or U1108 (N_1108,N_524,N_254);
nor U1109 (N_1109,In_581,N_517);
or U1110 (N_1110,In_216,In_104);
nor U1111 (N_1111,N_309,N_987);
and U1112 (N_1112,N_661,N_786);
and U1113 (N_1113,In_500,N_572);
xnor U1114 (N_1114,In_967,In_1695);
or U1115 (N_1115,In_1883,In_1436);
and U1116 (N_1116,In_1607,N_616);
and U1117 (N_1117,In_652,In_278);
nand U1118 (N_1118,N_507,In_174);
xnor U1119 (N_1119,N_821,N_727);
nor U1120 (N_1120,In_645,In_1072);
and U1121 (N_1121,N_902,In_127);
nand U1122 (N_1122,N_938,N_885);
nor U1123 (N_1123,In_1168,N_794);
and U1124 (N_1124,N_950,N_962);
nand U1125 (N_1125,N_856,In_1880);
or U1126 (N_1126,N_791,In_1150);
nor U1127 (N_1127,In_1565,In_792);
nand U1128 (N_1128,N_162,In_529);
nor U1129 (N_1129,N_481,N_862);
xnor U1130 (N_1130,In_1489,N_208);
nand U1131 (N_1131,N_880,In_1438);
xor U1132 (N_1132,In_1935,N_995);
or U1133 (N_1133,N_541,N_202);
and U1134 (N_1134,N_970,N_983);
xnor U1135 (N_1135,N_303,In_90);
or U1136 (N_1136,In_1250,N_573);
nand U1137 (N_1137,N_287,N_933);
and U1138 (N_1138,In_1153,In_1816);
nand U1139 (N_1139,N_753,N_85);
nand U1140 (N_1140,N_988,N_823);
nand U1141 (N_1141,In_995,In_317);
xnor U1142 (N_1142,N_518,N_711);
xor U1143 (N_1143,N_835,N_628);
nand U1144 (N_1144,In_1683,N_603);
xnor U1145 (N_1145,N_548,N_795);
nor U1146 (N_1146,In_462,N_485);
xnor U1147 (N_1147,In_286,N_871);
or U1148 (N_1148,In_999,N_629);
or U1149 (N_1149,N_930,N_192);
nand U1150 (N_1150,N_971,In_592);
nand U1151 (N_1151,N_736,N_527);
xnor U1152 (N_1152,In_1455,N_81);
and U1153 (N_1153,In_597,N_762);
xnor U1154 (N_1154,N_929,N_785);
or U1155 (N_1155,N_244,N_956);
and U1156 (N_1156,N_637,N_919);
nand U1157 (N_1157,N_750,In_220);
xor U1158 (N_1158,In_1973,N_829);
and U1159 (N_1159,N_766,N_847);
or U1160 (N_1160,N_86,N_872);
and U1161 (N_1161,N_728,In_1599);
xor U1162 (N_1162,In_771,In_1010);
or U1163 (N_1163,In_514,In_375);
or U1164 (N_1164,In_1915,In_1832);
and U1165 (N_1165,In_473,N_359);
nor U1166 (N_1166,In_1381,N_915);
nand U1167 (N_1167,In_1961,In_1383);
nand U1168 (N_1168,N_808,N_272);
or U1169 (N_1169,In_538,N_770);
nor U1170 (N_1170,In_1398,N_422);
or U1171 (N_1171,N_657,N_107);
or U1172 (N_1172,In_554,N_664);
and U1173 (N_1173,N_146,In_1796);
xnor U1174 (N_1174,In_962,In_1953);
nor U1175 (N_1175,N_402,In_1791);
and U1176 (N_1176,N_186,In_647);
nor U1177 (N_1177,In_545,N_854);
nand U1178 (N_1178,In_1159,N_158);
nand U1179 (N_1179,N_879,In_1735);
and U1180 (N_1180,N_897,In_1651);
or U1181 (N_1181,N_943,In_191);
xor U1182 (N_1182,In_1267,N_963);
nand U1183 (N_1183,In_696,In_1707);
xor U1184 (N_1184,N_836,In_1938);
xnor U1185 (N_1185,In_755,N_968);
nand U1186 (N_1186,N_955,In_1312);
nor U1187 (N_1187,In_1620,In_1340);
nand U1188 (N_1188,N_865,N_561);
xnor U1189 (N_1189,N_855,In_1231);
and U1190 (N_1190,N_746,In_369);
and U1191 (N_1191,In_422,N_355);
and U1192 (N_1192,N_853,In_1907);
and U1193 (N_1193,N_673,N_239);
nand U1194 (N_1194,N_837,In_260);
nor U1195 (N_1195,N_317,N_796);
and U1196 (N_1196,N_774,N_898);
and U1197 (N_1197,N_11,N_271);
nor U1198 (N_1198,N_935,N_252);
nor U1199 (N_1199,In_1119,In_1893);
xor U1200 (N_1200,N_745,In_15);
nor U1201 (N_1201,In_1287,N_265);
nand U1202 (N_1202,N_109,N_870);
and U1203 (N_1203,In_982,In_1266);
or U1204 (N_1204,N_802,In_1246);
nor U1205 (N_1205,In_1629,In_763);
nand U1206 (N_1206,N_20,In_1831);
or U1207 (N_1207,N_681,N_947);
nor U1208 (N_1208,N_353,N_147);
xnor U1209 (N_1209,N_833,In_467);
nand U1210 (N_1210,In_1458,In_593);
xor U1211 (N_1211,In_1534,N_675);
and U1212 (N_1212,N_136,N_100);
or U1213 (N_1213,N_488,N_476);
or U1214 (N_1214,In_1671,In_1517);
xnor U1215 (N_1215,In_371,In_1452);
xor U1216 (N_1216,In_1860,N_442);
xor U1217 (N_1217,N_775,In_1459);
nand U1218 (N_1218,N_436,In_29);
and U1219 (N_1219,N_194,N_542);
xnor U1220 (N_1220,N_761,N_619);
nor U1221 (N_1221,N_557,N_764);
nor U1222 (N_1222,N_325,N_822);
xnor U1223 (N_1223,In_959,In_1684);
nor U1224 (N_1224,N_560,In_636);
and U1225 (N_1225,In_377,N_516);
or U1226 (N_1226,N_860,N_866);
xor U1227 (N_1227,In_347,In_1326);
or U1228 (N_1228,N_546,In_617);
nor U1229 (N_1229,N_876,N_246);
and U1230 (N_1230,N_994,N_15);
nand U1231 (N_1231,In_760,In_1418);
or U1232 (N_1232,N_486,In_544);
xnor U1233 (N_1233,In_1555,In_1419);
and U1234 (N_1234,N_740,In_512);
nand U1235 (N_1235,N_351,In_534);
nand U1236 (N_1236,N_688,N_600);
nor U1237 (N_1237,N_887,N_969);
nor U1238 (N_1238,N_861,N_691);
xor U1239 (N_1239,N_450,N_502);
xor U1240 (N_1240,N_177,In_1057);
or U1241 (N_1241,In_600,N_104);
or U1242 (N_1242,N_268,N_617);
and U1243 (N_1243,N_444,In_433);
and U1244 (N_1244,In_1712,In_1087);
or U1245 (N_1245,N_849,N_397);
and U1246 (N_1246,N_33,In_1008);
xor U1247 (N_1247,N_314,In_791);
and U1248 (N_1248,In_574,N_590);
nor U1249 (N_1249,N_597,In_270);
and U1250 (N_1250,In_1492,N_479);
xor U1251 (N_1251,N_709,N_986);
or U1252 (N_1252,N_306,N_1082);
nand U1253 (N_1253,In_1522,N_1130);
or U1254 (N_1254,In_766,In_1604);
nor U1255 (N_1255,N_321,N_1047);
and U1256 (N_1256,N_912,In_1967);
nand U1257 (N_1257,N_807,N_1145);
xor U1258 (N_1258,N_168,In_1221);
xnor U1259 (N_1259,N_633,N_864);
nor U1260 (N_1260,N_984,N_599);
or U1261 (N_1261,N_941,N_1232);
or U1262 (N_1262,N_1179,N_1111);
xor U1263 (N_1263,N_379,N_714);
nand U1264 (N_1264,N_831,N_1188);
and U1265 (N_1265,In_1575,In_1615);
xnor U1266 (N_1266,N_1131,In_477);
or U1267 (N_1267,In_571,N_738);
nand U1268 (N_1268,N_323,N_553);
and U1269 (N_1269,In_1520,N_300);
xnor U1270 (N_1270,In_1909,N_1108);
nor U1271 (N_1271,N_1033,N_1199);
nor U1272 (N_1272,N_94,N_839);
xnor U1273 (N_1273,N_55,N_1072);
nand U1274 (N_1274,In_981,N_1168);
and U1275 (N_1275,N_999,N_1016);
or U1276 (N_1276,N_895,N_1248);
nand U1277 (N_1277,In_1211,N_1240);
xnor U1278 (N_1278,In_1790,In_1731);
xnor U1279 (N_1279,In_320,In_1659);
nor U1280 (N_1280,N_1156,In_1308);
nand U1281 (N_1281,N_1022,N_1230);
nand U1282 (N_1282,In_839,N_1162);
nor U1283 (N_1283,N_580,In_1143);
nor U1284 (N_1284,N_1216,In_782);
and U1285 (N_1285,N_768,N_1134);
nand U1286 (N_1286,N_813,N_1133);
and U1287 (N_1287,In_1840,N_896);
or U1288 (N_1288,In_1606,N_515);
nor U1289 (N_1289,N_674,N_461);
xnor U1290 (N_1290,N_1083,N_281);
xor U1291 (N_1291,N_544,In_684);
xor U1292 (N_1292,In_957,In_1978);
and U1293 (N_1293,N_1245,N_16);
and U1294 (N_1294,N_1193,N_689);
and U1295 (N_1295,N_1106,N_1170);
nor U1296 (N_1296,N_193,N_820);
nand U1297 (N_1297,N_1023,N_1005);
nand U1298 (N_1298,In_368,N_153);
or U1299 (N_1299,In_855,N_595);
nor U1300 (N_1300,In_1034,In_178);
or U1301 (N_1301,In_1351,N_982);
or U1302 (N_1302,N_1122,N_1173);
nor U1303 (N_1303,N_1097,In_1600);
nand U1304 (N_1304,N_1178,In_27);
or U1305 (N_1305,N_772,N_1004);
nand U1306 (N_1306,N_513,N_413);
and U1307 (N_1307,In_131,N_178);
or U1308 (N_1308,N_1217,N_932);
or U1309 (N_1309,N_843,N_1086);
nand U1310 (N_1310,N_1049,N_453);
or U1311 (N_1311,In_1303,N_558);
or U1312 (N_1312,In_1102,N_145);
or U1313 (N_1313,In_306,In_715);
nor U1314 (N_1314,N_1075,N_1109);
and U1315 (N_1315,N_1092,N_1114);
or U1316 (N_1316,N_779,In_842);
or U1317 (N_1317,N_526,N_564);
nor U1318 (N_1318,N_926,N_1195);
nor U1319 (N_1319,In_1466,N_1222);
and U1320 (N_1320,N_407,N_1206);
and U1321 (N_1321,N_345,In_1582);
xnor U1322 (N_1322,N_977,N_1045);
or U1323 (N_1323,In_1835,In_261);
nor U1324 (N_1324,N_1159,In_1608);
or U1325 (N_1325,In_524,N_1095);
nand U1326 (N_1326,N_464,N_1078);
and U1327 (N_1327,In_1971,In_1092);
nor U1328 (N_1328,N_1201,In_606);
nand U1329 (N_1329,In_200,N_1040);
or U1330 (N_1330,In_1721,N_974);
nand U1331 (N_1331,N_570,N_981);
or U1332 (N_1332,N_543,N_1196);
xor U1333 (N_1333,N_948,N_782);
nor U1334 (N_1334,In_493,N_650);
xnor U1335 (N_1335,N_457,N_1001);
and U1336 (N_1336,In_1451,N_922);
nand U1337 (N_1337,In_45,N_1090);
or U1338 (N_1338,N_722,N_592);
and U1339 (N_1339,N_1129,N_918);
nor U1340 (N_1340,N_1154,N_806);
nor U1341 (N_1341,In_476,N_771);
nor U1342 (N_1342,N_635,N_1091);
xnor U1343 (N_1343,N_1017,N_1115);
and U1344 (N_1344,N_1198,N_196);
nand U1345 (N_1345,N_900,In_1933);
nand U1346 (N_1346,N_1175,In_579);
xor U1347 (N_1347,In_1093,N_1057);
nor U1348 (N_1348,N_723,N_725);
nand U1349 (N_1349,In_944,N_439);
xnor U1350 (N_1350,In_1944,N_416);
and U1351 (N_1351,N_1180,N_381);
nor U1352 (N_1352,N_368,In_1643);
xor U1353 (N_1353,In_1649,N_1066);
xnor U1354 (N_1354,N_1050,N_1241);
and U1355 (N_1355,N_817,N_211);
and U1356 (N_1356,In_411,In_783);
nand U1357 (N_1357,N_1080,N_421);
and U1358 (N_1358,N_1079,N_195);
and U1359 (N_1359,N_907,In_1255);
nor U1360 (N_1360,N_1026,In_916);
xor U1361 (N_1361,N_1074,N_706);
nor U1362 (N_1362,N_1085,In_1771);
or U1363 (N_1363,In_254,N_906);
xor U1364 (N_1364,N_696,N_1152);
and U1365 (N_1365,In_1485,In_911);
xnor U1366 (N_1366,N_618,N_1010);
or U1367 (N_1367,In_80,In_1138);
xor U1368 (N_1368,N_747,N_939);
or U1369 (N_1369,N_756,N_207);
nor U1370 (N_1370,In_407,In_946);
xnor U1371 (N_1371,N_1117,N_1103);
or U1372 (N_1372,N_1064,N_315);
nand U1373 (N_1373,N_863,In_820);
or U1374 (N_1374,In_1720,N_925);
and U1375 (N_1375,N_298,N_921);
xor U1376 (N_1376,N_262,In_802);
xnor U1377 (N_1377,N_1031,N_1204);
xnor U1378 (N_1378,N_1249,N_1120);
nor U1379 (N_1379,N_1096,N_1144);
nor U1380 (N_1380,N_1044,N_474);
and U1381 (N_1381,N_337,N_878);
nand U1382 (N_1382,N_672,In_115);
nand U1383 (N_1383,N_965,In_1208);
or U1384 (N_1384,In_1772,N_601);
nand U1385 (N_1385,N_1116,In_1963);
nand U1386 (N_1386,N_1028,N_972);
xor U1387 (N_1387,N_1006,N_662);
xor U1388 (N_1388,N_1185,N_993);
nand U1389 (N_1389,N_1073,N_1052);
nor U1390 (N_1390,In_555,N_1148);
nand U1391 (N_1391,N_1228,In_352);
and U1392 (N_1392,In_374,N_818);
nor U1393 (N_1393,In_1742,N_500);
nand U1394 (N_1394,N_1246,N_1166);
xnor U1395 (N_1395,N_1140,N_841);
and U1396 (N_1396,N_1211,N_763);
and U1397 (N_1397,N_1226,N_441);
or U1398 (N_1398,N_1142,In_290);
and U1399 (N_1399,N_1242,N_1183);
or U1400 (N_1400,N_1042,N_905);
or U1401 (N_1401,In_404,In_440);
nor U1402 (N_1402,N_1099,N_1181);
nand U1403 (N_1403,N_1169,N_1186);
and U1404 (N_1404,N_800,In_1320);
nor U1405 (N_1405,N_1055,N_1190);
or U1406 (N_1406,N_498,N_990);
or U1407 (N_1407,N_754,In_1833);
and U1408 (N_1408,N_804,N_307);
xor U1409 (N_1409,N_975,N_705);
and U1410 (N_1410,N_528,N_749);
nor U1411 (N_1411,N_538,N_505);
nand U1412 (N_1412,N_1110,N_842);
nor U1413 (N_1413,In_1480,In_406);
xnor U1414 (N_1414,N_992,N_1219);
or U1415 (N_1415,In_1362,N_1032);
nand U1416 (N_1416,N_399,In_1668);
nand U1417 (N_1417,N_776,N_1127);
nand U1418 (N_1418,In_1107,N_1012);
nor U1419 (N_1419,N_419,N_653);
nor U1420 (N_1420,N_953,In_93);
nand U1421 (N_1421,N_1089,N_931);
and U1422 (N_1422,N_378,N_1236);
nor U1423 (N_1423,In_1113,N_1107);
or U1424 (N_1424,N_1149,N_382);
and U1425 (N_1425,N_36,N_1136);
nand U1426 (N_1426,In_877,N_1084);
or U1427 (N_1427,N_1202,N_901);
nor U1428 (N_1428,N_1141,N_914);
or U1429 (N_1429,N_1003,N_559);
nor U1430 (N_1430,N_699,N_1112);
nor U1431 (N_1431,In_1670,N_1172);
or U1432 (N_1432,N_1194,N_679);
or U1433 (N_1433,N_1247,N_1157);
nor U1434 (N_1434,N_923,N_1205);
or U1435 (N_1435,N_859,N_892);
nand U1436 (N_1436,In_1146,N_1087);
or U1437 (N_1437,N_1203,N_1015);
or U1438 (N_1438,N_1243,N_367);
xnor U1439 (N_1439,N_1121,In_1134);
and U1440 (N_1440,N_469,In_1443);
nor U1441 (N_1441,N_707,N_556);
nand U1442 (N_1442,N_1177,N_1176);
nand U1443 (N_1443,N_1174,In_280);
nor U1444 (N_1444,In_102,In_1429);
xnor U1445 (N_1445,In_1002,N_888);
nor U1446 (N_1446,In_977,N_602);
nor U1447 (N_1447,In_1936,In_44);
and U1448 (N_1448,N_98,N_394);
xor U1449 (N_1449,N_1014,In_1952);
nor U1450 (N_1450,In_585,N_1046);
nand U1451 (N_1451,N_1123,In_900);
xnor U1452 (N_1452,N_844,N_1182);
nand U1453 (N_1453,In_1463,In_1839);
nand U1454 (N_1454,N_659,N_1126);
xor U1455 (N_1455,N_1207,N_825);
and U1456 (N_1456,In_1108,N_1065);
or U1457 (N_1457,N_1125,N_959);
nor U1458 (N_1458,N_1009,N_1008);
or U1459 (N_1459,In_1856,N_793);
xnor U1460 (N_1460,N_1061,N_868);
nor U1461 (N_1461,N_1034,N_827);
nor U1462 (N_1462,N_1036,In_305);
or U1463 (N_1463,N_814,In_564);
nor U1464 (N_1464,In_1469,N_1100);
xnor U1465 (N_1465,N_1143,N_942);
or U1466 (N_1466,N_352,N_249);
nand U1467 (N_1467,N_80,N_719);
and U1468 (N_1468,In_1120,N_1020);
xnor U1469 (N_1469,In_1588,In_624);
nand U1470 (N_1470,N_781,In_1559);
or U1471 (N_1471,N_1164,In_702);
xnor U1472 (N_1472,N_1118,In_908);
nand U1473 (N_1473,In_1147,N_385);
and U1474 (N_1474,N_425,N_1231);
nor U1475 (N_1475,N_801,N_1038);
and U1476 (N_1476,In_61,In_1813);
or U1477 (N_1477,N_979,N_1160);
nor U1478 (N_1478,N_1102,N_140);
and U1479 (N_1479,N_1124,N_1013);
and U1480 (N_1480,N_997,N_1088);
or U1481 (N_1481,N_693,N_1209);
nand U1482 (N_1482,N_92,N_765);
xnor U1483 (N_1483,N_812,N_1150);
and U1484 (N_1484,N_1237,N_1235);
or U1485 (N_1485,N_891,N_520);
nor U1486 (N_1486,N_400,In_1324);
nand U1487 (N_1487,N_1225,N_1002);
and U1488 (N_1488,In_1626,N_1229);
nand U1489 (N_1489,N_1210,N_57);
or U1490 (N_1490,N_631,N_819);
nand U1491 (N_1491,N_632,In_958);
or U1492 (N_1492,In_812,N_389);
xor U1493 (N_1493,In_258,N_1054);
or U1494 (N_1494,N_467,N_1223);
xor U1495 (N_1495,N_704,In_530);
xnor U1496 (N_1496,N_1068,N_780);
and U1497 (N_1497,N_1024,N_1077);
xor U1498 (N_1498,N_1011,N_549);
nand U1499 (N_1499,N_1138,In_1566);
nand U1500 (N_1500,N_683,N_1367);
nor U1501 (N_1501,N_649,N_1424);
or U1502 (N_1502,In_235,In_1593);
xor U1503 (N_1503,N_438,N_1213);
nor U1504 (N_1504,N_574,N_1030);
and U1505 (N_1505,N_1289,N_1317);
xor U1506 (N_1506,N_815,N_752);
xnor U1507 (N_1507,In_1937,N_1406);
nor U1508 (N_1508,N_1362,In_666);
or U1509 (N_1509,N_1490,N_373);
or U1510 (N_1510,N_1187,N_1270);
and U1511 (N_1511,N_911,N_1264);
and U1512 (N_1512,N_1266,N_1200);
nor U1513 (N_1513,N_1376,N_1421);
nand U1514 (N_1514,N_1304,N_1007);
xor U1515 (N_1515,N_1293,N_1056);
nor U1516 (N_1516,N_1352,N_1340);
nand U1517 (N_1517,N_1286,N_751);
xnor U1518 (N_1518,In_1746,N_996);
and U1519 (N_1519,N_1262,N_1416);
nand U1520 (N_1520,In_1809,N_1476);
xnor U1521 (N_1521,N_1462,N_1184);
nor U1522 (N_1522,N_1482,N_1439);
and U1523 (N_1523,N_1335,N_1487);
xor U1524 (N_1524,N_1301,N_65);
and U1525 (N_1525,N_1390,N_1290);
or U1526 (N_1526,N_149,N_1239);
and U1527 (N_1527,N_1428,N_620);
nor U1528 (N_1528,N_1358,N_1330);
and U1529 (N_1529,N_1444,N_1161);
and U1530 (N_1530,N_1491,N_1244);
and U1531 (N_1531,N_1324,N_1051);
nand U1532 (N_1532,N_1283,N_1468);
nor U1533 (N_1533,N_1039,N_1474);
xor U1534 (N_1534,N_1062,In_378);
nand U1535 (N_1535,N_1385,N_587);
or U1536 (N_1536,N_1450,In_1169);
nor U1537 (N_1537,N_1167,N_458);
and U1538 (N_1538,N_1261,N_1437);
nor U1539 (N_1539,N_1018,N_985);
nor U1540 (N_1540,N_1191,N_1325);
or U1541 (N_1541,N_858,N_1105);
and U1542 (N_1542,N_940,N_1446);
or U1543 (N_1543,N_1430,N_311);
xor U1544 (N_1544,N_978,N_1479);
or U1545 (N_1545,N_1292,N_1272);
nor U1546 (N_1546,N_1274,N_1067);
or U1547 (N_1547,In_1408,N_1360);
or U1548 (N_1548,N_1025,N_946);
nor U1549 (N_1549,N_1392,N_1321);
and U1550 (N_1550,N_1461,In_943);
and U1551 (N_1551,N_51,N_1275);
and U1552 (N_1552,N_290,In_1941);
nor U1553 (N_1553,In_824,N_1492);
nand U1554 (N_1554,N_1346,N_1485);
and U1555 (N_1555,N_292,N_1258);
and U1556 (N_1556,In_1863,N_1280);
nand U1557 (N_1557,In_402,N_1238);
or U1558 (N_1558,N_1401,N_1267);
and U1559 (N_1559,N_742,N_1147);
nor U1560 (N_1560,N_1396,N_1171);
xnor U1561 (N_1561,In_841,N_1254);
nor U1562 (N_1562,N_1441,In_1889);
and U1563 (N_1563,N_1494,N_1497);
or U1564 (N_1564,N_1000,N_1489);
nand U1565 (N_1565,N_1282,N_1155);
nor U1566 (N_1566,N_1053,N_758);
nor U1567 (N_1567,N_944,N_1336);
or U1568 (N_1568,N_957,N_1460);
nand U1569 (N_1569,N_1398,N_1364);
nand U1570 (N_1570,N_1347,N_1305);
nand U1571 (N_1571,N_954,In_1786);
and U1572 (N_1572,N_247,N_1415);
or U1573 (N_1573,N_967,N_1448);
xor U1574 (N_1574,N_1281,In_1165);
or U1575 (N_1575,N_1456,N_1297);
xnor U1576 (N_1576,N_1455,N_759);
xnor U1577 (N_1577,In_499,N_1343);
or U1578 (N_1578,N_1119,N_1291);
or U1579 (N_1579,N_349,In_595);
or U1580 (N_1580,N_1383,N_1417);
and U1581 (N_1581,N_1334,N_1273);
and U1582 (N_1582,N_1356,N_284);
and U1583 (N_1583,N_1158,N_1379);
xor U1584 (N_1584,N_1377,N_1329);
and U1585 (N_1585,N_529,N_1477);
and U1586 (N_1586,N_1309,In_1286);
or U1587 (N_1587,In_1925,N_1464);
or U1588 (N_1588,N_1483,N_1372);
and U1589 (N_1589,N_875,N_1279);
nor U1590 (N_1590,N_1069,N_44);
xnor U1591 (N_1591,In_891,N_1451);
nor U1592 (N_1592,In_862,N_420);
nand U1593 (N_1593,N_790,N_512);
nand U1594 (N_1594,N_838,N_1374);
and U1595 (N_1595,N_1313,N_1373);
xnor U1596 (N_1596,N_1486,N_1197);
nor U1597 (N_1597,In_801,N_1423);
xnor U1598 (N_1598,In_219,In_166);
nand U1599 (N_1599,N_1370,In_190);
nor U1600 (N_1600,N_1440,N_1308);
nor U1601 (N_1601,In_648,In_489);
nor U1602 (N_1602,N_1499,N_1354);
nor U1603 (N_1603,N_1422,N_1378);
nor U1604 (N_1604,N_1471,In_1758);
nand U1605 (N_1605,N_1412,N_1447);
or U1606 (N_1606,N_873,N_1063);
and U1607 (N_1607,N_1250,N_1113);
nand U1608 (N_1608,N_1041,N_565);
or U1609 (N_1609,N_1382,N_1255);
nor U1610 (N_1610,N_591,N_1420);
or U1611 (N_1611,In_1049,N_1463);
nand U1612 (N_1612,N_1333,In_1178);
nor U1613 (N_1613,In_1203,N_1350);
xor U1614 (N_1614,N_1218,N_1408);
xor U1615 (N_1615,N_1263,N_1331);
or U1616 (N_1616,N_1429,N_1189);
xnor U1617 (N_1617,N_640,N_1480);
or U1618 (N_1618,N_642,N_417);
nand U1619 (N_1619,N_1251,N_525);
or U1620 (N_1620,N_1233,N_1434);
and U1621 (N_1621,In_1688,N_1214);
and U1622 (N_1622,N_1453,N_1137);
xor U1623 (N_1623,N_1081,In_1428);
or U1624 (N_1624,In_525,N_1278);
xnor U1625 (N_1625,N_1470,N_424);
xor U1626 (N_1626,In_917,N_1443);
or U1627 (N_1627,N_1227,N_1284);
nor U1628 (N_1628,N_466,N_1027);
xnor U1629 (N_1629,N_1436,N_1271);
or U1630 (N_1630,N_845,N_1320);
xor U1631 (N_1631,N_1224,N_1493);
nor U1632 (N_1632,N_1365,N_577);
xor U1633 (N_1633,In_1112,N_1132);
and U1634 (N_1634,N_1043,N_1466);
xor U1635 (N_1635,N_1475,N_834);
nor U1636 (N_1636,N_639,N_189);
nand U1637 (N_1637,N_908,N_1488);
nand U1638 (N_1638,N_1288,N_1393);
xor U1639 (N_1639,N_1410,N_1498);
and U1640 (N_1640,N_1318,N_1345);
nand U1641 (N_1641,N_1151,N_1265);
nor U1642 (N_1642,N_626,N_1391);
nand U1643 (N_1643,N_1234,N_1035);
or U1644 (N_1644,N_1426,N_1357);
xnor U1645 (N_1645,N_1029,N_384);
and U1646 (N_1646,N_431,N_648);
or U1647 (N_1647,N_1326,N_1071);
nand U1648 (N_1648,N_1298,N_184);
xnor U1649 (N_1649,N_643,N_1019);
or U1650 (N_1650,N_869,N_1432);
nand U1651 (N_1651,N_1319,N_1277);
and U1652 (N_1652,N_1253,In_932);
or U1653 (N_1653,N_1394,N_1413);
nor U1654 (N_1654,N_1403,In_415);
or U1655 (N_1655,N_88,N_1467);
nand U1656 (N_1656,N_1449,N_1355);
nor U1657 (N_1657,N_1388,N_1359);
xnor U1658 (N_1658,In_947,N_1060);
or U1659 (N_1659,N_1427,N_1306);
nand U1660 (N_1660,In_1449,N_1276);
and U1661 (N_1661,N_503,N_1307);
xnor U1662 (N_1662,N_282,N_1215);
xor U1663 (N_1663,In_370,N_1348);
nor U1664 (N_1664,N_235,N_1296);
nor U1665 (N_1665,N_798,N_1294);
or U1666 (N_1666,N_1349,In_758);
nand U1667 (N_1667,N_1295,In_1986);
nand U1668 (N_1668,N_1310,N_1351);
nand U1669 (N_1669,In_1642,N_1104);
nand U1670 (N_1670,N_225,N_1386);
nor U1671 (N_1671,N_877,N_883);
or U1672 (N_1672,In_1063,N_720);
xor U1673 (N_1673,N_1478,N_1472);
and U1674 (N_1674,N_1419,N_789);
nor U1675 (N_1675,N_1058,N_1220);
nor U1676 (N_1676,N_989,N_447);
or U1677 (N_1677,N_830,N_1404);
nand U1678 (N_1678,N_1135,N_1369);
nand U1679 (N_1679,N_788,N_1363);
nand U1680 (N_1680,N_1153,N_1381);
nand U1681 (N_1681,In_1052,N_191);
xnor U1682 (N_1682,N_1344,N_1400);
nand U1683 (N_1683,N_1314,N_1311);
xor U1684 (N_1684,N_1375,N_1315);
xor U1685 (N_1685,In_548,N_449);
xor U1686 (N_1686,N_1021,N_375);
and U1687 (N_1687,N_1452,N_1192);
nand U1688 (N_1688,N_1312,In_1654);
or U1689 (N_1689,N_1128,N_1212);
nor U1690 (N_1690,N_1361,In_472);
or U1691 (N_1691,In_1931,N_1384);
and U1692 (N_1692,N_1322,In_1806);
xor U1693 (N_1693,N_1442,N_1208);
nor U1694 (N_1694,In_705,N_1405);
and U1695 (N_1695,In_57,N_1414);
and U1696 (N_1696,N_739,N_1407);
and U1697 (N_1697,N_1465,N_1303);
or U1698 (N_1698,N_1287,In_864);
xor U1699 (N_1699,In_100,N_1328);
or U1700 (N_1700,N_1146,N_1418);
or U1701 (N_1701,N_1469,N_1048);
and U1702 (N_1702,N_1059,N_767);
or U1703 (N_1703,N_1454,N_522);
xnor U1704 (N_1704,N_200,N_1425);
nor U1705 (N_1705,N_1397,N_803);
nand U1706 (N_1706,N_773,N_14);
or U1707 (N_1707,N_1332,In_789);
nor U1708 (N_1708,N_96,N_1402);
or U1709 (N_1709,N_904,In_515);
or U1710 (N_1710,N_1285,N_1484);
nand U1711 (N_1711,N_777,N_1094);
or U1712 (N_1712,N_1496,N_1327);
xor U1713 (N_1713,N_328,In_1393);
nor U1714 (N_1714,N_213,N_1409);
or U1715 (N_1715,N_1323,In_642);
nand U1716 (N_1716,N_493,N_1380);
nor U1717 (N_1717,N_1268,In_1584);
and U1718 (N_1718,N_1338,N_1252);
or U1719 (N_1719,N_1371,N_1098);
or U1720 (N_1720,N_1457,N_934);
or U1721 (N_1721,N_1260,N_1259);
xor U1722 (N_1722,N_1395,N_769);
or U1723 (N_1723,N_1411,N_1093);
nand U1724 (N_1724,N_1445,N_1353);
nor U1725 (N_1725,N_484,N_1337);
nand U1726 (N_1726,N_1302,N_1037);
or U1727 (N_1727,In_759,N_889);
xor U1728 (N_1728,N_1256,N_1070);
and U1729 (N_1729,N_409,In_1974);
and U1730 (N_1730,N_890,N_646);
and U1731 (N_1731,N_1366,N_1368);
or U1732 (N_1732,In_1343,N_1221);
nand U1733 (N_1733,N_608,N_1458);
xor U1734 (N_1734,N_1473,N_1459);
nor U1735 (N_1735,N_1269,N_1339);
nor U1736 (N_1736,N_1438,N_1435);
and U1737 (N_1737,N_1139,N_1341);
or U1738 (N_1738,In_183,N_1076);
or U1739 (N_1739,N_1431,N_1257);
xnor U1740 (N_1740,N_288,N_1165);
or U1741 (N_1741,N_1163,N_221);
nand U1742 (N_1742,N_215,N_678);
nand U1743 (N_1743,N_1101,N_1300);
nand U1744 (N_1744,N_1389,N_1433);
and U1745 (N_1745,N_783,In_1309);
or U1746 (N_1746,N_1387,N_1495);
nand U1747 (N_1747,N_1316,N_1399);
xnor U1748 (N_1748,N_778,N_1481);
nor U1749 (N_1749,N_1342,N_1299);
nand U1750 (N_1750,N_1684,N_1694);
nand U1751 (N_1751,N_1644,N_1594);
or U1752 (N_1752,N_1743,N_1507);
or U1753 (N_1753,N_1725,N_1606);
xor U1754 (N_1754,N_1653,N_1565);
and U1755 (N_1755,N_1666,N_1629);
nor U1756 (N_1756,N_1664,N_1723);
nand U1757 (N_1757,N_1575,N_1554);
and U1758 (N_1758,N_1624,N_1505);
nand U1759 (N_1759,N_1718,N_1609);
xnor U1760 (N_1760,N_1673,N_1553);
xor U1761 (N_1761,N_1611,N_1667);
nor U1762 (N_1762,N_1628,N_1742);
nand U1763 (N_1763,N_1707,N_1548);
xnor U1764 (N_1764,N_1523,N_1520);
nor U1765 (N_1765,N_1541,N_1540);
or U1766 (N_1766,N_1598,N_1516);
or U1767 (N_1767,N_1517,N_1619);
xor U1768 (N_1768,N_1732,N_1552);
xor U1769 (N_1769,N_1646,N_1643);
nand U1770 (N_1770,N_1680,N_1519);
xor U1771 (N_1771,N_1682,N_1692);
nand U1772 (N_1772,N_1669,N_1648);
or U1773 (N_1773,N_1687,N_1538);
nand U1774 (N_1774,N_1581,N_1634);
and U1775 (N_1775,N_1522,N_1588);
and U1776 (N_1776,N_1524,N_1592);
and U1777 (N_1777,N_1702,N_1597);
nand U1778 (N_1778,N_1572,N_1593);
and U1779 (N_1779,N_1740,N_1733);
and U1780 (N_1780,N_1675,N_1662);
nand U1781 (N_1781,N_1734,N_1659);
nor U1782 (N_1782,N_1508,N_1615);
or U1783 (N_1783,N_1570,N_1567);
or U1784 (N_1784,N_1591,N_1603);
nor U1785 (N_1785,N_1748,N_1510);
xnor U1786 (N_1786,N_1627,N_1712);
or U1787 (N_1787,N_1713,N_1551);
or U1788 (N_1788,N_1642,N_1559);
and U1789 (N_1789,N_1504,N_1542);
nor U1790 (N_1790,N_1547,N_1549);
and U1791 (N_1791,N_1660,N_1728);
or U1792 (N_1792,N_1599,N_1543);
and U1793 (N_1793,N_1525,N_1530);
or U1794 (N_1794,N_1717,N_1651);
nor U1795 (N_1795,N_1539,N_1671);
and U1796 (N_1796,N_1584,N_1537);
or U1797 (N_1797,N_1561,N_1512);
nand U1798 (N_1798,N_1557,N_1566);
nor U1799 (N_1799,N_1722,N_1700);
and U1800 (N_1800,N_1737,N_1689);
or U1801 (N_1801,N_1558,N_1635);
and U1802 (N_1802,N_1589,N_1502);
nor U1803 (N_1803,N_1511,N_1564);
nand U1804 (N_1804,N_1645,N_1656);
or U1805 (N_1805,N_1587,N_1500);
and U1806 (N_1806,N_1726,N_1562);
and U1807 (N_1807,N_1583,N_1716);
or U1808 (N_1808,N_1714,N_1605);
nor U1809 (N_1809,N_1681,N_1623);
nand U1810 (N_1810,N_1631,N_1617);
and U1811 (N_1811,N_1657,N_1715);
nand U1812 (N_1812,N_1556,N_1585);
or U1813 (N_1813,N_1665,N_1576);
nor U1814 (N_1814,N_1730,N_1678);
nor U1815 (N_1815,N_1749,N_1699);
or U1816 (N_1816,N_1695,N_1744);
and U1817 (N_1817,N_1720,N_1649);
nor U1818 (N_1818,N_1688,N_1625);
nor U1819 (N_1819,N_1683,N_1618);
nand U1820 (N_1820,N_1602,N_1672);
nand U1821 (N_1821,N_1641,N_1626);
and U1822 (N_1822,N_1677,N_1632);
or U1823 (N_1823,N_1580,N_1703);
nor U1824 (N_1824,N_1735,N_1674);
nand U1825 (N_1825,N_1620,N_1721);
and U1826 (N_1826,N_1705,N_1710);
nand U1827 (N_1827,N_1698,N_1661);
or U1828 (N_1828,N_1696,N_1515);
and U1829 (N_1829,N_1630,N_1637);
or U1830 (N_1830,N_1697,N_1600);
and U1831 (N_1831,N_1555,N_1724);
xor U1832 (N_1832,N_1532,N_1747);
nand U1833 (N_1833,N_1650,N_1638);
or U1834 (N_1834,N_1739,N_1704);
and U1835 (N_1835,N_1526,N_1569);
nand U1836 (N_1836,N_1663,N_1521);
or U1837 (N_1837,N_1652,N_1708);
xor U1838 (N_1838,N_1745,N_1729);
nand U1839 (N_1839,N_1518,N_1514);
or U1840 (N_1840,N_1595,N_1527);
and U1841 (N_1841,N_1686,N_1690);
xnor U1842 (N_1842,N_1590,N_1693);
nand U1843 (N_1843,N_1550,N_1613);
xnor U1844 (N_1844,N_1563,N_1582);
and U1845 (N_1845,N_1528,N_1578);
xnor U1846 (N_1846,N_1531,N_1501);
nor U1847 (N_1847,N_1655,N_1612);
nand U1848 (N_1848,N_1621,N_1544);
nor U1849 (N_1849,N_1679,N_1736);
or U1850 (N_1850,N_1640,N_1610);
and U1851 (N_1851,N_1711,N_1506);
or U1852 (N_1852,N_1685,N_1647);
and U1853 (N_1853,N_1533,N_1654);
and U1854 (N_1854,N_1639,N_1738);
or U1855 (N_1855,N_1574,N_1614);
or U1856 (N_1856,N_1676,N_1535);
xnor U1857 (N_1857,N_1568,N_1571);
or U1858 (N_1858,N_1622,N_1706);
or U1859 (N_1859,N_1579,N_1636);
and U1860 (N_1860,N_1560,N_1607);
or U1861 (N_1861,N_1746,N_1616);
xnor U1862 (N_1862,N_1701,N_1691);
xnor U1863 (N_1863,N_1536,N_1601);
nor U1864 (N_1864,N_1503,N_1596);
and U1865 (N_1865,N_1545,N_1633);
nor U1866 (N_1866,N_1513,N_1731);
nand U1867 (N_1867,N_1709,N_1658);
nor U1868 (N_1868,N_1668,N_1529);
nand U1869 (N_1869,N_1577,N_1534);
and U1870 (N_1870,N_1608,N_1546);
or U1871 (N_1871,N_1509,N_1719);
nand U1872 (N_1872,N_1604,N_1586);
nand U1873 (N_1873,N_1573,N_1670);
nor U1874 (N_1874,N_1741,N_1727);
or U1875 (N_1875,N_1738,N_1522);
nand U1876 (N_1876,N_1579,N_1528);
or U1877 (N_1877,N_1506,N_1500);
nand U1878 (N_1878,N_1549,N_1507);
xor U1879 (N_1879,N_1663,N_1727);
and U1880 (N_1880,N_1632,N_1518);
nand U1881 (N_1881,N_1542,N_1735);
nand U1882 (N_1882,N_1630,N_1674);
nand U1883 (N_1883,N_1566,N_1709);
and U1884 (N_1884,N_1587,N_1693);
xnor U1885 (N_1885,N_1630,N_1603);
nor U1886 (N_1886,N_1697,N_1688);
nor U1887 (N_1887,N_1622,N_1651);
and U1888 (N_1888,N_1687,N_1659);
xnor U1889 (N_1889,N_1620,N_1624);
and U1890 (N_1890,N_1595,N_1583);
nand U1891 (N_1891,N_1642,N_1644);
xnor U1892 (N_1892,N_1653,N_1678);
or U1893 (N_1893,N_1625,N_1552);
xor U1894 (N_1894,N_1688,N_1519);
nand U1895 (N_1895,N_1748,N_1653);
nor U1896 (N_1896,N_1513,N_1678);
nand U1897 (N_1897,N_1585,N_1738);
nor U1898 (N_1898,N_1617,N_1542);
xnor U1899 (N_1899,N_1743,N_1613);
nor U1900 (N_1900,N_1558,N_1726);
nor U1901 (N_1901,N_1742,N_1679);
xor U1902 (N_1902,N_1506,N_1672);
xnor U1903 (N_1903,N_1585,N_1631);
or U1904 (N_1904,N_1584,N_1690);
nand U1905 (N_1905,N_1648,N_1737);
nor U1906 (N_1906,N_1714,N_1721);
xnor U1907 (N_1907,N_1698,N_1745);
nand U1908 (N_1908,N_1529,N_1698);
nand U1909 (N_1909,N_1666,N_1541);
nor U1910 (N_1910,N_1691,N_1606);
or U1911 (N_1911,N_1507,N_1653);
and U1912 (N_1912,N_1581,N_1549);
nor U1913 (N_1913,N_1726,N_1580);
nand U1914 (N_1914,N_1548,N_1567);
xor U1915 (N_1915,N_1515,N_1665);
and U1916 (N_1916,N_1710,N_1630);
xnor U1917 (N_1917,N_1573,N_1531);
or U1918 (N_1918,N_1580,N_1568);
xor U1919 (N_1919,N_1747,N_1739);
nand U1920 (N_1920,N_1572,N_1513);
nand U1921 (N_1921,N_1625,N_1730);
nor U1922 (N_1922,N_1671,N_1611);
and U1923 (N_1923,N_1668,N_1710);
nand U1924 (N_1924,N_1576,N_1718);
xnor U1925 (N_1925,N_1644,N_1619);
and U1926 (N_1926,N_1644,N_1626);
or U1927 (N_1927,N_1610,N_1699);
or U1928 (N_1928,N_1575,N_1680);
and U1929 (N_1929,N_1731,N_1688);
or U1930 (N_1930,N_1582,N_1681);
nand U1931 (N_1931,N_1720,N_1586);
nor U1932 (N_1932,N_1556,N_1567);
xor U1933 (N_1933,N_1714,N_1532);
or U1934 (N_1934,N_1568,N_1601);
nor U1935 (N_1935,N_1584,N_1634);
xnor U1936 (N_1936,N_1546,N_1704);
and U1937 (N_1937,N_1733,N_1716);
or U1938 (N_1938,N_1672,N_1675);
nand U1939 (N_1939,N_1652,N_1723);
xor U1940 (N_1940,N_1515,N_1707);
nor U1941 (N_1941,N_1685,N_1680);
and U1942 (N_1942,N_1611,N_1579);
nor U1943 (N_1943,N_1682,N_1553);
nand U1944 (N_1944,N_1656,N_1547);
nand U1945 (N_1945,N_1700,N_1565);
nand U1946 (N_1946,N_1662,N_1520);
nand U1947 (N_1947,N_1713,N_1524);
or U1948 (N_1948,N_1625,N_1550);
and U1949 (N_1949,N_1521,N_1559);
nor U1950 (N_1950,N_1543,N_1749);
or U1951 (N_1951,N_1722,N_1584);
or U1952 (N_1952,N_1668,N_1524);
and U1953 (N_1953,N_1642,N_1537);
or U1954 (N_1954,N_1573,N_1593);
and U1955 (N_1955,N_1654,N_1660);
nand U1956 (N_1956,N_1562,N_1598);
or U1957 (N_1957,N_1721,N_1532);
nor U1958 (N_1958,N_1713,N_1607);
and U1959 (N_1959,N_1578,N_1601);
nor U1960 (N_1960,N_1655,N_1650);
nor U1961 (N_1961,N_1693,N_1532);
and U1962 (N_1962,N_1725,N_1536);
nor U1963 (N_1963,N_1544,N_1505);
and U1964 (N_1964,N_1632,N_1601);
xor U1965 (N_1965,N_1591,N_1676);
xor U1966 (N_1966,N_1506,N_1544);
and U1967 (N_1967,N_1660,N_1579);
xor U1968 (N_1968,N_1588,N_1557);
xor U1969 (N_1969,N_1729,N_1518);
or U1970 (N_1970,N_1619,N_1518);
and U1971 (N_1971,N_1519,N_1682);
and U1972 (N_1972,N_1609,N_1522);
or U1973 (N_1973,N_1679,N_1618);
nand U1974 (N_1974,N_1681,N_1569);
xnor U1975 (N_1975,N_1682,N_1691);
or U1976 (N_1976,N_1737,N_1599);
nor U1977 (N_1977,N_1727,N_1724);
or U1978 (N_1978,N_1509,N_1539);
nor U1979 (N_1979,N_1694,N_1654);
nor U1980 (N_1980,N_1547,N_1552);
and U1981 (N_1981,N_1749,N_1583);
nand U1982 (N_1982,N_1706,N_1617);
nor U1983 (N_1983,N_1706,N_1503);
nand U1984 (N_1984,N_1521,N_1611);
nor U1985 (N_1985,N_1552,N_1630);
nor U1986 (N_1986,N_1572,N_1649);
xnor U1987 (N_1987,N_1561,N_1747);
or U1988 (N_1988,N_1552,N_1747);
nor U1989 (N_1989,N_1667,N_1562);
nand U1990 (N_1990,N_1567,N_1632);
or U1991 (N_1991,N_1541,N_1692);
nor U1992 (N_1992,N_1694,N_1517);
nand U1993 (N_1993,N_1565,N_1567);
and U1994 (N_1994,N_1617,N_1521);
nand U1995 (N_1995,N_1565,N_1687);
and U1996 (N_1996,N_1611,N_1699);
or U1997 (N_1997,N_1505,N_1696);
or U1998 (N_1998,N_1741,N_1630);
and U1999 (N_1999,N_1529,N_1691);
xor U2000 (N_2000,N_1851,N_1782);
and U2001 (N_2001,N_1925,N_1928);
nor U2002 (N_2002,N_1856,N_1770);
and U2003 (N_2003,N_1860,N_1984);
nand U2004 (N_2004,N_1803,N_1861);
or U2005 (N_2005,N_1800,N_1854);
and U2006 (N_2006,N_1793,N_1980);
nor U2007 (N_2007,N_1963,N_1957);
nor U2008 (N_2008,N_1761,N_1781);
and U2009 (N_2009,N_1874,N_1972);
nor U2010 (N_2010,N_1763,N_1758);
nor U2011 (N_2011,N_1838,N_1864);
nor U2012 (N_2012,N_1978,N_1853);
xor U2013 (N_2013,N_1900,N_1869);
xnor U2014 (N_2014,N_1934,N_1959);
xor U2015 (N_2015,N_1767,N_1756);
and U2016 (N_2016,N_1780,N_1943);
and U2017 (N_2017,N_1941,N_1919);
xnor U2018 (N_2018,N_1776,N_1893);
and U2019 (N_2019,N_1983,N_1786);
nor U2020 (N_2020,N_1995,N_1891);
or U2021 (N_2021,N_1842,N_1839);
or U2022 (N_2022,N_1956,N_1792);
nand U2023 (N_2023,N_1923,N_1931);
or U2024 (N_2024,N_1977,N_1989);
nor U2025 (N_2025,N_1762,N_1911);
nor U2026 (N_2026,N_1933,N_1929);
nand U2027 (N_2027,N_1914,N_1917);
and U2028 (N_2028,N_1942,N_1915);
nand U2029 (N_2029,N_1750,N_1766);
nor U2030 (N_2030,N_1817,N_1990);
xor U2031 (N_2031,N_1909,N_1831);
or U2032 (N_2032,N_1952,N_1787);
nand U2033 (N_2033,N_1849,N_1932);
or U2034 (N_2034,N_1798,N_1808);
nor U2035 (N_2035,N_1958,N_1960);
xor U2036 (N_2036,N_1898,N_1961);
and U2037 (N_2037,N_1829,N_1826);
nor U2038 (N_2038,N_1788,N_1754);
or U2039 (N_2039,N_1884,N_1807);
nand U2040 (N_2040,N_1821,N_1975);
nor U2041 (N_2041,N_1982,N_1913);
nand U2042 (N_2042,N_1843,N_1771);
xnor U2043 (N_2043,N_1901,N_1920);
nand U2044 (N_2044,N_1847,N_1889);
or U2045 (N_2045,N_1946,N_1938);
nor U2046 (N_2046,N_1918,N_1992);
and U2047 (N_2047,N_1773,N_1947);
or U2048 (N_2048,N_1962,N_1924);
xor U2049 (N_2049,N_1797,N_1882);
nand U2050 (N_2050,N_1791,N_1812);
xor U2051 (N_2051,N_1954,N_1769);
nor U2052 (N_2052,N_1795,N_1885);
nand U2053 (N_2053,N_1796,N_1944);
xnor U2054 (N_2054,N_1772,N_1815);
xor U2055 (N_2055,N_1810,N_1970);
or U2056 (N_2056,N_1804,N_1921);
or U2057 (N_2057,N_1840,N_1835);
xor U2058 (N_2058,N_1953,N_1996);
or U2059 (N_2059,N_1937,N_1836);
and U2060 (N_2060,N_1862,N_1899);
or U2061 (N_2061,N_1852,N_1896);
or U2062 (N_2062,N_1828,N_1955);
nand U2063 (N_2063,N_1866,N_1872);
nand U2064 (N_2064,N_1827,N_1875);
xor U2065 (N_2065,N_1892,N_1988);
nand U2066 (N_2066,N_1824,N_1912);
or U2067 (N_2067,N_1846,N_1908);
and U2068 (N_2068,N_1877,N_1755);
and U2069 (N_2069,N_1816,N_1813);
nand U2070 (N_2070,N_1876,N_1858);
and U2071 (N_2071,N_1751,N_1855);
xnor U2072 (N_2072,N_1823,N_1834);
and U2073 (N_2073,N_1859,N_1880);
nor U2074 (N_2074,N_1865,N_1979);
nor U2075 (N_2075,N_1799,N_1878);
nand U2076 (N_2076,N_1895,N_1777);
nand U2077 (N_2077,N_1886,N_1819);
or U2078 (N_2078,N_1775,N_1789);
or U2079 (N_2079,N_1969,N_1805);
nor U2080 (N_2080,N_1890,N_1973);
or U2081 (N_2081,N_1910,N_1950);
nor U2082 (N_2082,N_1820,N_1993);
nor U2083 (N_2083,N_1974,N_1935);
nor U2084 (N_2084,N_1906,N_1811);
nor U2085 (N_2085,N_1922,N_1879);
nand U2086 (N_2086,N_1873,N_1774);
and U2087 (N_2087,N_1987,N_1916);
and U2088 (N_2088,N_1863,N_1848);
nand U2089 (N_2089,N_1867,N_1940);
or U2090 (N_2090,N_1936,N_1902);
and U2091 (N_2091,N_1965,N_1991);
nand U2092 (N_2092,N_1759,N_1841);
nand U2093 (N_2093,N_1794,N_1997);
nor U2094 (N_2094,N_1926,N_1814);
and U2095 (N_2095,N_1753,N_1844);
nand U2096 (N_2096,N_1968,N_1966);
nand U2097 (N_2097,N_1985,N_1883);
or U2098 (N_2098,N_1783,N_1888);
xnor U2099 (N_2099,N_1850,N_1949);
nor U2100 (N_2100,N_1778,N_1830);
and U2101 (N_2101,N_1967,N_1971);
nand U2102 (N_2102,N_1785,N_1976);
xnor U2103 (N_2103,N_1832,N_1857);
and U2104 (N_2104,N_1802,N_1768);
nand U2105 (N_2105,N_1871,N_1927);
nand U2106 (N_2106,N_1806,N_1994);
and U2107 (N_2107,N_1903,N_1845);
nor U2108 (N_2108,N_1764,N_1951);
or U2109 (N_2109,N_1981,N_1809);
nand U2110 (N_2110,N_1801,N_1870);
and U2111 (N_2111,N_1905,N_1887);
and U2112 (N_2112,N_1948,N_1986);
xor U2113 (N_2113,N_1939,N_1999);
nand U2114 (N_2114,N_1760,N_1945);
and U2115 (N_2115,N_1894,N_1779);
and U2116 (N_2116,N_1833,N_1904);
xnor U2117 (N_2117,N_1784,N_1964);
nor U2118 (N_2118,N_1825,N_1998);
nor U2119 (N_2119,N_1752,N_1881);
nor U2120 (N_2120,N_1822,N_1837);
and U2121 (N_2121,N_1930,N_1868);
and U2122 (N_2122,N_1897,N_1790);
xor U2123 (N_2123,N_1765,N_1907);
nand U2124 (N_2124,N_1757,N_1818);
xnor U2125 (N_2125,N_1774,N_1800);
nand U2126 (N_2126,N_1954,N_1808);
xnor U2127 (N_2127,N_1972,N_1764);
xnor U2128 (N_2128,N_1802,N_1913);
xnor U2129 (N_2129,N_1844,N_1817);
or U2130 (N_2130,N_1821,N_1969);
nand U2131 (N_2131,N_1965,N_1913);
and U2132 (N_2132,N_1998,N_1890);
or U2133 (N_2133,N_1754,N_1849);
and U2134 (N_2134,N_1774,N_1950);
nor U2135 (N_2135,N_1987,N_1897);
xor U2136 (N_2136,N_1892,N_1767);
and U2137 (N_2137,N_1841,N_1973);
nand U2138 (N_2138,N_1874,N_1993);
nor U2139 (N_2139,N_1928,N_1791);
and U2140 (N_2140,N_1910,N_1836);
xnor U2141 (N_2141,N_1788,N_1973);
xor U2142 (N_2142,N_1968,N_1987);
nand U2143 (N_2143,N_1813,N_1846);
nand U2144 (N_2144,N_1761,N_1776);
and U2145 (N_2145,N_1842,N_1893);
and U2146 (N_2146,N_1849,N_1855);
xor U2147 (N_2147,N_1913,N_1940);
nor U2148 (N_2148,N_1851,N_1966);
nand U2149 (N_2149,N_1987,N_1954);
and U2150 (N_2150,N_1849,N_1850);
nor U2151 (N_2151,N_1848,N_1942);
and U2152 (N_2152,N_1896,N_1929);
or U2153 (N_2153,N_1796,N_1883);
xnor U2154 (N_2154,N_1966,N_1769);
and U2155 (N_2155,N_1984,N_1850);
and U2156 (N_2156,N_1819,N_1798);
nand U2157 (N_2157,N_1825,N_1982);
and U2158 (N_2158,N_1824,N_1884);
or U2159 (N_2159,N_1783,N_1918);
nor U2160 (N_2160,N_1904,N_1872);
or U2161 (N_2161,N_1957,N_1842);
nand U2162 (N_2162,N_1903,N_1949);
and U2163 (N_2163,N_1978,N_1847);
xor U2164 (N_2164,N_1840,N_1988);
and U2165 (N_2165,N_1779,N_1878);
nand U2166 (N_2166,N_1934,N_1884);
nand U2167 (N_2167,N_1751,N_1934);
or U2168 (N_2168,N_1942,N_1988);
nor U2169 (N_2169,N_1997,N_1958);
or U2170 (N_2170,N_1832,N_1994);
xnor U2171 (N_2171,N_1751,N_1995);
nand U2172 (N_2172,N_1753,N_1781);
and U2173 (N_2173,N_1858,N_1828);
or U2174 (N_2174,N_1806,N_1927);
xor U2175 (N_2175,N_1921,N_1820);
and U2176 (N_2176,N_1796,N_1956);
nand U2177 (N_2177,N_1897,N_1840);
nand U2178 (N_2178,N_1950,N_1941);
nand U2179 (N_2179,N_1858,N_1973);
nand U2180 (N_2180,N_1944,N_1886);
xnor U2181 (N_2181,N_1773,N_1833);
nor U2182 (N_2182,N_1780,N_1800);
nand U2183 (N_2183,N_1949,N_1912);
xnor U2184 (N_2184,N_1810,N_1820);
or U2185 (N_2185,N_1908,N_1817);
nor U2186 (N_2186,N_1946,N_1797);
and U2187 (N_2187,N_1803,N_1923);
nor U2188 (N_2188,N_1765,N_1800);
or U2189 (N_2189,N_1905,N_1933);
and U2190 (N_2190,N_1941,N_1925);
or U2191 (N_2191,N_1972,N_1800);
and U2192 (N_2192,N_1772,N_1826);
nor U2193 (N_2193,N_1818,N_1872);
xor U2194 (N_2194,N_1778,N_1999);
nand U2195 (N_2195,N_1831,N_1976);
nand U2196 (N_2196,N_1914,N_1906);
nand U2197 (N_2197,N_1917,N_1898);
nor U2198 (N_2198,N_1810,N_1923);
nor U2199 (N_2199,N_1801,N_1973);
nand U2200 (N_2200,N_1817,N_1862);
xor U2201 (N_2201,N_1866,N_1838);
and U2202 (N_2202,N_1956,N_1762);
and U2203 (N_2203,N_1993,N_1962);
or U2204 (N_2204,N_1917,N_1821);
and U2205 (N_2205,N_1981,N_1982);
nor U2206 (N_2206,N_1827,N_1750);
xor U2207 (N_2207,N_1893,N_1947);
nor U2208 (N_2208,N_1786,N_1818);
and U2209 (N_2209,N_1840,N_1909);
and U2210 (N_2210,N_1830,N_1849);
nor U2211 (N_2211,N_1874,N_1766);
nor U2212 (N_2212,N_1994,N_1909);
nand U2213 (N_2213,N_1911,N_1796);
nand U2214 (N_2214,N_1790,N_1880);
nor U2215 (N_2215,N_1968,N_1909);
nor U2216 (N_2216,N_1962,N_1777);
xor U2217 (N_2217,N_1979,N_1934);
nand U2218 (N_2218,N_1974,N_1861);
nor U2219 (N_2219,N_1840,N_1963);
xor U2220 (N_2220,N_1921,N_1983);
and U2221 (N_2221,N_1964,N_1831);
nor U2222 (N_2222,N_1914,N_1910);
nor U2223 (N_2223,N_1764,N_1860);
nor U2224 (N_2224,N_1798,N_1824);
nor U2225 (N_2225,N_1957,N_1894);
nand U2226 (N_2226,N_1836,N_1933);
nand U2227 (N_2227,N_1885,N_1845);
nor U2228 (N_2228,N_1812,N_1940);
and U2229 (N_2229,N_1969,N_1923);
or U2230 (N_2230,N_1960,N_1956);
and U2231 (N_2231,N_1756,N_1861);
and U2232 (N_2232,N_1968,N_1854);
xnor U2233 (N_2233,N_1805,N_1940);
and U2234 (N_2234,N_1862,N_1751);
xor U2235 (N_2235,N_1867,N_1887);
or U2236 (N_2236,N_1833,N_1966);
or U2237 (N_2237,N_1784,N_1992);
and U2238 (N_2238,N_1923,N_1939);
xor U2239 (N_2239,N_1869,N_1758);
xnor U2240 (N_2240,N_1954,N_1960);
or U2241 (N_2241,N_1934,N_1994);
or U2242 (N_2242,N_1973,N_1945);
or U2243 (N_2243,N_1860,N_1811);
nor U2244 (N_2244,N_1830,N_1844);
nand U2245 (N_2245,N_1901,N_1986);
xor U2246 (N_2246,N_1832,N_1974);
nand U2247 (N_2247,N_1750,N_1991);
nor U2248 (N_2248,N_1958,N_1769);
nor U2249 (N_2249,N_1757,N_1882);
and U2250 (N_2250,N_2097,N_2153);
nand U2251 (N_2251,N_2088,N_2247);
or U2252 (N_2252,N_2172,N_2244);
and U2253 (N_2253,N_2152,N_2140);
or U2254 (N_2254,N_2132,N_2234);
xor U2255 (N_2255,N_2191,N_2025);
nor U2256 (N_2256,N_2120,N_2056);
xnor U2257 (N_2257,N_2134,N_2066);
nor U2258 (N_2258,N_2116,N_2080);
or U2259 (N_2259,N_2170,N_2161);
nand U2260 (N_2260,N_2019,N_2195);
or U2261 (N_2261,N_2249,N_2053);
nor U2262 (N_2262,N_2210,N_2227);
xor U2263 (N_2263,N_2198,N_2118);
or U2264 (N_2264,N_2067,N_2110);
nand U2265 (N_2265,N_2197,N_2069);
and U2266 (N_2266,N_2165,N_2000);
or U2267 (N_2267,N_2219,N_2222);
and U2268 (N_2268,N_2087,N_2157);
nand U2269 (N_2269,N_2204,N_2005);
or U2270 (N_2270,N_2237,N_2171);
nand U2271 (N_2271,N_2178,N_2107);
xnor U2272 (N_2272,N_2201,N_2190);
or U2273 (N_2273,N_2183,N_2109);
or U2274 (N_2274,N_2021,N_2163);
and U2275 (N_2275,N_2052,N_2187);
and U2276 (N_2276,N_2168,N_2126);
xor U2277 (N_2277,N_2054,N_2013);
nand U2278 (N_2278,N_2081,N_2100);
or U2279 (N_2279,N_2167,N_2214);
or U2280 (N_2280,N_2131,N_2226);
nand U2281 (N_2281,N_2112,N_2068);
xnor U2282 (N_2282,N_2001,N_2185);
xor U2283 (N_2283,N_2155,N_2159);
or U2284 (N_2284,N_2039,N_2216);
nor U2285 (N_2285,N_2209,N_2221);
xnor U2286 (N_2286,N_2149,N_2138);
nand U2287 (N_2287,N_2236,N_2049);
xnor U2288 (N_2288,N_2030,N_2015);
xnor U2289 (N_2289,N_2042,N_2012);
or U2290 (N_2290,N_2213,N_2230);
or U2291 (N_2291,N_2215,N_2032);
or U2292 (N_2292,N_2202,N_2023);
nor U2293 (N_2293,N_2123,N_2114);
or U2294 (N_2294,N_2060,N_2045);
nand U2295 (N_2295,N_2093,N_2246);
or U2296 (N_2296,N_2016,N_2229);
or U2297 (N_2297,N_2156,N_2113);
nor U2298 (N_2298,N_2184,N_2206);
or U2299 (N_2299,N_2051,N_2104);
nand U2300 (N_2300,N_2004,N_2175);
and U2301 (N_2301,N_2011,N_2091);
and U2302 (N_2302,N_2099,N_2078);
and U2303 (N_2303,N_2029,N_2141);
nand U2304 (N_2304,N_2079,N_2173);
nand U2305 (N_2305,N_2063,N_2151);
and U2306 (N_2306,N_2127,N_2007);
xor U2307 (N_2307,N_2228,N_2074);
or U2308 (N_2308,N_2139,N_2203);
xor U2309 (N_2309,N_2121,N_2010);
nand U2310 (N_2310,N_2235,N_2128);
nor U2311 (N_2311,N_2096,N_2147);
or U2312 (N_2312,N_2090,N_2111);
nor U2313 (N_2313,N_2137,N_2022);
xnor U2314 (N_2314,N_2008,N_2208);
or U2315 (N_2315,N_2084,N_2014);
and U2316 (N_2316,N_2129,N_2142);
and U2317 (N_2317,N_2031,N_2046);
nand U2318 (N_2318,N_2166,N_2240);
nor U2319 (N_2319,N_2224,N_2106);
nand U2320 (N_2320,N_2154,N_2164);
or U2321 (N_2321,N_2232,N_2061);
xor U2322 (N_2322,N_2076,N_2055);
xor U2323 (N_2323,N_2059,N_2122);
or U2324 (N_2324,N_2125,N_2233);
nand U2325 (N_2325,N_2223,N_2217);
and U2326 (N_2326,N_2133,N_2071);
nor U2327 (N_2327,N_2057,N_2200);
xnor U2328 (N_2328,N_2115,N_2144);
and U2329 (N_2329,N_2026,N_2082);
and U2330 (N_2330,N_2072,N_2146);
or U2331 (N_2331,N_2103,N_2189);
nand U2332 (N_2332,N_2192,N_2186);
nand U2333 (N_2333,N_2033,N_2003);
xnor U2334 (N_2334,N_2058,N_2047);
or U2335 (N_2335,N_2083,N_2024);
or U2336 (N_2336,N_2070,N_2242);
nand U2337 (N_2337,N_2064,N_2037);
xor U2338 (N_2338,N_2245,N_2017);
or U2339 (N_2339,N_2196,N_2188);
nor U2340 (N_2340,N_2199,N_2098);
nand U2341 (N_2341,N_2136,N_2181);
nand U2342 (N_2342,N_2092,N_2009);
nor U2343 (N_2343,N_2048,N_2027);
or U2344 (N_2344,N_2040,N_2105);
and U2345 (N_2345,N_2150,N_2124);
or U2346 (N_2346,N_2119,N_2205);
nand U2347 (N_2347,N_2176,N_2050);
xor U2348 (N_2348,N_2135,N_2160);
xor U2349 (N_2349,N_2212,N_2041);
nand U2350 (N_2350,N_2034,N_2225);
or U2351 (N_2351,N_2038,N_2179);
and U2352 (N_2352,N_2094,N_2145);
xnor U2353 (N_2353,N_2073,N_2035);
and U2354 (N_2354,N_2194,N_2043);
xor U2355 (N_2355,N_2044,N_2095);
xnor U2356 (N_2356,N_2180,N_2102);
or U2357 (N_2357,N_2089,N_2158);
or U2358 (N_2358,N_2248,N_2075);
and U2359 (N_2359,N_2174,N_2108);
and U2360 (N_2360,N_2086,N_2238);
and U2361 (N_2361,N_2239,N_2220);
and U2362 (N_2362,N_2177,N_2117);
nand U2363 (N_2363,N_2028,N_2218);
nor U2364 (N_2364,N_2169,N_2148);
nand U2365 (N_2365,N_2207,N_2006);
nand U2366 (N_2366,N_2036,N_2101);
and U2367 (N_2367,N_2020,N_2211);
and U2368 (N_2368,N_2065,N_2231);
xnor U2369 (N_2369,N_2085,N_2018);
nand U2370 (N_2370,N_2162,N_2130);
and U2371 (N_2371,N_2243,N_2062);
xor U2372 (N_2372,N_2182,N_2241);
xnor U2373 (N_2373,N_2077,N_2143);
nand U2374 (N_2374,N_2002,N_2193);
nor U2375 (N_2375,N_2102,N_2021);
nor U2376 (N_2376,N_2108,N_2169);
and U2377 (N_2377,N_2247,N_2187);
nor U2378 (N_2378,N_2007,N_2017);
and U2379 (N_2379,N_2235,N_2218);
nor U2380 (N_2380,N_2017,N_2228);
nand U2381 (N_2381,N_2110,N_2198);
xnor U2382 (N_2382,N_2141,N_2160);
nand U2383 (N_2383,N_2175,N_2073);
nor U2384 (N_2384,N_2020,N_2180);
nor U2385 (N_2385,N_2205,N_2192);
and U2386 (N_2386,N_2130,N_2241);
or U2387 (N_2387,N_2032,N_2210);
nor U2388 (N_2388,N_2004,N_2183);
nand U2389 (N_2389,N_2043,N_2148);
nand U2390 (N_2390,N_2103,N_2025);
xnor U2391 (N_2391,N_2024,N_2058);
xor U2392 (N_2392,N_2207,N_2040);
nand U2393 (N_2393,N_2238,N_2119);
nor U2394 (N_2394,N_2187,N_2156);
and U2395 (N_2395,N_2129,N_2070);
or U2396 (N_2396,N_2183,N_2014);
nor U2397 (N_2397,N_2029,N_2055);
nand U2398 (N_2398,N_2110,N_2037);
xnor U2399 (N_2399,N_2118,N_2202);
or U2400 (N_2400,N_2185,N_2216);
xnor U2401 (N_2401,N_2206,N_2242);
or U2402 (N_2402,N_2040,N_2117);
nor U2403 (N_2403,N_2030,N_2041);
or U2404 (N_2404,N_2179,N_2213);
xnor U2405 (N_2405,N_2212,N_2172);
and U2406 (N_2406,N_2236,N_2149);
xor U2407 (N_2407,N_2018,N_2149);
nor U2408 (N_2408,N_2155,N_2193);
xnor U2409 (N_2409,N_2054,N_2164);
and U2410 (N_2410,N_2094,N_2193);
nor U2411 (N_2411,N_2041,N_2042);
or U2412 (N_2412,N_2166,N_2162);
nand U2413 (N_2413,N_2225,N_2130);
nor U2414 (N_2414,N_2200,N_2180);
nand U2415 (N_2415,N_2153,N_2140);
xor U2416 (N_2416,N_2210,N_2246);
nor U2417 (N_2417,N_2125,N_2195);
nand U2418 (N_2418,N_2104,N_2189);
and U2419 (N_2419,N_2099,N_2037);
nor U2420 (N_2420,N_2171,N_2020);
xnor U2421 (N_2421,N_2048,N_2066);
and U2422 (N_2422,N_2074,N_2154);
nand U2423 (N_2423,N_2039,N_2004);
nand U2424 (N_2424,N_2234,N_2114);
or U2425 (N_2425,N_2157,N_2166);
nand U2426 (N_2426,N_2020,N_2121);
or U2427 (N_2427,N_2109,N_2019);
nor U2428 (N_2428,N_2030,N_2014);
or U2429 (N_2429,N_2041,N_2141);
or U2430 (N_2430,N_2036,N_2243);
and U2431 (N_2431,N_2134,N_2059);
xor U2432 (N_2432,N_2104,N_2128);
and U2433 (N_2433,N_2071,N_2185);
and U2434 (N_2434,N_2102,N_2062);
or U2435 (N_2435,N_2228,N_2166);
or U2436 (N_2436,N_2003,N_2032);
or U2437 (N_2437,N_2180,N_2244);
nor U2438 (N_2438,N_2128,N_2233);
xnor U2439 (N_2439,N_2069,N_2034);
and U2440 (N_2440,N_2219,N_2101);
and U2441 (N_2441,N_2078,N_2094);
xor U2442 (N_2442,N_2127,N_2042);
nand U2443 (N_2443,N_2243,N_2159);
nor U2444 (N_2444,N_2118,N_2062);
xor U2445 (N_2445,N_2111,N_2036);
nand U2446 (N_2446,N_2227,N_2145);
xnor U2447 (N_2447,N_2065,N_2092);
nand U2448 (N_2448,N_2166,N_2124);
and U2449 (N_2449,N_2006,N_2096);
nor U2450 (N_2450,N_2131,N_2213);
and U2451 (N_2451,N_2078,N_2206);
xor U2452 (N_2452,N_2145,N_2071);
and U2453 (N_2453,N_2126,N_2232);
nor U2454 (N_2454,N_2187,N_2121);
nand U2455 (N_2455,N_2059,N_2217);
or U2456 (N_2456,N_2125,N_2086);
nand U2457 (N_2457,N_2019,N_2217);
nor U2458 (N_2458,N_2048,N_2042);
or U2459 (N_2459,N_2121,N_2101);
nor U2460 (N_2460,N_2216,N_2178);
nand U2461 (N_2461,N_2245,N_2239);
or U2462 (N_2462,N_2131,N_2168);
and U2463 (N_2463,N_2241,N_2137);
nor U2464 (N_2464,N_2120,N_2134);
or U2465 (N_2465,N_2027,N_2086);
or U2466 (N_2466,N_2210,N_2075);
xor U2467 (N_2467,N_2048,N_2008);
nor U2468 (N_2468,N_2022,N_2016);
nor U2469 (N_2469,N_2024,N_2120);
xor U2470 (N_2470,N_2014,N_2160);
xnor U2471 (N_2471,N_2017,N_2186);
and U2472 (N_2472,N_2198,N_2079);
or U2473 (N_2473,N_2018,N_2141);
and U2474 (N_2474,N_2087,N_2238);
or U2475 (N_2475,N_2051,N_2096);
nor U2476 (N_2476,N_2239,N_2106);
nor U2477 (N_2477,N_2242,N_2033);
and U2478 (N_2478,N_2225,N_2074);
or U2479 (N_2479,N_2044,N_2012);
and U2480 (N_2480,N_2144,N_2019);
xor U2481 (N_2481,N_2060,N_2004);
xor U2482 (N_2482,N_2195,N_2098);
or U2483 (N_2483,N_2058,N_2108);
nand U2484 (N_2484,N_2216,N_2187);
and U2485 (N_2485,N_2246,N_2078);
and U2486 (N_2486,N_2244,N_2230);
or U2487 (N_2487,N_2025,N_2036);
and U2488 (N_2488,N_2147,N_2205);
or U2489 (N_2489,N_2173,N_2093);
nor U2490 (N_2490,N_2027,N_2058);
xnor U2491 (N_2491,N_2111,N_2212);
nand U2492 (N_2492,N_2043,N_2211);
and U2493 (N_2493,N_2102,N_2217);
nor U2494 (N_2494,N_2228,N_2036);
or U2495 (N_2495,N_2119,N_2052);
nand U2496 (N_2496,N_2200,N_2066);
xnor U2497 (N_2497,N_2184,N_2106);
or U2498 (N_2498,N_2039,N_2201);
nand U2499 (N_2499,N_2122,N_2180);
and U2500 (N_2500,N_2378,N_2373);
or U2501 (N_2501,N_2448,N_2474);
nand U2502 (N_2502,N_2421,N_2430);
or U2503 (N_2503,N_2301,N_2258);
and U2504 (N_2504,N_2289,N_2307);
and U2505 (N_2505,N_2436,N_2253);
nor U2506 (N_2506,N_2438,N_2445);
or U2507 (N_2507,N_2452,N_2406);
nand U2508 (N_2508,N_2374,N_2275);
and U2509 (N_2509,N_2370,N_2252);
or U2510 (N_2510,N_2493,N_2280);
nand U2511 (N_2511,N_2371,N_2322);
nor U2512 (N_2512,N_2376,N_2291);
nor U2513 (N_2513,N_2480,N_2335);
or U2514 (N_2514,N_2302,N_2329);
nand U2515 (N_2515,N_2467,N_2295);
xor U2516 (N_2516,N_2409,N_2267);
and U2517 (N_2517,N_2380,N_2265);
and U2518 (N_2518,N_2484,N_2417);
nor U2519 (N_2519,N_2387,N_2412);
nand U2520 (N_2520,N_2328,N_2435);
nor U2521 (N_2521,N_2457,N_2444);
nand U2522 (N_2522,N_2405,N_2486);
and U2523 (N_2523,N_2282,N_2394);
or U2524 (N_2524,N_2303,N_2375);
xor U2525 (N_2525,N_2433,N_2365);
and U2526 (N_2526,N_2477,N_2447);
xor U2527 (N_2527,N_2422,N_2407);
or U2528 (N_2528,N_2494,N_2296);
or U2529 (N_2529,N_2345,N_2449);
xor U2530 (N_2530,N_2250,N_2453);
or U2531 (N_2531,N_2498,N_2260);
nor U2532 (N_2532,N_2451,N_2465);
and U2533 (N_2533,N_2355,N_2325);
nand U2534 (N_2534,N_2393,N_2276);
nor U2535 (N_2535,N_2473,N_2483);
xnor U2536 (N_2536,N_2326,N_2496);
and U2537 (N_2537,N_2344,N_2368);
or U2538 (N_2538,N_2333,N_2261);
nor U2539 (N_2539,N_2270,N_2372);
and U2540 (N_2540,N_2278,N_2454);
nand U2541 (N_2541,N_2497,N_2460);
and U2542 (N_2542,N_2426,N_2470);
and U2543 (N_2543,N_2492,N_2471);
nand U2544 (N_2544,N_2311,N_2415);
nor U2545 (N_2545,N_2424,N_2411);
xnor U2546 (N_2546,N_2300,N_2434);
xor U2547 (N_2547,N_2459,N_2277);
xor U2548 (N_2548,N_2298,N_2410);
xor U2549 (N_2549,N_2455,N_2396);
or U2550 (N_2550,N_2356,N_2456);
nor U2551 (N_2551,N_2429,N_2257);
nand U2552 (N_2552,N_2281,N_2461);
xnor U2553 (N_2553,N_2305,N_2262);
nand U2554 (N_2554,N_2330,N_2408);
or U2555 (N_2555,N_2418,N_2366);
xnor U2556 (N_2556,N_2468,N_2428);
or U2557 (N_2557,N_2463,N_2342);
nor U2558 (N_2558,N_2363,N_2313);
xnor U2559 (N_2559,N_2398,N_2495);
or U2560 (N_2560,N_2316,N_2327);
or U2561 (N_2561,N_2287,N_2332);
nor U2562 (N_2562,N_2478,N_2391);
nand U2563 (N_2563,N_2353,N_2420);
or U2564 (N_2564,N_2476,N_2264);
or U2565 (N_2565,N_2279,N_2401);
nand U2566 (N_2566,N_2399,N_2472);
xnor U2567 (N_2567,N_2377,N_2272);
or U2568 (N_2568,N_2425,N_2299);
and U2569 (N_2569,N_2427,N_2343);
or U2570 (N_2570,N_2285,N_2334);
xor U2571 (N_2571,N_2336,N_2259);
nand U2572 (N_2572,N_2382,N_2308);
or U2573 (N_2573,N_2349,N_2331);
and U2574 (N_2574,N_2318,N_2297);
and U2575 (N_2575,N_2266,N_2364);
nand U2576 (N_2576,N_2251,N_2439);
nand U2577 (N_2577,N_2323,N_2284);
or U2578 (N_2578,N_2306,N_2283);
nand U2579 (N_2579,N_2271,N_2414);
or U2580 (N_2580,N_2317,N_2350);
xnor U2581 (N_2581,N_2319,N_2274);
xnor U2582 (N_2582,N_2419,N_2400);
or U2583 (N_2583,N_2360,N_2475);
and U2584 (N_2584,N_2385,N_2383);
and U2585 (N_2585,N_2464,N_2392);
xor U2586 (N_2586,N_2443,N_2390);
nor U2587 (N_2587,N_2432,N_2381);
nor U2588 (N_2588,N_2403,N_2304);
nor U2589 (N_2589,N_2446,N_2481);
and U2590 (N_2590,N_2389,N_2369);
nor U2591 (N_2591,N_2379,N_2294);
or U2592 (N_2592,N_2273,N_2359);
and U2593 (N_2593,N_2362,N_2466);
nand U2594 (N_2594,N_2339,N_2367);
nand U2595 (N_2595,N_2440,N_2491);
xnor U2596 (N_2596,N_2315,N_2416);
or U2597 (N_2597,N_2487,N_2288);
nor U2598 (N_2598,N_2450,N_2337);
nor U2599 (N_2599,N_2395,N_2346);
nor U2600 (N_2600,N_2479,N_2351);
nand U2601 (N_2601,N_2357,N_2286);
xor U2602 (N_2602,N_2352,N_2269);
and U2603 (N_2603,N_2321,N_2485);
or U2604 (N_2604,N_2388,N_2482);
and U2605 (N_2605,N_2340,N_2489);
nand U2606 (N_2606,N_2293,N_2254);
nor U2607 (N_2607,N_2458,N_2290);
xnor U2608 (N_2608,N_2469,N_2386);
nor U2609 (N_2609,N_2324,N_2413);
or U2610 (N_2610,N_2488,N_2314);
xnor U2611 (N_2611,N_2442,N_2404);
xnor U2612 (N_2612,N_2423,N_2341);
or U2613 (N_2613,N_2499,N_2268);
nor U2614 (N_2614,N_2256,N_2431);
and U2615 (N_2615,N_2338,N_2320);
or U2616 (N_2616,N_2354,N_2255);
and U2617 (N_2617,N_2292,N_2361);
and U2618 (N_2618,N_2263,N_2490);
and U2619 (N_2619,N_2312,N_2309);
and U2620 (N_2620,N_2441,N_2310);
and U2621 (N_2621,N_2384,N_2402);
nor U2622 (N_2622,N_2437,N_2347);
and U2623 (N_2623,N_2358,N_2348);
or U2624 (N_2624,N_2462,N_2397);
nor U2625 (N_2625,N_2351,N_2295);
nand U2626 (N_2626,N_2294,N_2290);
or U2627 (N_2627,N_2496,N_2451);
xnor U2628 (N_2628,N_2290,N_2417);
nand U2629 (N_2629,N_2397,N_2295);
or U2630 (N_2630,N_2336,N_2480);
nor U2631 (N_2631,N_2409,N_2469);
or U2632 (N_2632,N_2459,N_2252);
nand U2633 (N_2633,N_2451,N_2375);
and U2634 (N_2634,N_2393,N_2294);
xnor U2635 (N_2635,N_2441,N_2274);
or U2636 (N_2636,N_2423,N_2409);
nor U2637 (N_2637,N_2286,N_2310);
xor U2638 (N_2638,N_2255,N_2325);
or U2639 (N_2639,N_2260,N_2444);
nand U2640 (N_2640,N_2337,N_2408);
nand U2641 (N_2641,N_2366,N_2402);
nand U2642 (N_2642,N_2474,N_2327);
or U2643 (N_2643,N_2411,N_2474);
xnor U2644 (N_2644,N_2449,N_2291);
and U2645 (N_2645,N_2272,N_2380);
nand U2646 (N_2646,N_2487,N_2412);
nand U2647 (N_2647,N_2256,N_2384);
nor U2648 (N_2648,N_2352,N_2399);
xnor U2649 (N_2649,N_2324,N_2361);
nor U2650 (N_2650,N_2440,N_2457);
nand U2651 (N_2651,N_2341,N_2470);
nor U2652 (N_2652,N_2375,N_2472);
nor U2653 (N_2653,N_2405,N_2497);
or U2654 (N_2654,N_2419,N_2469);
xnor U2655 (N_2655,N_2287,N_2394);
or U2656 (N_2656,N_2397,N_2289);
and U2657 (N_2657,N_2346,N_2401);
or U2658 (N_2658,N_2339,N_2259);
and U2659 (N_2659,N_2439,N_2267);
or U2660 (N_2660,N_2495,N_2353);
nand U2661 (N_2661,N_2321,N_2333);
or U2662 (N_2662,N_2499,N_2338);
nand U2663 (N_2663,N_2449,N_2483);
nor U2664 (N_2664,N_2287,N_2457);
or U2665 (N_2665,N_2386,N_2308);
xnor U2666 (N_2666,N_2346,N_2469);
nand U2667 (N_2667,N_2270,N_2262);
nand U2668 (N_2668,N_2260,N_2378);
xor U2669 (N_2669,N_2380,N_2457);
and U2670 (N_2670,N_2319,N_2485);
xnor U2671 (N_2671,N_2292,N_2420);
nor U2672 (N_2672,N_2319,N_2374);
xnor U2673 (N_2673,N_2427,N_2335);
and U2674 (N_2674,N_2348,N_2412);
nand U2675 (N_2675,N_2418,N_2454);
nand U2676 (N_2676,N_2371,N_2478);
or U2677 (N_2677,N_2358,N_2441);
and U2678 (N_2678,N_2382,N_2451);
or U2679 (N_2679,N_2370,N_2478);
xor U2680 (N_2680,N_2334,N_2373);
nor U2681 (N_2681,N_2432,N_2431);
or U2682 (N_2682,N_2308,N_2446);
nand U2683 (N_2683,N_2419,N_2451);
and U2684 (N_2684,N_2284,N_2392);
xor U2685 (N_2685,N_2379,N_2451);
nor U2686 (N_2686,N_2346,N_2440);
nor U2687 (N_2687,N_2313,N_2480);
xnor U2688 (N_2688,N_2436,N_2356);
and U2689 (N_2689,N_2447,N_2289);
or U2690 (N_2690,N_2364,N_2251);
or U2691 (N_2691,N_2483,N_2268);
nand U2692 (N_2692,N_2301,N_2331);
and U2693 (N_2693,N_2280,N_2314);
and U2694 (N_2694,N_2418,N_2388);
nor U2695 (N_2695,N_2334,N_2279);
and U2696 (N_2696,N_2382,N_2305);
or U2697 (N_2697,N_2316,N_2349);
nor U2698 (N_2698,N_2306,N_2447);
and U2699 (N_2699,N_2453,N_2374);
or U2700 (N_2700,N_2444,N_2459);
nand U2701 (N_2701,N_2469,N_2280);
xor U2702 (N_2702,N_2291,N_2283);
or U2703 (N_2703,N_2290,N_2346);
and U2704 (N_2704,N_2398,N_2367);
nand U2705 (N_2705,N_2402,N_2377);
and U2706 (N_2706,N_2359,N_2282);
nor U2707 (N_2707,N_2393,N_2366);
nor U2708 (N_2708,N_2471,N_2286);
nor U2709 (N_2709,N_2409,N_2412);
xor U2710 (N_2710,N_2478,N_2401);
and U2711 (N_2711,N_2371,N_2449);
nor U2712 (N_2712,N_2494,N_2429);
nor U2713 (N_2713,N_2450,N_2361);
nor U2714 (N_2714,N_2490,N_2307);
nor U2715 (N_2715,N_2312,N_2275);
xor U2716 (N_2716,N_2436,N_2417);
or U2717 (N_2717,N_2498,N_2318);
nor U2718 (N_2718,N_2291,N_2427);
nand U2719 (N_2719,N_2255,N_2413);
xor U2720 (N_2720,N_2352,N_2360);
nand U2721 (N_2721,N_2374,N_2426);
nor U2722 (N_2722,N_2451,N_2335);
and U2723 (N_2723,N_2479,N_2252);
and U2724 (N_2724,N_2425,N_2434);
nor U2725 (N_2725,N_2366,N_2372);
or U2726 (N_2726,N_2376,N_2367);
and U2727 (N_2727,N_2250,N_2399);
nor U2728 (N_2728,N_2256,N_2317);
xor U2729 (N_2729,N_2332,N_2462);
or U2730 (N_2730,N_2307,N_2486);
or U2731 (N_2731,N_2358,N_2347);
or U2732 (N_2732,N_2483,N_2335);
or U2733 (N_2733,N_2269,N_2469);
or U2734 (N_2734,N_2445,N_2487);
or U2735 (N_2735,N_2403,N_2405);
xor U2736 (N_2736,N_2422,N_2250);
nor U2737 (N_2737,N_2389,N_2439);
or U2738 (N_2738,N_2332,N_2330);
and U2739 (N_2739,N_2331,N_2460);
nor U2740 (N_2740,N_2390,N_2333);
nor U2741 (N_2741,N_2444,N_2427);
nor U2742 (N_2742,N_2261,N_2263);
xor U2743 (N_2743,N_2453,N_2427);
or U2744 (N_2744,N_2494,N_2411);
and U2745 (N_2745,N_2428,N_2354);
and U2746 (N_2746,N_2416,N_2256);
xor U2747 (N_2747,N_2350,N_2341);
nor U2748 (N_2748,N_2264,N_2347);
xor U2749 (N_2749,N_2381,N_2429);
xnor U2750 (N_2750,N_2501,N_2683);
nand U2751 (N_2751,N_2615,N_2636);
xor U2752 (N_2752,N_2572,N_2703);
xor U2753 (N_2753,N_2570,N_2708);
and U2754 (N_2754,N_2706,N_2730);
or U2755 (N_2755,N_2722,N_2532);
and U2756 (N_2756,N_2569,N_2548);
or U2757 (N_2757,N_2607,N_2596);
or U2758 (N_2758,N_2540,N_2566);
nor U2759 (N_2759,N_2676,N_2561);
nand U2760 (N_2760,N_2654,N_2662);
xnor U2761 (N_2761,N_2579,N_2687);
or U2762 (N_2762,N_2633,N_2527);
nand U2763 (N_2763,N_2549,N_2692);
and U2764 (N_2764,N_2659,N_2724);
and U2765 (N_2765,N_2719,N_2592);
and U2766 (N_2766,N_2515,N_2520);
and U2767 (N_2767,N_2559,N_2550);
and U2768 (N_2768,N_2589,N_2747);
xnor U2769 (N_2769,N_2737,N_2510);
xor U2770 (N_2770,N_2732,N_2564);
nor U2771 (N_2771,N_2547,N_2630);
and U2772 (N_2772,N_2695,N_2707);
and U2773 (N_2773,N_2541,N_2715);
nor U2774 (N_2774,N_2641,N_2598);
nor U2775 (N_2775,N_2728,N_2552);
nor U2776 (N_2776,N_2524,N_2593);
and U2777 (N_2777,N_2500,N_2698);
xor U2778 (N_2778,N_2702,N_2642);
and U2779 (N_2779,N_2583,N_2678);
xnor U2780 (N_2780,N_2689,N_2666);
nor U2781 (N_2781,N_2535,N_2723);
xor U2782 (N_2782,N_2656,N_2647);
nand U2783 (N_2783,N_2512,N_2617);
xor U2784 (N_2784,N_2660,N_2643);
nor U2785 (N_2785,N_2694,N_2578);
nand U2786 (N_2786,N_2717,N_2712);
and U2787 (N_2787,N_2628,N_2551);
xnor U2788 (N_2788,N_2612,N_2721);
nand U2789 (N_2789,N_2517,N_2711);
nor U2790 (N_2790,N_2710,N_2667);
xor U2791 (N_2791,N_2544,N_2685);
nor U2792 (N_2792,N_2634,N_2704);
or U2793 (N_2793,N_2701,N_2690);
nand U2794 (N_2794,N_2713,N_2502);
xor U2795 (N_2795,N_2584,N_2522);
nand U2796 (N_2796,N_2684,N_2665);
or U2797 (N_2797,N_2679,N_2650);
or U2798 (N_2798,N_2626,N_2733);
xnor U2799 (N_2799,N_2590,N_2597);
nand U2800 (N_2800,N_2623,N_2681);
nor U2801 (N_2801,N_2649,N_2503);
xnor U2802 (N_2802,N_2748,N_2591);
and U2803 (N_2803,N_2652,N_2506);
nor U2804 (N_2804,N_2675,N_2677);
or U2805 (N_2805,N_2619,N_2720);
nor U2806 (N_2806,N_2582,N_2726);
and U2807 (N_2807,N_2668,N_2575);
or U2808 (N_2808,N_2514,N_2568);
and U2809 (N_2809,N_2571,N_2709);
or U2810 (N_2810,N_2622,N_2587);
and U2811 (N_2811,N_2727,N_2577);
nor U2812 (N_2812,N_2671,N_2627);
nand U2813 (N_2813,N_2658,N_2739);
and U2814 (N_2814,N_2505,N_2686);
nor U2815 (N_2815,N_2504,N_2530);
or U2816 (N_2816,N_2508,N_2743);
nor U2817 (N_2817,N_2543,N_2537);
xor U2818 (N_2818,N_2714,N_2554);
xnor U2819 (N_2819,N_2638,N_2734);
or U2820 (N_2820,N_2576,N_2538);
or U2821 (N_2821,N_2509,N_2688);
and U2822 (N_2822,N_2624,N_2664);
xor U2823 (N_2823,N_2574,N_2725);
or U2824 (N_2824,N_2608,N_2542);
xnor U2825 (N_2825,N_2699,N_2605);
and U2826 (N_2826,N_2744,N_2610);
nor U2827 (N_2827,N_2657,N_2663);
nand U2828 (N_2828,N_2588,N_2594);
or U2829 (N_2829,N_2556,N_2516);
and U2830 (N_2830,N_2742,N_2735);
and U2831 (N_2831,N_2738,N_2640);
and U2832 (N_2832,N_2629,N_2533);
or U2833 (N_2833,N_2661,N_2613);
nand U2834 (N_2834,N_2511,N_2562);
xnor U2835 (N_2835,N_2632,N_2606);
xor U2836 (N_2836,N_2609,N_2696);
xor U2837 (N_2837,N_2534,N_2580);
nor U2838 (N_2838,N_2651,N_2741);
xnor U2839 (N_2839,N_2653,N_2518);
nand U2840 (N_2840,N_2546,N_2565);
xor U2841 (N_2841,N_2674,N_2637);
or U2842 (N_2842,N_2560,N_2697);
nor U2843 (N_2843,N_2693,N_2655);
xor U2844 (N_2844,N_2620,N_2746);
or U2845 (N_2845,N_2603,N_2585);
or U2846 (N_2846,N_2700,N_2595);
xor U2847 (N_2847,N_2736,N_2600);
and U2848 (N_2848,N_2602,N_2639);
xor U2849 (N_2849,N_2729,N_2731);
or U2850 (N_2850,N_2555,N_2519);
nor U2851 (N_2851,N_2604,N_2507);
xnor U2852 (N_2852,N_2586,N_2545);
and U2853 (N_2853,N_2648,N_2558);
or U2854 (N_2854,N_2557,N_2749);
and U2855 (N_2855,N_2567,N_2616);
nand U2856 (N_2856,N_2621,N_2618);
or U2857 (N_2857,N_2581,N_2745);
and U2858 (N_2858,N_2644,N_2513);
and U2859 (N_2859,N_2669,N_2523);
and U2860 (N_2860,N_2529,N_2526);
nand U2861 (N_2861,N_2525,N_2635);
nor U2862 (N_2862,N_2673,N_2716);
nor U2863 (N_2863,N_2611,N_2691);
xnor U2864 (N_2864,N_2645,N_2705);
and U2865 (N_2865,N_2646,N_2528);
nand U2866 (N_2866,N_2718,N_2601);
or U2867 (N_2867,N_2599,N_2625);
and U2868 (N_2868,N_2680,N_2539);
xor U2869 (N_2869,N_2682,N_2521);
nand U2870 (N_2870,N_2631,N_2672);
or U2871 (N_2871,N_2670,N_2536);
or U2872 (N_2872,N_2614,N_2563);
nor U2873 (N_2873,N_2553,N_2573);
and U2874 (N_2874,N_2531,N_2740);
nand U2875 (N_2875,N_2568,N_2734);
and U2876 (N_2876,N_2620,N_2607);
nor U2877 (N_2877,N_2633,N_2665);
nand U2878 (N_2878,N_2567,N_2724);
or U2879 (N_2879,N_2555,N_2713);
nor U2880 (N_2880,N_2668,N_2744);
xnor U2881 (N_2881,N_2701,N_2619);
nand U2882 (N_2882,N_2707,N_2508);
nand U2883 (N_2883,N_2506,N_2707);
xor U2884 (N_2884,N_2567,N_2742);
and U2885 (N_2885,N_2521,N_2546);
and U2886 (N_2886,N_2579,N_2703);
or U2887 (N_2887,N_2708,N_2667);
xnor U2888 (N_2888,N_2527,N_2589);
or U2889 (N_2889,N_2511,N_2722);
and U2890 (N_2890,N_2633,N_2518);
or U2891 (N_2891,N_2568,N_2724);
xor U2892 (N_2892,N_2629,N_2714);
or U2893 (N_2893,N_2566,N_2538);
or U2894 (N_2894,N_2684,N_2577);
and U2895 (N_2895,N_2620,N_2739);
nor U2896 (N_2896,N_2605,N_2541);
nand U2897 (N_2897,N_2670,N_2627);
xor U2898 (N_2898,N_2664,N_2644);
nand U2899 (N_2899,N_2500,N_2580);
xnor U2900 (N_2900,N_2534,N_2635);
or U2901 (N_2901,N_2526,N_2701);
nand U2902 (N_2902,N_2641,N_2688);
or U2903 (N_2903,N_2585,N_2572);
nand U2904 (N_2904,N_2601,N_2709);
xor U2905 (N_2905,N_2607,N_2695);
and U2906 (N_2906,N_2502,N_2586);
or U2907 (N_2907,N_2648,N_2687);
xnor U2908 (N_2908,N_2618,N_2593);
or U2909 (N_2909,N_2650,N_2741);
or U2910 (N_2910,N_2645,N_2578);
nand U2911 (N_2911,N_2611,N_2580);
xor U2912 (N_2912,N_2680,N_2620);
or U2913 (N_2913,N_2733,N_2655);
nand U2914 (N_2914,N_2716,N_2623);
and U2915 (N_2915,N_2703,N_2687);
or U2916 (N_2916,N_2633,N_2635);
and U2917 (N_2917,N_2588,N_2715);
nor U2918 (N_2918,N_2598,N_2549);
and U2919 (N_2919,N_2505,N_2722);
nand U2920 (N_2920,N_2680,N_2716);
nand U2921 (N_2921,N_2572,N_2715);
and U2922 (N_2922,N_2588,N_2700);
or U2923 (N_2923,N_2512,N_2557);
nor U2924 (N_2924,N_2512,N_2518);
nor U2925 (N_2925,N_2523,N_2578);
and U2926 (N_2926,N_2619,N_2664);
or U2927 (N_2927,N_2583,N_2615);
and U2928 (N_2928,N_2562,N_2708);
and U2929 (N_2929,N_2639,N_2677);
and U2930 (N_2930,N_2604,N_2732);
nor U2931 (N_2931,N_2518,N_2733);
nor U2932 (N_2932,N_2635,N_2665);
xnor U2933 (N_2933,N_2674,N_2570);
nand U2934 (N_2934,N_2705,N_2695);
xor U2935 (N_2935,N_2523,N_2576);
nand U2936 (N_2936,N_2699,N_2738);
xor U2937 (N_2937,N_2529,N_2680);
nand U2938 (N_2938,N_2716,N_2500);
or U2939 (N_2939,N_2611,N_2643);
nand U2940 (N_2940,N_2546,N_2705);
and U2941 (N_2941,N_2567,N_2500);
or U2942 (N_2942,N_2638,N_2596);
or U2943 (N_2943,N_2734,N_2687);
nor U2944 (N_2944,N_2692,N_2656);
nand U2945 (N_2945,N_2562,N_2636);
nand U2946 (N_2946,N_2628,N_2607);
nor U2947 (N_2947,N_2554,N_2506);
and U2948 (N_2948,N_2501,N_2587);
or U2949 (N_2949,N_2538,N_2612);
nor U2950 (N_2950,N_2592,N_2555);
xor U2951 (N_2951,N_2551,N_2531);
xor U2952 (N_2952,N_2653,N_2717);
and U2953 (N_2953,N_2654,N_2695);
nor U2954 (N_2954,N_2718,N_2556);
nand U2955 (N_2955,N_2616,N_2723);
nand U2956 (N_2956,N_2577,N_2593);
and U2957 (N_2957,N_2504,N_2619);
nor U2958 (N_2958,N_2615,N_2553);
and U2959 (N_2959,N_2511,N_2514);
nor U2960 (N_2960,N_2558,N_2504);
nor U2961 (N_2961,N_2579,N_2639);
nand U2962 (N_2962,N_2630,N_2583);
nor U2963 (N_2963,N_2608,N_2679);
and U2964 (N_2964,N_2657,N_2516);
xnor U2965 (N_2965,N_2631,N_2544);
and U2966 (N_2966,N_2730,N_2518);
and U2967 (N_2967,N_2653,N_2602);
and U2968 (N_2968,N_2669,N_2728);
or U2969 (N_2969,N_2634,N_2590);
or U2970 (N_2970,N_2553,N_2578);
xor U2971 (N_2971,N_2585,N_2651);
xnor U2972 (N_2972,N_2527,N_2659);
and U2973 (N_2973,N_2615,N_2554);
nand U2974 (N_2974,N_2686,N_2628);
xnor U2975 (N_2975,N_2732,N_2580);
nor U2976 (N_2976,N_2596,N_2598);
xor U2977 (N_2977,N_2511,N_2592);
or U2978 (N_2978,N_2677,N_2578);
nor U2979 (N_2979,N_2690,N_2671);
nand U2980 (N_2980,N_2562,N_2597);
or U2981 (N_2981,N_2636,N_2585);
and U2982 (N_2982,N_2697,N_2684);
xor U2983 (N_2983,N_2624,N_2738);
and U2984 (N_2984,N_2713,N_2535);
nand U2985 (N_2985,N_2530,N_2737);
nor U2986 (N_2986,N_2596,N_2730);
xnor U2987 (N_2987,N_2638,N_2745);
and U2988 (N_2988,N_2650,N_2692);
nor U2989 (N_2989,N_2706,N_2583);
nand U2990 (N_2990,N_2731,N_2674);
nand U2991 (N_2991,N_2612,N_2665);
nor U2992 (N_2992,N_2704,N_2656);
or U2993 (N_2993,N_2566,N_2680);
xor U2994 (N_2994,N_2639,N_2589);
or U2995 (N_2995,N_2715,N_2678);
or U2996 (N_2996,N_2746,N_2741);
xnor U2997 (N_2997,N_2659,N_2704);
and U2998 (N_2998,N_2605,N_2543);
nand U2999 (N_2999,N_2588,N_2699);
nor U3000 (N_3000,N_2839,N_2758);
nor U3001 (N_3001,N_2955,N_2876);
nand U3002 (N_3002,N_2789,N_2852);
and U3003 (N_3003,N_2919,N_2815);
or U3004 (N_3004,N_2980,N_2984);
and U3005 (N_3005,N_2996,N_2885);
or U3006 (N_3006,N_2987,N_2752);
nand U3007 (N_3007,N_2840,N_2882);
and U3008 (N_3008,N_2872,N_2765);
xnor U3009 (N_3009,N_2766,N_2799);
xor U3010 (N_3010,N_2925,N_2797);
xnor U3011 (N_3011,N_2909,N_2930);
nand U3012 (N_3012,N_2782,N_2786);
and U3013 (N_3013,N_2953,N_2954);
nor U3014 (N_3014,N_2802,N_2798);
nor U3015 (N_3015,N_2877,N_2785);
nor U3016 (N_3016,N_2776,N_2905);
and U3017 (N_3017,N_2933,N_2975);
or U3018 (N_3018,N_2948,N_2808);
xnor U3019 (N_3019,N_2844,N_2801);
xor U3020 (N_3020,N_2965,N_2757);
nor U3021 (N_3021,N_2938,N_2795);
nand U3022 (N_3022,N_2762,N_2773);
nand U3023 (N_3023,N_2884,N_2849);
or U3024 (N_3024,N_2780,N_2932);
nand U3025 (N_3025,N_2914,N_2959);
xor U3026 (N_3026,N_2855,N_2866);
or U3027 (N_3027,N_2807,N_2770);
nand U3028 (N_3028,N_2829,N_2993);
nand U3029 (N_3029,N_2822,N_2875);
or U3030 (N_3030,N_2833,N_2800);
or U3031 (N_3031,N_2806,N_2767);
xnor U3032 (N_3032,N_2810,N_2777);
or U3033 (N_3033,N_2994,N_2768);
nand U3034 (N_3034,N_2856,N_2963);
nand U3035 (N_3035,N_2887,N_2957);
or U3036 (N_3036,N_2937,N_2899);
xnor U3037 (N_3037,N_2972,N_2790);
nor U3038 (N_3038,N_2900,N_2968);
nor U3039 (N_3039,N_2854,N_2897);
nor U3040 (N_3040,N_2778,N_2843);
and U3041 (N_3041,N_2969,N_2956);
nor U3042 (N_3042,N_2772,N_2929);
nor U3043 (N_3043,N_2988,N_2788);
nor U3044 (N_3044,N_2967,N_2936);
nor U3045 (N_3045,N_2845,N_2754);
nand U3046 (N_3046,N_2809,N_2986);
nand U3047 (N_3047,N_2763,N_2970);
xnor U3048 (N_3048,N_2881,N_2761);
or U3049 (N_3049,N_2838,N_2853);
nor U3050 (N_3050,N_2858,N_2962);
xor U3051 (N_3051,N_2862,N_2983);
nand U3052 (N_3052,N_2913,N_2979);
nor U3053 (N_3053,N_2831,N_2835);
nand U3054 (N_3054,N_2784,N_2868);
or U3055 (N_3055,N_2977,N_2819);
xor U3056 (N_3056,N_2901,N_2774);
nand U3057 (N_3057,N_2997,N_2902);
or U3058 (N_3058,N_2935,N_2817);
and U3059 (N_3059,N_2952,N_2958);
and U3060 (N_3060,N_2787,N_2863);
nand U3061 (N_3061,N_2878,N_2926);
and U3062 (N_3062,N_2803,N_2945);
and U3063 (N_3063,N_2793,N_2889);
nor U3064 (N_3064,N_2794,N_2883);
nand U3065 (N_3065,N_2976,N_2944);
and U3066 (N_3066,N_2851,N_2904);
or U3067 (N_3067,N_2923,N_2960);
xor U3068 (N_3068,N_2850,N_2898);
and U3069 (N_3069,N_2918,N_2792);
nor U3070 (N_3070,N_2907,N_2814);
and U3071 (N_3071,N_2949,N_2992);
nor U3072 (N_3072,N_2771,N_2827);
or U3073 (N_3073,N_2890,N_2874);
nor U3074 (N_3074,N_2865,N_2846);
or U3075 (N_3075,N_2998,N_2871);
nand U3076 (N_3076,N_2895,N_2891);
or U3077 (N_3077,N_2981,N_2880);
and U3078 (N_3078,N_2805,N_2886);
nor U3079 (N_3079,N_2927,N_2811);
and U3080 (N_3080,N_2775,N_2873);
nand U3081 (N_3081,N_2859,N_2911);
or U3082 (N_3082,N_2824,N_2928);
and U3083 (N_3083,N_2922,N_2857);
nand U3084 (N_3084,N_2783,N_2946);
xnor U3085 (N_3085,N_2828,N_2924);
and U3086 (N_3086,N_2908,N_2756);
nand U3087 (N_3087,N_2941,N_2751);
nor U3088 (N_3088,N_2759,N_2921);
xnor U3089 (N_3089,N_2903,N_2834);
xnor U3090 (N_3090,N_2879,N_2985);
nand U3091 (N_3091,N_2951,N_2760);
nor U3092 (N_3092,N_2942,N_2982);
nand U3093 (N_3093,N_2978,N_2818);
xnor U3094 (N_3094,N_2915,N_2820);
nand U3095 (N_3095,N_2779,N_2961);
xor U3096 (N_3096,N_2825,N_2860);
nor U3097 (N_3097,N_2964,N_2750);
or U3098 (N_3098,N_2943,N_2931);
or U3099 (N_3099,N_2869,N_2755);
nor U3100 (N_3100,N_2995,N_2892);
nand U3101 (N_3101,N_2893,N_2950);
nand U3102 (N_3102,N_2781,N_2912);
and U3103 (N_3103,N_2841,N_2847);
xnor U3104 (N_3104,N_2848,N_2990);
nor U3105 (N_3105,N_2826,N_2830);
xnor U3106 (N_3106,N_2769,N_2947);
and U3107 (N_3107,N_2764,N_2864);
and U3108 (N_3108,N_2939,N_2906);
nand U3109 (N_3109,N_2796,N_2974);
or U3110 (N_3110,N_2813,N_2940);
or U3111 (N_3111,N_2753,N_2999);
or U3112 (N_3112,N_2971,N_2966);
and U3113 (N_3113,N_2842,N_2989);
or U3114 (N_3114,N_2888,N_2823);
nand U3115 (N_3115,N_2861,N_2910);
nand U3116 (N_3116,N_2934,N_2917);
and U3117 (N_3117,N_2791,N_2894);
and U3118 (N_3118,N_2896,N_2812);
nor U3119 (N_3119,N_2991,N_2816);
nor U3120 (N_3120,N_2804,N_2916);
and U3121 (N_3121,N_2973,N_2920);
or U3122 (N_3122,N_2837,N_2832);
nor U3123 (N_3123,N_2821,N_2867);
and U3124 (N_3124,N_2870,N_2836);
nor U3125 (N_3125,N_2860,N_2780);
and U3126 (N_3126,N_2752,N_2768);
or U3127 (N_3127,N_2831,N_2872);
and U3128 (N_3128,N_2835,N_2940);
nor U3129 (N_3129,N_2870,N_2859);
nor U3130 (N_3130,N_2761,N_2777);
nor U3131 (N_3131,N_2961,N_2807);
xnor U3132 (N_3132,N_2936,N_2991);
nand U3133 (N_3133,N_2761,N_2843);
nand U3134 (N_3134,N_2943,N_2756);
and U3135 (N_3135,N_2888,N_2851);
xor U3136 (N_3136,N_2850,N_2979);
nand U3137 (N_3137,N_2958,N_2851);
xnor U3138 (N_3138,N_2985,N_2955);
nand U3139 (N_3139,N_2758,N_2765);
nor U3140 (N_3140,N_2769,N_2760);
xor U3141 (N_3141,N_2779,N_2782);
xnor U3142 (N_3142,N_2882,N_2901);
or U3143 (N_3143,N_2975,N_2945);
nand U3144 (N_3144,N_2841,N_2997);
nor U3145 (N_3145,N_2923,N_2842);
xnor U3146 (N_3146,N_2965,N_2771);
or U3147 (N_3147,N_2805,N_2907);
or U3148 (N_3148,N_2963,N_2767);
and U3149 (N_3149,N_2821,N_2890);
and U3150 (N_3150,N_2798,N_2780);
nand U3151 (N_3151,N_2885,N_2755);
nor U3152 (N_3152,N_2993,N_2956);
nor U3153 (N_3153,N_2894,N_2859);
or U3154 (N_3154,N_2883,N_2840);
nand U3155 (N_3155,N_2894,N_2921);
nand U3156 (N_3156,N_2932,N_2996);
nor U3157 (N_3157,N_2796,N_2977);
nand U3158 (N_3158,N_2880,N_2875);
and U3159 (N_3159,N_2812,N_2852);
and U3160 (N_3160,N_2836,N_2834);
nand U3161 (N_3161,N_2815,N_2762);
and U3162 (N_3162,N_2941,N_2995);
and U3163 (N_3163,N_2826,N_2837);
xor U3164 (N_3164,N_2862,N_2914);
and U3165 (N_3165,N_2871,N_2873);
nand U3166 (N_3166,N_2970,N_2867);
nand U3167 (N_3167,N_2807,N_2852);
and U3168 (N_3168,N_2927,N_2848);
nand U3169 (N_3169,N_2868,N_2811);
nor U3170 (N_3170,N_2944,N_2986);
or U3171 (N_3171,N_2777,N_2898);
or U3172 (N_3172,N_2795,N_2797);
or U3173 (N_3173,N_2875,N_2881);
or U3174 (N_3174,N_2911,N_2963);
nand U3175 (N_3175,N_2825,N_2999);
nand U3176 (N_3176,N_2796,N_2887);
nand U3177 (N_3177,N_2948,N_2984);
nor U3178 (N_3178,N_2912,N_2964);
and U3179 (N_3179,N_2813,N_2885);
nor U3180 (N_3180,N_2889,N_2904);
nand U3181 (N_3181,N_2751,N_2771);
xor U3182 (N_3182,N_2848,N_2806);
nand U3183 (N_3183,N_2818,N_2988);
and U3184 (N_3184,N_2856,N_2772);
nand U3185 (N_3185,N_2985,N_2862);
xor U3186 (N_3186,N_2881,N_2990);
nor U3187 (N_3187,N_2905,N_2915);
xnor U3188 (N_3188,N_2933,N_2778);
or U3189 (N_3189,N_2761,N_2772);
or U3190 (N_3190,N_2941,N_2850);
nand U3191 (N_3191,N_2759,N_2981);
nor U3192 (N_3192,N_2754,N_2846);
nor U3193 (N_3193,N_2819,N_2866);
nand U3194 (N_3194,N_2985,N_2928);
xor U3195 (N_3195,N_2841,N_2935);
or U3196 (N_3196,N_2923,N_2858);
nor U3197 (N_3197,N_2767,N_2940);
nand U3198 (N_3198,N_2876,N_2844);
nor U3199 (N_3199,N_2845,N_2843);
xnor U3200 (N_3200,N_2900,N_2862);
nor U3201 (N_3201,N_2848,N_2763);
nor U3202 (N_3202,N_2902,N_2876);
xor U3203 (N_3203,N_2861,N_2984);
xor U3204 (N_3204,N_2965,N_2989);
xnor U3205 (N_3205,N_2753,N_2876);
xnor U3206 (N_3206,N_2756,N_2788);
nor U3207 (N_3207,N_2798,N_2807);
xor U3208 (N_3208,N_2929,N_2949);
nor U3209 (N_3209,N_2933,N_2757);
xor U3210 (N_3210,N_2783,N_2793);
and U3211 (N_3211,N_2938,N_2920);
nor U3212 (N_3212,N_2920,N_2813);
or U3213 (N_3213,N_2977,N_2783);
and U3214 (N_3214,N_2892,N_2813);
or U3215 (N_3215,N_2763,N_2827);
nor U3216 (N_3216,N_2973,N_2850);
nor U3217 (N_3217,N_2948,N_2892);
xnor U3218 (N_3218,N_2872,N_2993);
nor U3219 (N_3219,N_2801,N_2805);
nand U3220 (N_3220,N_2991,N_2902);
xnor U3221 (N_3221,N_2778,N_2856);
and U3222 (N_3222,N_2830,N_2759);
nor U3223 (N_3223,N_2978,N_2923);
or U3224 (N_3224,N_2753,N_2968);
nand U3225 (N_3225,N_2855,N_2967);
xor U3226 (N_3226,N_2965,N_2970);
and U3227 (N_3227,N_2968,N_2986);
and U3228 (N_3228,N_2838,N_2789);
or U3229 (N_3229,N_2884,N_2796);
or U3230 (N_3230,N_2845,N_2974);
and U3231 (N_3231,N_2883,N_2886);
or U3232 (N_3232,N_2772,N_2857);
and U3233 (N_3233,N_2976,N_2789);
nor U3234 (N_3234,N_2978,N_2972);
xnor U3235 (N_3235,N_2939,N_2882);
or U3236 (N_3236,N_2979,N_2867);
and U3237 (N_3237,N_2983,N_2974);
nor U3238 (N_3238,N_2956,N_2884);
or U3239 (N_3239,N_2979,N_2924);
or U3240 (N_3240,N_2822,N_2860);
xor U3241 (N_3241,N_2933,N_2983);
and U3242 (N_3242,N_2983,N_2889);
nor U3243 (N_3243,N_2853,N_2817);
xnor U3244 (N_3244,N_2904,N_2968);
nand U3245 (N_3245,N_2907,N_2800);
nor U3246 (N_3246,N_2785,N_2750);
nor U3247 (N_3247,N_2829,N_2998);
nand U3248 (N_3248,N_2781,N_2986);
and U3249 (N_3249,N_2993,N_2781);
and U3250 (N_3250,N_3231,N_3068);
and U3251 (N_3251,N_3205,N_3196);
xor U3252 (N_3252,N_3005,N_3041);
or U3253 (N_3253,N_3207,N_3108);
or U3254 (N_3254,N_3082,N_3209);
or U3255 (N_3255,N_3114,N_3055);
or U3256 (N_3256,N_3084,N_3248);
xor U3257 (N_3257,N_3092,N_3034);
and U3258 (N_3258,N_3160,N_3139);
nor U3259 (N_3259,N_3039,N_3140);
xnor U3260 (N_3260,N_3045,N_3053);
or U3261 (N_3261,N_3064,N_3003);
nand U3262 (N_3262,N_3130,N_3019);
nand U3263 (N_3263,N_3177,N_3184);
or U3264 (N_3264,N_3200,N_3129);
or U3265 (N_3265,N_3069,N_3116);
or U3266 (N_3266,N_3168,N_3101);
xor U3267 (N_3267,N_3199,N_3020);
nor U3268 (N_3268,N_3011,N_3193);
or U3269 (N_3269,N_3047,N_3010);
xor U3270 (N_3270,N_3042,N_3035);
nand U3271 (N_3271,N_3171,N_3172);
xor U3272 (N_3272,N_3127,N_3179);
nand U3273 (N_3273,N_3178,N_3164);
nand U3274 (N_3274,N_3033,N_3049);
nand U3275 (N_3275,N_3208,N_3137);
nand U3276 (N_3276,N_3183,N_3211);
xnor U3277 (N_3277,N_3221,N_3070);
xor U3278 (N_3278,N_3192,N_3220);
or U3279 (N_3279,N_3066,N_3214);
or U3280 (N_3280,N_3223,N_3028);
or U3281 (N_3281,N_3012,N_3075);
nand U3282 (N_3282,N_3191,N_3097);
xnor U3283 (N_3283,N_3198,N_3222);
or U3284 (N_3284,N_3001,N_3176);
nor U3285 (N_3285,N_3229,N_3190);
or U3286 (N_3286,N_3225,N_3206);
or U3287 (N_3287,N_3115,N_3197);
and U3288 (N_3288,N_3203,N_3113);
nor U3289 (N_3289,N_3046,N_3030);
and U3290 (N_3290,N_3210,N_3133);
or U3291 (N_3291,N_3175,N_3057);
and U3292 (N_3292,N_3050,N_3161);
or U3293 (N_3293,N_3119,N_3150);
or U3294 (N_3294,N_3093,N_3156);
nand U3295 (N_3295,N_3189,N_3100);
or U3296 (N_3296,N_3226,N_3106);
or U3297 (N_3297,N_3105,N_3083);
and U3298 (N_3298,N_3152,N_3123);
xor U3299 (N_3299,N_3024,N_3134);
or U3300 (N_3300,N_3163,N_3102);
nand U3301 (N_3301,N_3023,N_3228);
or U3302 (N_3302,N_3195,N_3167);
or U3303 (N_3303,N_3219,N_3096);
xnor U3304 (N_3304,N_3058,N_3224);
xnor U3305 (N_3305,N_3107,N_3235);
xnor U3306 (N_3306,N_3144,N_3218);
nand U3307 (N_3307,N_3087,N_3015);
nand U3308 (N_3308,N_3146,N_3165);
xor U3309 (N_3309,N_3056,N_3073);
or U3310 (N_3310,N_3004,N_3088);
or U3311 (N_3311,N_3240,N_3180);
or U3312 (N_3312,N_3040,N_3006);
xnor U3313 (N_3313,N_3060,N_3154);
or U3314 (N_3314,N_3076,N_3090);
nor U3315 (N_3315,N_3079,N_3249);
xnor U3316 (N_3316,N_3246,N_3008);
nor U3317 (N_3317,N_3048,N_3120);
or U3318 (N_3318,N_3109,N_3149);
nor U3319 (N_3319,N_3065,N_3018);
or U3320 (N_3320,N_3014,N_3086);
nand U3321 (N_3321,N_3043,N_3021);
xor U3322 (N_3322,N_3170,N_3081);
or U3323 (N_3323,N_3091,N_3245);
nand U3324 (N_3324,N_3121,N_3017);
xnor U3325 (N_3325,N_3099,N_3051);
nor U3326 (N_3326,N_3032,N_3009);
or U3327 (N_3327,N_3212,N_3232);
or U3328 (N_3328,N_3131,N_3244);
and U3329 (N_3329,N_3238,N_3182);
or U3330 (N_3330,N_3063,N_3242);
nand U3331 (N_3331,N_3078,N_3243);
and U3332 (N_3332,N_3126,N_3094);
nor U3333 (N_3333,N_3071,N_3132);
or U3334 (N_3334,N_3111,N_3110);
xnor U3335 (N_3335,N_3204,N_3061);
and U3336 (N_3336,N_3054,N_3128);
nand U3337 (N_3337,N_3026,N_3241);
nand U3338 (N_3338,N_3234,N_3044);
nand U3339 (N_3339,N_3000,N_3080);
nor U3340 (N_3340,N_3072,N_3216);
nor U3341 (N_3341,N_3142,N_3153);
xor U3342 (N_3342,N_3162,N_3202);
nor U3343 (N_3343,N_3155,N_3141);
xnor U3344 (N_3344,N_3052,N_3118);
nor U3345 (N_3345,N_3159,N_3239);
and U3346 (N_3346,N_3157,N_3098);
nand U3347 (N_3347,N_3125,N_3077);
nand U3348 (N_3348,N_3217,N_3215);
nor U3349 (N_3349,N_3213,N_3143);
xnor U3350 (N_3350,N_3201,N_3074);
xor U3351 (N_3351,N_3122,N_3145);
xnor U3352 (N_3352,N_3166,N_3029);
and U3353 (N_3353,N_3036,N_3031);
xor U3354 (N_3354,N_3188,N_3135);
or U3355 (N_3355,N_3169,N_3187);
nor U3356 (N_3356,N_3138,N_3002);
and U3357 (N_3357,N_3147,N_3233);
or U3358 (N_3358,N_3185,N_3059);
nand U3359 (N_3359,N_3016,N_3117);
and U3360 (N_3360,N_3027,N_3104);
nand U3361 (N_3361,N_3067,N_3173);
xor U3362 (N_3362,N_3124,N_3237);
nor U3363 (N_3363,N_3230,N_3037);
xor U3364 (N_3364,N_3236,N_3158);
nor U3365 (N_3365,N_3151,N_3112);
xor U3366 (N_3366,N_3025,N_3013);
or U3367 (N_3367,N_3022,N_3148);
and U3368 (N_3368,N_3085,N_3089);
xor U3369 (N_3369,N_3007,N_3103);
and U3370 (N_3370,N_3181,N_3136);
or U3371 (N_3371,N_3194,N_3227);
nand U3372 (N_3372,N_3038,N_3186);
and U3373 (N_3373,N_3174,N_3247);
nand U3374 (N_3374,N_3062,N_3095);
nand U3375 (N_3375,N_3159,N_3191);
nor U3376 (N_3376,N_3062,N_3134);
or U3377 (N_3377,N_3089,N_3173);
or U3378 (N_3378,N_3051,N_3082);
nor U3379 (N_3379,N_3032,N_3103);
xor U3380 (N_3380,N_3100,N_3050);
or U3381 (N_3381,N_3166,N_3240);
nor U3382 (N_3382,N_3167,N_3160);
nor U3383 (N_3383,N_3118,N_3096);
or U3384 (N_3384,N_3232,N_3031);
or U3385 (N_3385,N_3013,N_3161);
nor U3386 (N_3386,N_3185,N_3104);
or U3387 (N_3387,N_3204,N_3246);
and U3388 (N_3388,N_3002,N_3020);
xor U3389 (N_3389,N_3207,N_3152);
nand U3390 (N_3390,N_3073,N_3047);
nor U3391 (N_3391,N_3071,N_3033);
xnor U3392 (N_3392,N_3086,N_3009);
nand U3393 (N_3393,N_3235,N_3171);
and U3394 (N_3394,N_3120,N_3249);
or U3395 (N_3395,N_3152,N_3142);
nor U3396 (N_3396,N_3059,N_3036);
nand U3397 (N_3397,N_3010,N_3249);
nand U3398 (N_3398,N_3049,N_3004);
and U3399 (N_3399,N_3218,N_3074);
xor U3400 (N_3400,N_3065,N_3105);
and U3401 (N_3401,N_3159,N_3162);
xnor U3402 (N_3402,N_3150,N_3172);
or U3403 (N_3403,N_3141,N_3138);
nand U3404 (N_3404,N_3065,N_3238);
and U3405 (N_3405,N_3069,N_3182);
xor U3406 (N_3406,N_3063,N_3173);
nand U3407 (N_3407,N_3183,N_3075);
or U3408 (N_3408,N_3233,N_3182);
nor U3409 (N_3409,N_3128,N_3167);
and U3410 (N_3410,N_3105,N_3214);
nand U3411 (N_3411,N_3087,N_3029);
nand U3412 (N_3412,N_3192,N_3053);
nor U3413 (N_3413,N_3218,N_3197);
xnor U3414 (N_3414,N_3238,N_3203);
or U3415 (N_3415,N_3219,N_3236);
nor U3416 (N_3416,N_3079,N_3240);
or U3417 (N_3417,N_3248,N_3200);
xor U3418 (N_3418,N_3216,N_3047);
xor U3419 (N_3419,N_3066,N_3023);
and U3420 (N_3420,N_3038,N_3190);
nor U3421 (N_3421,N_3209,N_3114);
nor U3422 (N_3422,N_3097,N_3131);
nor U3423 (N_3423,N_3023,N_3007);
nor U3424 (N_3424,N_3190,N_3042);
nor U3425 (N_3425,N_3194,N_3198);
or U3426 (N_3426,N_3171,N_3084);
nand U3427 (N_3427,N_3213,N_3174);
and U3428 (N_3428,N_3130,N_3143);
nand U3429 (N_3429,N_3165,N_3116);
nor U3430 (N_3430,N_3036,N_3116);
and U3431 (N_3431,N_3111,N_3193);
nand U3432 (N_3432,N_3045,N_3191);
nor U3433 (N_3433,N_3249,N_3223);
nand U3434 (N_3434,N_3039,N_3217);
xnor U3435 (N_3435,N_3232,N_3220);
nand U3436 (N_3436,N_3107,N_3212);
or U3437 (N_3437,N_3244,N_3174);
and U3438 (N_3438,N_3099,N_3085);
and U3439 (N_3439,N_3132,N_3072);
nor U3440 (N_3440,N_3154,N_3102);
xor U3441 (N_3441,N_3106,N_3189);
or U3442 (N_3442,N_3223,N_3154);
xor U3443 (N_3443,N_3200,N_3050);
nand U3444 (N_3444,N_3023,N_3240);
xnor U3445 (N_3445,N_3132,N_3098);
nor U3446 (N_3446,N_3012,N_3205);
nand U3447 (N_3447,N_3160,N_3013);
xnor U3448 (N_3448,N_3157,N_3195);
or U3449 (N_3449,N_3021,N_3085);
xor U3450 (N_3450,N_3071,N_3123);
nor U3451 (N_3451,N_3081,N_3038);
and U3452 (N_3452,N_3139,N_3244);
xor U3453 (N_3453,N_3045,N_3120);
nor U3454 (N_3454,N_3139,N_3065);
nand U3455 (N_3455,N_3063,N_3026);
and U3456 (N_3456,N_3145,N_3159);
nor U3457 (N_3457,N_3052,N_3077);
nand U3458 (N_3458,N_3216,N_3207);
or U3459 (N_3459,N_3075,N_3006);
or U3460 (N_3460,N_3056,N_3155);
or U3461 (N_3461,N_3026,N_3204);
nand U3462 (N_3462,N_3109,N_3044);
and U3463 (N_3463,N_3138,N_3235);
nand U3464 (N_3464,N_3014,N_3032);
or U3465 (N_3465,N_3227,N_3190);
nor U3466 (N_3466,N_3061,N_3023);
or U3467 (N_3467,N_3001,N_3190);
or U3468 (N_3468,N_3023,N_3045);
nor U3469 (N_3469,N_3107,N_3089);
nand U3470 (N_3470,N_3061,N_3094);
xor U3471 (N_3471,N_3082,N_3112);
xor U3472 (N_3472,N_3062,N_3208);
or U3473 (N_3473,N_3119,N_3117);
nor U3474 (N_3474,N_3006,N_3034);
nor U3475 (N_3475,N_3237,N_3125);
nor U3476 (N_3476,N_3102,N_3040);
or U3477 (N_3477,N_3128,N_3241);
and U3478 (N_3478,N_3235,N_3119);
and U3479 (N_3479,N_3029,N_3007);
xor U3480 (N_3480,N_3229,N_3168);
and U3481 (N_3481,N_3154,N_3012);
and U3482 (N_3482,N_3102,N_3194);
xor U3483 (N_3483,N_3180,N_3023);
and U3484 (N_3484,N_3143,N_3003);
or U3485 (N_3485,N_3141,N_3224);
xnor U3486 (N_3486,N_3193,N_3115);
and U3487 (N_3487,N_3102,N_3156);
nor U3488 (N_3488,N_3207,N_3083);
xnor U3489 (N_3489,N_3087,N_3068);
and U3490 (N_3490,N_3201,N_3124);
nand U3491 (N_3491,N_3224,N_3181);
nor U3492 (N_3492,N_3152,N_3039);
or U3493 (N_3493,N_3233,N_3249);
and U3494 (N_3494,N_3010,N_3235);
or U3495 (N_3495,N_3049,N_3218);
nor U3496 (N_3496,N_3134,N_3053);
xnor U3497 (N_3497,N_3079,N_3147);
nor U3498 (N_3498,N_3029,N_3079);
xor U3499 (N_3499,N_3039,N_3177);
nand U3500 (N_3500,N_3306,N_3365);
and U3501 (N_3501,N_3399,N_3449);
xnor U3502 (N_3502,N_3491,N_3357);
nor U3503 (N_3503,N_3451,N_3418);
xnor U3504 (N_3504,N_3356,N_3408);
or U3505 (N_3505,N_3286,N_3396);
nand U3506 (N_3506,N_3334,N_3280);
xor U3507 (N_3507,N_3499,N_3293);
nand U3508 (N_3508,N_3482,N_3426);
and U3509 (N_3509,N_3327,N_3300);
xnor U3510 (N_3510,N_3481,N_3381);
and U3511 (N_3511,N_3360,N_3320);
and U3512 (N_3512,N_3270,N_3439);
nor U3513 (N_3513,N_3317,N_3350);
nor U3514 (N_3514,N_3427,N_3269);
xnor U3515 (N_3515,N_3376,N_3315);
or U3516 (N_3516,N_3337,N_3263);
nand U3517 (N_3517,N_3453,N_3390);
or U3518 (N_3518,N_3304,N_3340);
nand U3519 (N_3519,N_3415,N_3323);
nor U3520 (N_3520,N_3438,N_3478);
nor U3521 (N_3521,N_3310,N_3412);
nor U3522 (N_3522,N_3308,N_3281);
nand U3523 (N_3523,N_3452,N_3384);
or U3524 (N_3524,N_3490,N_3431);
xor U3525 (N_3525,N_3256,N_3328);
or U3526 (N_3526,N_3380,N_3254);
and U3527 (N_3527,N_3257,N_3339);
xor U3528 (N_3528,N_3329,N_3421);
nor U3529 (N_3529,N_3285,N_3348);
nand U3530 (N_3530,N_3423,N_3302);
xor U3531 (N_3531,N_3265,N_3261);
and U3532 (N_3532,N_3435,N_3311);
or U3533 (N_3533,N_3312,N_3367);
and U3534 (N_3534,N_3252,N_3400);
and U3535 (N_3535,N_3494,N_3255);
and U3536 (N_3536,N_3375,N_3343);
nand U3537 (N_3537,N_3370,N_3402);
or U3538 (N_3538,N_3457,N_3250);
and U3539 (N_3539,N_3366,N_3467);
xor U3540 (N_3540,N_3424,N_3294);
nor U3541 (N_3541,N_3338,N_3383);
xnor U3542 (N_3542,N_3448,N_3336);
nor U3543 (N_3543,N_3479,N_3260);
or U3544 (N_3544,N_3474,N_3473);
and U3545 (N_3545,N_3434,N_3283);
or U3546 (N_3546,N_3301,N_3437);
and U3547 (N_3547,N_3444,N_3291);
or U3548 (N_3548,N_3272,N_3489);
nand U3549 (N_3549,N_3287,N_3268);
nand U3550 (N_3550,N_3330,N_3361);
and U3551 (N_3551,N_3450,N_3472);
xnor U3552 (N_3552,N_3429,N_3305);
or U3553 (N_3553,N_3468,N_3321);
or U3554 (N_3554,N_3397,N_3319);
nand U3555 (N_3555,N_3284,N_3395);
and U3556 (N_3556,N_3441,N_3498);
xnor U3557 (N_3557,N_3295,N_3352);
xnor U3558 (N_3558,N_3440,N_3409);
xor U3559 (N_3559,N_3391,N_3347);
xor U3560 (N_3560,N_3369,N_3379);
and U3561 (N_3561,N_3278,N_3465);
or U3562 (N_3562,N_3407,N_3303);
nand U3563 (N_3563,N_3388,N_3483);
xnor U3564 (N_3564,N_3460,N_3344);
and U3565 (N_3565,N_3298,N_3410);
nand U3566 (N_3566,N_3401,N_3493);
nand U3567 (N_3567,N_3386,N_3414);
or U3568 (N_3568,N_3349,N_3309);
xor U3569 (N_3569,N_3325,N_3442);
and U3570 (N_3570,N_3436,N_3363);
and U3571 (N_3571,N_3345,N_3471);
nand U3572 (N_3572,N_3413,N_3458);
nor U3573 (N_3573,N_3258,N_3353);
or U3574 (N_3574,N_3372,N_3267);
or U3575 (N_3575,N_3378,N_3475);
and U3576 (N_3576,N_3282,N_3264);
or U3577 (N_3577,N_3411,N_3389);
nor U3578 (N_3578,N_3359,N_3447);
or U3579 (N_3579,N_3420,N_3368);
or U3580 (N_3580,N_3394,N_3314);
or U3581 (N_3581,N_3496,N_3346);
and U3582 (N_3582,N_3406,N_3289);
xor U3583 (N_3583,N_3433,N_3371);
xor U3584 (N_3584,N_3279,N_3432);
and U3585 (N_3585,N_3492,N_3251);
nor U3586 (N_3586,N_3477,N_3292);
xnor U3587 (N_3587,N_3404,N_3488);
nor U3588 (N_3588,N_3335,N_3377);
and U3589 (N_3589,N_3425,N_3480);
nor U3590 (N_3590,N_3373,N_3290);
xnor U3591 (N_3591,N_3318,N_3484);
xor U3592 (N_3592,N_3277,N_3342);
or U3593 (N_3593,N_3351,N_3341);
xor U3594 (N_3594,N_3297,N_3313);
nor U3595 (N_3595,N_3445,N_3495);
nor U3596 (N_3596,N_3461,N_3463);
nand U3597 (N_3597,N_3274,N_3466);
and U3598 (N_3598,N_3398,N_3273);
nor U3599 (N_3599,N_3455,N_3382);
xnor U3600 (N_3600,N_3331,N_3497);
nand U3601 (N_3601,N_3470,N_3259);
nor U3602 (N_3602,N_3476,N_3262);
nor U3603 (N_3603,N_3485,N_3469);
nor U3604 (N_3604,N_3387,N_3428);
nor U3605 (N_3605,N_3322,N_3276);
or U3606 (N_3606,N_3459,N_3419);
and U3607 (N_3607,N_3416,N_3296);
xnor U3608 (N_3608,N_3446,N_3403);
xor U3609 (N_3609,N_3307,N_3354);
and U3610 (N_3610,N_3486,N_3316);
nor U3611 (N_3611,N_3362,N_3443);
nor U3612 (N_3612,N_3358,N_3266);
nor U3613 (N_3613,N_3405,N_3299);
xor U3614 (N_3614,N_3324,N_3417);
xnor U3615 (N_3615,N_3332,N_3355);
or U3616 (N_3616,N_3333,N_3487);
and U3617 (N_3617,N_3462,N_3364);
or U3618 (N_3618,N_3430,N_3253);
nand U3619 (N_3619,N_3275,N_3374);
and U3620 (N_3620,N_3392,N_3271);
nor U3621 (N_3621,N_3422,N_3454);
or U3622 (N_3622,N_3456,N_3326);
xor U3623 (N_3623,N_3393,N_3385);
nor U3624 (N_3624,N_3464,N_3288);
or U3625 (N_3625,N_3414,N_3303);
xnor U3626 (N_3626,N_3331,N_3380);
and U3627 (N_3627,N_3284,N_3487);
nor U3628 (N_3628,N_3329,N_3393);
and U3629 (N_3629,N_3260,N_3498);
nand U3630 (N_3630,N_3335,N_3359);
nor U3631 (N_3631,N_3489,N_3467);
or U3632 (N_3632,N_3254,N_3480);
or U3633 (N_3633,N_3386,N_3256);
xnor U3634 (N_3634,N_3319,N_3394);
and U3635 (N_3635,N_3412,N_3340);
nor U3636 (N_3636,N_3434,N_3266);
or U3637 (N_3637,N_3308,N_3263);
nor U3638 (N_3638,N_3483,N_3430);
nor U3639 (N_3639,N_3491,N_3371);
or U3640 (N_3640,N_3320,N_3284);
xor U3641 (N_3641,N_3326,N_3476);
and U3642 (N_3642,N_3290,N_3463);
nor U3643 (N_3643,N_3456,N_3479);
nor U3644 (N_3644,N_3340,N_3437);
xor U3645 (N_3645,N_3470,N_3459);
and U3646 (N_3646,N_3270,N_3281);
xnor U3647 (N_3647,N_3374,N_3491);
and U3648 (N_3648,N_3318,N_3354);
xnor U3649 (N_3649,N_3325,N_3351);
and U3650 (N_3650,N_3261,N_3349);
xor U3651 (N_3651,N_3305,N_3289);
nand U3652 (N_3652,N_3253,N_3474);
or U3653 (N_3653,N_3463,N_3454);
or U3654 (N_3654,N_3253,N_3254);
or U3655 (N_3655,N_3277,N_3303);
or U3656 (N_3656,N_3374,N_3285);
and U3657 (N_3657,N_3489,N_3417);
nand U3658 (N_3658,N_3353,N_3274);
or U3659 (N_3659,N_3498,N_3302);
nor U3660 (N_3660,N_3263,N_3258);
xor U3661 (N_3661,N_3313,N_3366);
xor U3662 (N_3662,N_3275,N_3379);
nor U3663 (N_3663,N_3430,N_3415);
nand U3664 (N_3664,N_3361,N_3494);
and U3665 (N_3665,N_3354,N_3303);
and U3666 (N_3666,N_3385,N_3495);
and U3667 (N_3667,N_3265,N_3361);
xnor U3668 (N_3668,N_3472,N_3380);
nand U3669 (N_3669,N_3261,N_3404);
or U3670 (N_3670,N_3326,N_3458);
nand U3671 (N_3671,N_3462,N_3491);
nor U3672 (N_3672,N_3286,N_3372);
nand U3673 (N_3673,N_3495,N_3388);
or U3674 (N_3674,N_3475,N_3319);
or U3675 (N_3675,N_3301,N_3433);
and U3676 (N_3676,N_3285,N_3304);
nand U3677 (N_3677,N_3463,N_3439);
or U3678 (N_3678,N_3416,N_3337);
nor U3679 (N_3679,N_3285,N_3373);
nand U3680 (N_3680,N_3309,N_3396);
nor U3681 (N_3681,N_3307,N_3416);
nand U3682 (N_3682,N_3476,N_3309);
nand U3683 (N_3683,N_3309,N_3306);
or U3684 (N_3684,N_3412,N_3305);
xor U3685 (N_3685,N_3392,N_3482);
xnor U3686 (N_3686,N_3465,N_3352);
nand U3687 (N_3687,N_3252,N_3439);
nor U3688 (N_3688,N_3333,N_3497);
or U3689 (N_3689,N_3473,N_3353);
nand U3690 (N_3690,N_3439,N_3272);
xnor U3691 (N_3691,N_3322,N_3347);
and U3692 (N_3692,N_3410,N_3423);
or U3693 (N_3693,N_3484,N_3465);
nand U3694 (N_3694,N_3489,N_3369);
nand U3695 (N_3695,N_3300,N_3355);
or U3696 (N_3696,N_3397,N_3297);
nand U3697 (N_3697,N_3428,N_3354);
nor U3698 (N_3698,N_3480,N_3325);
or U3699 (N_3699,N_3343,N_3410);
xor U3700 (N_3700,N_3449,N_3276);
nand U3701 (N_3701,N_3456,N_3418);
and U3702 (N_3702,N_3483,N_3357);
and U3703 (N_3703,N_3404,N_3359);
or U3704 (N_3704,N_3498,N_3325);
nand U3705 (N_3705,N_3391,N_3253);
and U3706 (N_3706,N_3365,N_3373);
and U3707 (N_3707,N_3388,N_3296);
or U3708 (N_3708,N_3302,N_3401);
xor U3709 (N_3709,N_3365,N_3391);
nor U3710 (N_3710,N_3429,N_3252);
nor U3711 (N_3711,N_3339,N_3266);
nand U3712 (N_3712,N_3493,N_3260);
or U3713 (N_3713,N_3329,N_3407);
xnor U3714 (N_3714,N_3280,N_3324);
nor U3715 (N_3715,N_3420,N_3458);
nor U3716 (N_3716,N_3388,N_3390);
nand U3717 (N_3717,N_3431,N_3402);
nor U3718 (N_3718,N_3372,N_3449);
and U3719 (N_3719,N_3254,N_3387);
or U3720 (N_3720,N_3415,N_3491);
xnor U3721 (N_3721,N_3358,N_3480);
and U3722 (N_3722,N_3274,N_3459);
nand U3723 (N_3723,N_3392,N_3444);
xor U3724 (N_3724,N_3412,N_3416);
and U3725 (N_3725,N_3480,N_3409);
or U3726 (N_3726,N_3254,N_3283);
xor U3727 (N_3727,N_3366,N_3403);
nand U3728 (N_3728,N_3430,N_3375);
nor U3729 (N_3729,N_3329,N_3365);
or U3730 (N_3730,N_3457,N_3310);
nand U3731 (N_3731,N_3300,N_3354);
or U3732 (N_3732,N_3355,N_3393);
xor U3733 (N_3733,N_3322,N_3395);
nand U3734 (N_3734,N_3414,N_3339);
xnor U3735 (N_3735,N_3299,N_3378);
and U3736 (N_3736,N_3286,N_3454);
nand U3737 (N_3737,N_3349,N_3270);
nor U3738 (N_3738,N_3378,N_3428);
nor U3739 (N_3739,N_3477,N_3372);
nand U3740 (N_3740,N_3379,N_3286);
nand U3741 (N_3741,N_3485,N_3392);
nand U3742 (N_3742,N_3324,N_3388);
nand U3743 (N_3743,N_3326,N_3446);
or U3744 (N_3744,N_3372,N_3279);
nand U3745 (N_3745,N_3388,N_3293);
nor U3746 (N_3746,N_3418,N_3362);
and U3747 (N_3747,N_3340,N_3350);
and U3748 (N_3748,N_3427,N_3452);
or U3749 (N_3749,N_3404,N_3372);
xor U3750 (N_3750,N_3684,N_3577);
nor U3751 (N_3751,N_3576,N_3745);
nor U3752 (N_3752,N_3572,N_3672);
nor U3753 (N_3753,N_3639,N_3696);
or U3754 (N_3754,N_3574,N_3625);
nor U3755 (N_3755,N_3523,N_3561);
nor U3756 (N_3756,N_3553,N_3533);
and U3757 (N_3757,N_3727,N_3676);
or U3758 (N_3758,N_3517,N_3512);
and U3759 (N_3759,N_3604,N_3504);
or U3760 (N_3760,N_3532,N_3522);
nand U3761 (N_3761,N_3706,N_3620);
nand U3762 (N_3762,N_3560,N_3644);
and U3763 (N_3763,N_3642,N_3693);
nand U3764 (N_3764,N_3503,N_3691);
and U3765 (N_3765,N_3559,N_3749);
nand U3766 (N_3766,N_3632,N_3526);
nand U3767 (N_3767,N_3660,N_3654);
xor U3768 (N_3768,N_3636,N_3571);
nor U3769 (N_3769,N_3717,N_3597);
and U3770 (N_3770,N_3613,N_3712);
and U3771 (N_3771,N_3700,N_3617);
or U3772 (N_3772,N_3501,N_3568);
xnor U3773 (N_3773,N_3547,N_3554);
nor U3774 (N_3774,N_3508,N_3590);
nor U3775 (N_3775,N_3668,N_3701);
nor U3776 (N_3776,N_3669,N_3630);
nor U3777 (N_3777,N_3623,N_3742);
and U3778 (N_3778,N_3528,N_3578);
nor U3779 (N_3779,N_3656,N_3529);
nand U3780 (N_3780,N_3605,N_3626);
nand U3781 (N_3781,N_3521,N_3628);
or U3782 (N_3782,N_3720,N_3531);
and U3783 (N_3783,N_3702,N_3705);
xor U3784 (N_3784,N_3733,N_3519);
nand U3785 (N_3785,N_3562,N_3510);
xnor U3786 (N_3786,N_3549,N_3723);
xnor U3787 (N_3787,N_3743,N_3552);
nor U3788 (N_3788,N_3688,N_3714);
or U3789 (N_3789,N_3697,N_3643);
nor U3790 (N_3790,N_3581,N_3619);
nor U3791 (N_3791,N_3537,N_3587);
or U3792 (N_3792,N_3724,N_3544);
or U3793 (N_3793,N_3566,N_3542);
or U3794 (N_3794,N_3685,N_3711);
nand U3795 (N_3795,N_3558,N_3748);
nor U3796 (N_3796,N_3563,N_3538);
xnor U3797 (N_3797,N_3735,N_3592);
nand U3798 (N_3798,N_3591,N_3659);
xor U3799 (N_3799,N_3500,N_3683);
xnor U3800 (N_3800,N_3629,N_3565);
and U3801 (N_3801,N_3595,N_3556);
nor U3802 (N_3802,N_3730,N_3695);
or U3803 (N_3803,N_3618,N_3699);
nand U3804 (N_3804,N_3737,N_3648);
or U3805 (N_3805,N_3707,N_3543);
or U3806 (N_3806,N_3739,N_3663);
nand U3807 (N_3807,N_3575,N_3652);
nor U3808 (N_3808,N_3677,N_3525);
or U3809 (N_3809,N_3678,N_3715);
or U3810 (N_3810,N_3722,N_3627);
and U3811 (N_3811,N_3589,N_3602);
or U3812 (N_3812,N_3747,N_3585);
nor U3813 (N_3813,N_3738,N_3657);
nand U3814 (N_3814,N_3507,N_3545);
and U3815 (N_3815,N_3539,N_3640);
nor U3816 (N_3816,N_3582,N_3726);
or U3817 (N_3817,N_3694,N_3687);
or U3818 (N_3818,N_3725,N_3598);
or U3819 (N_3819,N_3596,N_3665);
xor U3820 (N_3820,N_3650,N_3634);
or U3821 (N_3821,N_3670,N_3713);
xnor U3822 (N_3822,N_3615,N_3740);
and U3823 (N_3823,N_3600,N_3505);
xnor U3824 (N_3824,N_3732,N_3734);
or U3825 (N_3825,N_3710,N_3664);
nand U3826 (N_3826,N_3631,N_3611);
or U3827 (N_3827,N_3610,N_3731);
and U3828 (N_3828,N_3520,N_3599);
nor U3829 (N_3829,N_3513,N_3511);
xor U3830 (N_3830,N_3703,N_3593);
nand U3831 (N_3831,N_3638,N_3588);
nand U3832 (N_3832,N_3682,N_3616);
and U3833 (N_3833,N_3709,N_3681);
or U3834 (N_3834,N_3579,N_3584);
nor U3835 (N_3835,N_3679,N_3603);
or U3836 (N_3836,N_3535,N_3515);
nor U3837 (N_3837,N_3608,N_3716);
nand U3838 (N_3838,N_3675,N_3708);
nand U3839 (N_3839,N_3534,N_3612);
and U3840 (N_3840,N_3651,N_3661);
or U3841 (N_3841,N_3633,N_3540);
nand U3842 (N_3842,N_3728,N_3671);
xnor U3843 (N_3843,N_3557,N_3530);
nand U3844 (N_3844,N_3516,N_3541);
and U3845 (N_3845,N_3551,N_3689);
or U3846 (N_3846,N_3570,N_3686);
or U3847 (N_3847,N_3614,N_3621);
or U3848 (N_3848,N_3666,N_3729);
nor U3849 (N_3849,N_3673,N_3680);
nand U3850 (N_3850,N_3536,N_3506);
nor U3851 (N_3851,N_3721,N_3692);
xnor U3852 (N_3852,N_3548,N_3647);
nand U3853 (N_3853,N_3655,N_3524);
xor U3854 (N_3854,N_3601,N_3569);
nand U3855 (N_3855,N_3502,N_3609);
xor U3856 (N_3856,N_3704,N_3649);
and U3857 (N_3857,N_3518,N_3624);
xnor U3858 (N_3858,N_3509,N_3637);
or U3859 (N_3859,N_3607,N_3736);
nand U3860 (N_3860,N_3573,N_3690);
xor U3861 (N_3861,N_3674,N_3514);
nand U3862 (N_3862,N_3698,N_3646);
xnor U3863 (N_3863,N_3555,N_3550);
or U3864 (N_3864,N_3658,N_3719);
xnor U3865 (N_3865,N_3586,N_3641);
nor U3866 (N_3866,N_3746,N_3662);
xnor U3867 (N_3867,N_3594,N_3667);
nand U3868 (N_3868,N_3580,N_3653);
nand U3869 (N_3869,N_3564,N_3741);
xor U3870 (N_3870,N_3744,N_3645);
nor U3871 (N_3871,N_3567,N_3527);
nor U3872 (N_3872,N_3546,N_3718);
or U3873 (N_3873,N_3583,N_3622);
nand U3874 (N_3874,N_3606,N_3635);
and U3875 (N_3875,N_3531,N_3520);
nand U3876 (N_3876,N_3539,N_3625);
and U3877 (N_3877,N_3721,N_3691);
or U3878 (N_3878,N_3651,N_3531);
xor U3879 (N_3879,N_3656,N_3520);
or U3880 (N_3880,N_3725,N_3602);
nand U3881 (N_3881,N_3583,N_3620);
or U3882 (N_3882,N_3654,N_3504);
nand U3883 (N_3883,N_3640,N_3692);
and U3884 (N_3884,N_3636,N_3589);
or U3885 (N_3885,N_3592,N_3544);
xor U3886 (N_3886,N_3623,N_3503);
xor U3887 (N_3887,N_3544,N_3531);
and U3888 (N_3888,N_3702,N_3607);
and U3889 (N_3889,N_3702,N_3658);
or U3890 (N_3890,N_3656,N_3734);
and U3891 (N_3891,N_3575,N_3749);
nor U3892 (N_3892,N_3677,N_3662);
nor U3893 (N_3893,N_3595,N_3588);
and U3894 (N_3894,N_3597,N_3609);
or U3895 (N_3895,N_3541,N_3605);
nand U3896 (N_3896,N_3702,N_3578);
nor U3897 (N_3897,N_3536,N_3609);
nor U3898 (N_3898,N_3522,N_3540);
or U3899 (N_3899,N_3688,N_3650);
nand U3900 (N_3900,N_3655,N_3514);
xor U3901 (N_3901,N_3523,N_3581);
or U3902 (N_3902,N_3562,N_3631);
and U3903 (N_3903,N_3658,N_3572);
or U3904 (N_3904,N_3626,N_3689);
xor U3905 (N_3905,N_3511,N_3706);
xor U3906 (N_3906,N_3743,N_3685);
or U3907 (N_3907,N_3564,N_3649);
or U3908 (N_3908,N_3739,N_3748);
nor U3909 (N_3909,N_3656,N_3560);
nor U3910 (N_3910,N_3643,N_3727);
nand U3911 (N_3911,N_3529,N_3523);
or U3912 (N_3912,N_3507,N_3656);
or U3913 (N_3913,N_3624,N_3718);
nor U3914 (N_3914,N_3697,N_3638);
and U3915 (N_3915,N_3711,N_3514);
nand U3916 (N_3916,N_3579,N_3537);
or U3917 (N_3917,N_3562,N_3577);
and U3918 (N_3918,N_3647,N_3543);
nor U3919 (N_3919,N_3594,N_3580);
xor U3920 (N_3920,N_3690,N_3695);
nor U3921 (N_3921,N_3686,N_3636);
xor U3922 (N_3922,N_3590,N_3545);
nor U3923 (N_3923,N_3624,N_3572);
nand U3924 (N_3924,N_3657,N_3512);
nor U3925 (N_3925,N_3705,N_3579);
or U3926 (N_3926,N_3576,N_3601);
xnor U3927 (N_3927,N_3625,N_3726);
or U3928 (N_3928,N_3626,N_3660);
xnor U3929 (N_3929,N_3582,N_3501);
or U3930 (N_3930,N_3738,N_3575);
nor U3931 (N_3931,N_3581,N_3622);
or U3932 (N_3932,N_3728,N_3610);
nand U3933 (N_3933,N_3514,N_3717);
or U3934 (N_3934,N_3711,N_3568);
and U3935 (N_3935,N_3627,N_3619);
xnor U3936 (N_3936,N_3700,N_3549);
and U3937 (N_3937,N_3720,N_3631);
nand U3938 (N_3938,N_3521,N_3602);
and U3939 (N_3939,N_3745,N_3662);
nor U3940 (N_3940,N_3649,N_3696);
nand U3941 (N_3941,N_3609,N_3591);
nand U3942 (N_3942,N_3618,N_3684);
and U3943 (N_3943,N_3619,N_3602);
nand U3944 (N_3944,N_3530,N_3615);
xnor U3945 (N_3945,N_3663,N_3601);
xor U3946 (N_3946,N_3666,N_3676);
and U3947 (N_3947,N_3588,N_3671);
nor U3948 (N_3948,N_3545,N_3617);
and U3949 (N_3949,N_3691,N_3554);
nor U3950 (N_3950,N_3720,N_3615);
nor U3951 (N_3951,N_3607,N_3628);
and U3952 (N_3952,N_3592,N_3655);
nand U3953 (N_3953,N_3559,N_3543);
nand U3954 (N_3954,N_3637,N_3727);
and U3955 (N_3955,N_3523,N_3637);
xnor U3956 (N_3956,N_3661,N_3518);
or U3957 (N_3957,N_3627,N_3683);
nand U3958 (N_3958,N_3648,N_3634);
or U3959 (N_3959,N_3609,N_3704);
or U3960 (N_3960,N_3708,N_3508);
or U3961 (N_3961,N_3605,N_3564);
or U3962 (N_3962,N_3667,N_3530);
and U3963 (N_3963,N_3597,N_3628);
xnor U3964 (N_3964,N_3697,N_3715);
and U3965 (N_3965,N_3703,N_3640);
nand U3966 (N_3966,N_3688,N_3586);
and U3967 (N_3967,N_3573,N_3649);
nand U3968 (N_3968,N_3644,N_3630);
or U3969 (N_3969,N_3645,N_3589);
and U3970 (N_3970,N_3598,N_3741);
or U3971 (N_3971,N_3718,N_3674);
or U3972 (N_3972,N_3523,N_3693);
nand U3973 (N_3973,N_3548,N_3542);
nor U3974 (N_3974,N_3568,N_3506);
nor U3975 (N_3975,N_3537,N_3730);
and U3976 (N_3976,N_3655,N_3574);
xor U3977 (N_3977,N_3717,N_3550);
nand U3978 (N_3978,N_3592,N_3692);
nor U3979 (N_3979,N_3607,N_3570);
or U3980 (N_3980,N_3593,N_3611);
and U3981 (N_3981,N_3637,N_3648);
nor U3982 (N_3982,N_3695,N_3747);
xor U3983 (N_3983,N_3577,N_3739);
or U3984 (N_3984,N_3551,N_3710);
nor U3985 (N_3985,N_3648,N_3589);
nor U3986 (N_3986,N_3713,N_3656);
xnor U3987 (N_3987,N_3601,N_3635);
nand U3988 (N_3988,N_3727,N_3558);
xnor U3989 (N_3989,N_3503,N_3531);
and U3990 (N_3990,N_3588,N_3723);
xnor U3991 (N_3991,N_3582,N_3525);
or U3992 (N_3992,N_3564,N_3532);
or U3993 (N_3993,N_3631,N_3525);
or U3994 (N_3994,N_3613,N_3664);
nand U3995 (N_3995,N_3515,N_3509);
xnor U3996 (N_3996,N_3580,N_3572);
nand U3997 (N_3997,N_3681,N_3734);
or U3998 (N_3998,N_3684,N_3578);
xor U3999 (N_3999,N_3550,N_3662);
and U4000 (N_4000,N_3901,N_3805);
nor U4001 (N_4001,N_3883,N_3772);
nand U4002 (N_4002,N_3868,N_3759);
nor U4003 (N_4003,N_3869,N_3779);
or U4004 (N_4004,N_3842,N_3782);
xor U4005 (N_4005,N_3963,N_3914);
or U4006 (N_4006,N_3845,N_3961);
and U4007 (N_4007,N_3995,N_3938);
nand U4008 (N_4008,N_3986,N_3804);
nor U4009 (N_4009,N_3895,N_3802);
xnor U4010 (N_4010,N_3829,N_3957);
nor U4011 (N_4011,N_3789,N_3989);
and U4012 (N_4012,N_3816,N_3786);
nand U4013 (N_4013,N_3858,N_3857);
nor U4014 (N_4014,N_3890,N_3960);
nor U4015 (N_4015,N_3867,N_3970);
nor U4016 (N_4016,N_3921,N_3937);
nor U4017 (N_4017,N_3771,N_3962);
or U4018 (N_4018,N_3971,N_3828);
or U4019 (N_4019,N_3835,N_3811);
and U4020 (N_4020,N_3856,N_3777);
nand U4021 (N_4021,N_3863,N_3958);
nand U4022 (N_4022,N_3841,N_3955);
xor U4023 (N_4023,N_3840,N_3791);
xor U4024 (N_4024,N_3815,N_3767);
nor U4025 (N_4025,N_3966,N_3753);
xor U4026 (N_4026,N_3803,N_3915);
xor U4027 (N_4027,N_3899,N_3874);
xor U4028 (N_4028,N_3846,N_3806);
nor U4029 (N_4029,N_3801,N_3999);
or U4030 (N_4030,N_3773,N_3973);
nor U4031 (N_4031,N_3768,N_3774);
xnor U4032 (N_4032,N_3953,N_3876);
xnor U4033 (N_4033,N_3821,N_3935);
nor U4034 (N_4034,N_3956,N_3794);
nor U4035 (N_4035,N_3847,N_3944);
xor U4036 (N_4036,N_3933,N_3952);
nand U4037 (N_4037,N_3752,N_3861);
or U4038 (N_4038,N_3780,N_3964);
nand U4039 (N_4039,N_3950,N_3954);
nand U4040 (N_4040,N_3755,N_3934);
xnor U4041 (N_4041,N_3884,N_3968);
or U4042 (N_4042,N_3996,N_3864);
nor U4043 (N_4043,N_3945,N_3891);
and U4044 (N_4044,N_3751,N_3987);
xnor U4045 (N_4045,N_3893,N_3758);
xor U4046 (N_4046,N_3946,N_3792);
and U4047 (N_4047,N_3939,N_3998);
nor U4048 (N_4048,N_3756,N_3888);
or U4049 (N_4049,N_3808,N_3942);
xnor U4050 (N_4050,N_3880,N_3783);
nand U4051 (N_4051,N_3831,N_3854);
xor U4052 (N_4052,N_3839,N_3807);
nor U4053 (N_4053,N_3983,N_3906);
nand U4054 (N_4054,N_3793,N_3787);
nor U4055 (N_4055,N_3838,N_3907);
xor U4056 (N_4056,N_3882,N_3905);
nor U4057 (N_4057,N_3902,N_3760);
or U4058 (N_4058,N_3993,N_3927);
or U4059 (N_4059,N_3965,N_3928);
nor U4060 (N_4060,N_3809,N_3775);
xnor U4061 (N_4061,N_3959,N_3866);
and U4062 (N_4062,N_3823,N_3862);
and U4063 (N_4063,N_3929,N_3900);
nand U4064 (N_4064,N_3799,N_3834);
and U4065 (N_4065,N_3810,N_3980);
and U4066 (N_4066,N_3877,N_3819);
xor U4067 (N_4067,N_3837,N_3788);
nand U4068 (N_4068,N_3879,N_3979);
or U4069 (N_4069,N_3912,N_3885);
and U4070 (N_4070,N_3776,N_3833);
xnor U4071 (N_4071,N_3827,N_3865);
and U4072 (N_4072,N_3814,N_3764);
nor U4073 (N_4073,N_3800,N_3784);
xor U4074 (N_4074,N_3992,N_3818);
xor U4075 (N_4075,N_3785,N_3894);
xor U4076 (N_4076,N_3919,N_3978);
nor U4077 (N_4077,N_3836,N_3860);
or U4078 (N_4078,N_3763,N_3930);
or U4079 (N_4079,N_3947,N_3896);
nor U4080 (N_4080,N_3982,N_3812);
nor U4081 (N_4081,N_3898,N_3813);
or U4082 (N_4082,N_3825,N_3972);
and U4083 (N_4083,N_3940,N_3798);
xnor U4084 (N_4084,N_3832,N_3850);
nor U4085 (N_4085,N_3994,N_3769);
nor U4086 (N_4086,N_3871,N_3889);
xnor U4087 (N_4087,N_3988,N_3909);
xor U4088 (N_4088,N_3881,N_3976);
xnor U4089 (N_4089,N_3826,N_3931);
or U4090 (N_4090,N_3797,N_3852);
or U4091 (N_4091,N_3897,N_3848);
xnor U4092 (N_4092,N_3873,N_3911);
nor U4093 (N_4093,N_3754,N_3853);
or U4094 (N_4094,N_3922,N_3761);
xor U4095 (N_4095,N_3851,N_3918);
nand U4096 (N_4096,N_3849,N_3981);
nand U4097 (N_4097,N_3843,N_3875);
nor U4098 (N_4098,N_3925,N_3997);
nor U4099 (N_4099,N_3917,N_3926);
nand U4100 (N_4100,N_3948,N_3778);
or U4101 (N_4101,N_3872,N_3913);
and U4102 (N_4102,N_3974,N_3781);
and U4103 (N_4103,N_3943,N_3967);
nor U4104 (N_4104,N_3924,N_3766);
nor U4105 (N_4105,N_3762,N_3844);
or U4106 (N_4106,N_3790,N_3969);
nor U4107 (N_4107,N_3975,N_3822);
or U4108 (N_4108,N_3870,N_3796);
nor U4109 (N_4109,N_3932,N_3951);
xnor U4110 (N_4110,N_3991,N_3878);
xor U4111 (N_4111,N_3830,N_3920);
nor U4112 (N_4112,N_3916,N_3908);
xor U4113 (N_4113,N_3903,N_3817);
nor U4114 (N_4114,N_3990,N_3770);
and U4115 (N_4115,N_3765,N_3949);
or U4116 (N_4116,N_3910,N_3886);
nand U4117 (N_4117,N_3887,N_3904);
and U4118 (N_4118,N_3936,N_3923);
or U4119 (N_4119,N_3977,N_3941);
or U4120 (N_4120,N_3985,N_3859);
nor U4121 (N_4121,N_3750,N_3824);
xnor U4122 (N_4122,N_3820,N_3795);
nand U4123 (N_4123,N_3892,N_3984);
nor U4124 (N_4124,N_3855,N_3757);
or U4125 (N_4125,N_3857,N_3922);
xor U4126 (N_4126,N_3953,N_3893);
nand U4127 (N_4127,N_3752,N_3822);
xnor U4128 (N_4128,N_3919,N_3962);
and U4129 (N_4129,N_3843,N_3901);
nand U4130 (N_4130,N_3914,N_3837);
xnor U4131 (N_4131,N_3984,N_3880);
nand U4132 (N_4132,N_3817,N_3803);
or U4133 (N_4133,N_3802,N_3847);
or U4134 (N_4134,N_3808,N_3809);
nor U4135 (N_4135,N_3957,N_3870);
and U4136 (N_4136,N_3838,N_3996);
nand U4137 (N_4137,N_3772,N_3830);
nand U4138 (N_4138,N_3891,N_3779);
nand U4139 (N_4139,N_3934,N_3977);
nor U4140 (N_4140,N_3827,N_3786);
or U4141 (N_4141,N_3949,N_3900);
xor U4142 (N_4142,N_3917,N_3763);
nor U4143 (N_4143,N_3972,N_3981);
or U4144 (N_4144,N_3768,N_3869);
or U4145 (N_4145,N_3924,N_3975);
or U4146 (N_4146,N_3982,N_3797);
xnor U4147 (N_4147,N_3865,N_3812);
and U4148 (N_4148,N_3910,N_3926);
or U4149 (N_4149,N_3844,N_3831);
nor U4150 (N_4150,N_3771,N_3795);
nand U4151 (N_4151,N_3974,N_3920);
nand U4152 (N_4152,N_3936,N_3776);
nor U4153 (N_4153,N_3945,N_3812);
or U4154 (N_4154,N_3759,N_3839);
nand U4155 (N_4155,N_3838,N_3937);
xor U4156 (N_4156,N_3953,N_3909);
xnor U4157 (N_4157,N_3790,N_3861);
nand U4158 (N_4158,N_3921,N_3903);
xor U4159 (N_4159,N_3828,N_3946);
or U4160 (N_4160,N_3857,N_3923);
xnor U4161 (N_4161,N_3883,N_3848);
or U4162 (N_4162,N_3982,N_3750);
nand U4163 (N_4163,N_3976,N_3873);
nand U4164 (N_4164,N_3840,N_3861);
xor U4165 (N_4165,N_3896,N_3763);
or U4166 (N_4166,N_3796,N_3897);
and U4167 (N_4167,N_3810,N_3865);
and U4168 (N_4168,N_3958,N_3966);
and U4169 (N_4169,N_3928,N_3838);
xnor U4170 (N_4170,N_3974,N_3937);
nor U4171 (N_4171,N_3869,N_3837);
nand U4172 (N_4172,N_3800,N_3780);
or U4173 (N_4173,N_3884,N_3847);
nand U4174 (N_4174,N_3869,N_3986);
nand U4175 (N_4175,N_3974,N_3847);
and U4176 (N_4176,N_3950,N_3828);
nand U4177 (N_4177,N_3915,N_3907);
or U4178 (N_4178,N_3803,N_3906);
or U4179 (N_4179,N_3965,N_3820);
and U4180 (N_4180,N_3848,N_3782);
xor U4181 (N_4181,N_3823,N_3951);
xnor U4182 (N_4182,N_3956,N_3872);
and U4183 (N_4183,N_3869,N_3780);
xor U4184 (N_4184,N_3920,N_3794);
and U4185 (N_4185,N_3928,N_3822);
nor U4186 (N_4186,N_3841,N_3885);
nand U4187 (N_4187,N_3992,N_3820);
and U4188 (N_4188,N_3823,N_3884);
nor U4189 (N_4189,N_3842,N_3902);
and U4190 (N_4190,N_3965,N_3956);
nor U4191 (N_4191,N_3950,N_3805);
nor U4192 (N_4192,N_3876,N_3769);
nand U4193 (N_4193,N_3907,N_3758);
nand U4194 (N_4194,N_3842,N_3767);
nor U4195 (N_4195,N_3928,N_3879);
xor U4196 (N_4196,N_3877,N_3902);
or U4197 (N_4197,N_3924,N_3961);
and U4198 (N_4198,N_3911,N_3999);
nor U4199 (N_4199,N_3863,N_3939);
nor U4200 (N_4200,N_3991,N_3844);
and U4201 (N_4201,N_3971,N_3910);
and U4202 (N_4202,N_3907,N_3914);
xnor U4203 (N_4203,N_3851,N_3839);
nor U4204 (N_4204,N_3814,N_3875);
nand U4205 (N_4205,N_3818,N_3814);
and U4206 (N_4206,N_3841,N_3994);
xor U4207 (N_4207,N_3823,N_3847);
nor U4208 (N_4208,N_3792,N_3822);
nand U4209 (N_4209,N_3850,N_3964);
or U4210 (N_4210,N_3835,N_3776);
xnor U4211 (N_4211,N_3849,N_3856);
or U4212 (N_4212,N_3821,N_3787);
and U4213 (N_4213,N_3866,N_3790);
nor U4214 (N_4214,N_3929,N_3955);
xor U4215 (N_4215,N_3853,N_3963);
xor U4216 (N_4216,N_3960,N_3834);
nor U4217 (N_4217,N_3992,N_3856);
or U4218 (N_4218,N_3994,N_3961);
xor U4219 (N_4219,N_3813,N_3809);
xor U4220 (N_4220,N_3849,N_3752);
nand U4221 (N_4221,N_3880,N_3893);
nor U4222 (N_4222,N_3882,N_3914);
and U4223 (N_4223,N_3885,N_3803);
nor U4224 (N_4224,N_3975,N_3957);
or U4225 (N_4225,N_3906,N_3915);
nor U4226 (N_4226,N_3965,N_3764);
xor U4227 (N_4227,N_3983,N_3944);
and U4228 (N_4228,N_3984,N_3936);
xor U4229 (N_4229,N_3984,N_3985);
nor U4230 (N_4230,N_3820,N_3972);
and U4231 (N_4231,N_3943,N_3849);
or U4232 (N_4232,N_3786,N_3888);
and U4233 (N_4233,N_3801,N_3905);
and U4234 (N_4234,N_3880,N_3803);
and U4235 (N_4235,N_3823,N_3927);
nor U4236 (N_4236,N_3838,N_3914);
or U4237 (N_4237,N_3915,N_3867);
or U4238 (N_4238,N_3998,N_3797);
and U4239 (N_4239,N_3899,N_3807);
or U4240 (N_4240,N_3924,N_3815);
nand U4241 (N_4241,N_3923,N_3762);
or U4242 (N_4242,N_3975,N_3916);
or U4243 (N_4243,N_3853,N_3857);
xnor U4244 (N_4244,N_3944,N_3776);
nand U4245 (N_4245,N_3753,N_3948);
or U4246 (N_4246,N_3816,N_3793);
xor U4247 (N_4247,N_3773,N_3852);
nor U4248 (N_4248,N_3965,N_3970);
nand U4249 (N_4249,N_3937,N_3934);
nand U4250 (N_4250,N_4113,N_4100);
or U4251 (N_4251,N_4073,N_4199);
nand U4252 (N_4252,N_4215,N_4224);
nand U4253 (N_4253,N_4020,N_4122);
xnor U4254 (N_4254,N_4174,N_4200);
and U4255 (N_4255,N_4127,N_4006);
nor U4256 (N_4256,N_4105,N_4208);
and U4257 (N_4257,N_4197,N_4172);
nand U4258 (N_4258,N_4019,N_4139);
xnor U4259 (N_4259,N_4158,N_4219);
nand U4260 (N_4260,N_4184,N_4231);
or U4261 (N_4261,N_4063,N_4159);
or U4262 (N_4262,N_4069,N_4039);
or U4263 (N_4263,N_4126,N_4007);
or U4264 (N_4264,N_4054,N_4015);
nor U4265 (N_4265,N_4226,N_4177);
nor U4266 (N_4266,N_4048,N_4025);
xor U4267 (N_4267,N_4027,N_4090);
and U4268 (N_4268,N_4143,N_4094);
nor U4269 (N_4269,N_4202,N_4028);
nand U4270 (N_4270,N_4001,N_4145);
nor U4271 (N_4271,N_4084,N_4044);
and U4272 (N_4272,N_4056,N_4120);
or U4273 (N_4273,N_4166,N_4012);
or U4274 (N_4274,N_4067,N_4107);
nand U4275 (N_4275,N_4157,N_4024);
nand U4276 (N_4276,N_4142,N_4065);
or U4277 (N_4277,N_4121,N_4013);
nand U4278 (N_4278,N_4130,N_4002);
nor U4279 (N_4279,N_4136,N_4232);
and U4280 (N_4280,N_4017,N_4185);
nor U4281 (N_4281,N_4086,N_4077);
and U4282 (N_4282,N_4099,N_4004);
or U4283 (N_4283,N_4156,N_4070);
and U4284 (N_4284,N_4179,N_4026);
nor U4285 (N_4285,N_4188,N_4233);
and U4286 (N_4286,N_4243,N_4194);
and U4287 (N_4287,N_4021,N_4047);
xor U4288 (N_4288,N_4018,N_4191);
nand U4289 (N_4289,N_4060,N_4124);
or U4290 (N_4290,N_4080,N_4128);
nor U4291 (N_4291,N_4169,N_4132);
or U4292 (N_4292,N_4138,N_4062);
nor U4293 (N_4293,N_4178,N_4153);
and U4294 (N_4294,N_4175,N_4152);
nand U4295 (N_4295,N_4170,N_4083);
nor U4296 (N_4296,N_4050,N_4049);
xor U4297 (N_4297,N_4244,N_4163);
nor U4298 (N_4298,N_4237,N_4076);
nand U4299 (N_4299,N_4149,N_4196);
nor U4300 (N_4300,N_4053,N_4003);
or U4301 (N_4301,N_4097,N_4221);
and U4302 (N_4302,N_4245,N_4195);
or U4303 (N_4303,N_4119,N_4095);
nor U4304 (N_4304,N_4239,N_4072);
xnor U4305 (N_4305,N_4168,N_4096);
and U4306 (N_4306,N_4059,N_4223);
and U4307 (N_4307,N_4043,N_4147);
and U4308 (N_4308,N_4182,N_4135);
nand U4309 (N_4309,N_4000,N_4148);
nand U4310 (N_4310,N_4220,N_4078);
xor U4311 (N_4311,N_4218,N_4209);
xor U4312 (N_4312,N_4206,N_4085);
or U4313 (N_4313,N_4108,N_4129);
nor U4314 (N_4314,N_4066,N_4204);
xnor U4315 (N_4315,N_4045,N_4167);
and U4316 (N_4316,N_4171,N_4133);
nand U4317 (N_4317,N_4187,N_4023);
nor U4318 (N_4318,N_4037,N_4150);
or U4319 (N_4319,N_4104,N_4229);
nand U4320 (N_4320,N_4248,N_4110);
nor U4321 (N_4321,N_4212,N_4058);
nor U4322 (N_4322,N_4033,N_4011);
nand U4323 (N_4323,N_4201,N_4040);
xor U4324 (N_4324,N_4140,N_4141);
nor U4325 (N_4325,N_4118,N_4041);
xnor U4326 (N_4326,N_4249,N_4176);
xor U4327 (N_4327,N_4186,N_4181);
or U4328 (N_4328,N_4225,N_4217);
xnor U4329 (N_4329,N_4082,N_4234);
and U4330 (N_4330,N_4115,N_4088);
nor U4331 (N_4331,N_4109,N_4101);
nand U4332 (N_4332,N_4098,N_4055);
xnor U4333 (N_4333,N_4022,N_4183);
nor U4334 (N_4334,N_4164,N_4134);
xnor U4335 (N_4335,N_4203,N_4222);
nor U4336 (N_4336,N_4093,N_4240);
xor U4337 (N_4337,N_4162,N_4144);
nor U4338 (N_4338,N_4035,N_4236);
nor U4339 (N_4339,N_4112,N_4125);
xor U4340 (N_4340,N_4198,N_4235);
and U4341 (N_4341,N_4061,N_4160);
nor U4342 (N_4342,N_4030,N_4106);
nand U4343 (N_4343,N_4068,N_4246);
xnor U4344 (N_4344,N_4036,N_4051);
xor U4345 (N_4345,N_4111,N_4089);
or U4346 (N_4346,N_4009,N_4034);
nor U4347 (N_4347,N_4008,N_4190);
nor U4348 (N_4348,N_4081,N_4213);
and U4349 (N_4349,N_4247,N_4074);
xnor U4350 (N_4350,N_4114,N_4146);
nand U4351 (N_4351,N_4238,N_4038);
xor U4352 (N_4352,N_4216,N_4207);
nor U4353 (N_4353,N_4042,N_4155);
nor U4354 (N_4354,N_4071,N_4210);
xor U4355 (N_4355,N_4241,N_4046);
nor U4356 (N_4356,N_4161,N_4154);
nor U4357 (N_4357,N_4193,N_4151);
xor U4358 (N_4358,N_4228,N_4005);
nand U4359 (N_4359,N_4092,N_4173);
and U4360 (N_4360,N_4064,N_4103);
xor U4361 (N_4361,N_4165,N_4057);
or U4362 (N_4362,N_4117,N_4010);
and U4363 (N_4363,N_4227,N_4032);
and U4364 (N_4364,N_4211,N_4087);
and U4365 (N_4365,N_4091,N_4116);
or U4366 (N_4366,N_4029,N_4131);
and U4367 (N_4367,N_4052,N_4205);
xnor U4368 (N_4368,N_4102,N_4230);
xor U4369 (N_4369,N_4192,N_4014);
xnor U4370 (N_4370,N_4180,N_4214);
nand U4371 (N_4371,N_4075,N_4031);
xnor U4372 (N_4372,N_4079,N_4016);
and U4373 (N_4373,N_4137,N_4123);
and U4374 (N_4374,N_4242,N_4189);
xnor U4375 (N_4375,N_4245,N_4209);
nor U4376 (N_4376,N_4188,N_4224);
and U4377 (N_4377,N_4168,N_4091);
xor U4378 (N_4378,N_4056,N_4077);
xor U4379 (N_4379,N_4055,N_4066);
nand U4380 (N_4380,N_4214,N_4098);
nor U4381 (N_4381,N_4249,N_4189);
nor U4382 (N_4382,N_4071,N_4012);
nor U4383 (N_4383,N_4099,N_4173);
or U4384 (N_4384,N_4015,N_4007);
nor U4385 (N_4385,N_4183,N_4210);
and U4386 (N_4386,N_4221,N_4016);
xor U4387 (N_4387,N_4122,N_4101);
nand U4388 (N_4388,N_4038,N_4151);
or U4389 (N_4389,N_4245,N_4088);
nand U4390 (N_4390,N_4072,N_4147);
nand U4391 (N_4391,N_4075,N_4188);
or U4392 (N_4392,N_4237,N_4232);
nor U4393 (N_4393,N_4187,N_4062);
or U4394 (N_4394,N_4047,N_4133);
or U4395 (N_4395,N_4076,N_4133);
nor U4396 (N_4396,N_4044,N_4175);
nand U4397 (N_4397,N_4142,N_4166);
xor U4398 (N_4398,N_4242,N_4062);
nor U4399 (N_4399,N_4219,N_4169);
nand U4400 (N_4400,N_4167,N_4148);
nor U4401 (N_4401,N_4166,N_4043);
xor U4402 (N_4402,N_4066,N_4031);
xor U4403 (N_4403,N_4203,N_4094);
nand U4404 (N_4404,N_4203,N_4227);
or U4405 (N_4405,N_4130,N_4091);
nor U4406 (N_4406,N_4133,N_4088);
nand U4407 (N_4407,N_4184,N_4020);
or U4408 (N_4408,N_4152,N_4180);
and U4409 (N_4409,N_4064,N_4087);
nor U4410 (N_4410,N_4105,N_4042);
xnor U4411 (N_4411,N_4247,N_4146);
nor U4412 (N_4412,N_4216,N_4225);
nand U4413 (N_4413,N_4029,N_4092);
xor U4414 (N_4414,N_4228,N_4045);
nor U4415 (N_4415,N_4010,N_4169);
and U4416 (N_4416,N_4221,N_4111);
and U4417 (N_4417,N_4022,N_4141);
and U4418 (N_4418,N_4013,N_4090);
or U4419 (N_4419,N_4211,N_4011);
nor U4420 (N_4420,N_4199,N_4188);
nor U4421 (N_4421,N_4195,N_4015);
xor U4422 (N_4422,N_4031,N_4182);
or U4423 (N_4423,N_4163,N_4240);
or U4424 (N_4424,N_4233,N_4227);
or U4425 (N_4425,N_4189,N_4201);
and U4426 (N_4426,N_4110,N_4207);
nor U4427 (N_4427,N_4002,N_4140);
or U4428 (N_4428,N_4098,N_4229);
and U4429 (N_4429,N_4167,N_4132);
nor U4430 (N_4430,N_4220,N_4203);
or U4431 (N_4431,N_4059,N_4037);
or U4432 (N_4432,N_4247,N_4135);
or U4433 (N_4433,N_4046,N_4168);
and U4434 (N_4434,N_4092,N_4147);
nand U4435 (N_4435,N_4110,N_4054);
and U4436 (N_4436,N_4070,N_4061);
and U4437 (N_4437,N_4044,N_4005);
or U4438 (N_4438,N_4083,N_4055);
xnor U4439 (N_4439,N_4246,N_4170);
nor U4440 (N_4440,N_4198,N_4242);
or U4441 (N_4441,N_4108,N_4145);
xnor U4442 (N_4442,N_4246,N_4051);
xnor U4443 (N_4443,N_4025,N_4002);
nand U4444 (N_4444,N_4164,N_4102);
nor U4445 (N_4445,N_4024,N_4091);
or U4446 (N_4446,N_4180,N_4205);
nand U4447 (N_4447,N_4145,N_4187);
and U4448 (N_4448,N_4172,N_4155);
xnor U4449 (N_4449,N_4119,N_4010);
nand U4450 (N_4450,N_4133,N_4115);
nand U4451 (N_4451,N_4061,N_4013);
xor U4452 (N_4452,N_4110,N_4242);
nand U4453 (N_4453,N_4084,N_4247);
and U4454 (N_4454,N_4111,N_4237);
xor U4455 (N_4455,N_4045,N_4126);
nor U4456 (N_4456,N_4180,N_4139);
xnor U4457 (N_4457,N_4093,N_4053);
and U4458 (N_4458,N_4153,N_4111);
nand U4459 (N_4459,N_4130,N_4078);
nand U4460 (N_4460,N_4159,N_4049);
nand U4461 (N_4461,N_4026,N_4063);
xor U4462 (N_4462,N_4219,N_4198);
and U4463 (N_4463,N_4089,N_4102);
nor U4464 (N_4464,N_4116,N_4183);
xnor U4465 (N_4465,N_4043,N_4003);
or U4466 (N_4466,N_4124,N_4096);
or U4467 (N_4467,N_4210,N_4184);
xnor U4468 (N_4468,N_4006,N_4106);
nand U4469 (N_4469,N_4117,N_4166);
nand U4470 (N_4470,N_4143,N_4034);
or U4471 (N_4471,N_4160,N_4027);
nor U4472 (N_4472,N_4015,N_4114);
nor U4473 (N_4473,N_4108,N_4163);
or U4474 (N_4474,N_4224,N_4022);
or U4475 (N_4475,N_4207,N_4146);
and U4476 (N_4476,N_4029,N_4208);
nor U4477 (N_4477,N_4035,N_4209);
xnor U4478 (N_4478,N_4169,N_4194);
or U4479 (N_4479,N_4037,N_4241);
and U4480 (N_4480,N_4129,N_4234);
nor U4481 (N_4481,N_4012,N_4084);
xor U4482 (N_4482,N_4227,N_4223);
xnor U4483 (N_4483,N_4125,N_4167);
xor U4484 (N_4484,N_4247,N_4220);
or U4485 (N_4485,N_4148,N_4100);
and U4486 (N_4486,N_4212,N_4200);
nand U4487 (N_4487,N_4060,N_4183);
xor U4488 (N_4488,N_4090,N_4151);
xor U4489 (N_4489,N_4190,N_4131);
nand U4490 (N_4490,N_4145,N_4045);
and U4491 (N_4491,N_4108,N_4088);
nor U4492 (N_4492,N_4026,N_4119);
nand U4493 (N_4493,N_4105,N_4093);
nor U4494 (N_4494,N_4076,N_4115);
nor U4495 (N_4495,N_4146,N_4068);
and U4496 (N_4496,N_4177,N_4095);
or U4497 (N_4497,N_4039,N_4006);
nand U4498 (N_4498,N_4244,N_4122);
or U4499 (N_4499,N_4006,N_4032);
and U4500 (N_4500,N_4479,N_4474);
nor U4501 (N_4501,N_4369,N_4342);
or U4502 (N_4502,N_4300,N_4291);
or U4503 (N_4503,N_4256,N_4282);
nor U4504 (N_4504,N_4321,N_4433);
nor U4505 (N_4505,N_4453,N_4435);
nor U4506 (N_4506,N_4272,N_4396);
and U4507 (N_4507,N_4380,N_4460);
or U4508 (N_4508,N_4417,N_4304);
xnor U4509 (N_4509,N_4441,N_4326);
and U4510 (N_4510,N_4305,N_4400);
xnor U4511 (N_4511,N_4466,N_4381);
nand U4512 (N_4512,N_4260,N_4325);
or U4513 (N_4513,N_4347,N_4356);
nand U4514 (N_4514,N_4399,N_4492);
nor U4515 (N_4515,N_4440,N_4259);
nand U4516 (N_4516,N_4350,N_4254);
xnor U4517 (N_4517,N_4491,N_4255);
and U4518 (N_4518,N_4274,N_4404);
or U4519 (N_4519,N_4276,N_4478);
and U4520 (N_4520,N_4408,N_4384);
or U4521 (N_4521,N_4368,N_4425);
and U4522 (N_4522,N_4318,N_4377);
nor U4523 (N_4523,N_4261,N_4401);
or U4524 (N_4524,N_4270,N_4324);
nand U4525 (N_4525,N_4357,N_4486);
and U4526 (N_4526,N_4430,N_4407);
or U4527 (N_4527,N_4364,N_4482);
or U4528 (N_4528,N_4320,N_4286);
or U4529 (N_4529,N_4252,N_4372);
or U4530 (N_4530,N_4355,N_4340);
nand U4531 (N_4531,N_4424,N_4378);
nand U4532 (N_4532,N_4351,N_4299);
nor U4533 (N_4533,N_4386,N_4284);
nor U4534 (N_4534,N_4303,N_4343);
and U4535 (N_4535,N_4266,N_4497);
xnor U4536 (N_4536,N_4370,N_4337);
and U4537 (N_4537,N_4329,N_4308);
xor U4538 (N_4538,N_4289,N_4288);
or U4539 (N_4539,N_4450,N_4301);
or U4540 (N_4540,N_4297,N_4298);
nor U4541 (N_4541,N_4319,N_4280);
xnor U4542 (N_4542,N_4416,N_4432);
nor U4543 (N_4543,N_4315,N_4271);
nor U4544 (N_4544,N_4294,N_4346);
nand U4545 (N_4545,N_4473,N_4498);
nor U4546 (N_4546,N_4264,N_4338);
xor U4547 (N_4547,N_4339,N_4376);
nand U4548 (N_4548,N_4485,N_4461);
and U4549 (N_4549,N_4317,N_4327);
or U4550 (N_4550,N_4456,N_4402);
or U4551 (N_4551,N_4390,N_4349);
and U4552 (N_4552,N_4306,N_4487);
and U4553 (N_4553,N_4275,N_4458);
nand U4554 (N_4554,N_4354,N_4448);
nor U4555 (N_4555,N_4366,N_4421);
nor U4556 (N_4556,N_4419,N_4262);
and U4557 (N_4557,N_4316,N_4309);
xnor U4558 (N_4558,N_4287,N_4375);
and U4559 (N_4559,N_4468,N_4281);
or U4560 (N_4560,N_4341,N_4428);
nand U4561 (N_4561,N_4277,N_4423);
nand U4562 (N_4562,N_4267,N_4290);
xnor U4563 (N_4563,N_4385,N_4470);
nor U4564 (N_4564,N_4253,N_4352);
nor U4565 (N_4565,N_4457,N_4471);
nand U4566 (N_4566,N_4472,N_4314);
and U4567 (N_4567,N_4488,N_4394);
xor U4568 (N_4568,N_4462,N_4459);
or U4569 (N_4569,N_4363,N_4344);
xor U4570 (N_4570,N_4444,N_4383);
or U4571 (N_4571,N_4499,N_4361);
nand U4572 (N_4572,N_4265,N_4273);
or U4573 (N_4573,N_4463,N_4446);
nor U4574 (N_4574,N_4387,N_4269);
nor U4575 (N_4575,N_4345,N_4283);
xnor U4576 (N_4576,N_4334,N_4296);
or U4577 (N_4577,N_4483,N_4415);
nand U4578 (N_4578,N_4454,N_4335);
nand U4579 (N_4579,N_4452,N_4251);
and U4580 (N_4580,N_4250,N_4420);
nor U4581 (N_4581,N_4367,N_4469);
and U4582 (N_4582,N_4307,N_4494);
nand U4583 (N_4583,N_4403,N_4437);
nand U4584 (N_4584,N_4431,N_4475);
nor U4585 (N_4585,N_4449,N_4389);
xnor U4586 (N_4586,N_4310,N_4412);
nor U4587 (N_4587,N_4295,N_4429);
and U4588 (N_4588,N_4398,N_4484);
xor U4589 (N_4589,N_4302,N_4481);
nand U4590 (N_4590,N_4360,N_4395);
and U4591 (N_4591,N_4392,N_4292);
and U4592 (N_4592,N_4373,N_4332);
nor U4593 (N_4593,N_4257,N_4439);
nand U4594 (N_4594,N_4322,N_4382);
and U4595 (N_4595,N_4427,N_4358);
nor U4596 (N_4596,N_4413,N_4493);
nor U4597 (N_4597,N_4426,N_4362);
nand U4598 (N_4598,N_4371,N_4258);
nand U4599 (N_4599,N_4405,N_4268);
and U4600 (N_4600,N_4490,N_4455);
or U4601 (N_4601,N_4442,N_4336);
nor U4602 (N_4602,N_4359,N_4422);
nor U4603 (N_4603,N_4406,N_4328);
xor U4604 (N_4604,N_4391,N_4313);
nand U4605 (N_4605,N_4434,N_4323);
and U4606 (N_4606,N_4436,N_4379);
xnor U4607 (N_4607,N_4393,N_4331);
xor U4608 (N_4608,N_4465,N_4365);
or U4609 (N_4609,N_4464,N_4467);
or U4610 (N_4610,N_4312,N_4411);
and U4611 (N_4611,N_4414,N_4495);
nor U4612 (N_4612,N_4279,N_4333);
xnor U4613 (N_4613,N_4451,N_4278);
or U4614 (N_4614,N_4293,N_4447);
or U4615 (N_4615,N_4410,N_4330);
or U4616 (N_4616,N_4397,N_4311);
nor U4617 (N_4617,N_4409,N_4285);
xor U4618 (N_4618,N_4418,N_4496);
xnor U4619 (N_4619,N_4438,N_4443);
and U4620 (N_4620,N_4477,N_4480);
xnor U4621 (N_4621,N_4348,N_4353);
or U4622 (N_4622,N_4489,N_4374);
nand U4623 (N_4623,N_4263,N_4445);
nand U4624 (N_4624,N_4388,N_4476);
xor U4625 (N_4625,N_4493,N_4266);
nand U4626 (N_4626,N_4415,N_4457);
or U4627 (N_4627,N_4487,N_4448);
nor U4628 (N_4628,N_4434,N_4443);
nand U4629 (N_4629,N_4475,N_4439);
and U4630 (N_4630,N_4379,N_4496);
and U4631 (N_4631,N_4482,N_4435);
and U4632 (N_4632,N_4287,N_4428);
nor U4633 (N_4633,N_4250,N_4328);
or U4634 (N_4634,N_4474,N_4273);
nor U4635 (N_4635,N_4377,N_4454);
nand U4636 (N_4636,N_4450,N_4275);
and U4637 (N_4637,N_4281,N_4367);
nand U4638 (N_4638,N_4424,N_4495);
nand U4639 (N_4639,N_4278,N_4498);
nor U4640 (N_4640,N_4438,N_4369);
xnor U4641 (N_4641,N_4381,N_4487);
nand U4642 (N_4642,N_4259,N_4258);
nor U4643 (N_4643,N_4310,N_4468);
nand U4644 (N_4644,N_4479,N_4452);
nor U4645 (N_4645,N_4360,N_4389);
and U4646 (N_4646,N_4412,N_4465);
and U4647 (N_4647,N_4492,N_4398);
or U4648 (N_4648,N_4339,N_4362);
xnor U4649 (N_4649,N_4424,N_4310);
nor U4650 (N_4650,N_4289,N_4315);
and U4651 (N_4651,N_4331,N_4297);
or U4652 (N_4652,N_4441,N_4373);
and U4653 (N_4653,N_4300,N_4442);
and U4654 (N_4654,N_4287,N_4362);
or U4655 (N_4655,N_4368,N_4403);
nand U4656 (N_4656,N_4257,N_4483);
nand U4657 (N_4657,N_4489,N_4416);
nor U4658 (N_4658,N_4425,N_4328);
or U4659 (N_4659,N_4401,N_4290);
nand U4660 (N_4660,N_4474,N_4423);
nor U4661 (N_4661,N_4302,N_4474);
and U4662 (N_4662,N_4440,N_4430);
nor U4663 (N_4663,N_4351,N_4337);
xnor U4664 (N_4664,N_4431,N_4302);
or U4665 (N_4665,N_4494,N_4454);
nand U4666 (N_4666,N_4416,N_4288);
nor U4667 (N_4667,N_4312,N_4477);
and U4668 (N_4668,N_4488,N_4425);
nand U4669 (N_4669,N_4421,N_4299);
nand U4670 (N_4670,N_4358,N_4332);
xnor U4671 (N_4671,N_4445,N_4433);
nand U4672 (N_4672,N_4262,N_4267);
or U4673 (N_4673,N_4335,N_4416);
xnor U4674 (N_4674,N_4265,N_4294);
xor U4675 (N_4675,N_4285,N_4405);
xor U4676 (N_4676,N_4285,N_4425);
and U4677 (N_4677,N_4406,N_4431);
xor U4678 (N_4678,N_4468,N_4295);
and U4679 (N_4679,N_4403,N_4451);
nand U4680 (N_4680,N_4313,N_4329);
xnor U4681 (N_4681,N_4396,N_4298);
xor U4682 (N_4682,N_4256,N_4465);
xor U4683 (N_4683,N_4477,N_4460);
or U4684 (N_4684,N_4315,N_4272);
nand U4685 (N_4685,N_4357,N_4256);
and U4686 (N_4686,N_4412,N_4298);
nor U4687 (N_4687,N_4276,N_4394);
or U4688 (N_4688,N_4466,N_4388);
nand U4689 (N_4689,N_4306,N_4412);
nor U4690 (N_4690,N_4313,N_4452);
nor U4691 (N_4691,N_4377,N_4367);
and U4692 (N_4692,N_4313,N_4427);
nand U4693 (N_4693,N_4298,N_4321);
nor U4694 (N_4694,N_4452,N_4395);
or U4695 (N_4695,N_4279,N_4377);
and U4696 (N_4696,N_4339,N_4375);
nor U4697 (N_4697,N_4377,N_4475);
nor U4698 (N_4698,N_4287,N_4286);
or U4699 (N_4699,N_4354,N_4328);
or U4700 (N_4700,N_4297,N_4460);
or U4701 (N_4701,N_4257,N_4488);
nor U4702 (N_4702,N_4364,N_4340);
xor U4703 (N_4703,N_4463,N_4344);
xor U4704 (N_4704,N_4270,N_4463);
xor U4705 (N_4705,N_4445,N_4256);
xor U4706 (N_4706,N_4418,N_4383);
and U4707 (N_4707,N_4454,N_4455);
nand U4708 (N_4708,N_4434,N_4468);
and U4709 (N_4709,N_4326,N_4464);
nand U4710 (N_4710,N_4319,N_4251);
or U4711 (N_4711,N_4470,N_4458);
nand U4712 (N_4712,N_4342,N_4415);
nor U4713 (N_4713,N_4305,N_4349);
or U4714 (N_4714,N_4396,N_4359);
nand U4715 (N_4715,N_4346,N_4376);
and U4716 (N_4716,N_4413,N_4374);
nand U4717 (N_4717,N_4461,N_4342);
or U4718 (N_4718,N_4410,N_4279);
or U4719 (N_4719,N_4410,N_4493);
and U4720 (N_4720,N_4340,N_4444);
nand U4721 (N_4721,N_4482,N_4456);
xnor U4722 (N_4722,N_4378,N_4371);
nor U4723 (N_4723,N_4466,N_4351);
nand U4724 (N_4724,N_4362,N_4324);
xnor U4725 (N_4725,N_4255,N_4290);
xnor U4726 (N_4726,N_4313,N_4465);
nor U4727 (N_4727,N_4286,N_4360);
xnor U4728 (N_4728,N_4454,N_4375);
nand U4729 (N_4729,N_4389,N_4474);
nor U4730 (N_4730,N_4361,N_4424);
xor U4731 (N_4731,N_4435,N_4286);
nand U4732 (N_4732,N_4472,N_4399);
nand U4733 (N_4733,N_4346,N_4328);
xnor U4734 (N_4734,N_4348,N_4489);
xor U4735 (N_4735,N_4251,N_4460);
nand U4736 (N_4736,N_4488,N_4416);
and U4737 (N_4737,N_4437,N_4452);
nand U4738 (N_4738,N_4299,N_4348);
and U4739 (N_4739,N_4256,N_4302);
nand U4740 (N_4740,N_4373,N_4370);
nor U4741 (N_4741,N_4294,N_4304);
or U4742 (N_4742,N_4335,N_4377);
nor U4743 (N_4743,N_4334,N_4262);
nand U4744 (N_4744,N_4340,N_4406);
nor U4745 (N_4745,N_4400,N_4334);
nor U4746 (N_4746,N_4337,N_4341);
and U4747 (N_4747,N_4336,N_4348);
and U4748 (N_4748,N_4378,N_4483);
nand U4749 (N_4749,N_4293,N_4409);
and U4750 (N_4750,N_4602,N_4611);
or U4751 (N_4751,N_4685,N_4712);
nand U4752 (N_4752,N_4678,N_4671);
and U4753 (N_4753,N_4644,N_4572);
and U4754 (N_4754,N_4716,N_4717);
nand U4755 (N_4755,N_4512,N_4664);
or U4756 (N_4756,N_4709,N_4626);
or U4757 (N_4757,N_4704,N_4558);
or U4758 (N_4758,N_4625,N_4576);
or U4759 (N_4759,N_4503,N_4645);
nand U4760 (N_4760,N_4598,N_4615);
nand U4761 (N_4761,N_4525,N_4562);
xnor U4762 (N_4762,N_4532,N_4630);
nor U4763 (N_4763,N_4601,N_4698);
xnor U4764 (N_4764,N_4741,N_4680);
nand U4765 (N_4765,N_4560,N_4675);
or U4766 (N_4766,N_4731,N_4563);
xor U4767 (N_4767,N_4553,N_4662);
nor U4768 (N_4768,N_4573,N_4647);
xnor U4769 (N_4769,N_4679,N_4556);
xnor U4770 (N_4770,N_4642,N_4546);
nand U4771 (N_4771,N_4551,N_4591);
nor U4772 (N_4772,N_4708,N_4640);
nor U4773 (N_4773,N_4557,N_4508);
or U4774 (N_4774,N_4540,N_4739);
nor U4775 (N_4775,N_4550,N_4633);
or U4776 (N_4776,N_4606,N_4649);
xor U4777 (N_4777,N_4618,N_4722);
nand U4778 (N_4778,N_4746,N_4581);
and U4779 (N_4779,N_4693,N_4518);
and U4780 (N_4780,N_4736,N_4720);
and U4781 (N_4781,N_4669,N_4545);
and U4782 (N_4782,N_4531,N_4529);
xnor U4783 (N_4783,N_4578,N_4569);
xnor U4784 (N_4784,N_4723,N_4530);
xor U4785 (N_4785,N_4605,N_4730);
nand U4786 (N_4786,N_4665,N_4652);
and U4787 (N_4787,N_4747,N_4663);
or U4788 (N_4788,N_4537,N_4543);
nand U4789 (N_4789,N_4509,N_4710);
xor U4790 (N_4790,N_4570,N_4506);
nor U4791 (N_4791,N_4511,N_4707);
and U4792 (N_4792,N_4701,N_4660);
nand U4793 (N_4793,N_4728,N_4586);
xnor U4794 (N_4794,N_4564,N_4523);
and U4795 (N_4795,N_4691,N_4513);
and U4796 (N_4796,N_4634,N_4737);
nor U4797 (N_4797,N_4502,N_4734);
nand U4798 (N_4798,N_4619,N_4654);
nor U4799 (N_4799,N_4639,N_4585);
and U4800 (N_4800,N_4657,N_4745);
xnor U4801 (N_4801,N_4536,N_4603);
xnor U4802 (N_4802,N_4519,N_4700);
nand U4803 (N_4803,N_4686,N_4596);
nor U4804 (N_4804,N_4705,N_4735);
xor U4805 (N_4805,N_4588,N_4667);
or U4806 (N_4806,N_4677,N_4517);
xor U4807 (N_4807,N_4661,N_4539);
and U4808 (N_4808,N_4515,N_4547);
nor U4809 (N_4809,N_4706,N_4617);
xnor U4810 (N_4810,N_4582,N_4610);
or U4811 (N_4811,N_4594,N_4656);
or U4812 (N_4812,N_4621,N_4628);
nor U4813 (N_4813,N_4714,N_4697);
or U4814 (N_4814,N_4579,N_4505);
nor U4815 (N_4815,N_4533,N_4609);
nand U4816 (N_4816,N_4666,N_4524);
xor U4817 (N_4817,N_4718,N_4554);
nor U4818 (N_4818,N_4629,N_4528);
nor U4819 (N_4819,N_4672,N_4608);
nand U4820 (N_4820,N_4648,N_4583);
and U4821 (N_4821,N_4538,N_4552);
xor U4822 (N_4822,N_4544,N_4692);
or U4823 (N_4823,N_4719,N_4541);
and U4824 (N_4824,N_4616,N_4699);
or U4825 (N_4825,N_4743,N_4690);
or U4826 (N_4826,N_4565,N_4650);
nand U4827 (N_4827,N_4670,N_4548);
nor U4828 (N_4828,N_4729,N_4724);
xnor U4829 (N_4829,N_4643,N_4504);
nor U4830 (N_4830,N_4668,N_4674);
nand U4831 (N_4831,N_4721,N_4655);
nor U4832 (N_4832,N_4584,N_4627);
and U4833 (N_4833,N_4738,N_4561);
xnor U4834 (N_4834,N_4631,N_4636);
nor U4835 (N_4835,N_4744,N_4742);
and U4836 (N_4836,N_4571,N_4507);
or U4837 (N_4837,N_4549,N_4559);
nor U4838 (N_4838,N_4555,N_4695);
nor U4839 (N_4839,N_4614,N_4587);
xnor U4840 (N_4840,N_4658,N_4580);
or U4841 (N_4841,N_4501,N_4676);
nor U4842 (N_4842,N_4600,N_4567);
nor U4843 (N_4843,N_4715,N_4632);
xor U4844 (N_4844,N_4590,N_4542);
nor U4845 (N_4845,N_4620,N_4684);
nand U4846 (N_4846,N_4688,N_4592);
and U4847 (N_4847,N_4595,N_4589);
nor U4848 (N_4848,N_4651,N_4749);
nand U4849 (N_4849,N_4659,N_4575);
nand U4850 (N_4850,N_4607,N_4703);
xor U4851 (N_4851,N_4624,N_4622);
or U4852 (N_4852,N_4568,N_4534);
or U4853 (N_4853,N_4637,N_4500);
nand U4854 (N_4854,N_4604,N_4566);
xnor U4855 (N_4855,N_4516,N_4612);
xor U4856 (N_4856,N_4593,N_4748);
and U4857 (N_4857,N_4687,N_4727);
nand U4858 (N_4858,N_4682,N_4689);
xnor U4859 (N_4859,N_4733,N_4574);
nor U4860 (N_4860,N_4673,N_4522);
nand U4861 (N_4861,N_4646,N_4577);
and U4862 (N_4862,N_4713,N_4694);
nor U4863 (N_4863,N_4641,N_4711);
and U4864 (N_4864,N_4635,N_4613);
nand U4865 (N_4865,N_4520,N_4681);
xnor U4866 (N_4866,N_4521,N_4653);
or U4867 (N_4867,N_4535,N_4526);
xor U4868 (N_4868,N_4638,N_4623);
nor U4869 (N_4869,N_4740,N_4510);
xor U4870 (N_4870,N_4726,N_4514);
and U4871 (N_4871,N_4732,N_4597);
nand U4872 (N_4872,N_4527,N_4702);
xnor U4873 (N_4873,N_4683,N_4725);
and U4874 (N_4874,N_4599,N_4696);
or U4875 (N_4875,N_4540,N_4674);
or U4876 (N_4876,N_4514,N_4570);
or U4877 (N_4877,N_4562,N_4728);
xnor U4878 (N_4878,N_4520,N_4684);
and U4879 (N_4879,N_4745,N_4645);
xnor U4880 (N_4880,N_4629,N_4655);
nor U4881 (N_4881,N_4637,N_4534);
or U4882 (N_4882,N_4518,N_4656);
nand U4883 (N_4883,N_4635,N_4743);
xnor U4884 (N_4884,N_4555,N_4648);
or U4885 (N_4885,N_4572,N_4725);
and U4886 (N_4886,N_4647,N_4669);
nor U4887 (N_4887,N_4560,N_4654);
xor U4888 (N_4888,N_4672,N_4522);
and U4889 (N_4889,N_4742,N_4527);
nand U4890 (N_4890,N_4623,N_4540);
nand U4891 (N_4891,N_4749,N_4702);
nor U4892 (N_4892,N_4660,N_4528);
nor U4893 (N_4893,N_4675,N_4632);
and U4894 (N_4894,N_4660,N_4748);
nand U4895 (N_4895,N_4671,N_4528);
xnor U4896 (N_4896,N_4641,N_4713);
or U4897 (N_4897,N_4556,N_4518);
nor U4898 (N_4898,N_4500,N_4593);
nand U4899 (N_4899,N_4595,N_4511);
nand U4900 (N_4900,N_4661,N_4597);
xor U4901 (N_4901,N_4660,N_4669);
and U4902 (N_4902,N_4694,N_4726);
nor U4903 (N_4903,N_4655,N_4553);
nor U4904 (N_4904,N_4687,N_4631);
nor U4905 (N_4905,N_4585,N_4506);
and U4906 (N_4906,N_4721,N_4593);
or U4907 (N_4907,N_4739,N_4686);
nor U4908 (N_4908,N_4545,N_4571);
nor U4909 (N_4909,N_4743,N_4730);
nand U4910 (N_4910,N_4700,N_4638);
nor U4911 (N_4911,N_4556,N_4730);
nand U4912 (N_4912,N_4566,N_4542);
and U4913 (N_4913,N_4718,N_4587);
nand U4914 (N_4914,N_4671,N_4585);
nor U4915 (N_4915,N_4523,N_4673);
nand U4916 (N_4916,N_4515,N_4583);
or U4917 (N_4917,N_4680,N_4682);
or U4918 (N_4918,N_4608,N_4500);
and U4919 (N_4919,N_4543,N_4723);
xnor U4920 (N_4920,N_4744,N_4605);
nor U4921 (N_4921,N_4645,N_4570);
or U4922 (N_4922,N_4748,N_4726);
xor U4923 (N_4923,N_4641,N_4502);
and U4924 (N_4924,N_4517,N_4698);
nor U4925 (N_4925,N_4588,N_4515);
xor U4926 (N_4926,N_4504,N_4730);
nand U4927 (N_4927,N_4591,N_4636);
or U4928 (N_4928,N_4630,N_4627);
nand U4929 (N_4929,N_4685,N_4523);
nor U4930 (N_4930,N_4561,N_4743);
and U4931 (N_4931,N_4503,N_4566);
xnor U4932 (N_4932,N_4614,N_4627);
and U4933 (N_4933,N_4652,N_4688);
nor U4934 (N_4934,N_4596,N_4679);
xor U4935 (N_4935,N_4741,N_4731);
and U4936 (N_4936,N_4712,N_4510);
and U4937 (N_4937,N_4657,N_4701);
xor U4938 (N_4938,N_4553,N_4561);
nor U4939 (N_4939,N_4580,N_4727);
and U4940 (N_4940,N_4575,N_4688);
nand U4941 (N_4941,N_4639,N_4542);
xnor U4942 (N_4942,N_4568,N_4528);
nand U4943 (N_4943,N_4521,N_4714);
and U4944 (N_4944,N_4654,N_4675);
or U4945 (N_4945,N_4749,N_4584);
or U4946 (N_4946,N_4723,N_4748);
nor U4947 (N_4947,N_4744,N_4714);
nand U4948 (N_4948,N_4635,N_4651);
xnor U4949 (N_4949,N_4549,N_4591);
xnor U4950 (N_4950,N_4574,N_4735);
xor U4951 (N_4951,N_4562,N_4647);
nor U4952 (N_4952,N_4619,N_4596);
nand U4953 (N_4953,N_4633,N_4746);
xor U4954 (N_4954,N_4690,N_4604);
or U4955 (N_4955,N_4542,N_4520);
and U4956 (N_4956,N_4520,N_4563);
or U4957 (N_4957,N_4526,N_4708);
and U4958 (N_4958,N_4568,N_4623);
or U4959 (N_4959,N_4549,N_4553);
nand U4960 (N_4960,N_4644,N_4636);
nand U4961 (N_4961,N_4568,N_4650);
nand U4962 (N_4962,N_4575,N_4576);
nand U4963 (N_4963,N_4516,N_4629);
nor U4964 (N_4964,N_4513,N_4576);
or U4965 (N_4965,N_4597,N_4703);
nor U4966 (N_4966,N_4675,N_4645);
nor U4967 (N_4967,N_4513,N_4695);
or U4968 (N_4968,N_4655,N_4536);
xnor U4969 (N_4969,N_4698,N_4720);
or U4970 (N_4970,N_4543,N_4560);
and U4971 (N_4971,N_4500,N_4738);
or U4972 (N_4972,N_4573,N_4739);
nor U4973 (N_4973,N_4619,N_4742);
and U4974 (N_4974,N_4594,N_4575);
nor U4975 (N_4975,N_4698,N_4640);
nand U4976 (N_4976,N_4673,N_4692);
nand U4977 (N_4977,N_4546,N_4718);
xor U4978 (N_4978,N_4669,N_4705);
xor U4979 (N_4979,N_4544,N_4672);
or U4980 (N_4980,N_4574,N_4614);
xnor U4981 (N_4981,N_4502,N_4733);
and U4982 (N_4982,N_4625,N_4739);
xor U4983 (N_4983,N_4572,N_4653);
xor U4984 (N_4984,N_4660,N_4532);
and U4985 (N_4985,N_4639,N_4707);
nand U4986 (N_4986,N_4709,N_4712);
and U4987 (N_4987,N_4726,N_4554);
and U4988 (N_4988,N_4665,N_4702);
and U4989 (N_4989,N_4651,N_4535);
xnor U4990 (N_4990,N_4646,N_4641);
xor U4991 (N_4991,N_4578,N_4538);
or U4992 (N_4992,N_4529,N_4683);
or U4993 (N_4993,N_4577,N_4746);
xnor U4994 (N_4994,N_4681,N_4527);
or U4995 (N_4995,N_4524,N_4623);
or U4996 (N_4996,N_4688,N_4553);
or U4997 (N_4997,N_4593,N_4624);
nand U4998 (N_4998,N_4580,N_4636);
xor U4999 (N_4999,N_4545,N_4582);
and U5000 (N_5000,N_4770,N_4885);
and U5001 (N_5001,N_4769,N_4812);
xor U5002 (N_5002,N_4760,N_4789);
and U5003 (N_5003,N_4937,N_4849);
and U5004 (N_5004,N_4883,N_4992);
xnor U5005 (N_5005,N_4975,N_4833);
xor U5006 (N_5006,N_4775,N_4831);
or U5007 (N_5007,N_4822,N_4906);
nor U5008 (N_5008,N_4844,N_4820);
and U5009 (N_5009,N_4862,N_4797);
nor U5010 (N_5010,N_4819,N_4949);
nand U5011 (N_5011,N_4889,N_4825);
nand U5012 (N_5012,N_4936,N_4841);
and U5013 (N_5013,N_4787,N_4805);
nand U5014 (N_5014,N_4791,N_4972);
nor U5015 (N_5015,N_4919,N_4907);
nor U5016 (N_5016,N_4998,N_4839);
nand U5017 (N_5017,N_4943,N_4955);
xor U5018 (N_5018,N_4980,N_4873);
nor U5019 (N_5019,N_4814,N_4781);
nand U5020 (N_5020,N_4855,N_4934);
nand U5021 (N_5021,N_4864,N_4804);
xor U5022 (N_5022,N_4989,N_4891);
or U5023 (N_5023,N_4903,N_4914);
nor U5024 (N_5024,N_4939,N_4821);
nor U5025 (N_5025,N_4778,N_4963);
nor U5026 (N_5026,N_4995,N_4986);
xor U5027 (N_5027,N_4878,N_4780);
and U5028 (N_5028,N_4913,N_4897);
and U5029 (N_5029,N_4796,N_4852);
or U5030 (N_5030,N_4857,N_4771);
and U5031 (N_5031,N_4793,N_4872);
nand U5032 (N_5032,N_4886,N_4868);
nand U5033 (N_5033,N_4846,N_4899);
xnor U5034 (N_5034,N_4764,N_4880);
and U5035 (N_5035,N_4921,N_4948);
nor U5036 (N_5036,N_4794,N_4884);
nor U5037 (N_5037,N_4959,N_4984);
and U5038 (N_5038,N_4946,N_4993);
or U5039 (N_5039,N_4938,N_4920);
or U5040 (N_5040,N_4942,N_4837);
and U5041 (N_5041,N_4973,N_4836);
nand U5042 (N_5042,N_4982,N_4991);
xor U5043 (N_5043,N_4815,N_4843);
nand U5044 (N_5044,N_4790,N_4887);
and U5045 (N_5045,N_4924,N_4823);
nor U5046 (N_5046,N_4828,N_4751);
nand U5047 (N_5047,N_4900,N_4768);
and U5048 (N_5048,N_4757,N_4809);
nor U5049 (N_5049,N_4990,N_4935);
nand U5050 (N_5050,N_4803,N_4850);
nor U5051 (N_5051,N_4902,N_4853);
and U5052 (N_5052,N_4918,N_4896);
xor U5053 (N_5053,N_4956,N_4786);
and U5054 (N_5054,N_4763,N_4863);
or U5055 (N_5055,N_4783,N_4867);
nor U5056 (N_5056,N_4871,N_4890);
nand U5057 (N_5057,N_4964,N_4944);
xor U5058 (N_5058,N_4818,N_4877);
xnor U5059 (N_5059,N_4826,N_4970);
xor U5060 (N_5060,N_4908,N_4917);
or U5061 (N_5061,N_4951,N_4881);
nand U5062 (N_5062,N_4997,N_4926);
or U5063 (N_5063,N_4807,N_4999);
xor U5064 (N_5064,N_4953,N_4952);
nand U5065 (N_5065,N_4824,N_4861);
or U5066 (N_5066,N_4892,N_4945);
and U5067 (N_5067,N_4947,N_4830);
nor U5068 (N_5068,N_4750,N_4865);
or U5069 (N_5069,N_4759,N_4869);
or U5070 (N_5070,N_4829,N_4974);
xor U5071 (N_5071,N_4772,N_4859);
nand U5072 (N_5072,N_4933,N_4761);
and U5073 (N_5073,N_4785,N_4879);
or U5074 (N_5074,N_4976,N_4876);
or U5075 (N_5075,N_4983,N_4792);
xor U5076 (N_5076,N_4842,N_4838);
or U5077 (N_5077,N_4985,N_4898);
or U5078 (N_5078,N_4755,N_4860);
nand U5079 (N_5079,N_4988,N_4777);
nand U5080 (N_5080,N_4977,N_4782);
nand U5081 (N_5081,N_4911,N_4758);
nand U5082 (N_5082,N_4813,N_4774);
or U5083 (N_5083,N_4962,N_4895);
nand U5084 (N_5084,N_4932,N_4784);
nand U5085 (N_5085,N_4776,N_4929);
xnor U5086 (N_5086,N_4882,N_4806);
nor U5087 (N_5087,N_4971,N_4870);
or U5088 (N_5088,N_4752,N_4979);
nand U5089 (N_5089,N_4874,N_4957);
nand U5090 (N_5090,N_4795,N_4847);
xnor U5091 (N_5091,N_4856,N_4910);
xor U5092 (N_5092,N_4912,N_4969);
xor U5093 (N_5093,N_4923,N_4940);
or U5094 (N_5094,N_4779,N_4909);
nand U5095 (N_5095,N_4840,N_4773);
or U5096 (N_5096,N_4834,N_4893);
nor U5097 (N_5097,N_4987,N_4765);
nand U5098 (N_5098,N_4767,N_4845);
nand U5099 (N_5099,N_4916,N_4858);
and U5100 (N_5100,N_4762,N_4808);
or U5101 (N_5101,N_4799,N_4922);
nand U5102 (N_5102,N_4978,N_4958);
or U5103 (N_5103,N_4753,N_4816);
nor U5104 (N_5104,N_4788,N_4854);
nand U5105 (N_5105,N_4800,N_4866);
and U5106 (N_5106,N_4801,N_4927);
and U5107 (N_5107,N_4901,N_4811);
nand U5108 (N_5108,N_4954,N_4925);
and U5109 (N_5109,N_4996,N_4798);
or U5110 (N_5110,N_4968,N_4967);
or U5111 (N_5111,N_4802,N_4915);
xnor U5112 (N_5112,N_4994,N_4960);
nand U5113 (N_5113,N_4931,N_4766);
xnor U5114 (N_5114,N_4894,N_4817);
nor U5115 (N_5115,N_4756,N_4928);
xor U5116 (N_5116,N_4835,N_4981);
nand U5117 (N_5117,N_4848,N_4961);
xnor U5118 (N_5118,N_4851,N_4832);
nand U5119 (N_5119,N_4888,N_4754);
xor U5120 (N_5120,N_4875,N_4810);
xor U5121 (N_5121,N_4905,N_4966);
nor U5122 (N_5122,N_4904,N_4827);
nand U5123 (N_5123,N_4941,N_4930);
xor U5124 (N_5124,N_4965,N_4950);
or U5125 (N_5125,N_4877,N_4895);
xnor U5126 (N_5126,N_4847,N_4932);
xnor U5127 (N_5127,N_4894,N_4761);
or U5128 (N_5128,N_4920,N_4895);
nor U5129 (N_5129,N_4750,N_4801);
xor U5130 (N_5130,N_4879,N_4813);
nor U5131 (N_5131,N_4813,N_4836);
xnor U5132 (N_5132,N_4844,N_4866);
and U5133 (N_5133,N_4829,N_4919);
nand U5134 (N_5134,N_4781,N_4788);
nor U5135 (N_5135,N_4994,N_4814);
nand U5136 (N_5136,N_4809,N_4894);
nand U5137 (N_5137,N_4828,N_4976);
xnor U5138 (N_5138,N_4823,N_4977);
nor U5139 (N_5139,N_4870,N_4832);
nand U5140 (N_5140,N_4999,N_4988);
nor U5141 (N_5141,N_4774,N_4960);
nand U5142 (N_5142,N_4892,N_4905);
nand U5143 (N_5143,N_4802,N_4791);
nor U5144 (N_5144,N_4879,N_4811);
and U5145 (N_5145,N_4787,N_4984);
or U5146 (N_5146,N_4784,N_4778);
xnor U5147 (N_5147,N_4782,N_4795);
or U5148 (N_5148,N_4942,N_4892);
or U5149 (N_5149,N_4851,N_4769);
and U5150 (N_5150,N_4903,N_4937);
xnor U5151 (N_5151,N_4989,N_4924);
and U5152 (N_5152,N_4940,N_4794);
and U5153 (N_5153,N_4845,N_4994);
nor U5154 (N_5154,N_4936,N_4800);
or U5155 (N_5155,N_4770,N_4962);
or U5156 (N_5156,N_4905,N_4865);
and U5157 (N_5157,N_4914,N_4839);
nor U5158 (N_5158,N_4822,N_4905);
nor U5159 (N_5159,N_4919,N_4822);
and U5160 (N_5160,N_4976,N_4926);
or U5161 (N_5161,N_4876,N_4793);
or U5162 (N_5162,N_4996,N_4931);
or U5163 (N_5163,N_4840,N_4877);
or U5164 (N_5164,N_4962,N_4822);
xnor U5165 (N_5165,N_4964,N_4758);
xor U5166 (N_5166,N_4976,N_4774);
xor U5167 (N_5167,N_4807,N_4935);
nand U5168 (N_5168,N_4785,N_4765);
or U5169 (N_5169,N_4938,N_4966);
nor U5170 (N_5170,N_4936,N_4833);
xnor U5171 (N_5171,N_4964,N_4771);
nor U5172 (N_5172,N_4959,N_4901);
nor U5173 (N_5173,N_4905,N_4967);
or U5174 (N_5174,N_4811,N_4947);
xor U5175 (N_5175,N_4903,N_4890);
xor U5176 (N_5176,N_4807,N_4907);
nand U5177 (N_5177,N_4810,N_4835);
nand U5178 (N_5178,N_4875,N_4898);
and U5179 (N_5179,N_4788,N_4757);
nand U5180 (N_5180,N_4991,N_4870);
nor U5181 (N_5181,N_4783,N_4918);
nand U5182 (N_5182,N_4989,N_4912);
nor U5183 (N_5183,N_4873,N_4856);
nand U5184 (N_5184,N_4915,N_4936);
or U5185 (N_5185,N_4921,N_4958);
and U5186 (N_5186,N_4889,N_4940);
and U5187 (N_5187,N_4886,N_4961);
xor U5188 (N_5188,N_4954,N_4819);
nand U5189 (N_5189,N_4897,N_4915);
and U5190 (N_5190,N_4890,N_4994);
or U5191 (N_5191,N_4987,N_4793);
xnor U5192 (N_5192,N_4778,N_4989);
nor U5193 (N_5193,N_4952,N_4913);
nand U5194 (N_5194,N_4809,N_4869);
nand U5195 (N_5195,N_4800,N_4858);
nand U5196 (N_5196,N_4969,N_4989);
nor U5197 (N_5197,N_4852,N_4826);
nor U5198 (N_5198,N_4921,N_4865);
nand U5199 (N_5199,N_4894,N_4787);
nand U5200 (N_5200,N_4901,N_4822);
xor U5201 (N_5201,N_4856,N_4782);
nand U5202 (N_5202,N_4895,N_4917);
xor U5203 (N_5203,N_4822,N_4913);
xor U5204 (N_5204,N_4765,N_4827);
or U5205 (N_5205,N_4810,N_4967);
xnor U5206 (N_5206,N_4988,N_4782);
xor U5207 (N_5207,N_4775,N_4985);
or U5208 (N_5208,N_4751,N_4902);
and U5209 (N_5209,N_4909,N_4801);
nand U5210 (N_5210,N_4807,N_4804);
nand U5211 (N_5211,N_4817,N_4776);
xnor U5212 (N_5212,N_4908,N_4760);
and U5213 (N_5213,N_4836,N_4817);
nor U5214 (N_5214,N_4894,N_4783);
xnor U5215 (N_5215,N_4992,N_4790);
xnor U5216 (N_5216,N_4984,N_4752);
nand U5217 (N_5217,N_4884,N_4910);
or U5218 (N_5218,N_4973,N_4812);
xnor U5219 (N_5219,N_4944,N_4991);
or U5220 (N_5220,N_4761,N_4920);
nor U5221 (N_5221,N_4789,N_4888);
and U5222 (N_5222,N_4862,N_4759);
xnor U5223 (N_5223,N_4752,N_4788);
nand U5224 (N_5224,N_4775,N_4837);
or U5225 (N_5225,N_4805,N_4950);
xor U5226 (N_5226,N_4864,N_4962);
nand U5227 (N_5227,N_4852,N_4776);
or U5228 (N_5228,N_4961,N_4841);
and U5229 (N_5229,N_4906,N_4798);
and U5230 (N_5230,N_4791,N_4860);
or U5231 (N_5231,N_4915,N_4968);
and U5232 (N_5232,N_4849,N_4847);
nand U5233 (N_5233,N_4962,N_4844);
or U5234 (N_5234,N_4853,N_4906);
nor U5235 (N_5235,N_4861,N_4794);
xnor U5236 (N_5236,N_4793,N_4881);
and U5237 (N_5237,N_4979,N_4866);
nor U5238 (N_5238,N_4921,N_4754);
nor U5239 (N_5239,N_4813,N_4797);
nor U5240 (N_5240,N_4767,N_4849);
nor U5241 (N_5241,N_4960,N_4997);
nand U5242 (N_5242,N_4938,N_4929);
nand U5243 (N_5243,N_4842,N_4965);
and U5244 (N_5244,N_4926,N_4794);
nor U5245 (N_5245,N_4914,N_4910);
nor U5246 (N_5246,N_4848,N_4912);
nand U5247 (N_5247,N_4847,N_4771);
or U5248 (N_5248,N_4860,N_4824);
xor U5249 (N_5249,N_4777,N_4863);
nand U5250 (N_5250,N_5196,N_5000);
or U5251 (N_5251,N_5017,N_5170);
nand U5252 (N_5252,N_5155,N_5180);
nand U5253 (N_5253,N_5200,N_5206);
and U5254 (N_5254,N_5095,N_5187);
or U5255 (N_5255,N_5043,N_5157);
nor U5256 (N_5256,N_5243,N_5171);
and U5257 (N_5257,N_5124,N_5209);
nand U5258 (N_5258,N_5228,N_5247);
and U5259 (N_5259,N_5093,N_5211);
xnor U5260 (N_5260,N_5229,N_5060);
xor U5261 (N_5261,N_5055,N_5057);
or U5262 (N_5262,N_5245,N_5241);
or U5263 (N_5263,N_5233,N_5064);
nor U5264 (N_5264,N_5040,N_5129);
xnor U5265 (N_5265,N_5005,N_5092);
xnor U5266 (N_5266,N_5199,N_5079);
xnor U5267 (N_5267,N_5238,N_5136);
and U5268 (N_5268,N_5028,N_5069);
or U5269 (N_5269,N_5194,N_5003);
xor U5270 (N_5270,N_5094,N_5022);
nor U5271 (N_5271,N_5117,N_5018);
nor U5272 (N_5272,N_5008,N_5048);
nor U5273 (N_5273,N_5183,N_5220);
xor U5274 (N_5274,N_5097,N_5162);
nand U5275 (N_5275,N_5009,N_5120);
nor U5276 (N_5276,N_5218,N_5154);
xor U5277 (N_5277,N_5002,N_5163);
xor U5278 (N_5278,N_5016,N_5042);
nor U5279 (N_5279,N_5148,N_5110);
or U5280 (N_5280,N_5121,N_5081);
xor U5281 (N_5281,N_5177,N_5054);
nor U5282 (N_5282,N_5212,N_5135);
nand U5283 (N_5283,N_5026,N_5032);
nor U5284 (N_5284,N_5029,N_5050);
or U5285 (N_5285,N_5234,N_5207);
nor U5286 (N_5286,N_5244,N_5045);
nand U5287 (N_5287,N_5172,N_5138);
or U5288 (N_5288,N_5116,N_5039);
or U5289 (N_5289,N_5226,N_5181);
nor U5290 (N_5290,N_5202,N_5031);
and U5291 (N_5291,N_5114,N_5023);
nand U5292 (N_5292,N_5041,N_5070);
xnor U5293 (N_5293,N_5239,N_5127);
xor U5294 (N_5294,N_5053,N_5144);
xor U5295 (N_5295,N_5061,N_5109);
or U5296 (N_5296,N_5046,N_5189);
and U5297 (N_5297,N_5131,N_5006);
nand U5298 (N_5298,N_5160,N_5025);
nand U5299 (N_5299,N_5221,N_5216);
nand U5300 (N_5300,N_5165,N_5176);
and U5301 (N_5301,N_5237,N_5240);
nand U5302 (N_5302,N_5132,N_5084);
and U5303 (N_5303,N_5049,N_5063);
and U5304 (N_5304,N_5013,N_5075);
or U5305 (N_5305,N_5178,N_5108);
nand U5306 (N_5306,N_5098,N_5012);
nor U5307 (N_5307,N_5133,N_5100);
nand U5308 (N_5308,N_5224,N_5166);
or U5309 (N_5309,N_5204,N_5037);
nand U5310 (N_5310,N_5066,N_5236);
nor U5311 (N_5311,N_5231,N_5150);
nor U5312 (N_5312,N_5091,N_5134);
nor U5313 (N_5313,N_5174,N_5085);
xnor U5314 (N_5314,N_5077,N_5158);
nand U5315 (N_5315,N_5137,N_5130);
or U5316 (N_5316,N_5198,N_5020);
nand U5317 (N_5317,N_5071,N_5188);
or U5318 (N_5318,N_5047,N_5036);
or U5319 (N_5319,N_5147,N_5011);
nor U5320 (N_5320,N_5225,N_5125);
and U5321 (N_5321,N_5089,N_5159);
xor U5322 (N_5322,N_5118,N_5068);
or U5323 (N_5323,N_5019,N_5190);
or U5324 (N_5324,N_5219,N_5111);
or U5325 (N_5325,N_5038,N_5021);
nor U5326 (N_5326,N_5222,N_5248);
nand U5327 (N_5327,N_5030,N_5223);
xor U5328 (N_5328,N_5208,N_5001);
and U5329 (N_5329,N_5086,N_5227);
xnor U5330 (N_5330,N_5007,N_5193);
nor U5331 (N_5331,N_5076,N_5195);
and U5332 (N_5332,N_5151,N_5249);
and U5333 (N_5333,N_5024,N_5088);
and U5334 (N_5334,N_5062,N_5210);
nor U5335 (N_5335,N_5103,N_5182);
nand U5336 (N_5336,N_5142,N_5126);
nor U5337 (N_5337,N_5192,N_5052);
and U5338 (N_5338,N_5168,N_5106);
nand U5339 (N_5339,N_5156,N_5027);
nor U5340 (N_5340,N_5232,N_5051);
or U5341 (N_5341,N_5149,N_5230);
nor U5342 (N_5342,N_5179,N_5078);
nand U5343 (N_5343,N_5067,N_5105);
or U5344 (N_5344,N_5122,N_5015);
and U5345 (N_5345,N_5072,N_5123);
nor U5346 (N_5346,N_5087,N_5112);
xor U5347 (N_5347,N_5104,N_5090);
nand U5348 (N_5348,N_5191,N_5185);
nand U5349 (N_5349,N_5139,N_5065);
and U5350 (N_5350,N_5102,N_5099);
nor U5351 (N_5351,N_5004,N_5044);
and U5352 (N_5352,N_5217,N_5203);
nand U5353 (N_5353,N_5034,N_5101);
nor U5354 (N_5354,N_5115,N_5153);
xnor U5355 (N_5355,N_5215,N_5058);
nor U5356 (N_5356,N_5073,N_5056);
xor U5357 (N_5357,N_5083,N_5113);
nor U5358 (N_5358,N_5033,N_5161);
nor U5359 (N_5359,N_5143,N_5214);
nor U5360 (N_5360,N_5184,N_5152);
nor U5361 (N_5361,N_5213,N_5186);
or U5362 (N_5362,N_5242,N_5128);
or U5363 (N_5363,N_5173,N_5119);
nor U5364 (N_5364,N_5197,N_5164);
or U5365 (N_5365,N_5141,N_5169);
nor U5366 (N_5366,N_5167,N_5014);
or U5367 (N_5367,N_5145,N_5035);
nor U5368 (N_5368,N_5010,N_5205);
and U5369 (N_5369,N_5074,N_5146);
xor U5370 (N_5370,N_5175,N_5096);
nand U5371 (N_5371,N_5059,N_5082);
or U5372 (N_5372,N_5235,N_5140);
nor U5373 (N_5373,N_5107,N_5246);
nor U5374 (N_5374,N_5201,N_5080);
nand U5375 (N_5375,N_5184,N_5031);
or U5376 (N_5376,N_5244,N_5066);
or U5377 (N_5377,N_5173,N_5162);
or U5378 (N_5378,N_5176,N_5046);
or U5379 (N_5379,N_5204,N_5244);
xnor U5380 (N_5380,N_5047,N_5201);
xnor U5381 (N_5381,N_5062,N_5237);
xnor U5382 (N_5382,N_5129,N_5221);
xnor U5383 (N_5383,N_5124,N_5128);
xor U5384 (N_5384,N_5249,N_5227);
nor U5385 (N_5385,N_5015,N_5215);
xnor U5386 (N_5386,N_5161,N_5217);
and U5387 (N_5387,N_5051,N_5081);
nand U5388 (N_5388,N_5207,N_5082);
xnor U5389 (N_5389,N_5038,N_5125);
and U5390 (N_5390,N_5216,N_5102);
nor U5391 (N_5391,N_5010,N_5097);
and U5392 (N_5392,N_5139,N_5229);
or U5393 (N_5393,N_5045,N_5167);
nand U5394 (N_5394,N_5152,N_5191);
or U5395 (N_5395,N_5247,N_5080);
nand U5396 (N_5396,N_5109,N_5237);
nand U5397 (N_5397,N_5148,N_5247);
nand U5398 (N_5398,N_5032,N_5190);
nand U5399 (N_5399,N_5225,N_5037);
and U5400 (N_5400,N_5000,N_5182);
or U5401 (N_5401,N_5138,N_5182);
and U5402 (N_5402,N_5159,N_5143);
or U5403 (N_5403,N_5105,N_5077);
and U5404 (N_5404,N_5167,N_5028);
and U5405 (N_5405,N_5176,N_5183);
nand U5406 (N_5406,N_5065,N_5129);
or U5407 (N_5407,N_5045,N_5175);
xnor U5408 (N_5408,N_5077,N_5052);
and U5409 (N_5409,N_5001,N_5125);
nor U5410 (N_5410,N_5000,N_5229);
nand U5411 (N_5411,N_5047,N_5247);
nand U5412 (N_5412,N_5031,N_5173);
and U5413 (N_5413,N_5023,N_5151);
or U5414 (N_5414,N_5007,N_5138);
nor U5415 (N_5415,N_5128,N_5003);
nor U5416 (N_5416,N_5002,N_5123);
xnor U5417 (N_5417,N_5086,N_5029);
xor U5418 (N_5418,N_5002,N_5016);
nor U5419 (N_5419,N_5234,N_5139);
or U5420 (N_5420,N_5084,N_5216);
or U5421 (N_5421,N_5008,N_5087);
xor U5422 (N_5422,N_5087,N_5086);
nand U5423 (N_5423,N_5154,N_5208);
nand U5424 (N_5424,N_5158,N_5042);
nand U5425 (N_5425,N_5013,N_5104);
and U5426 (N_5426,N_5010,N_5131);
nand U5427 (N_5427,N_5080,N_5166);
nor U5428 (N_5428,N_5097,N_5012);
nand U5429 (N_5429,N_5157,N_5133);
xor U5430 (N_5430,N_5156,N_5004);
nor U5431 (N_5431,N_5102,N_5201);
nand U5432 (N_5432,N_5225,N_5200);
and U5433 (N_5433,N_5249,N_5209);
nor U5434 (N_5434,N_5163,N_5123);
or U5435 (N_5435,N_5210,N_5085);
nor U5436 (N_5436,N_5221,N_5065);
and U5437 (N_5437,N_5118,N_5108);
or U5438 (N_5438,N_5038,N_5003);
and U5439 (N_5439,N_5157,N_5186);
and U5440 (N_5440,N_5049,N_5103);
nor U5441 (N_5441,N_5089,N_5129);
and U5442 (N_5442,N_5133,N_5195);
or U5443 (N_5443,N_5070,N_5145);
or U5444 (N_5444,N_5157,N_5228);
and U5445 (N_5445,N_5217,N_5052);
nand U5446 (N_5446,N_5052,N_5128);
nor U5447 (N_5447,N_5098,N_5160);
xnor U5448 (N_5448,N_5244,N_5059);
and U5449 (N_5449,N_5015,N_5114);
xor U5450 (N_5450,N_5077,N_5249);
nand U5451 (N_5451,N_5028,N_5052);
or U5452 (N_5452,N_5206,N_5149);
xnor U5453 (N_5453,N_5128,N_5217);
nand U5454 (N_5454,N_5194,N_5058);
xnor U5455 (N_5455,N_5205,N_5137);
and U5456 (N_5456,N_5195,N_5035);
or U5457 (N_5457,N_5030,N_5178);
nor U5458 (N_5458,N_5218,N_5071);
and U5459 (N_5459,N_5095,N_5062);
nor U5460 (N_5460,N_5001,N_5154);
xor U5461 (N_5461,N_5122,N_5055);
nor U5462 (N_5462,N_5142,N_5058);
or U5463 (N_5463,N_5089,N_5007);
xor U5464 (N_5464,N_5075,N_5043);
and U5465 (N_5465,N_5079,N_5119);
nor U5466 (N_5466,N_5038,N_5211);
or U5467 (N_5467,N_5149,N_5061);
xnor U5468 (N_5468,N_5200,N_5018);
nor U5469 (N_5469,N_5234,N_5117);
or U5470 (N_5470,N_5242,N_5139);
and U5471 (N_5471,N_5068,N_5021);
nand U5472 (N_5472,N_5062,N_5143);
xnor U5473 (N_5473,N_5093,N_5140);
nand U5474 (N_5474,N_5172,N_5106);
and U5475 (N_5475,N_5098,N_5132);
nand U5476 (N_5476,N_5075,N_5025);
nor U5477 (N_5477,N_5160,N_5159);
nor U5478 (N_5478,N_5039,N_5216);
nor U5479 (N_5479,N_5132,N_5145);
nand U5480 (N_5480,N_5181,N_5008);
nand U5481 (N_5481,N_5071,N_5074);
xnor U5482 (N_5482,N_5138,N_5052);
nor U5483 (N_5483,N_5163,N_5249);
or U5484 (N_5484,N_5130,N_5027);
nand U5485 (N_5485,N_5172,N_5125);
nand U5486 (N_5486,N_5064,N_5101);
xnor U5487 (N_5487,N_5217,N_5142);
and U5488 (N_5488,N_5092,N_5068);
xnor U5489 (N_5489,N_5214,N_5124);
or U5490 (N_5490,N_5208,N_5123);
nand U5491 (N_5491,N_5006,N_5038);
nor U5492 (N_5492,N_5009,N_5047);
and U5493 (N_5493,N_5081,N_5230);
nand U5494 (N_5494,N_5134,N_5239);
nor U5495 (N_5495,N_5150,N_5059);
and U5496 (N_5496,N_5125,N_5059);
xnor U5497 (N_5497,N_5212,N_5197);
nand U5498 (N_5498,N_5031,N_5054);
or U5499 (N_5499,N_5076,N_5221);
nor U5500 (N_5500,N_5329,N_5440);
or U5501 (N_5501,N_5393,N_5316);
or U5502 (N_5502,N_5277,N_5274);
or U5503 (N_5503,N_5463,N_5281);
or U5504 (N_5504,N_5388,N_5362);
nand U5505 (N_5505,N_5372,N_5443);
xor U5506 (N_5506,N_5264,N_5377);
nor U5507 (N_5507,N_5400,N_5498);
nor U5508 (N_5508,N_5252,N_5358);
or U5509 (N_5509,N_5475,N_5438);
and U5510 (N_5510,N_5477,N_5251);
or U5511 (N_5511,N_5413,N_5367);
xor U5512 (N_5512,N_5276,N_5387);
xnor U5513 (N_5513,N_5455,N_5320);
xnor U5514 (N_5514,N_5467,N_5315);
nand U5515 (N_5515,N_5352,N_5497);
and U5516 (N_5516,N_5254,N_5312);
nand U5517 (N_5517,N_5349,N_5479);
xor U5518 (N_5518,N_5426,N_5336);
and U5519 (N_5519,N_5285,N_5326);
xor U5520 (N_5520,N_5404,N_5442);
or U5521 (N_5521,N_5273,N_5271);
and U5522 (N_5522,N_5472,N_5476);
xnor U5523 (N_5523,N_5395,N_5392);
or U5524 (N_5524,N_5489,N_5366);
nand U5525 (N_5525,N_5257,N_5499);
and U5526 (N_5526,N_5373,N_5286);
nand U5527 (N_5527,N_5408,N_5494);
nor U5528 (N_5528,N_5363,N_5449);
and U5529 (N_5529,N_5385,N_5324);
nand U5530 (N_5530,N_5396,N_5347);
nand U5531 (N_5531,N_5275,N_5411);
xnor U5532 (N_5532,N_5290,N_5266);
nand U5533 (N_5533,N_5345,N_5348);
nand U5534 (N_5534,N_5343,N_5441);
or U5535 (N_5535,N_5350,N_5459);
and U5536 (N_5536,N_5323,N_5368);
and U5537 (N_5537,N_5485,N_5325);
and U5538 (N_5538,N_5268,N_5452);
nor U5539 (N_5539,N_5280,N_5296);
nand U5540 (N_5540,N_5436,N_5302);
xnor U5541 (N_5541,N_5383,N_5306);
and U5542 (N_5542,N_5311,N_5431);
xor U5543 (N_5543,N_5256,N_5425);
nand U5544 (N_5544,N_5424,N_5468);
and U5545 (N_5545,N_5305,N_5308);
xnor U5546 (N_5546,N_5356,N_5279);
xnor U5547 (N_5547,N_5297,N_5420);
nor U5548 (N_5548,N_5293,N_5483);
and U5549 (N_5549,N_5430,N_5374);
xnor U5550 (N_5550,N_5493,N_5351);
nor U5551 (N_5551,N_5407,N_5331);
nor U5552 (N_5552,N_5321,N_5454);
nand U5553 (N_5553,N_5355,N_5389);
or U5554 (N_5554,N_5429,N_5380);
nor U5555 (N_5555,N_5370,N_5282);
nor U5556 (N_5556,N_5284,N_5446);
or U5557 (N_5557,N_5381,N_5402);
nand U5558 (N_5558,N_5319,N_5287);
xor U5559 (N_5559,N_5405,N_5437);
nand U5560 (N_5560,N_5397,N_5342);
nand U5561 (N_5561,N_5416,N_5480);
or U5562 (N_5562,N_5469,N_5291);
or U5563 (N_5563,N_5435,N_5414);
nand U5564 (N_5564,N_5258,N_5341);
nor U5565 (N_5565,N_5327,N_5272);
or U5566 (N_5566,N_5394,N_5265);
and U5567 (N_5567,N_5482,N_5486);
or U5568 (N_5568,N_5300,N_5461);
nor U5569 (N_5569,N_5492,N_5322);
nand U5570 (N_5570,N_5354,N_5432);
nor U5571 (N_5571,N_5375,N_5371);
xnor U5572 (N_5572,N_5299,N_5295);
nor U5573 (N_5573,N_5401,N_5448);
nor U5574 (N_5574,N_5270,N_5445);
or U5575 (N_5575,N_5386,N_5376);
and U5576 (N_5576,N_5439,N_5317);
nor U5577 (N_5577,N_5384,N_5269);
nand U5578 (N_5578,N_5466,N_5487);
and U5579 (N_5579,N_5398,N_5481);
and U5580 (N_5580,N_5309,N_5382);
or U5581 (N_5581,N_5450,N_5457);
or U5582 (N_5582,N_5422,N_5412);
nor U5583 (N_5583,N_5250,N_5490);
nand U5584 (N_5584,N_5390,N_5346);
xnor U5585 (N_5585,N_5417,N_5267);
xnor U5586 (N_5586,N_5314,N_5460);
nor U5587 (N_5587,N_5318,N_5391);
or U5588 (N_5588,N_5337,N_5462);
nand U5589 (N_5589,N_5361,N_5263);
xor U5590 (N_5590,N_5334,N_5495);
nor U5591 (N_5591,N_5303,N_5427);
xnor U5592 (N_5592,N_5474,N_5338);
or U5593 (N_5593,N_5353,N_5419);
nand U5594 (N_5594,N_5288,N_5464);
or U5595 (N_5595,N_5340,N_5453);
and U5596 (N_5596,N_5360,N_5301);
xor U5597 (N_5597,N_5415,N_5434);
nand U5598 (N_5598,N_5458,N_5289);
nor U5599 (N_5599,N_5421,N_5339);
or U5600 (N_5600,N_5328,N_5488);
or U5601 (N_5601,N_5444,N_5473);
and U5602 (N_5602,N_5451,N_5478);
nand U5603 (N_5603,N_5409,N_5260);
xor U5604 (N_5604,N_5335,N_5310);
xor U5605 (N_5605,N_5294,N_5261);
xnor U5606 (N_5606,N_5304,N_5399);
or U5607 (N_5607,N_5379,N_5428);
or U5608 (N_5608,N_5253,N_5496);
or U5609 (N_5609,N_5357,N_5344);
nor U5610 (N_5610,N_5298,N_5491);
nor U5611 (N_5611,N_5406,N_5465);
and U5612 (N_5612,N_5278,N_5484);
xor U5613 (N_5613,N_5332,N_5471);
nand U5614 (N_5614,N_5292,N_5333);
and U5615 (N_5615,N_5313,N_5259);
and U5616 (N_5616,N_5447,N_5364);
and U5617 (N_5617,N_5456,N_5378);
or U5618 (N_5618,N_5283,N_5330);
or U5619 (N_5619,N_5403,N_5369);
or U5620 (N_5620,N_5418,N_5359);
xnor U5621 (N_5621,N_5307,N_5255);
nand U5622 (N_5622,N_5433,N_5423);
xor U5623 (N_5623,N_5365,N_5262);
nand U5624 (N_5624,N_5410,N_5470);
nand U5625 (N_5625,N_5494,N_5262);
nor U5626 (N_5626,N_5441,N_5391);
xnor U5627 (N_5627,N_5473,N_5312);
and U5628 (N_5628,N_5492,N_5377);
nand U5629 (N_5629,N_5487,N_5447);
nand U5630 (N_5630,N_5367,N_5443);
or U5631 (N_5631,N_5264,N_5410);
nor U5632 (N_5632,N_5381,N_5324);
or U5633 (N_5633,N_5370,N_5329);
nor U5634 (N_5634,N_5418,N_5481);
xnor U5635 (N_5635,N_5340,N_5439);
or U5636 (N_5636,N_5447,N_5302);
nand U5637 (N_5637,N_5447,N_5347);
or U5638 (N_5638,N_5270,N_5395);
nand U5639 (N_5639,N_5254,N_5447);
or U5640 (N_5640,N_5446,N_5448);
xor U5641 (N_5641,N_5292,N_5273);
or U5642 (N_5642,N_5433,N_5334);
or U5643 (N_5643,N_5350,N_5364);
and U5644 (N_5644,N_5461,N_5441);
and U5645 (N_5645,N_5478,N_5434);
nor U5646 (N_5646,N_5400,N_5446);
or U5647 (N_5647,N_5263,N_5464);
xnor U5648 (N_5648,N_5350,N_5305);
and U5649 (N_5649,N_5261,N_5350);
and U5650 (N_5650,N_5285,N_5363);
xnor U5651 (N_5651,N_5406,N_5482);
and U5652 (N_5652,N_5475,N_5337);
and U5653 (N_5653,N_5438,N_5373);
nor U5654 (N_5654,N_5349,N_5350);
and U5655 (N_5655,N_5498,N_5357);
or U5656 (N_5656,N_5320,N_5280);
and U5657 (N_5657,N_5334,N_5448);
nor U5658 (N_5658,N_5330,N_5302);
xnor U5659 (N_5659,N_5451,N_5300);
and U5660 (N_5660,N_5287,N_5410);
xor U5661 (N_5661,N_5421,N_5250);
xnor U5662 (N_5662,N_5447,N_5432);
nor U5663 (N_5663,N_5475,N_5425);
nor U5664 (N_5664,N_5373,N_5465);
nor U5665 (N_5665,N_5435,N_5473);
nor U5666 (N_5666,N_5392,N_5418);
and U5667 (N_5667,N_5262,N_5461);
and U5668 (N_5668,N_5444,N_5308);
and U5669 (N_5669,N_5263,N_5252);
nor U5670 (N_5670,N_5461,N_5452);
xnor U5671 (N_5671,N_5474,N_5436);
nor U5672 (N_5672,N_5275,N_5370);
and U5673 (N_5673,N_5295,N_5475);
xor U5674 (N_5674,N_5388,N_5421);
nor U5675 (N_5675,N_5294,N_5304);
or U5676 (N_5676,N_5395,N_5401);
and U5677 (N_5677,N_5282,N_5298);
xor U5678 (N_5678,N_5370,N_5292);
and U5679 (N_5679,N_5488,N_5449);
nand U5680 (N_5680,N_5408,N_5424);
xor U5681 (N_5681,N_5397,N_5339);
or U5682 (N_5682,N_5327,N_5489);
or U5683 (N_5683,N_5268,N_5481);
xor U5684 (N_5684,N_5359,N_5320);
or U5685 (N_5685,N_5322,N_5346);
nand U5686 (N_5686,N_5353,N_5493);
nor U5687 (N_5687,N_5360,N_5294);
nand U5688 (N_5688,N_5360,N_5261);
nand U5689 (N_5689,N_5368,N_5308);
xnor U5690 (N_5690,N_5318,N_5411);
xor U5691 (N_5691,N_5459,N_5396);
xor U5692 (N_5692,N_5277,N_5379);
and U5693 (N_5693,N_5286,N_5495);
xor U5694 (N_5694,N_5457,N_5264);
xnor U5695 (N_5695,N_5454,N_5463);
or U5696 (N_5696,N_5389,N_5483);
xor U5697 (N_5697,N_5472,N_5364);
and U5698 (N_5698,N_5269,N_5437);
xnor U5699 (N_5699,N_5409,N_5280);
or U5700 (N_5700,N_5356,N_5405);
xor U5701 (N_5701,N_5454,N_5362);
nand U5702 (N_5702,N_5278,N_5416);
xor U5703 (N_5703,N_5328,N_5282);
xnor U5704 (N_5704,N_5274,N_5370);
xnor U5705 (N_5705,N_5487,N_5334);
nor U5706 (N_5706,N_5298,N_5255);
nor U5707 (N_5707,N_5454,N_5469);
xnor U5708 (N_5708,N_5274,N_5331);
xnor U5709 (N_5709,N_5499,N_5443);
nand U5710 (N_5710,N_5418,N_5299);
xnor U5711 (N_5711,N_5471,N_5465);
or U5712 (N_5712,N_5262,N_5350);
or U5713 (N_5713,N_5431,N_5447);
or U5714 (N_5714,N_5435,N_5464);
xnor U5715 (N_5715,N_5265,N_5267);
nor U5716 (N_5716,N_5348,N_5264);
or U5717 (N_5717,N_5443,N_5305);
nor U5718 (N_5718,N_5281,N_5478);
xor U5719 (N_5719,N_5349,N_5297);
nor U5720 (N_5720,N_5283,N_5492);
and U5721 (N_5721,N_5455,N_5423);
or U5722 (N_5722,N_5262,N_5361);
or U5723 (N_5723,N_5298,N_5326);
nand U5724 (N_5724,N_5452,N_5340);
xor U5725 (N_5725,N_5333,N_5260);
nand U5726 (N_5726,N_5388,N_5489);
and U5727 (N_5727,N_5354,N_5491);
nand U5728 (N_5728,N_5259,N_5444);
and U5729 (N_5729,N_5429,N_5412);
or U5730 (N_5730,N_5416,N_5321);
and U5731 (N_5731,N_5312,N_5459);
nand U5732 (N_5732,N_5400,N_5416);
nand U5733 (N_5733,N_5394,N_5337);
xor U5734 (N_5734,N_5395,N_5309);
or U5735 (N_5735,N_5415,N_5315);
nor U5736 (N_5736,N_5386,N_5282);
xor U5737 (N_5737,N_5405,N_5333);
and U5738 (N_5738,N_5451,N_5450);
or U5739 (N_5739,N_5473,N_5362);
or U5740 (N_5740,N_5310,N_5497);
xnor U5741 (N_5741,N_5455,N_5322);
and U5742 (N_5742,N_5482,N_5457);
nor U5743 (N_5743,N_5256,N_5409);
and U5744 (N_5744,N_5368,N_5299);
nand U5745 (N_5745,N_5312,N_5286);
xor U5746 (N_5746,N_5461,N_5293);
or U5747 (N_5747,N_5262,N_5458);
nand U5748 (N_5748,N_5427,N_5361);
and U5749 (N_5749,N_5331,N_5420);
nor U5750 (N_5750,N_5628,N_5714);
nand U5751 (N_5751,N_5716,N_5705);
or U5752 (N_5752,N_5603,N_5747);
or U5753 (N_5753,N_5601,N_5561);
and U5754 (N_5754,N_5510,N_5579);
or U5755 (N_5755,N_5643,N_5547);
or U5756 (N_5756,N_5686,N_5504);
xor U5757 (N_5757,N_5653,N_5548);
or U5758 (N_5758,N_5597,N_5644);
nor U5759 (N_5759,N_5718,N_5719);
nand U5760 (N_5760,N_5632,N_5604);
nand U5761 (N_5761,N_5618,N_5540);
nor U5762 (N_5762,N_5542,N_5676);
nand U5763 (N_5763,N_5672,N_5622);
and U5764 (N_5764,N_5728,N_5515);
nand U5765 (N_5765,N_5683,N_5512);
nor U5766 (N_5766,N_5602,N_5577);
or U5767 (N_5767,N_5664,N_5661);
xnor U5768 (N_5768,N_5662,N_5563);
or U5769 (N_5769,N_5569,N_5582);
xor U5770 (N_5770,N_5551,N_5543);
nand U5771 (N_5771,N_5518,N_5648);
and U5772 (N_5772,N_5699,N_5568);
xor U5773 (N_5773,N_5655,N_5533);
nand U5774 (N_5774,N_5591,N_5641);
nor U5775 (N_5775,N_5634,N_5721);
or U5776 (N_5776,N_5558,N_5640);
and U5777 (N_5777,N_5535,N_5710);
and U5778 (N_5778,N_5685,N_5682);
nor U5779 (N_5779,N_5521,N_5649);
xor U5780 (N_5780,N_5516,N_5555);
xnor U5781 (N_5781,N_5593,N_5623);
and U5782 (N_5782,N_5595,N_5736);
and U5783 (N_5783,N_5616,N_5665);
nor U5784 (N_5784,N_5566,N_5578);
xnor U5785 (N_5785,N_5584,N_5530);
and U5786 (N_5786,N_5556,N_5654);
nand U5787 (N_5787,N_5658,N_5549);
or U5788 (N_5788,N_5734,N_5743);
and U5789 (N_5789,N_5608,N_5611);
and U5790 (N_5790,N_5739,N_5565);
nor U5791 (N_5791,N_5537,N_5738);
nor U5792 (N_5792,N_5712,N_5624);
or U5793 (N_5793,N_5646,N_5652);
or U5794 (N_5794,N_5633,N_5539);
nand U5795 (N_5795,N_5669,N_5717);
nor U5796 (N_5796,N_5694,N_5706);
nor U5797 (N_5797,N_5725,N_5726);
xnor U5798 (N_5798,N_5745,N_5749);
xnor U5799 (N_5799,N_5557,N_5687);
nor U5800 (N_5800,N_5528,N_5713);
and U5801 (N_5801,N_5519,N_5615);
xnor U5802 (N_5802,N_5677,N_5585);
nor U5803 (N_5803,N_5703,N_5627);
or U5804 (N_5804,N_5586,N_5552);
and U5805 (N_5805,N_5659,N_5681);
and U5806 (N_5806,N_5517,N_5746);
and U5807 (N_5807,N_5503,N_5571);
and U5808 (N_5808,N_5511,N_5607);
nand U5809 (N_5809,N_5554,N_5668);
and U5810 (N_5810,N_5570,N_5576);
nand U5811 (N_5811,N_5696,N_5700);
xor U5812 (N_5812,N_5625,N_5698);
or U5813 (N_5813,N_5724,N_5708);
nand U5814 (N_5814,N_5619,N_5574);
or U5815 (N_5815,N_5520,N_5567);
nand U5816 (N_5816,N_5707,N_5667);
nand U5817 (N_5817,N_5553,N_5651);
or U5818 (N_5818,N_5678,N_5740);
xor U5819 (N_5819,N_5513,N_5505);
and U5820 (N_5820,N_5580,N_5663);
xor U5821 (N_5821,N_5723,N_5671);
or U5822 (N_5822,N_5701,N_5502);
or U5823 (N_5823,N_5660,N_5729);
or U5824 (N_5824,N_5536,N_5524);
or U5825 (N_5825,N_5523,N_5605);
nor U5826 (N_5826,N_5656,N_5506);
and U5827 (N_5827,N_5732,N_5684);
or U5828 (N_5828,N_5610,N_5720);
nand U5829 (N_5829,N_5645,N_5629);
xor U5830 (N_5830,N_5722,N_5617);
or U5831 (N_5831,N_5500,N_5679);
or U5832 (N_5832,N_5709,N_5742);
xnor U5833 (N_5833,N_5748,N_5635);
nor U5834 (N_5834,N_5744,N_5650);
and U5835 (N_5835,N_5598,N_5638);
nand U5836 (N_5836,N_5509,N_5559);
xnor U5837 (N_5837,N_5546,N_5613);
nor U5838 (N_5838,N_5564,N_5702);
nand U5839 (N_5839,N_5639,N_5592);
nor U5840 (N_5840,N_5545,N_5733);
or U5841 (N_5841,N_5680,N_5606);
and U5842 (N_5842,N_5590,N_5689);
nor U5843 (N_5843,N_5507,N_5501);
xnor U5844 (N_5844,N_5614,N_5527);
xnor U5845 (N_5845,N_5531,N_5731);
nor U5846 (N_5846,N_5636,N_5538);
and U5847 (N_5847,N_5691,N_5673);
and U5848 (N_5848,N_5589,N_5514);
nor U5849 (N_5849,N_5508,N_5550);
nand U5850 (N_5850,N_5637,N_5572);
and U5851 (N_5851,N_5711,N_5599);
and U5852 (N_5852,N_5688,N_5541);
or U5853 (N_5853,N_5631,N_5544);
nand U5854 (N_5854,N_5692,N_5587);
xnor U5855 (N_5855,N_5596,N_5626);
and U5856 (N_5856,N_5612,N_5588);
nand U5857 (N_5857,N_5642,N_5609);
and U5858 (N_5858,N_5522,N_5573);
xnor U5859 (N_5859,N_5670,N_5675);
xor U5860 (N_5860,N_5737,N_5697);
xnor U5861 (N_5861,N_5560,N_5704);
nand U5862 (N_5862,N_5715,N_5693);
or U5863 (N_5863,N_5647,N_5657);
xor U5864 (N_5864,N_5562,N_5630);
or U5865 (N_5865,N_5526,N_5529);
nand U5866 (N_5866,N_5534,N_5575);
and U5867 (N_5867,N_5735,N_5674);
nor U5868 (N_5868,N_5600,N_5581);
nand U5869 (N_5869,N_5525,N_5695);
nor U5870 (N_5870,N_5730,N_5583);
and U5871 (N_5871,N_5666,N_5621);
or U5872 (N_5872,N_5620,N_5532);
xor U5873 (N_5873,N_5690,N_5594);
nand U5874 (N_5874,N_5727,N_5741);
xor U5875 (N_5875,N_5650,N_5563);
nand U5876 (N_5876,N_5664,N_5513);
xor U5877 (N_5877,N_5660,N_5634);
nor U5878 (N_5878,N_5676,N_5654);
and U5879 (N_5879,N_5534,N_5734);
nand U5880 (N_5880,N_5550,N_5668);
or U5881 (N_5881,N_5511,N_5691);
xor U5882 (N_5882,N_5606,N_5728);
xnor U5883 (N_5883,N_5681,N_5732);
xor U5884 (N_5884,N_5550,N_5642);
nor U5885 (N_5885,N_5523,N_5710);
or U5886 (N_5886,N_5606,N_5718);
xor U5887 (N_5887,N_5648,N_5699);
nor U5888 (N_5888,N_5605,N_5630);
xnor U5889 (N_5889,N_5698,N_5636);
and U5890 (N_5890,N_5724,N_5655);
nor U5891 (N_5891,N_5721,N_5603);
nor U5892 (N_5892,N_5525,N_5726);
and U5893 (N_5893,N_5725,N_5628);
and U5894 (N_5894,N_5598,N_5568);
and U5895 (N_5895,N_5739,N_5683);
xnor U5896 (N_5896,N_5561,N_5571);
xor U5897 (N_5897,N_5567,N_5694);
nand U5898 (N_5898,N_5604,N_5694);
xor U5899 (N_5899,N_5642,N_5624);
and U5900 (N_5900,N_5654,N_5543);
or U5901 (N_5901,N_5699,N_5640);
nor U5902 (N_5902,N_5629,N_5672);
xnor U5903 (N_5903,N_5713,N_5591);
nand U5904 (N_5904,N_5581,N_5737);
xnor U5905 (N_5905,N_5540,N_5578);
nand U5906 (N_5906,N_5697,N_5692);
or U5907 (N_5907,N_5522,N_5576);
nand U5908 (N_5908,N_5708,N_5590);
and U5909 (N_5909,N_5556,N_5738);
nor U5910 (N_5910,N_5520,N_5509);
or U5911 (N_5911,N_5699,N_5601);
nor U5912 (N_5912,N_5688,N_5571);
nand U5913 (N_5913,N_5618,N_5680);
or U5914 (N_5914,N_5613,N_5640);
or U5915 (N_5915,N_5589,N_5500);
and U5916 (N_5916,N_5659,N_5676);
or U5917 (N_5917,N_5566,N_5571);
xnor U5918 (N_5918,N_5564,N_5673);
xor U5919 (N_5919,N_5628,N_5596);
nor U5920 (N_5920,N_5670,N_5734);
nor U5921 (N_5921,N_5633,N_5715);
nand U5922 (N_5922,N_5667,N_5622);
and U5923 (N_5923,N_5564,N_5654);
and U5924 (N_5924,N_5741,N_5695);
xnor U5925 (N_5925,N_5507,N_5586);
and U5926 (N_5926,N_5710,N_5542);
xnor U5927 (N_5927,N_5684,N_5663);
xnor U5928 (N_5928,N_5566,N_5510);
or U5929 (N_5929,N_5692,N_5630);
nor U5930 (N_5930,N_5713,N_5619);
and U5931 (N_5931,N_5567,N_5742);
and U5932 (N_5932,N_5630,N_5699);
or U5933 (N_5933,N_5718,N_5509);
and U5934 (N_5934,N_5731,N_5622);
xnor U5935 (N_5935,N_5662,N_5607);
nor U5936 (N_5936,N_5735,N_5550);
nor U5937 (N_5937,N_5590,N_5548);
xnor U5938 (N_5938,N_5617,N_5606);
or U5939 (N_5939,N_5697,N_5585);
nand U5940 (N_5940,N_5636,N_5609);
nor U5941 (N_5941,N_5748,N_5693);
nor U5942 (N_5942,N_5683,N_5678);
nor U5943 (N_5943,N_5687,N_5733);
nand U5944 (N_5944,N_5600,N_5611);
or U5945 (N_5945,N_5638,N_5578);
or U5946 (N_5946,N_5574,N_5715);
xor U5947 (N_5947,N_5634,N_5713);
and U5948 (N_5948,N_5512,N_5511);
nand U5949 (N_5949,N_5592,N_5515);
nand U5950 (N_5950,N_5690,N_5544);
or U5951 (N_5951,N_5506,N_5700);
nor U5952 (N_5952,N_5658,N_5570);
nor U5953 (N_5953,N_5634,N_5700);
or U5954 (N_5954,N_5557,N_5748);
and U5955 (N_5955,N_5648,N_5659);
or U5956 (N_5956,N_5689,N_5554);
or U5957 (N_5957,N_5532,N_5719);
nor U5958 (N_5958,N_5735,N_5702);
xnor U5959 (N_5959,N_5537,N_5530);
nand U5960 (N_5960,N_5609,N_5718);
or U5961 (N_5961,N_5600,N_5617);
or U5962 (N_5962,N_5657,N_5519);
and U5963 (N_5963,N_5671,N_5524);
nand U5964 (N_5964,N_5736,N_5502);
and U5965 (N_5965,N_5522,N_5736);
nand U5966 (N_5966,N_5681,N_5677);
nand U5967 (N_5967,N_5538,N_5734);
and U5968 (N_5968,N_5742,N_5636);
nor U5969 (N_5969,N_5541,N_5538);
and U5970 (N_5970,N_5539,N_5598);
and U5971 (N_5971,N_5688,N_5648);
xnor U5972 (N_5972,N_5736,N_5662);
or U5973 (N_5973,N_5501,N_5656);
xor U5974 (N_5974,N_5646,N_5533);
nand U5975 (N_5975,N_5584,N_5679);
or U5976 (N_5976,N_5626,N_5570);
nor U5977 (N_5977,N_5734,N_5668);
or U5978 (N_5978,N_5715,N_5615);
nor U5979 (N_5979,N_5736,N_5704);
nor U5980 (N_5980,N_5689,N_5664);
xor U5981 (N_5981,N_5536,N_5529);
nor U5982 (N_5982,N_5560,N_5642);
and U5983 (N_5983,N_5621,N_5534);
nand U5984 (N_5984,N_5687,N_5610);
nor U5985 (N_5985,N_5593,N_5701);
and U5986 (N_5986,N_5629,N_5554);
nand U5987 (N_5987,N_5502,N_5644);
nor U5988 (N_5988,N_5569,N_5519);
nand U5989 (N_5989,N_5683,N_5575);
xor U5990 (N_5990,N_5599,N_5680);
nor U5991 (N_5991,N_5555,N_5517);
and U5992 (N_5992,N_5591,N_5647);
or U5993 (N_5993,N_5530,N_5679);
xor U5994 (N_5994,N_5655,N_5526);
nand U5995 (N_5995,N_5708,N_5561);
xnor U5996 (N_5996,N_5570,N_5516);
and U5997 (N_5997,N_5621,N_5604);
or U5998 (N_5998,N_5576,N_5558);
nor U5999 (N_5999,N_5600,N_5642);
nor U6000 (N_6000,N_5826,N_5972);
xor U6001 (N_6001,N_5994,N_5815);
and U6002 (N_6002,N_5985,N_5997);
nor U6003 (N_6003,N_5772,N_5872);
or U6004 (N_6004,N_5845,N_5974);
xnor U6005 (N_6005,N_5860,N_5912);
and U6006 (N_6006,N_5876,N_5906);
and U6007 (N_6007,N_5907,N_5802);
nor U6008 (N_6008,N_5920,N_5937);
xnor U6009 (N_6009,N_5883,N_5797);
xor U6010 (N_6010,N_5840,N_5804);
and U6011 (N_6011,N_5889,N_5771);
or U6012 (N_6012,N_5969,N_5773);
nand U6013 (N_6013,N_5793,N_5824);
or U6014 (N_6014,N_5759,N_5975);
and U6015 (N_6015,N_5885,N_5816);
or U6016 (N_6016,N_5808,N_5925);
nand U6017 (N_6017,N_5904,N_5818);
nand U6018 (N_6018,N_5962,N_5943);
nand U6019 (N_6019,N_5865,N_5813);
nand U6020 (N_6020,N_5799,N_5891);
xor U6021 (N_6021,N_5774,N_5950);
nand U6022 (N_6022,N_5814,N_5961);
xnor U6023 (N_6023,N_5896,N_5981);
xnor U6024 (N_6024,N_5977,N_5778);
xor U6025 (N_6025,N_5834,N_5982);
nor U6026 (N_6026,N_5916,N_5780);
nor U6027 (N_6027,N_5957,N_5949);
nor U6028 (N_6028,N_5871,N_5867);
or U6029 (N_6029,N_5991,N_5837);
nand U6030 (N_6030,N_5788,N_5852);
xnor U6031 (N_6031,N_5844,N_5958);
xnor U6032 (N_6032,N_5767,N_5864);
nand U6033 (N_6033,N_5944,N_5953);
nand U6034 (N_6034,N_5888,N_5817);
and U6035 (N_6035,N_5850,N_5785);
and U6036 (N_6036,N_5890,N_5929);
or U6037 (N_6037,N_5976,N_5805);
xor U6038 (N_6038,N_5849,N_5789);
nor U6039 (N_6039,N_5870,N_5938);
or U6040 (N_6040,N_5952,N_5819);
or U6041 (N_6041,N_5931,N_5971);
or U6042 (N_6042,N_5756,N_5866);
or U6043 (N_6043,N_5956,N_5966);
or U6044 (N_6044,N_5884,N_5963);
and U6045 (N_6045,N_5859,N_5783);
or U6046 (N_6046,N_5893,N_5915);
nor U6047 (N_6047,N_5921,N_5766);
xor U6048 (N_6048,N_5758,N_5892);
nor U6049 (N_6049,N_5954,N_5782);
or U6050 (N_6050,N_5869,N_5959);
and U6051 (N_6051,N_5762,N_5894);
and U6052 (N_6052,N_5903,N_5847);
or U6053 (N_6053,N_5951,N_5830);
nor U6054 (N_6054,N_5911,N_5812);
nand U6055 (N_6055,N_5790,N_5923);
xnor U6056 (N_6056,N_5993,N_5828);
and U6057 (N_6057,N_5947,N_5922);
nor U6058 (N_6058,N_5902,N_5820);
nand U6059 (N_6059,N_5935,N_5996);
xnor U6060 (N_6060,N_5900,N_5768);
xor U6061 (N_6061,N_5980,N_5833);
nand U6062 (N_6062,N_5765,N_5861);
xor U6063 (N_6063,N_5795,N_5887);
or U6064 (N_6064,N_5965,N_5913);
xor U6065 (N_6065,N_5933,N_5809);
nand U6066 (N_6066,N_5851,N_5945);
and U6067 (N_6067,N_5946,N_5770);
and U6068 (N_6068,N_5811,N_5978);
xnor U6069 (N_6069,N_5769,N_5881);
nor U6070 (N_6070,N_5886,N_5761);
xnor U6071 (N_6071,N_5853,N_5827);
nand U6072 (N_6072,N_5763,N_5800);
or U6073 (N_6073,N_5939,N_5908);
or U6074 (N_6074,N_5968,N_5786);
xor U6075 (N_6075,N_5750,N_5899);
nor U6076 (N_6076,N_5995,N_5926);
nand U6077 (N_6077,N_5858,N_5901);
and U6078 (N_6078,N_5843,N_5874);
xor U6079 (N_6079,N_5753,N_5989);
nor U6080 (N_6080,N_5835,N_5999);
nor U6081 (N_6081,N_5895,N_5764);
nor U6082 (N_6082,N_5964,N_5777);
or U6083 (N_6083,N_5787,N_5807);
nor U6084 (N_6084,N_5781,N_5948);
nand U6085 (N_6085,N_5910,N_5846);
nor U6086 (N_6086,N_5988,N_5941);
xor U6087 (N_6087,N_5942,N_5897);
xor U6088 (N_6088,N_5751,N_5822);
or U6089 (N_6089,N_5979,N_5936);
or U6090 (N_6090,N_5986,N_5810);
nand U6091 (N_6091,N_5854,N_5905);
xnor U6092 (N_6092,N_5967,N_5877);
or U6093 (N_6093,N_5924,N_5868);
xnor U6094 (N_6094,N_5779,N_5841);
or U6095 (N_6095,N_5882,N_5878);
nand U6096 (N_6096,N_5960,N_5970);
xor U6097 (N_6097,N_5825,N_5776);
xnor U6098 (N_6098,N_5990,N_5752);
nor U6099 (N_6099,N_5919,N_5839);
xor U6100 (N_6100,N_5998,N_5940);
nor U6101 (N_6101,N_5879,N_5775);
and U6102 (N_6102,N_5898,N_5757);
nor U6103 (N_6103,N_5928,N_5798);
or U6104 (N_6104,N_5984,N_5842);
xnor U6105 (N_6105,N_5875,N_5909);
or U6106 (N_6106,N_5856,N_5792);
and U6107 (N_6107,N_5932,N_5927);
nor U6108 (N_6108,N_5857,N_5755);
nand U6109 (N_6109,N_5801,N_5832);
nand U6110 (N_6110,N_5855,N_5829);
or U6111 (N_6111,N_5880,N_5930);
nand U6112 (N_6112,N_5873,N_5803);
nand U6113 (N_6113,N_5983,N_5823);
nand U6114 (N_6114,N_5838,N_5918);
nand U6115 (N_6115,N_5955,N_5862);
and U6116 (N_6116,N_5987,N_5796);
or U6117 (N_6117,N_5754,N_5784);
nor U6118 (N_6118,N_5760,N_5848);
nand U6119 (N_6119,N_5794,N_5831);
xnor U6120 (N_6120,N_5821,N_5917);
nand U6121 (N_6121,N_5973,N_5914);
nor U6122 (N_6122,N_5836,N_5992);
xor U6123 (N_6123,N_5806,N_5791);
xor U6124 (N_6124,N_5934,N_5863);
and U6125 (N_6125,N_5832,N_5999);
nand U6126 (N_6126,N_5984,N_5855);
nand U6127 (N_6127,N_5846,N_5752);
nand U6128 (N_6128,N_5944,N_5937);
nor U6129 (N_6129,N_5829,N_5807);
and U6130 (N_6130,N_5958,N_5995);
xnor U6131 (N_6131,N_5884,N_5752);
xnor U6132 (N_6132,N_5915,N_5932);
nor U6133 (N_6133,N_5865,N_5855);
nor U6134 (N_6134,N_5994,N_5774);
xnor U6135 (N_6135,N_5856,N_5942);
and U6136 (N_6136,N_5819,N_5999);
nand U6137 (N_6137,N_5938,N_5806);
and U6138 (N_6138,N_5968,N_5808);
or U6139 (N_6139,N_5767,N_5831);
xor U6140 (N_6140,N_5787,N_5917);
nor U6141 (N_6141,N_5924,N_5968);
xor U6142 (N_6142,N_5946,N_5780);
nor U6143 (N_6143,N_5972,N_5750);
or U6144 (N_6144,N_5873,N_5842);
xor U6145 (N_6145,N_5801,N_5843);
xnor U6146 (N_6146,N_5849,N_5819);
nor U6147 (N_6147,N_5865,N_5759);
nand U6148 (N_6148,N_5929,N_5834);
xnor U6149 (N_6149,N_5900,N_5821);
or U6150 (N_6150,N_5766,N_5758);
xnor U6151 (N_6151,N_5752,N_5861);
xor U6152 (N_6152,N_5910,N_5915);
nor U6153 (N_6153,N_5771,N_5983);
xor U6154 (N_6154,N_5965,N_5967);
xor U6155 (N_6155,N_5897,N_5829);
or U6156 (N_6156,N_5928,N_5960);
nor U6157 (N_6157,N_5932,N_5973);
or U6158 (N_6158,N_5981,N_5952);
nand U6159 (N_6159,N_5786,N_5847);
and U6160 (N_6160,N_5936,N_5889);
or U6161 (N_6161,N_5921,N_5959);
and U6162 (N_6162,N_5913,N_5782);
xor U6163 (N_6163,N_5969,N_5975);
and U6164 (N_6164,N_5916,N_5920);
nor U6165 (N_6165,N_5845,N_5892);
nor U6166 (N_6166,N_5832,N_5866);
and U6167 (N_6167,N_5977,N_5804);
or U6168 (N_6168,N_5902,N_5920);
xor U6169 (N_6169,N_5897,N_5826);
or U6170 (N_6170,N_5913,N_5905);
or U6171 (N_6171,N_5914,N_5988);
xnor U6172 (N_6172,N_5945,N_5828);
nand U6173 (N_6173,N_5772,N_5965);
xor U6174 (N_6174,N_5929,N_5985);
or U6175 (N_6175,N_5825,N_5945);
nor U6176 (N_6176,N_5840,N_5918);
nor U6177 (N_6177,N_5948,N_5844);
nand U6178 (N_6178,N_5967,N_5780);
and U6179 (N_6179,N_5966,N_5867);
or U6180 (N_6180,N_5797,N_5993);
xnor U6181 (N_6181,N_5952,N_5919);
xnor U6182 (N_6182,N_5791,N_5840);
and U6183 (N_6183,N_5894,N_5795);
or U6184 (N_6184,N_5761,N_5929);
nor U6185 (N_6185,N_5977,N_5992);
nand U6186 (N_6186,N_5829,N_5903);
nor U6187 (N_6187,N_5765,N_5907);
and U6188 (N_6188,N_5903,N_5930);
xor U6189 (N_6189,N_5851,N_5984);
nor U6190 (N_6190,N_5840,N_5829);
or U6191 (N_6191,N_5910,N_5902);
nand U6192 (N_6192,N_5995,N_5908);
xnor U6193 (N_6193,N_5908,N_5946);
nor U6194 (N_6194,N_5867,N_5888);
and U6195 (N_6195,N_5773,N_5884);
nor U6196 (N_6196,N_5984,N_5870);
and U6197 (N_6197,N_5840,N_5790);
or U6198 (N_6198,N_5982,N_5763);
and U6199 (N_6199,N_5909,N_5771);
xnor U6200 (N_6200,N_5871,N_5927);
nand U6201 (N_6201,N_5914,N_5875);
or U6202 (N_6202,N_5812,N_5983);
and U6203 (N_6203,N_5988,N_5962);
nor U6204 (N_6204,N_5883,N_5838);
or U6205 (N_6205,N_5802,N_5904);
and U6206 (N_6206,N_5841,N_5973);
nand U6207 (N_6207,N_5795,N_5984);
and U6208 (N_6208,N_5932,N_5993);
nor U6209 (N_6209,N_5989,N_5986);
nand U6210 (N_6210,N_5951,N_5842);
nor U6211 (N_6211,N_5903,N_5897);
or U6212 (N_6212,N_5849,N_5899);
xnor U6213 (N_6213,N_5805,N_5958);
nor U6214 (N_6214,N_5894,N_5938);
nand U6215 (N_6215,N_5923,N_5910);
and U6216 (N_6216,N_5893,N_5763);
or U6217 (N_6217,N_5778,N_5938);
or U6218 (N_6218,N_5762,N_5917);
nand U6219 (N_6219,N_5771,N_5961);
or U6220 (N_6220,N_5850,N_5977);
nor U6221 (N_6221,N_5853,N_5839);
and U6222 (N_6222,N_5823,N_5921);
or U6223 (N_6223,N_5750,N_5943);
or U6224 (N_6224,N_5877,N_5837);
nand U6225 (N_6225,N_5795,N_5780);
or U6226 (N_6226,N_5985,N_5944);
xor U6227 (N_6227,N_5837,N_5791);
xor U6228 (N_6228,N_5761,N_5999);
and U6229 (N_6229,N_5877,N_5920);
and U6230 (N_6230,N_5962,N_5874);
xnor U6231 (N_6231,N_5774,N_5963);
nor U6232 (N_6232,N_5856,N_5842);
nor U6233 (N_6233,N_5867,N_5799);
xor U6234 (N_6234,N_5983,N_5961);
and U6235 (N_6235,N_5989,N_5917);
xnor U6236 (N_6236,N_5896,N_5906);
and U6237 (N_6237,N_5782,N_5937);
nand U6238 (N_6238,N_5914,N_5989);
and U6239 (N_6239,N_5885,N_5904);
xor U6240 (N_6240,N_5806,N_5941);
and U6241 (N_6241,N_5921,N_5883);
xor U6242 (N_6242,N_5909,N_5984);
or U6243 (N_6243,N_5800,N_5881);
nand U6244 (N_6244,N_5912,N_5772);
nor U6245 (N_6245,N_5830,N_5985);
nor U6246 (N_6246,N_5809,N_5876);
nor U6247 (N_6247,N_5929,N_5910);
xnor U6248 (N_6248,N_5987,N_5885);
nor U6249 (N_6249,N_5866,N_5953);
or U6250 (N_6250,N_6092,N_6086);
or U6251 (N_6251,N_6084,N_6141);
nand U6252 (N_6252,N_6157,N_6011);
nor U6253 (N_6253,N_6033,N_6179);
or U6254 (N_6254,N_6211,N_6074);
or U6255 (N_6255,N_6122,N_6216);
xor U6256 (N_6256,N_6151,N_6055);
nor U6257 (N_6257,N_6109,N_6002);
or U6258 (N_6258,N_6104,N_6144);
nand U6259 (N_6259,N_6045,N_6110);
or U6260 (N_6260,N_6245,N_6191);
nor U6261 (N_6261,N_6244,N_6215);
nor U6262 (N_6262,N_6066,N_6154);
xor U6263 (N_6263,N_6003,N_6108);
or U6264 (N_6264,N_6030,N_6209);
or U6265 (N_6265,N_6016,N_6146);
nand U6266 (N_6266,N_6249,N_6035);
and U6267 (N_6267,N_6198,N_6130);
and U6268 (N_6268,N_6168,N_6203);
or U6269 (N_6269,N_6170,N_6153);
or U6270 (N_6270,N_6222,N_6037);
nand U6271 (N_6271,N_6043,N_6004);
nor U6272 (N_6272,N_6202,N_6226);
or U6273 (N_6273,N_6248,N_6132);
or U6274 (N_6274,N_6046,N_6021);
or U6275 (N_6275,N_6199,N_6161);
or U6276 (N_6276,N_6178,N_6176);
and U6277 (N_6277,N_6220,N_6050);
xor U6278 (N_6278,N_6128,N_6026);
nand U6279 (N_6279,N_6027,N_6242);
xor U6280 (N_6280,N_6081,N_6177);
or U6281 (N_6281,N_6113,N_6166);
xor U6282 (N_6282,N_6133,N_6064);
and U6283 (N_6283,N_6195,N_6227);
nor U6284 (N_6284,N_6228,N_6075);
nand U6285 (N_6285,N_6067,N_6038);
or U6286 (N_6286,N_6138,N_6159);
and U6287 (N_6287,N_6029,N_6208);
or U6288 (N_6288,N_6160,N_6097);
and U6289 (N_6289,N_6156,N_6241);
or U6290 (N_6290,N_6076,N_6047);
xnor U6291 (N_6291,N_6167,N_6082);
or U6292 (N_6292,N_6096,N_6193);
xor U6293 (N_6293,N_6012,N_6162);
or U6294 (N_6294,N_6182,N_6186);
nor U6295 (N_6295,N_6148,N_6196);
nor U6296 (N_6296,N_6124,N_6164);
xnor U6297 (N_6297,N_6225,N_6083);
nand U6298 (N_6298,N_6210,N_6140);
nand U6299 (N_6299,N_6173,N_6224);
nor U6300 (N_6300,N_6219,N_6247);
xor U6301 (N_6301,N_6185,N_6078);
and U6302 (N_6302,N_6090,N_6013);
and U6303 (N_6303,N_6042,N_6152);
xnor U6304 (N_6304,N_6040,N_6201);
nor U6305 (N_6305,N_6031,N_6136);
nand U6306 (N_6306,N_6054,N_6213);
and U6307 (N_6307,N_6184,N_6022);
xnor U6308 (N_6308,N_6005,N_6073);
xnor U6309 (N_6309,N_6006,N_6231);
xnor U6310 (N_6310,N_6172,N_6024);
or U6311 (N_6311,N_6181,N_6023);
nand U6312 (N_6312,N_6014,N_6150);
nand U6313 (N_6313,N_6008,N_6165);
and U6314 (N_6314,N_6062,N_6189);
xor U6315 (N_6315,N_6127,N_6072);
and U6316 (N_6316,N_6137,N_6221);
and U6317 (N_6317,N_6180,N_6129);
or U6318 (N_6318,N_6095,N_6143);
xnor U6319 (N_6319,N_6060,N_6218);
xor U6320 (N_6320,N_6106,N_6183);
nor U6321 (N_6321,N_6036,N_6206);
nand U6322 (N_6322,N_6214,N_6102);
nor U6323 (N_6323,N_6171,N_6069);
nor U6324 (N_6324,N_6053,N_6194);
nor U6325 (N_6325,N_6119,N_6085);
or U6326 (N_6326,N_6229,N_6020);
nand U6327 (N_6327,N_6238,N_6116);
nand U6328 (N_6328,N_6091,N_6028);
xor U6329 (N_6329,N_6117,N_6175);
nand U6330 (N_6330,N_6099,N_6158);
xor U6331 (N_6331,N_6058,N_6061);
nor U6332 (N_6332,N_6115,N_6098);
nor U6333 (N_6333,N_6131,N_6192);
or U6334 (N_6334,N_6240,N_6243);
nand U6335 (N_6335,N_6039,N_6212);
or U6336 (N_6336,N_6080,N_6049);
xnor U6337 (N_6337,N_6155,N_6123);
xor U6338 (N_6338,N_6089,N_6112);
or U6339 (N_6339,N_6190,N_6057);
and U6340 (N_6340,N_6139,N_6149);
xor U6341 (N_6341,N_6032,N_6163);
and U6342 (N_6342,N_6125,N_6087);
nor U6343 (N_6343,N_6048,N_6235);
and U6344 (N_6344,N_6114,N_6007);
or U6345 (N_6345,N_6105,N_6118);
or U6346 (N_6346,N_6111,N_6134);
nand U6347 (N_6347,N_6010,N_6056);
nor U6348 (N_6348,N_6088,N_6217);
xnor U6349 (N_6349,N_6174,N_6051);
xor U6350 (N_6350,N_6093,N_6120);
nand U6351 (N_6351,N_6052,N_6207);
xor U6352 (N_6352,N_6200,N_6001);
xor U6353 (N_6353,N_6009,N_6041);
nand U6354 (N_6354,N_6236,N_6100);
nor U6355 (N_6355,N_6018,N_6232);
nor U6356 (N_6356,N_6188,N_6063);
xor U6357 (N_6357,N_6187,N_6142);
nor U6358 (N_6358,N_6103,N_6234);
nor U6359 (N_6359,N_6147,N_6107);
xor U6360 (N_6360,N_6121,N_6017);
or U6361 (N_6361,N_6233,N_6019);
and U6362 (N_6362,N_6094,N_6204);
or U6363 (N_6363,N_6065,N_6135);
or U6364 (N_6364,N_6077,N_6079);
or U6365 (N_6365,N_6071,N_6025);
or U6366 (N_6366,N_6070,N_6101);
nand U6367 (N_6367,N_6015,N_6000);
or U6368 (N_6368,N_6246,N_6145);
xor U6369 (N_6369,N_6126,N_6223);
nand U6370 (N_6370,N_6169,N_6237);
xnor U6371 (N_6371,N_6230,N_6197);
nand U6372 (N_6372,N_6059,N_6034);
xnor U6373 (N_6373,N_6239,N_6068);
nand U6374 (N_6374,N_6044,N_6205);
and U6375 (N_6375,N_6155,N_6032);
and U6376 (N_6376,N_6029,N_6118);
nand U6377 (N_6377,N_6234,N_6201);
nor U6378 (N_6378,N_6116,N_6163);
and U6379 (N_6379,N_6187,N_6123);
or U6380 (N_6380,N_6040,N_6022);
xnor U6381 (N_6381,N_6249,N_6010);
nand U6382 (N_6382,N_6080,N_6113);
xnor U6383 (N_6383,N_6194,N_6091);
or U6384 (N_6384,N_6149,N_6204);
or U6385 (N_6385,N_6068,N_6187);
nor U6386 (N_6386,N_6136,N_6154);
nand U6387 (N_6387,N_6014,N_6079);
or U6388 (N_6388,N_6056,N_6058);
and U6389 (N_6389,N_6063,N_6246);
and U6390 (N_6390,N_6109,N_6102);
nand U6391 (N_6391,N_6085,N_6144);
or U6392 (N_6392,N_6206,N_6021);
and U6393 (N_6393,N_6071,N_6092);
nor U6394 (N_6394,N_6081,N_6143);
xnor U6395 (N_6395,N_6073,N_6132);
or U6396 (N_6396,N_6230,N_6165);
nor U6397 (N_6397,N_6189,N_6012);
or U6398 (N_6398,N_6106,N_6002);
nor U6399 (N_6399,N_6181,N_6092);
nor U6400 (N_6400,N_6016,N_6149);
xor U6401 (N_6401,N_6150,N_6000);
and U6402 (N_6402,N_6171,N_6224);
nand U6403 (N_6403,N_6175,N_6106);
or U6404 (N_6404,N_6184,N_6144);
nor U6405 (N_6405,N_6203,N_6217);
and U6406 (N_6406,N_6123,N_6066);
nand U6407 (N_6407,N_6189,N_6144);
nand U6408 (N_6408,N_6034,N_6011);
nor U6409 (N_6409,N_6210,N_6016);
or U6410 (N_6410,N_6213,N_6158);
or U6411 (N_6411,N_6152,N_6173);
xor U6412 (N_6412,N_6010,N_6018);
or U6413 (N_6413,N_6195,N_6072);
or U6414 (N_6414,N_6080,N_6199);
or U6415 (N_6415,N_6022,N_6079);
nand U6416 (N_6416,N_6247,N_6013);
nor U6417 (N_6417,N_6118,N_6021);
or U6418 (N_6418,N_6191,N_6152);
or U6419 (N_6419,N_6165,N_6236);
nor U6420 (N_6420,N_6157,N_6010);
or U6421 (N_6421,N_6144,N_6187);
xnor U6422 (N_6422,N_6070,N_6172);
and U6423 (N_6423,N_6183,N_6152);
nor U6424 (N_6424,N_6170,N_6084);
and U6425 (N_6425,N_6247,N_6023);
nand U6426 (N_6426,N_6144,N_6006);
xnor U6427 (N_6427,N_6004,N_6208);
nor U6428 (N_6428,N_6240,N_6124);
nand U6429 (N_6429,N_6023,N_6232);
nor U6430 (N_6430,N_6040,N_6224);
nor U6431 (N_6431,N_6116,N_6241);
xor U6432 (N_6432,N_6078,N_6172);
and U6433 (N_6433,N_6060,N_6131);
and U6434 (N_6434,N_6130,N_6063);
xor U6435 (N_6435,N_6101,N_6213);
nand U6436 (N_6436,N_6206,N_6078);
nand U6437 (N_6437,N_6040,N_6163);
xor U6438 (N_6438,N_6181,N_6172);
and U6439 (N_6439,N_6108,N_6096);
nor U6440 (N_6440,N_6017,N_6183);
and U6441 (N_6441,N_6004,N_6166);
and U6442 (N_6442,N_6022,N_6055);
nand U6443 (N_6443,N_6151,N_6060);
or U6444 (N_6444,N_6080,N_6135);
nand U6445 (N_6445,N_6002,N_6086);
nand U6446 (N_6446,N_6000,N_6104);
nor U6447 (N_6447,N_6106,N_6243);
or U6448 (N_6448,N_6182,N_6011);
or U6449 (N_6449,N_6079,N_6233);
nor U6450 (N_6450,N_6155,N_6172);
xnor U6451 (N_6451,N_6059,N_6242);
nor U6452 (N_6452,N_6221,N_6143);
or U6453 (N_6453,N_6201,N_6153);
nand U6454 (N_6454,N_6143,N_6135);
xor U6455 (N_6455,N_6153,N_6093);
xor U6456 (N_6456,N_6081,N_6153);
or U6457 (N_6457,N_6202,N_6215);
or U6458 (N_6458,N_6116,N_6199);
xnor U6459 (N_6459,N_6144,N_6202);
or U6460 (N_6460,N_6049,N_6092);
nand U6461 (N_6461,N_6012,N_6221);
or U6462 (N_6462,N_6107,N_6183);
xor U6463 (N_6463,N_6043,N_6185);
xnor U6464 (N_6464,N_6226,N_6223);
and U6465 (N_6465,N_6120,N_6091);
xnor U6466 (N_6466,N_6185,N_6109);
nor U6467 (N_6467,N_6119,N_6104);
nor U6468 (N_6468,N_6023,N_6218);
nand U6469 (N_6469,N_6069,N_6025);
and U6470 (N_6470,N_6110,N_6000);
and U6471 (N_6471,N_6037,N_6210);
nand U6472 (N_6472,N_6122,N_6003);
nand U6473 (N_6473,N_6062,N_6100);
nand U6474 (N_6474,N_6120,N_6045);
or U6475 (N_6475,N_6088,N_6056);
and U6476 (N_6476,N_6153,N_6135);
or U6477 (N_6477,N_6197,N_6108);
xnor U6478 (N_6478,N_6015,N_6006);
or U6479 (N_6479,N_6039,N_6144);
and U6480 (N_6480,N_6239,N_6082);
xnor U6481 (N_6481,N_6029,N_6238);
or U6482 (N_6482,N_6077,N_6226);
nor U6483 (N_6483,N_6032,N_6135);
nand U6484 (N_6484,N_6167,N_6221);
nor U6485 (N_6485,N_6071,N_6121);
or U6486 (N_6486,N_6162,N_6218);
nor U6487 (N_6487,N_6118,N_6035);
xnor U6488 (N_6488,N_6150,N_6121);
nand U6489 (N_6489,N_6214,N_6233);
or U6490 (N_6490,N_6104,N_6041);
nor U6491 (N_6491,N_6077,N_6214);
nand U6492 (N_6492,N_6106,N_6132);
xor U6493 (N_6493,N_6068,N_6096);
and U6494 (N_6494,N_6004,N_6200);
nor U6495 (N_6495,N_6093,N_6019);
nand U6496 (N_6496,N_6118,N_6038);
nor U6497 (N_6497,N_6164,N_6240);
xor U6498 (N_6498,N_6162,N_6198);
nand U6499 (N_6499,N_6199,N_6052);
xor U6500 (N_6500,N_6470,N_6328);
or U6501 (N_6501,N_6451,N_6413);
nand U6502 (N_6502,N_6344,N_6392);
or U6503 (N_6503,N_6296,N_6271);
nor U6504 (N_6504,N_6486,N_6410);
nor U6505 (N_6505,N_6387,N_6313);
or U6506 (N_6506,N_6363,N_6411);
or U6507 (N_6507,N_6304,N_6311);
xor U6508 (N_6508,N_6417,N_6260);
nand U6509 (N_6509,N_6258,N_6330);
or U6510 (N_6510,N_6341,N_6376);
or U6511 (N_6511,N_6444,N_6337);
and U6512 (N_6512,N_6397,N_6450);
nor U6513 (N_6513,N_6400,N_6358);
and U6514 (N_6514,N_6329,N_6463);
and U6515 (N_6515,N_6307,N_6415);
or U6516 (N_6516,N_6472,N_6266);
or U6517 (N_6517,N_6374,N_6382);
nor U6518 (N_6518,N_6416,N_6488);
nand U6519 (N_6519,N_6436,N_6331);
or U6520 (N_6520,N_6487,N_6403);
or U6521 (N_6521,N_6325,N_6425);
xnor U6522 (N_6522,N_6385,N_6435);
nand U6523 (N_6523,N_6345,N_6390);
nand U6524 (N_6524,N_6437,N_6303);
nand U6525 (N_6525,N_6377,N_6332);
or U6526 (N_6526,N_6365,N_6373);
nand U6527 (N_6527,N_6484,N_6432);
nand U6528 (N_6528,N_6280,N_6367);
nand U6529 (N_6529,N_6379,N_6490);
and U6530 (N_6530,N_6368,N_6485);
and U6531 (N_6531,N_6306,N_6499);
or U6532 (N_6532,N_6380,N_6476);
nand U6533 (N_6533,N_6265,N_6336);
nand U6534 (N_6534,N_6312,N_6441);
nand U6535 (N_6535,N_6346,N_6347);
xnor U6536 (N_6536,N_6464,N_6443);
nor U6537 (N_6537,N_6278,N_6474);
nor U6538 (N_6538,N_6272,N_6497);
and U6539 (N_6539,N_6388,N_6357);
nor U6540 (N_6540,N_6354,N_6339);
xnor U6541 (N_6541,N_6355,N_6316);
and U6542 (N_6542,N_6335,N_6324);
nand U6543 (N_6543,N_6458,N_6319);
or U6544 (N_6544,N_6273,N_6279);
or U6545 (N_6545,N_6250,N_6391);
and U6546 (N_6546,N_6338,N_6478);
nand U6547 (N_6547,N_6283,N_6323);
or U6548 (N_6548,N_6466,N_6461);
nor U6549 (N_6549,N_6428,N_6465);
nor U6550 (N_6550,N_6327,N_6442);
and U6551 (N_6551,N_6251,N_6493);
and U6552 (N_6552,N_6492,N_6456);
xnor U6553 (N_6553,N_6291,N_6429);
and U6554 (N_6554,N_6395,N_6427);
and U6555 (N_6555,N_6262,N_6356);
or U6556 (N_6556,N_6453,N_6375);
and U6557 (N_6557,N_6407,N_6412);
nor U6558 (N_6558,N_6275,N_6322);
xor U6559 (N_6559,N_6301,N_6438);
or U6560 (N_6560,N_6287,N_6398);
nand U6561 (N_6561,N_6420,N_6360);
and U6562 (N_6562,N_6292,N_6393);
or U6563 (N_6563,N_6372,N_6383);
or U6564 (N_6564,N_6270,N_6255);
xnor U6565 (N_6565,N_6289,N_6361);
or U6566 (N_6566,N_6252,N_6264);
nor U6567 (N_6567,N_6261,N_6369);
and U6568 (N_6568,N_6419,N_6396);
and U6569 (N_6569,N_6268,N_6310);
and U6570 (N_6570,N_6263,N_6481);
xnor U6571 (N_6571,N_6334,N_6406);
xnor U6572 (N_6572,N_6256,N_6371);
xnor U6573 (N_6573,N_6321,N_6290);
nor U6574 (N_6574,N_6299,N_6495);
nand U6575 (N_6575,N_6494,N_6317);
nand U6576 (N_6576,N_6479,N_6424);
nand U6577 (N_6577,N_6286,N_6343);
and U6578 (N_6578,N_6457,N_6452);
or U6579 (N_6579,N_6440,N_6293);
nor U6580 (N_6580,N_6480,N_6364);
nor U6581 (N_6581,N_6381,N_6342);
nor U6582 (N_6582,N_6352,N_6433);
nor U6583 (N_6583,N_6455,N_6350);
nor U6584 (N_6584,N_6288,N_6315);
or U6585 (N_6585,N_6446,N_6314);
nand U6586 (N_6586,N_6370,N_6431);
xnor U6587 (N_6587,N_6447,N_6454);
nor U6588 (N_6588,N_6402,N_6302);
nand U6589 (N_6589,N_6309,N_6473);
and U6590 (N_6590,N_6468,N_6426);
xor U6591 (N_6591,N_6274,N_6409);
or U6592 (N_6592,N_6351,N_6257);
nor U6593 (N_6593,N_6477,N_6253);
nand U6594 (N_6594,N_6445,N_6418);
xor U6595 (N_6595,N_6267,N_6399);
or U6596 (N_6596,N_6469,N_6491);
nand U6597 (N_6597,N_6483,N_6300);
xor U6598 (N_6598,N_6496,N_6348);
and U6599 (N_6599,N_6439,N_6308);
and U6600 (N_6600,N_6366,N_6333);
nor U6601 (N_6601,N_6359,N_6318);
or U6602 (N_6602,N_6405,N_6269);
xor U6603 (N_6603,N_6422,N_6460);
and U6604 (N_6604,N_6389,N_6414);
xnor U6605 (N_6605,N_6340,N_6281);
and U6606 (N_6606,N_6386,N_6294);
nor U6607 (N_6607,N_6475,N_6430);
and U6608 (N_6608,N_6284,N_6362);
nor U6609 (N_6609,N_6282,N_6320);
nor U6610 (N_6610,N_6448,N_6423);
and U6611 (N_6611,N_6449,N_6394);
or U6612 (N_6612,N_6489,N_6498);
or U6613 (N_6613,N_6434,N_6276);
or U6614 (N_6614,N_6482,N_6471);
or U6615 (N_6615,N_6408,N_6353);
or U6616 (N_6616,N_6459,N_6384);
or U6617 (N_6617,N_6467,N_6326);
nand U6618 (N_6618,N_6254,N_6349);
or U6619 (N_6619,N_6305,N_6401);
xor U6620 (N_6620,N_6259,N_6404);
nand U6621 (N_6621,N_6421,N_6378);
nand U6622 (N_6622,N_6285,N_6297);
xnor U6623 (N_6623,N_6277,N_6298);
and U6624 (N_6624,N_6462,N_6295);
or U6625 (N_6625,N_6357,N_6389);
nor U6626 (N_6626,N_6402,N_6448);
and U6627 (N_6627,N_6346,N_6252);
or U6628 (N_6628,N_6496,N_6351);
nand U6629 (N_6629,N_6409,N_6411);
and U6630 (N_6630,N_6405,N_6332);
or U6631 (N_6631,N_6485,N_6396);
and U6632 (N_6632,N_6410,N_6298);
xnor U6633 (N_6633,N_6421,N_6292);
nor U6634 (N_6634,N_6278,N_6476);
or U6635 (N_6635,N_6409,N_6268);
or U6636 (N_6636,N_6255,N_6318);
xnor U6637 (N_6637,N_6321,N_6316);
nor U6638 (N_6638,N_6394,N_6379);
nor U6639 (N_6639,N_6428,N_6301);
or U6640 (N_6640,N_6320,N_6428);
or U6641 (N_6641,N_6417,N_6463);
or U6642 (N_6642,N_6456,N_6419);
xor U6643 (N_6643,N_6263,N_6427);
nand U6644 (N_6644,N_6391,N_6412);
nor U6645 (N_6645,N_6422,N_6379);
xnor U6646 (N_6646,N_6254,N_6303);
or U6647 (N_6647,N_6369,N_6278);
and U6648 (N_6648,N_6413,N_6473);
nor U6649 (N_6649,N_6276,N_6280);
xor U6650 (N_6650,N_6251,N_6300);
and U6651 (N_6651,N_6418,N_6268);
xor U6652 (N_6652,N_6473,N_6391);
and U6653 (N_6653,N_6337,N_6363);
xnor U6654 (N_6654,N_6425,N_6345);
nand U6655 (N_6655,N_6321,N_6366);
or U6656 (N_6656,N_6390,N_6480);
nor U6657 (N_6657,N_6344,N_6444);
and U6658 (N_6658,N_6437,N_6375);
nand U6659 (N_6659,N_6450,N_6441);
or U6660 (N_6660,N_6346,N_6447);
nor U6661 (N_6661,N_6275,N_6479);
nor U6662 (N_6662,N_6352,N_6310);
or U6663 (N_6663,N_6453,N_6391);
or U6664 (N_6664,N_6451,N_6355);
xnor U6665 (N_6665,N_6382,N_6272);
nand U6666 (N_6666,N_6411,N_6458);
and U6667 (N_6667,N_6314,N_6265);
nand U6668 (N_6668,N_6304,N_6375);
or U6669 (N_6669,N_6378,N_6468);
nor U6670 (N_6670,N_6435,N_6397);
xnor U6671 (N_6671,N_6495,N_6388);
nor U6672 (N_6672,N_6410,N_6267);
or U6673 (N_6673,N_6308,N_6256);
nor U6674 (N_6674,N_6275,N_6384);
xnor U6675 (N_6675,N_6397,N_6341);
nand U6676 (N_6676,N_6420,N_6391);
nand U6677 (N_6677,N_6451,N_6387);
nand U6678 (N_6678,N_6337,N_6336);
or U6679 (N_6679,N_6409,N_6348);
or U6680 (N_6680,N_6369,N_6407);
nand U6681 (N_6681,N_6382,N_6431);
and U6682 (N_6682,N_6453,N_6394);
and U6683 (N_6683,N_6317,N_6300);
and U6684 (N_6684,N_6467,N_6358);
nand U6685 (N_6685,N_6396,N_6479);
xor U6686 (N_6686,N_6333,N_6372);
and U6687 (N_6687,N_6457,N_6396);
nand U6688 (N_6688,N_6469,N_6380);
nor U6689 (N_6689,N_6457,N_6296);
xor U6690 (N_6690,N_6440,N_6304);
nor U6691 (N_6691,N_6312,N_6326);
xor U6692 (N_6692,N_6388,N_6458);
nand U6693 (N_6693,N_6415,N_6350);
and U6694 (N_6694,N_6461,N_6307);
nand U6695 (N_6695,N_6413,N_6393);
nand U6696 (N_6696,N_6437,N_6499);
nor U6697 (N_6697,N_6257,N_6359);
xnor U6698 (N_6698,N_6391,N_6352);
xor U6699 (N_6699,N_6280,N_6333);
and U6700 (N_6700,N_6351,N_6273);
and U6701 (N_6701,N_6388,N_6377);
nor U6702 (N_6702,N_6389,N_6431);
xor U6703 (N_6703,N_6437,N_6357);
xnor U6704 (N_6704,N_6280,N_6281);
and U6705 (N_6705,N_6371,N_6343);
and U6706 (N_6706,N_6432,N_6440);
nor U6707 (N_6707,N_6273,N_6385);
nor U6708 (N_6708,N_6306,N_6343);
or U6709 (N_6709,N_6258,N_6267);
nand U6710 (N_6710,N_6348,N_6362);
and U6711 (N_6711,N_6323,N_6451);
and U6712 (N_6712,N_6349,N_6358);
xor U6713 (N_6713,N_6417,N_6282);
or U6714 (N_6714,N_6271,N_6371);
or U6715 (N_6715,N_6261,N_6319);
nor U6716 (N_6716,N_6407,N_6357);
nand U6717 (N_6717,N_6333,N_6317);
xor U6718 (N_6718,N_6317,N_6280);
nor U6719 (N_6719,N_6441,N_6438);
xnor U6720 (N_6720,N_6483,N_6424);
nand U6721 (N_6721,N_6412,N_6394);
xor U6722 (N_6722,N_6496,N_6403);
nand U6723 (N_6723,N_6450,N_6499);
xor U6724 (N_6724,N_6454,N_6259);
nand U6725 (N_6725,N_6273,N_6426);
xor U6726 (N_6726,N_6425,N_6426);
xor U6727 (N_6727,N_6371,N_6471);
xor U6728 (N_6728,N_6293,N_6314);
and U6729 (N_6729,N_6383,N_6278);
nand U6730 (N_6730,N_6318,N_6467);
xnor U6731 (N_6731,N_6424,N_6368);
xor U6732 (N_6732,N_6445,N_6484);
nand U6733 (N_6733,N_6321,N_6365);
xor U6734 (N_6734,N_6426,N_6451);
and U6735 (N_6735,N_6390,N_6425);
or U6736 (N_6736,N_6448,N_6298);
and U6737 (N_6737,N_6375,N_6488);
or U6738 (N_6738,N_6413,N_6411);
or U6739 (N_6739,N_6322,N_6423);
xor U6740 (N_6740,N_6449,N_6295);
xor U6741 (N_6741,N_6255,N_6470);
nor U6742 (N_6742,N_6281,N_6422);
or U6743 (N_6743,N_6446,N_6458);
or U6744 (N_6744,N_6462,N_6460);
nor U6745 (N_6745,N_6362,N_6309);
nor U6746 (N_6746,N_6356,N_6258);
and U6747 (N_6747,N_6283,N_6435);
or U6748 (N_6748,N_6419,N_6310);
xnor U6749 (N_6749,N_6313,N_6431);
xor U6750 (N_6750,N_6500,N_6543);
or U6751 (N_6751,N_6680,N_6551);
nor U6752 (N_6752,N_6579,N_6661);
nor U6753 (N_6753,N_6523,N_6559);
and U6754 (N_6754,N_6657,N_6652);
and U6755 (N_6755,N_6541,N_6624);
or U6756 (N_6756,N_6524,N_6571);
or U6757 (N_6757,N_6689,N_6504);
or U6758 (N_6758,N_6679,N_6632);
or U6759 (N_6759,N_6691,N_6690);
nand U6760 (N_6760,N_6717,N_6711);
and U6761 (N_6761,N_6605,N_6641);
nor U6762 (N_6762,N_6615,N_6710);
xor U6763 (N_6763,N_6638,N_6586);
nor U6764 (N_6764,N_6598,N_6702);
and U6765 (N_6765,N_6516,N_6533);
and U6766 (N_6766,N_6606,N_6589);
and U6767 (N_6767,N_6709,N_6723);
nand U6768 (N_6768,N_6655,N_6728);
nor U6769 (N_6769,N_6739,N_6526);
nand U6770 (N_6770,N_6603,N_6736);
nand U6771 (N_6771,N_6614,N_6570);
and U6772 (N_6772,N_6629,N_6740);
xnor U6773 (N_6773,N_6677,N_6540);
or U6774 (N_6774,N_6686,N_6715);
nand U6775 (N_6775,N_6577,N_6721);
xor U6776 (N_6776,N_6597,N_6631);
xnor U6777 (N_6777,N_6590,N_6654);
nor U6778 (N_6778,N_6720,N_6694);
nor U6779 (N_6779,N_6563,N_6507);
nor U6780 (N_6780,N_6749,N_6644);
and U6781 (N_6781,N_6576,N_6648);
or U6782 (N_6782,N_6688,N_6515);
nor U6783 (N_6783,N_6707,N_6668);
and U6784 (N_6784,N_6678,N_6512);
xor U6785 (N_6785,N_6514,N_6672);
xnor U6786 (N_6786,N_6556,N_6685);
nor U6787 (N_6787,N_6660,N_6633);
nor U6788 (N_6788,N_6663,N_6664);
nand U6789 (N_6789,N_6608,N_6636);
nor U6790 (N_6790,N_6534,N_6503);
nand U6791 (N_6791,N_6506,N_6596);
or U6792 (N_6792,N_6716,N_6670);
and U6793 (N_6793,N_6646,N_6675);
nor U6794 (N_6794,N_6746,N_6741);
or U6795 (N_6795,N_6613,N_6650);
or U6796 (N_6796,N_6669,N_6725);
and U6797 (N_6797,N_6607,N_6713);
nor U6798 (N_6798,N_6546,N_6682);
or U6799 (N_6799,N_6553,N_6628);
or U6800 (N_6800,N_6568,N_6616);
or U6801 (N_6801,N_6537,N_6671);
or U6802 (N_6802,N_6642,N_6529);
nor U6803 (N_6803,N_6639,N_6738);
and U6804 (N_6804,N_6530,N_6735);
and U6805 (N_6805,N_6531,N_6592);
or U6806 (N_6806,N_6547,N_6649);
nand U6807 (N_6807,N_6706,N_6593);
and U6808 (N_6808,N_6674,N_6712);
nand U6809 (N_6809,N_6595,N_6532);
nor U6810 (N_6810,N_6548,N_6714);
and U6811 (N_6811,N_6525,N_6698);
or U6812 (N_6812,N_6703,N_6519);
and U6813 (N_6813,N_6722,N_6604);
xor U6814 (N_6814,N_6584,N_6748);
nand U6815 (N_6815,N_6665,N_6666);
or U6816 (N_6816,N_6501,N_6742);
nor U6817 (N_6817,N_6585,N_6704);
or U6818 (N_6818,N_6620,N_6520);
and U6819 (N_6819,N_6574,N_6509);
nor U6820 (N_6820,N_6719,N_6699);
and U6821 (N_6821,N_6676,N_6730);
nand U6822 (N_6822,N_6695,N_6625);
nand U6823 (N_6823,N_6518,N_6692);
and U6824 (N_6824,N_6696,N_6609);
xnor U6825 (N_6825,N_6542,N_6673);
or U6826 (N_6826,N_6508,N_6659);
xnor U6827 (N_6827,N_6581,N_6617);
and U6828 (N_6828,N_6647,N_6573);
or U6829 (N_6829,N_6627,N_6656);
xor U6830 (N_6830,N_6505,N_6718);
and U6831 (N_6831,N_6634,N_6502);
nand U6832 (N_6832,N_6562,N_6591);
nand U6833 (N_6833,N_6727,N_6550);
and U6834 (N_6834,N_6536,N_6557);
nor U6835 (N_6835,N_6635,N_6681);
or U6836 (N_6836,N_6560,N_6693);
and U6837 (N_6837,N_6732,N_6697);
nand U6838 (N_6838,N_6619,N_6667);
and U6839 (N_6839,N_6527,N_6561);
nand U6840 (N_6840,N_6658,N_6601);
or U6841 (N_6841,N_6588,N_6731);
nor U6842 (N_6842,N_6626,N_6569);
nand U6843 (N_6843,N_6521,N_6567);
or U6844 (N_6844,N_6610,N_6564);
nand U6845 (N_6845,N_6621,N_6683);
xnor U6846 (N_6846,N_6575,N_6555);
or U6847 (N_6847,N_6552,N_6544);
and U6848 (N_6848,N_6708,N_6511);
or U6849 (N_6849,N_6611,N_6622);
or U6850 (N_6850,N_6687,N_6640);
or U6851 (N_6851,N_6701,N_6545);
and U6852 (N_6852,N_6572,N_6517);
nor U6853 (N_6853,N_6747,N_6643);
nor U6854 (N_6854,N_6724,N_6558);
nor U6855 (N_6855,N_6744,N_6583);
nor U6856 (N_6856,N_6637,N_6726);
xnor U6857 (N_6857,N_6587,N_6729);
and U6858 (N_6858,N_6700,N_6743);
nor U6859 (N_6859,N_6565,N_6612);
nor U6860 (N_6860,N_6705,N_6522);
or U6861 (N_6861,N_6684,N_6513);
and U6862 (N_6862,N_6745,N_6535);
or U6863 (N_6863,N_6602,N_6580);
nor U6864 (N_6864,N_6510,N_6734);
nand U6865 (N_6865,N_6645,N_6600);
nand U6866 (N_6866,N_6549,N_6599);
nand U6867 (N_6867,N_6618,N_6582);
xnor U6868 (N_6868,N_6733,N_6528);
nor U6869 (N_6869,N_6623,N_6651);
xor U6870 (N_6870,N_6630,N_6737);
and U6871 (N_6871,N_6566,N_6554);
nand U6872 (N_6872,N_6662,N_6578);
xor U6873 (N_6873,N_6539,N_6538);
or U6874 (N_6874,N_6594,N_6653);
and U6875 (N_6875,N_6697,N_6679);
xor U6876 (N_6876,N_6583,N_6627);
and U6877 (N_6877,N_6685,N_6705);
and U6878 (N_6878,N_6712,N_6635);
nor U6879 (N_6879,N_6711,N_6618);
xor U6880 (N_6880,N_6615,N_6676);
nand U6881 (N_6881,N_6749,N_6650);
nand U6882 (N_6882,N_6503,N_6690);
nand U6883 (N_6883,N_6601,N_6729);
xor U6884 (N_6884,N_6650,N_6557);
and U6885 (N_6885,N_6742,N_6505);
nor U6886 (N_6886,N_6623,N_6614);
or U6887 (N_6887,N_6513,N_6711);
and U6888 (N_6888,N_6679,N_6500);
xnor U6889 (N_6889,N_6512,N_6663);
and U6890 (N_6890,N_6547,N_6519);
and U6891 (N_6891,N_6700,N_6590);
nor U6892 (N_6892,N_6536,N_6594);
and U6893 (N_6893,N_6585,N_6668);
nor U6894 (N_6894,N_6562,N_6698);
and U6895 (N_6895,N_6514,N_6505);
nand U6896 (N_6896,N_6614,N_6580);
xnor U6897 (N_6897,N_6502,N_6545);
or U6898 (N_6898,N_6713,N_6637);
and U6899 (N_6899,N_6567,N_6691);
xor U6900 (N_6900,N_6620,N_6512);
and U6901 (N_6901,N_6525,N_6731);
or U6902 (N_6902,N_6700,N_6623);
nor U6903 (N_6903,N_6668,N_6506);
or U6904 (N_6904,N_6625,N_6648);
xor U6905 (N_6905,N_6698,N_6670);
and U6906 (N_6906,N_6501,N_6620);
nor U6907 (N_6907,N_6737,N_6621);
nor U6908 (N_6908,N_6672,N_6710);
nor U6909 (N_6909,N_6616,N_6656);
and U6910 (N_6910,N_6607,N_6613);
and U6911 (N_6911,N_6569,N_6676);
nand U6912 (N_6912,N_6705,N_6616);
and U6913 (N_6913,N_6566,N_6544);
nor U6914 (N_6914,N_6500,N_6626);
nand U6915 (N_6915,N_6651,N_6661);
and U6916 (N_6916,N_6749,N_6668);
xnor U6917 (N_6917,N_6534,N_6674);
nor U6918 (N_6918,N_6601,N_6502);
nand U6919 (N_6919,N_6522,N_6519);
or U6920 (N_6920,N_6561,N_6530);
nor U6921 (N_6921,N_6547,N_6591);
or U6922 (N_6922,N_6641,N_6681);
nor U6923 (N_6923,N_6623,N_6609);
xor U6924 (N_6924,N_6609,N_6647);
or U6925 (N_6925,N_6646,N_6503);
nand U6926 (N_6926,N_6742,N_6597);
and U6927 (N_6927,N_6606,N_6691);
nor U6928 (N_6928,N_6585,N_6543);
nand U6929 (N_6929,N_6510,N_6741);
xor U6930 (N_6930,N_6739,N_6679);
nor U6931 (N_6931,N_6744,N_6737);
xnor U6932 (N_6932,N_6601,N_6597);
nor U6933 (N_6933,N_6531,N_6676);
nand U6934 (N_6934,N_6533,N_6670);
xor U6935 (N_6935,N_6511,N_6500);
xor U6936 (N_6936,N_6687,N_6543);
xor U6937 (N_6937,N_6592,N_6522);
nand U6938 (N_6938,N_6678,N_6580);
xnor U6939 (N_6939,N_6525,N_6628);
nand U6940 (N_6940,N_6529,N_6598);
nor U6941 (N_6941,N_6701,N_6639);
nor U6942 (N_6942,N_6580,N_6597);
nand U6943 (N_6943,N_6624,N_6699);
or U6944 (N_6944,N_6577,N_6603);
xnor U6945 (N_6945,N_6559,N_6719);
nand U6946 (N_6946,N_6742,N_6664);
nand U6947 (N_6947,N_6633,N_6675);
nand U6948 (N_6948,N_6664,N_6636);
and U6949 (N_6949,N_6648,N_6538);
and U6950 (N_6950,N_6603,N_6598);
nor U6951 (N_6951,N_6561,N_6661);
xor U6952 (N_6952,N_6686,N_6717);
xnor U6953 (N_6953,N_6606,N_6699);
and U6954 (N_6954,N_6546,N_6539);
nand U6955 (N_6955,N_6559,N_6557);
or U6956 (N_6956,N_6716,N_6561);
and U6957 (N_6957,N_6584,N_6685);
or U6958 (N_6958,N_6586,N_6682);
xor U6959 (N_6959,N_6548,N_6566);
xnor U6960 (N_6960,N_6616,N_6588);
nor U6961 (N_6961,N_6674,N_6578);
nand U6962 (N_6962,N_6619,N_6720);
nand U6963 (N_6963,N_6651,N_6555);
nor U6964 (N_6964,N_6565,N_6596);
or U6965 (N_6965,N_6526,N_6566);
nand U6966 (N_6966,N_6711,N_6526);
xor U6967 (N_6967,N_6563,N_6616);
nand U6968 (N_6968,N_6581,N_6685);
or U6969 (N_6969,N_6513,N_6563);
nand U6970 (N_6970,N_6631,N_6542);
nand U6971 (N_6971,N_6547,N_6605);
xnor U6972 (N_6972,N_6612,N_6741);
nand U6973 (N_6973,N_6612,N_6700);
and U6974 (N_6974,N_6742,N_6618);
xor U6975 (N_6975,N_6748,N_6627);
and U6976 (N_6976,N_6682,N_6604);
nor U6977 (N_6977,N_6558,N_6542);
and U6978 (N_6978,N_6501,N_6663);
nand U6979 (N_6979,N_6674,N_6598);
nor U6980 (N_6980,N_6548,N_6635);
and U6981 (N_6981,N_6577,N_6609);
or U6982 (N_6982,N_6673,N_6703);
xnor U6983 (N_6983,N_6623,N_6718);
or U6984 (N_6984,N_6606,N_6659);
nand U6985 (N_6985,N_6583,N_6504);
or U6986 (N_6986,N_6534,N_6739);
and U6987 (N_6987,N_6567,N_6591);
and U6988 (N_6988,N_6591,N_6696);
and U6989 (N_6989,N_6515,N_6716);
nor U6990 (N_6990,N_6727,N_6637);
nand U6991 (N_6991,N_6598,N_6707);
and U6992 (N_6992,N_6679,N_6724);
xor U6993 (N_6993,N_6500,N_6649);
xnor U6994 (N_6994,N_6695,N_6741);
nand U6995 (N_6995,N_6593,N_6551);
xor U6996 (N_6996,N_6625,N_6568);
and U6997 (N_6997,N_6739,N_6522);
or U6998 (N_6998,N_6618,N_6732);
or U6999 (N_6999,N_6562,N_6530);
and U7000 (N_7000,N_6863,N_6856);
or U7001 (N_7001,N_6936,N_6806);
or U7002 (N_7002,N_6908,N_6797);
nand U7003 (N_7003,N_6795,N_6851);
and U7004 (N_7004,N_6864,N_6932);
and U7005 (N_7005,N_6910,N_6794);
or U7006 (N_7006,N_6967,N_6764);
nand U7007 (N_7007,N_6954,N_6841);
nor U7008 (N_7008,N_6986,N_6876);
or U7009 (N_7009,N_6884,N_6957);
and U7010 (N_7010,N_6962,N_6828);
nor U7011 (N_7011,N_6919,N_6879);
nand U7012 (N_7012,N_6818,N_6784);
and U7013 (N_7013,N_6773,N_6801);
xor U7014 (N_7014,N_6903,N_6781);
and U7015 (N_7015,N_6855,N_6783);
nand U7016 (N_7016,N_6940,N_6949);
xor U7017 (N_7017,N_6933,N_6771);
nand U7018 (N_7018,N_6946,N_6812);
nor U7019 (N_7019,N_6937,N_6975);
nand U7020 (N_7020,N_6819,N_6898);
nand U7021 (N_7021,N_6897,N_6815);
and U7022 (N_7022,N_6899,N_6950);
xor U7023 (N_7023,N_6878,N_6750);
and U7024 (N_7024,N_6869,N_6770);
nand U7025 (N_7025,N_6843,N_6961);
nor U7026 (N_7026,N_6798,N_6942);
and U7027 (N_7027,N_6772,N_6906);
or U7028 (N_7028,N_6846,N_6861);
and U7029 (N_7029,N_6960,N_6998);
xnor U7030 (N_7030,N_6928,N_6862);
and U7031 (N_7031,N_6965,N_6912);
xor U7032 (N_7032,N_6787,N_6814);
or U7033 (N_7033,N_6973,N_6766);
nor U7034 (N_7034,N_6823,N_6977);
xor U7035 (N_7035,N_6844,N_6845);
or U7036 (N_7036,N_6907,N_6935);
nand U7037 (N_7037,N_6881,N_6829);
nor U7038 (N_7038,N_6997,N_6836);
xnor U7039 (N_7039,N_6969,N_6927);
or U7040 (N_7040,N_6785,N_6892);
or U7041 (N_7041,N_6758,N_6759);
nand U7042 (N_7042,N_6917,N_6947);
nand U7043 (N_7043,N_6870,N_6800);
and U7044 (N_7044,N_6796,N_6993);
and U7045 (N_7045,N_6754,N_6871);
and U7046 (N_7046,N_6808,N_6921);
or U7047 (N_7047,N_6788,N_6945);
or U7048 (N_7048,N_6761,N_6914);
and U7049 (N_7049,N_6887,N_6989);
xor U7050 (N_7050,N_6813,N_6832);
nand U7051 (N_7051,N_6756,N_6775);
xnor U7052 (N_7052,N_6779,N_6753);
xnor U7053 (N_7053,N_6952,N_6924);
or U7054 (N_7054,N_6847,N_6987);
or U7055 (N_7055,N_6971,N_6896);
xor U7056 (N_7056,N_6979,N_6956);
or U7057 (N_7057,N_6874,N_6765);
and U7058 (N_7058,N_6763,N_6951);
nor U7059 (N_7059,N_6891,N_6976);
nor U7060 (N_7060,N_6833,N_6838);
and U7061 (N_7061,N_6982,N_6966);
nor U7062 (N_7062,N_6918,N_6939);
or U7063 (N_7063,N_6840,N_6824);
nand U7064 (N_7064,N_6983,N_6854);
or U7065 (N_7065,N_6880,N_6826);
xnor U7066 (N_7066,N_6882,N_6981);
nand U7067 (N_7067,N_6852,N_6886);
xor U7068 (N_7068,N_6755,N_6901);
xor U7069 (N_7069,N_6790,N_6842);
xnor U7070 (N_7070,N_6804,N_6799);
nor U7071 (N_7071,N_6978,N_6831);
nand U7072 (N_7072,N_6889,N_6980);
and U7073 (N_7073,N_6768,N_6866);
xnor U7074 (N_7074,N_6858,N_6778);
xor U7075 (N_7075,N_6791,N_6948);
nor U7076 (N_7076,N_6849,N_6964);
nand U7077 (N_7077,N_6894,N_6857);
nand U7078 (N_7078,N_6968,N_6873);
or U7079 (N_7079,N_6991,N_6895);
and U7080 (N_7080,N_6913,N_6835);
xor U7081 (N_7081,N_6958,N_6920);
and U7082 (N_7082,N_6850,N_6931);
nand U7083 (N_7083,N_6959,N_6995);
nand U7084 (N_7084,N_6926,N_6807);
xnor U7085 (N_7085,N_6974,N_6834);
xnor U7086 (N_7086,N_6789,N_6777);
or U7087 (N_7087,N_6751,N_6792);
nand U7088 (N_7088,N_6848,N_6963);
and U7089 (N_7089,N_6930,N_6827);
and U7090 (N_7090,N_6994,N_6817);
nor U7091 (N_7091,N_6905,N_6923);
nor U7092 (N_7092,N_6902,N_6820);
nor U7093 (N_7093,N_6769,N_6875);
xnor U7094 (N_7094,N_6816,N_6934);
nor U7095 (N_7095,N_6865,N_6985);
xnor U7096 (N_7096,N_6970,N_6872);
nand U7097 (N_7097,N_6830,N_6810);
or U7098 (N_7098,N_6859,N_6955);
nor U7099 (N_7099,N_6953,N_6988);
and U7100 (N_7100,N_6776,N_6883);
nand U7101 (N_7101,N_6825,N_6941);
and U7102 (N_7102,N_6888,N_6944);
or U7103 (N_7103,N_6760,N_6909);
and U7104 (N_7104,N_6809,N_6893);
xnor U7105 (N_7105,N_6868,N_6984);
nand U7106 (N_7106,N_6922,N_6821);
nand U7107 (N_7107,N_6811,N_6999);
nand U7108 (N_7108,N_6767,N_6802);
xnor U7109 (N_7109,N_6943,N_6853);
and U7110 (N_7110,N_6877,N_6752);
xor U7111 (N_7111,N_6786,N_6762);
and U7112 (N_7112,N_6911,N_6837);
nand U7113 (N_7113,N_6885,N_6793);
and U7114 (N_7114,N_6929,N_6780);
or U7115 (N_7115,N_6782,N_6867);
nand U7116 (N_7116,N_6992,N_6925);
or U7117 (N_7117,N_6990,N_6805);
or U7118 (N_7118,N_6938,N_6774);
nand U7119 (N_7119,N_6996,N_6839);
xnor U7120 (N_7120,N_6915,N_6972);
nor U7121 (N_7121,N_6904,N_6900);
nor U7122 (N_7122,N_6890,N_6822);
nand U7123 (N_7123,N_6803,N_6916);
nor U7124 (N_7124,N_6860,N_6757);
nand U7125 (N_7125,N_6926,N_6915);
xor U7126 (N_7126,N_6879,N_6963);
nor U7127 (N_7127,N_6816,N_6889);
nor U7128 (N_7128,N_6811,N_6855);
or U7129 (N_7129,N_6829,N_6858);
or U7130 (N_7130,N_6757,N_6769);
nand U7131 (N_7131,N_6872,N_6905);
nand U7132 (N_7132,N_6780,N_6940);
and U7133 (N_7133,N_6755,N_6853);
xnor U7134 (N_7134,N_6783,N_6822);
and U7135 (N_7135,N_6846,N_6842);
and U7136 (N_7136,N_6895,N_6913);
and U7137 (N_7137,N_6952,N_6916);
and U7138 (N_7138,N_6983,N_6891);
or U7139 (N_7139,N_6883,N_6840);
xnor U7140 (N_7140,N_6928,N_6896);
or U7141 (N_7141,N_6864,N_6848);
nor U7142 (N_7142,N_6942,N_6884);
xor U7143 (N_7143,N_6759,N_6972);
or U7144 (N_7144,N_6780,N_6992);
and U7145 (N_7145,N_6920,N_6793);
xnor U7146 (N_7146,N_6913,N_6787);
or U7147 (N_7147,N_6852,N_6877);
xnor U7148 (N_7148,N_6780,N_6903);
xnor U7149 (N_7149,N_6794,N_6994);
xor U7150 (N_7150,N_6818,N_6997);
or U7151 (N_7151,N_6944,N_6997);
nand U7152 (N_7152,N_6965,N_6922);
xnor U7153 (N_7153,N_6861,N_6987);
xnor U7154 (N_7154,N_6793,N_6966);
nor U7155 (N_7155,N_6815,N_6838);
xnor U7156 (N_7156,N_6758,N_6832);
nor U7157 (N_7157,N_6927,N_6987);
xor U7158 (N_7158,N_6864,N_6776);
nor U7159 (N_7159,N_6820,N_6876);
and U7160 (N_7160,N_6766,N_6758);
or U7161 (N_7161,N_6853,N_6994);
nand U7162 (N_7162,N_6858,N_6974);
nand U7163 (N_7163,N_6948,N_6814);
nor U7164 (N_7164,N_6765,N_6814);
or U7165 (N_7165,N_6903,N_6809);
nor U7166 (N_7166,N_6819,N_6859);
and U7167 (N_7167,N_6932,N_6850);
nand U7168 (N_7168,N_6931,N_6989);
xnor U7169 (N_7169,N_6768,N_6890);
or U7170 (N_7170,N_6841,N_6986);
xnor U7171 (N_7171,N_6805,N_6911);
nor U7172 (N_7172,N_6967,N_6940);
nor U7173 (N_7173,N_6847,N_6978);
nor U7174 (N_7174,N_6786,N_6861);
nor U7175 (N_7175,N_6835,N_6938);
or U7176 (N_7176,N_6839,N_6856);
nand U7177 (N_7177,N_6967,N_6891);
and U7178 (N_7178,N_6951,N_6983);
and U7179 (N_7179,N_6943,N_6959);
and U7180 (N_7180,N_6807,N_6868);
and U7181 (N_7181,N_6761,N_6849);
nand U7182 (N_7182,N_6856,N_6920);
or U7183 (N_7183,N_6921,N_6947);
nand U7184 (N_7184,N_6752,N_6966);
or U7185 (N_7185,N_6782,N_6950);
and U7186 (N_7186,N_6944,N_6993);
nor U7187 (N_7187,N_6791,N_6905);
and U7188 (N_7188,N_6872,N_6824);
and U7189 (N_7189,N_6858,N_6933);
nand U7190 (N_7190,N_6955,N_6811);
nand U7191 (N_7191,N_6827,N_6826);
xor U7192 (N_7192,N_6853,N_6750);
nand U7193 (N_7193,N_6826,N_6889);
and U7194 (N_7194,N_6939,N_6927);
or U7195 (N_7195,N_6936,N_6850);
or U7196 (N_7196,N_6864,N_6816);
or U7197 (N_7197,N_6906,N_6811);
xnor U7198 (N_7198,N_6950,N_6808);
nand U7199 (N_7199,N_6959,N_6795);
nand U7200 (N_7200,N_6782,N_6830);
nand U7201 (N_7201,N_6967,N_6813);
nand U7202 (N_7202,N_6861,N_6803);
xor U7203 (N_7203,N_6946,N_6943);
xnor U7204 (N_7204,N_6899,N_6857);
and U7205 (N_7205,N_6771,N_6832);
nor U7206 (N_7206,N_6934,N_6961);
and U7207 (N_7207,N_6973,N_6781);
nor U7208 (N_7208,N_6795,N_6775);
nor U7209 (N_7209,N_6810,N_6837);
and U7210 (N_7210,N_6969,N_6955);
nor U7211 (N_7211,N_6834,N_6835);
or U7212 (N_7212,N_6945,N_6972);
and U7213 (N_7213,N_6760,N_6838);
and U7214 (N_7214,N_6913,N_6885);
and U7215 (N_7215,N_6784,N_6870);
nor U7216 (N_7216,N_6771,N_6858);
or U7217 (N_7217,N_6770,N_6946);
and U7218 (N_7218,N_6804,N_6966);
or U7219 (N_7219,N_6761,N_6852);
nor U7220 (N_7220,N_6808,N_6892);
nor U7221 (N_7221,N_6793,N_6825);
or U7222 (N_7222,N_6868,N_6869);
or U7223 (N_7223,N_6784,N_6956);
nor U7224 (N_7224,N_6980,N_6952);
or U7225 (N_7225,N_6886,N_6820);
or U7226 (N_7226,N_6785,N_6833);
xor U7227 (N_7227,N_6760,N_6906);
xor U7228 (N_7228,N_6802,N_6877);
xor U7229 (N_7229,N_6943,N_6753);
nand U7230 (N_7230,N_6964,N_6806);
or U7231 (N_7231,N_6919,N_6952);
or U7232 (N_7232,N_6996,N_6753);
nor U7233 (N_7233,N_6935,N_6928);
nand U7234 (N_7234,N_6866,N_6957);
nor U7235 (N_7235,N_6879,N_6870);
xor U7236 (N_7236,N_6821,N_6957);
nor U7237 (N_7237,N_6988,N_6876);
nand U7238 (N_7238,N_6998,N_6877);
or U7239 (N_7239,N_6870,N_6853);
xor U7240 (N_7240,N_6846,N_6751);
nor U7241 (N_7241,N_6858,N_6927);
xor U7242 (N_7242,N_6939,N_6848);
and U7243 (N_7243,N_6773,N_6793);
and U7244 (N_7244,N_6784,N_6770);
nand U7245 (N_7245,N_6833,N_6897);
or U7246 (N_7246,N_6766,N_6931);
nor U7247 (N_7247,N_6905,N_6770);
nand U7248 (N_7248,N_6770,N_6826);
xnor U7249 (N_7249,N_6838,N_6961);
nor U7250 (N_7250,N_7172,N_7233);
nor U7251 (N_7251,N_7144,N_7055);
nand U7252 (N_7252,N_7028,N_7186);
nand U7253 (N_7253,N_7222,N_7036);
nor U7254 (N_7254,N_7127,N_7034);
xnor U7255 (N_7255,N_7185,N_7207);
nor U7256 (N_7256,N_7155,N_7130);
or U7257 (N_7257,N_7002,N_7202);
xnor U7258 (N_7258,N_7027,N_7069);
nor U7259 (N_7259,N_7158,N_7171);
or U7260 (N_7260,N_7248,N_7210);
nor U7261 (N_7261,N_7134,N_7166);
nor U7262 (N_7262,N_7225,N_7153);
and U7263 (N_7263,N_7215,N_7243);
and U7264 (N_7264,N_7173,N_7216);
or U7265 (N_7265,N_7198,N_7089);
nand U7266 (N_7266,N_7108,N_7204);
nor U7267 (N_7267,N_7132,N_7212);
and U7268 (N_7268,N_7227,N_7213);
and U7269 (N_7269,N_7109,N_7030);
or U7270 (N_7270,N_7119,N_7107);
nand U7271 (N_7271,N_7063,N_7240);
nand U7272 (N_7272,N_7062,N_7223);
xnor U7273 (N_7273,N_7190,N_7052);
and U7274 (N_7274,N_7131,N_7219);
nand U7275 (N_7275,N_7046,N_7082);
xnor U7276 (N_7276,N_7137,N_7050);
nor U7277 (N_7277,N_7023,N_7241);
or U7278 (N_7278,N_7182,N_7197);
nor U7279 (N_7279,N_7125,N_7018);
and U7280 (N_7280,N_7145,N_7101);
xor U7281 (N_7281,N_7175,N_7011);
nand U7282 (N_7282,N_7054,N_7168);
and U7283 (N_7283,N_7122,N_7151);
or U7284 (N_7284,N_7105,N_7010);
xnor U7285 (N_7285,N_7195,N_7091);
xnor U7286 (N_7286,N_7084,N_7013);
xnor U7287 (N_7287,N_7059,N_7060);
xor U7288 (N_7288,N_7188,N_7200);
nor U7289 (N_7289,N_7087,N_7029);
xnor U7290 (N_7290,N_7051,N_7096);
and U7291 (N_7291,N_7176,N_7019);
nor U7292 (N_7292,N_7043,N_7070);
or U7293 (N_7293,N_7114,N_7199);
or U7294 (N_7294,N_7037,N_7143);
nor U7295 (N_7295,N_7220,N_7041);
or U7296 (N_7296,N_7039,N_7135);
xor U7297 (N_7297,N_7174,N_7235);
nor U7298 (N_7298,N_7203,N_7071);
and U7299 (N_7299,N_7136,N_7249);
or U7300 (N_7300,N_7209,N_7061);
xnor U7301 (N_7301,N_7184,N_7066);
xor U7302 (N_7302,N_7040,N_7126);
and U7303 (N_7303,N_7008,N_7115);
nand U7304 (N_7304,N_7189,N_7129);
xor U7305 (N_7305,N_7149,N_7026);
or U7306 (N_7306,N_7057,N_7118);
xnor U7307 (N_7307,N_7120,N_7100);
nor U7308 (N_7308,N_7237,N_7160);
nand U7309 (N_7309,N_7232,N_7090);
xor U7310 (N_7310,N_7156,N_7191);
nand U7311 (N_7311,N_7242,N_7094);
nand U7312 (N_7312,N_7081,N_7234);
nor U7313 (N_7313,N_7077,N_7238);
nor U7314 (N_7314,N_7072,N_7229);
xor U7315 (N_7315,N_7086,N_7142);
nor U7316 (N_7316,N_7092,N_7009);
xnor U7317 (N_7317,N_7067,N_7102);
xnor U7318 (N_7318,N_7079,N_7110);
or U7319 (N_7319,N_7083,N_7206);
nor U7320 (N_7320,N_7074,N_7075);
or U7321 (N_7321,N_7247,N_7139);
or U7322 (N_7322,N_7228,N_7245);
xor U7323 (N_7323,N_7231,N_7169);
and U7324 (N_7324,N_7147,N_7183);
nor U7325 (N_7325,N_7048,N_7159);
or U7326 (N_7326,N_7016,N_7214);
nand U7327 (N_7327,N_7058,N_7116);
nor U7328 (N_7328,N_7022,N_7020);
and U7329 (N_7329,N_7146,N_7244);
or U7330 (N_7330,N_7236,N_7049);
nand U7331 (N_7331,N_7194,N_7167);
or U7332 (N_7332,N_7113,N_7117);
xor U7333 (N_7333,N_7162,N_7128);
nor U7334 (N_7334,N_7000,N_7047);
xnor U7335 (N_7335,N_7150,N_7123);
xor U7336 (N_7336,N_7226,N_7133);
and U7337 (N_7337,N_7015,N_7140);
xnor U7338 (N_7338,N_7178,N_7103);
and U7339 (N_7339,N_7164,N_7095);
nor U7340 (N_7340,N_7106,N_7042);
and U7341 (N_7341,N_7068,N_7045);
or U7342 (N_7342,N_7161,N_7038);
or U7343 (N_7343,N_7138,N_7014);
nor U7344 (N_7344,N_7078,N_7080);
or U7345 (N_7345,N_7208,N_7239);
or U7346 (N_7346,N_7017,N_7007);
nand U7347 (N_7347,N_7031,N_7073);
or U7348 (N_7348,N_7217,N_7187);
or U7349 (N_7349,N_7025,N_7192);
nand U7350 (N_7350,N_7093,N_7154);
and U7351 (N_7351,N_7112,N_7224);
nand U7352 (N_7352,N_7004,N_7177);
nand U7353 (N_7353,N_7065,N_7076);
nand U7354 (N_7354,N_7003,N_7032);
nor U7355 (N_7355,N_7033,N_7124);
xor U7356 (N_7356,N_7035,N_7170);
nand U7357 (N_7357,N_7001,N_7021);
nor U7358 (N_7358,N_7053,N_7012);
xor U7359 (N_7359,N_7056,N_7201);
nand U7360 (N_7360,N_7121,N_7148);
nor U7361 (N_7361,N_7205,N_7246);
or U7362 (N_7362,N_7111,N_7097);
or U7363 (N_7363,N_7179,N_7005);
nand U7364 (N_7364,N_7165,N_7152);
and U7365 (N_7365,N_7180,N_7141);
nand U7366 (N_7366,N_7006,N_7196);
nand U7367 (N_7367,N_7157,N_7064);
and U7368 (N_7368,N_7211,N_7104);
nand U7369 (N_7369,N_7181,N_7024);
and U7370 (N_7370,N_7098,N_7221);
and U7371 (N_7371,N_7230,N_7163);
and U7372 (N_7372,N_7099,N_7218);
nand U7373 (N_7373,N_7085,N_7088);
nor U7374 (N_7374,N_7193,N_7044);
or U7375 (N_7375,N_7151,N_7104);
nand U7376 (N_7376,N_7011,N_7089);
nand U7377 (N_7377,N_7053,N_7227);
nand U7378 (N_7378,N_7232,N_7111);
xnor U7379 (N_7379,N_7091,N_7200);
and U7380 (N_7380,N_7240,N_7161);
nor U7381 (N_7381,N_7058,N_7109);
nand U7382 (N_7382,N_7007,N_7153);
nor U7383 (N_7383,N_7051,N_7189);
and U7384 (N_7384,N_7248,N_7147);
xor U7385 (N_7385,N_7228,N_7098);
or U7386 (N_7386,N_7233,N_7239);
and U7387 (N_7387,N_7174,N_7128);
xnor U7388 (N_7388,N_7063,N_7000);
xor U7389 (N_7389,N_7046,N_7167);
or U7390 (N_7390,N_7209,N_7092);
and U7391 (N_7391,N_7039,N_7220);
and U7392 (N_7392,N_7028,N_7231);
or U7393 (N_7393,N_7205,N_7133);
and U7394 (N_7394,N_7006,N_7189);
xor U7395 (N_7395,N_7048,N_7012);
nand U7396 (N_7396,N_7211,N_7111);
xnor U7397 (N_7397,N_7123,N_7063);
and U7398 (N_7398,N_7107,N_7141);
xor U7399 (N_7399,N_7164,N_7075);
nand U7400 (N_7400,N_7108,N_7036);
xor U7401 (N_7401,N_7196,N_7130);
nor U7402 (N_7402,N_7155,N_7218);
and U7403 (N_7403,N_7044,N_7136);
xor U7404 (N_7404,N_7244,N_7187);
nor U7405 (N_7405,N_7246,N_7115);
nor U7406 (N_7406,N_7055,N_7082);
and U7407 (N_7407,N_7163,N_7207);
nor U7408 (N_7408,N_7034,N_7091);
nand U7409 (N_7409,N_7211,N_7223);
or U7410 (N_7410,N_7019,N_7129);
nor U7411 (N_7411,N_7218,N_7189);
nor U7412 (N_7412,N_7195,N_7139);
and U7413 (N_7413,N_7224,N_7219);
xnor U7414 (N_7414,N_7057,N_7157);
xor U7415 (N_7415,N_7154,N_7084);
or U7416 (N_7416,N_7109,N_7140);
nand U7417 (N_7417,N_7060,N_7089);
and U7418 (N_7418,N_7052,N_7071);
and U7419 (N_7419,N_7138,N_7232);
nand U7420 (N_7420,N_7218,N_7045);
xor U7421 (N_7421,N_7208,N_7195);
nand U7422 (N_7422,N_7223,N_7209);
or U7423 (N_7423,N_7032,N_7031);
nor U7424 (N_7424,N_7162,N_7068);
nand U7425 (N_7425,N_7072,N_7166);
or U7426 (N_7426,N_7213,N_7217);
and U7427 (N_7427,N_7241,N_7071);
nor U7428 (N_7428,N_7007,N_7116);
nor U7429 (N_7429,N_7015,N_7064);
xnor U7430 (N_7430,N_7122,N_7231);
xor U7431 (N_7431,N_7034,N_7007);
and U7432 (N_7432,N_7142,N_7147);
or U7433 (N_7433,N_7123,N_7160);
xnor U7434 (N_7434,N_7194,N_7038);
nand U7435 (N_7435,N_7056,N_7046);
nand U7436 (N_7436,N_7100,N_7021);
nand U7437 (N_7437,N_7016,N_7213);
xor U7438 (N_7438,N_7133,N_7167);
and U7439 (N_7439,N_7100,N_7058);
nor U7440 (N_7440,N_7151,N_7222);
xor U7441 (N_7441,N_7114,N_7165);
nor U7442 (N_7442,N_7111,N_7086);
or U7443 (N_7443,N_7238,N_7200);
or U7444 (N_7444,N_7031,N_7095);
nand U7445 (N_7445,N_7169,N_7078);
and U7446 (N_7446,N_7151,N_7123);
or U7447 (N_7447,N_7009,N_7221);
xnor U7448 (N_7448,N_7037,N_7147);
xor U7449 (N_7449,N_7146,N_7181);
nand U7450 (N_7450,N_7163,N_7107);
nand U7451 (N_7451,N_7014,N_7166);
and U7452 (N_7452,N_7090,N_7248);
nand U7453 (N_7453,N_7080,N_7239);
nand U7454 (N_7454,N_7064,N_7034);
and U7455 (N_7455,N_7118,N_7065);
nand U7456 (N_7456,N_7026,N_7088);
and U7457 (N_7457,N_7148,N_7028);
nand U7458 (N_7458,N_7053,N_7197);
nor U7459 (N_7459,N_7055,N_7122);
nor U7460 (N_7460,N_7218,N_7165);
xor U7461 (N_7461,N_7145,N_7179);
nand U7462 (N_7462,N_7055,N_7047);
nand U7463 (N_7463,N_7184,N_7016);
and U7464 (N_7464,N_7178,N_7080);
nand U7465 (N_7465,N_7102,N_7018);
nor U7466 (N_7466,N_7104,N_7230);
or U7467 (N_7467,N_7065,N_7119);
or U7468 (N_7468,N_7220,N_7150);
xor U7469 (N_7469,N_7211,N_7177);
and U7470 (N_7470,N_7181,N_7147);
or U7471 (N_7471,N_7033,N_7051);
nand U7472 (N_7472,N_7001,N_7125);
xor U7473 (N_7473,N_7196,N_7025);
nand U7474 (N_7474,N_7015,N_7008);
and U7475 (N_7475,N_7019,N_7124);
xnor U7476 (N_7476,N_7057,N_7127);
nand U7477 (N_7477,N_7240,N_7154);
and U7478 (N_7478,N_7043,N_7080);
xnor U7479 (N_7479,N_7031,N_7215);
xnor U7480 (N_7480,N_7163,N_7007);
nand U7481 (N_7481,N_7223,N_7114);
and U7482 (N_7482,N_7103,N_7093);
and U7483 (N_7483,N_7222,N_7195);
xor U7484 (N_7484,N_7242,N_7083);
xnor U7485 (N_7485,N_7202,N_7032);
xnor U7486 (N_7486,N_7059,N_7092);
or U7487 (N_7487,N_7084,N_7246);
and U7488 (N_7488,N_7080,N_7190);
nand U7489 (N_7489,N_7242,N_7102);
nor U7490 (N_7490,N_7203,N_7127);
xor U7491 (N_7491,N_7092,N_7158);
nand U7492 (N_7492,N_7104,N_7041);
or U7493 (N_7493,N_7163,N_7030);
nor U7494 (N_7494,N_7061,N_7163);
nand U7495 (N_7495,N_7067,N_7215);
nor U7496 (N_7496,N_7219,N_7095);
and U7497 (N_7497,N_7064,N_7104);
and U7498 (N_7498,N_7217,N_7104);
or U7499 (N_7499,N_7031,N_7223);
xnor U7500 (N_7500,N_7299,N_7289);
nor U7501 (N_7501,N_7274,N_7281);
nor U7502 (N_7502,N_7444,N_7447);
nand U7503 (N_7503,N_7341,N_7431);
or U7504 (N_7504,N_7441,N_7414);
and U7505 (N_7505,N_7352,N_7458);
and U7506 (N_7506,N_7297,N_7305);
and U7507 (N_7507,N_7300,N_7307);
and U7508 (N_7508,N_7373,N_7379);
xor U7509 (N_7509,N_7446,N_7495);
or U7510 (N_7510,N_7287,N_7467);
xnor U7511 (N_7511,N_7426,N_7275);
or U7512 (N_7512,N_7321,N_7420);
nand U7513 (N_7513,N_7423,N_7437);
xnor U7514 (N_7514,N_7354,N_7417);
nor U7515 (N_7515,N_7416,N_7377);
or U7516 (N_7516,N_7427,N_7291);
nor U7517 (N_7517,N_7293,N_7366);
nor U7518 (N_7518,N_7466,N_7445);
nor U7519 (N_7519,N_7360,N_7484);
or U7520 (N_7520,N_7361,N_7311);
and U7521 (N_7521,N_7411,N_7255);
nand U7522 (N_7522,N_7481,N_7272);
nand U7523 (N_7523,N_7319,N_7451);
and U7524 (N_7524,N_7418,N_7348);
and U7525 (N_7525,N_7276,N_7488);
and U7526 (N_7526,N_7318,N_7372);
and U7527 (N_7527,N_7415,N_7455);
nor U7528 (N_7528,N_7256,N_7257);
nor U7529 (N_7529,N_7357,N_7324);
nor U7530 (N_7530,N_7286,N_7363);
and U7531 (N_7531,N_7489,N_7265);
xnor U7532 (N_7532,N_7302,N_7296);
and U7533 (N_7533,N_7421,N_7497);
xnor U7534 (N_7534,N_7351,N_7483);
xnor U7535 (N_7535,N_7252,N_7422);
and U7536 (N_7536,N_7261,N_7337);
and U7537 (N_7537,N_7380,N_7464);
nand U7538 (N_7538,N_7450,N_7314);
nand U7539 (N_7539,N_7432,N_7388);
nand U7540 (N_7540,N_7442,N_7453);
or U7541 (N_7541,N_7264,N_7387);
and U7542 (N_7542,N_7438,N_7457);
xnor U7543 (N_7543,N_7381,N_7374);
or U7544 (N_7544,N_7315,N_7350);
xnor U7545 (N_7545,N_7408,N_7413);
or U7546 (N_7546,N_7402,N_7498);
nor U7547 (N_7547,N_7294,N_7430);
xnor U7548 (N_7548,N_7303,N_7283);
nor U7549 (N_7549,N_7460,N_7340);
or U7550 (N_7550,N_7353,N_7344);
or U7551 (N_7551,N_7384,N_7449);
nand U7552 (N_7552,N_7269,N_7439);
nor U7553 (N_7553,N_7277,N_7270);
nand U7554 (N_7554,N_7273,N_7356);
xnor U7555 (N_7555,N_7371,N_7267);
nor U7556 (N_7556,N_7382,N_7399);
xor U7557 (N_7557,N_7262,N_7309);
xor U7558 (N_7558,N_7436,N_7428);
xnor U7559 (N_7559,N_7364,N_7469);
or U7560 (N_7560,N_7345,N_7346);
or U7561 (N_7561,N_7339,N_7260);
nor U7562 (N_7562,N_7429,N_7409);
xnor U7563 (N_7563,N_7288,N_7280);
or U7564 (N_7564,N_7312,N_7338);
nand U7565 (N_7565,N_7390,N_7347);
xnor U7566 (N_7566,N_7395,N_7478);
nand U7567 (N_7567,N_7448,N_7474);
and U7568 (N_7568,N_7285,N_7349);
nand U7569 (N_7569,N_7394,N_7365);
nand U7570 (N_7570,N_7326,N_7266);
xor U7571 (N_7571,N_7471,N_7391);
or U7572 (N_7572,N_7330,N_7492);
xor U7573 (N_7573,N_7325,N_7425);
and U7574 (N_7574,N_7486,N_7343);
or U7575 (N_7575,N_7462,N_7468);
nand U7576 (N_7576,N_7434,N_7459);
nand U7577 (N_7577,N_7412,N_7392);
nor U7578 (N_7578,N_7393,N_7298);
or U7579 (N_7579,N_7320,N_7494);
or U7580 (N_7580,N_7463,N_7403);
nand U7581 (N_7581,N_7383,N_7396);
nor U7582 (N_7582,N_7443,N_7473);
nor U7583 (N_7583,N_7499,N_7490);
xor U7584 (N_7584,N_7331,N_7477);
nor U7585 (N_7585,N_7358,N_7284);
or U7586 (N_7586,N_7342,N_7476);
nor U7587 (N_7587,N_7496,N_7355);
nor U7588 (N_7588,N_7475,N_7435);
nand U7589 (N_7589,N_7317,N_7323);
nand U7590 (N_7590,N_7322,N_7398);
or U7591 (N_7591,N_7310,N_7278);
xor U7592 (N_7592,N_7406,N_7452);
nor U7593 (N_7593,N_7279,N_7461);
nor U7594 (N_7594,N_7316,N_7250);
xnor U7595 (N_7595,N_7465,N_7359);
nand U7596 (N_7596,N_7405,N_7487);
xor U7597 (N_7597,N_7301,N_7410);
xor U7598 (N_7598,N_7386,N_7304);
xor U7599 (N_7599,N_7424,N_7268);
xor U7600 (N_7600,N_7389,N_7327);
nand U7601 (N_7601,N_7254,N_7368);
or U7602 (N_7602,N_7440,N_7329);
xnor U7603 (N_7603,N_7454,N_7400);
nor U7604 (N_7604,N_7328,N_7369);
xor U7605 (N_7605,N_7306,N_7282);
or U7606 (N_7606,N_7308,N_7433);
nand U7607 (N_7607,N_7378,N_7407);
nand U7608 (N_7608,N_7385,N_7401);
nor U7609 (N_7609,N_7259,N_7292);
or U7610 (N_7610,N_7470,N_7313);
and U7611 (N_7611,N_7485,N_7271);
nor U7612 (N_7612,N_7295,N_7370);
nor U7613 (N_7613,N_7251,N_7332);
or U7614 (N_7614,N_7419,N_7258);
or U7615 (N_7615,N_7335,N_7290);
xor U7616 (N_7616,N_7479,N_7336);
nor U7617 (N_7617,N_7375,N_7472);
and U7618 (N_7618,N_7376,N_7367);
and U7619 (N_7619,N_7253,N_7333);
or U7620 (N_7620,N_7491,N_7404);
or U7621 (N_7621,N_7334,N_7456);
or U7622 (N_7622,N_7480,N_7362);
xor U7623 (N_7623,N_7263,N_7482);
xor U7624 (N_7624,N_7493,N_7397);
or U7625 (N_7625,N_7478,N_7336);
or U7626 (N_7626,N_7357,N_7270);
and U7627 (N_7627,N_7402,N_7290);
nor U7628 (N_7628,N_7302,N_7389);
and U7629 (N_7629,N_7467,N_7376);
xnor U7630 (N_7630,N_7251,N_7492);
nor U7631 (N_7631,N_7335,N_7446);
nand U7632 (N_7632,N_7345,N_7293);
or U7633 (N_7633,N_7416,N_7251);
and U7634 (N_7634,N_7411,N_7261);
nor U7635 (N_7635,N_7338,N_7348);
nand U7636 (N_7636,N_7456,N_7296);
nand U7637 (N_7637,N_7300,N_7348);
xnor U7638 (N_7638,N_7428,N_7364);
nand U7639 (N_7639,N_7430,N_7480);
xor U7640 (N_7640,N_7474,N_7312);
and U7641 (N_7641,N_7498,N_7281);
or U7642 (N_7642,N_7470,N_7445);
or U7643 (N_7643,N_7454,N_7435);
and U7644 (N_7644,N_7258,N_7262);
and U7645 (N_7645,N_7348,N_7265);
xor U7646 (N_7646,N_7343,N_7422);
nand U7647 (N_7647,N_7311,N_7359);
nand U7648 (N_7648,N_7417,N_7498);
or U7649 (N_7649,N_7314,N_7480);
and U7650 (N_7650,N_7339,N_7257);
and U7651 (N_7651,N_7271,N_7391);
nor U7652 (N_7652,N_7306,N_7351);
xor U7653 (N_7653,N_7450,N_7259);
or U7654 (N_7654,N_7266,N_7260);
and U7655 (N_7655,N_7404,N_7311);
and U7656 (N_7656,N_7283,N_7368);
nor U7657 (N_7657,N_7433,N_7421);
and U7658 (N_7658,N_7327,N_7257);
xnor U7659 (N_7659,N_7337,N_7440);
nor U7660 (N_7660,N_7435,N_7264);
nand U7661 (N_7661,N_7402,N_7496);
nor U7662 (N_7662,N_7331,N_7279);
nand U7663 (N_7663,N_7492,N_7457);
or U7664 (N_7664,N_7304,N_7359);
and U7665 (N_7665,N_7438,N_7297);
and U7666 (N_7666,N_7457,N_7387);
and U7667 (N_7667,N_7283,N_7392);
or U7668 (N_7668,N_7291,N_7326);
xnor U7669 (N_7669,N_7427,N_7411);
nor U7670 (N_7670,N_7484,N_7367);
or U7671 (N_7671,N_7365,N_7460);
or U7672 (N_7672,N_7468,N_7370);
xnor U7673 (N_7673,N_7464,N_7393);
nor U7674 (N_7674,N_7490,N_7414);
xnor U7675 (N_7675,N_7308,N_7447);
and U7676 (N_7676,N_7460,N_7418);
nor U7677 (N_7677,N_7351,N_7337);
nand U7678 (N_7678,N_7482,N_7396);
or U7679 (N_7679,N_7322,N_7453);
nor U7680 (N_7680,N_7390,N_7337);
nand U7681 (N_7681,N_7434,N_7485);
nand U7682 (N_7682,N_7425,N_7252);
nor U7683 (N_7683,N_7362,N_7267);
xnor U7684 (N_7684,N_7336,N_7306);
nand U7685 (N_7685,N_7294,N_7408);
nand U7686 (N_7686,N_7455,N_7438);
xor U7687 (N_7687,N_7284,N_7357);
or U7688 (N_7688,N_7305,N_7417);
and U7689 (N_7689,N_7479,N_7490);
nand U7690 (N_7690,N_7339,N_7353);
nand U7691 (N_7691,N_7366,N_7425);
nor U7692 (N_7692,N_7362,N_7471);
nor U7693 (N_7693,N_7297,N_7292);
nor U7694 (N_7694,N_7349,N_7473);
xnor U7695 (N_7695,N_7479,N_7488);
xor U7696 (N_7696,N_7490,N_7309);
xor U7697 (N_7697,N_7494,N_7363);
xnor U7698 (N_7698,N_7273,N_7307);
nand U7699 (N_7699,N_7340,N_7363);
and U7700 (N_7700,N_7316,N_7306);
xor U7701 (N_7701,N_7472,N_7497);
or U7702 (N_7702,N_7273,N_7461);
and U7703 (N_7703,N_7323,N_7465);
nand U7704 (N_7704,N_7424,N_7383);
or U7705 (N_7705,N_7324,N_7379);
nor U7706 (N_7706,N_7311,N_7348);
nand U7707 (N_7707,N_7431,N_7401);
nor U7708 (N_7708,N_7462,N_7378);
nand U7709 (N_7709,N_7401,N_7425);
or U7710 (N_7710,N_7387,N_7468);
or U7711 (N_7711,N_7306,N_7285);
nor U7712 (N_7712,N_7490,N_7487);
or U7713 (N_7713,N_7372,N_7338);
nor U7714 (N_7714,N_7471,N_7469);
nand U7715 (N_7715,N_7414,N_7422);
nor U7716 (N_7716,N_7333,N_7476);
nor U7717 (N_7717,N_7473,N_7404);
and U7718 (N_7718,N_7323,N_7257);
nor U7719 (N_7719,N_7379,N_7309);
nor U7720 (N_7720,N_7320,N_7445);
xnor U7721 (N_7721,N_7359,N_7284);
xnor U7722 (N_7722,N_7302,N_7256);
nor U7723 (N_7723,N_7464,N_7398);
xnor U7724 (N_7724,N_7433,N_7385);
xnor U7725 (N_7725,N_7411,N_7426);
xnor U7726 (N_7726,N_7437,N_7289);
and U7727 (N_7727,N_7399,N_7317);
xnor U7728 (N_7728,N_7346,N_7426);
xor U7729 (N_7729,N_7457,N_7298);
and U7730 (N_7730,N_7459,N_7356);
and U7731 (N_7731,N_7473,N_7438);
and U7732 (N_7732,N_7356,N_7337);
or U7733 (N_7733,N_7424,N_7251);
nand U7734 (N_7734,N_7437,N_7367);
and U7735 (N_7735,N_7280,N_7460);
nor U7736 (N_7736,N_7283,N_7432);
or U7737 (N_7737,N_7417,N_7441);
xor U7738 (N_7738,N_7385,N_7354);
xor U7739 (N_7739,N_7499,N_7292);
nor U7740 (N_7740,N_7450,N_7262);
nand U7741 (N_7741,N_7420,N_7374);
or U7742 (N_7742,N_7307,N_7442);
nand U7743 (N_7743,N_7339,N_7350);
and U7744 (N_7744,N_7350,N_7255);
nor U7745 (N_7745,N_7393,N_7460);
and U7746 (N_7746,N_7461,N_7456);
or U7747 (N_7747,N_7442,N_7456);
or U7748 (N_7748,N_7466,N_7477);
or U7749 (N_7749,N_7270,N_7487);
nand U7750 (N_7750,N_7646,N_7736);
nand U7751 (N_7751,N_7529,N_7615);
or U7752 (N_7752,N_7732,N_7623);
or U7753 (N_7753,N_7639,N_7579);
nor U7754 (N_7754,N_7525,N_7590);
nor U7755 (N_7755,N_7747,N_7628);
nand U7756 (N_7756,N_7500,N_7541);
nor U7757 (N_7757,N_7511,N_7563);
or U7758 (N_7758,N_7620,N_7575);
xnor U7759 (N_7759,N_7567,N_7634);
or U7760 (N_7760,N_7692,N_7560);
and U7761 (N_7761,N_7721,N_7506);
or U7762 (N_7762,N_7656,N_7641);
and U7763 (N_7763,N_7509,N_7657);
or U7764 (N_7764,N_7740,N_7562);
and U7765 (N_7765,N_7696,N_7532);
and U7766 (N_7766,N_7561,N_7543);
xor U7767 (N_7767,N_7688,N_7717);
nor U7768 (N_7768,N_7501,N_7533);
nor U7769 (N_7769,N_7719,N_7573);
or U7770 (N_7770,N_7733,N_7699);
and U7771 (N_7771,N_7606,N_7654);
or U7772 (N_7772,N_7691,N_7706);
or U7773 (N_7773,N_7693,N_7664);
nor U7774 (N_7774,N_7528,N_7516);
nand U7775 (N_7775,N_7743,N_7748);
nor U7776 (N_7776,N_7652,N_7546);
and U7777 (N_7777,N_7660,N_7683);
and U7778 (N_7778,N_7724,N_7678);
or U7779 (N_7779,N_7520,N_7666);
nand U7780 (N_7780,N_7582,N_7645);
nand U7781 (N_7781,N_7596,N_7648);
and U7782 (N_7782,N_7745,N_7653);
nor U7783 (N_7783,N_7507,N_7526);
nand U7784 (N_7784,N_7588,N_7597);
and U7785 (N_7785,N_7714,N_7744);
nor U7786 (N_7786,N_7647,N_7749);
or U7787 (N_7787,N_7594,N_7508);
nand U7788 (N_7788,N_7536,N_7662);
xor U7789 (N_7789,N_7503,N_7576);
nand U7790 (N_7790,N_7504,N_7684);
nand U7791 (N_7791,N_7604,N_7517);
nand U7792 (N_7792,N_7672,N_7589);
and U7793 (N_7793,N_7668,N_7535);
nand U7794 (N_7794,N_7627,N_7534);
nor U7795 (N_7795,N_7711,N_7669);
xnor U7796 (N_7796,N_7544,N_7713);
or U7797 (N_7797,N_7554,N_7559);
or U7798 (N_7798,N_7605,N_7515);
and U7799 (N_7799,N_7549,N_7607);
and U7800 (N_7800,N_7734,N_7695);
and U7801 (N_7801,N_7551,N_7531);
and U7802 (N_7802,N_7524,N_7737);
and U7803 (N_7803,N_7651,N_7626);
nand U7804 (N_7804,N_7568,N_7587);
or U7805 (N_7805,N_7742,N_7694);
or U7806 (N_7806,N_7581,N_7540);
nand U7807 (N_7807,N_7512,N_7655);
xnor U7808 (N_7808,N_7722,N_7697);
or U7809 (N_7809,N_7636,N_7704);
nor U7810 (N_7810,N_7618,N_7595);
or U7811 (N_7811,N_7518,N_7608);
and U7812 (N_7812,N_7601,N_7710);
nand U7813 (N_7813,N_7505,N_7539);
nand U7814 (N_7814,N_7550,N_7632);
or U7815 (N_7815,N_7616,N_7663);
or U7816 (N_7816,N_7730,N_7661);
or U7817 (N_7817,N_7557,N_7591);
xnor U7818 (N_7818,N_7746,N_7671);
or U7819 (N_7819,N_7705,N_7552);
xor U7820 (N_7820,N_7726,N_7675);
xnor U7821 (N_7821,N_7545,N_7708);
nor U7822 (N_7822,N_7592,N_7553);
xnor U7823 (N_7823,N_7580,N_7718);
and U7824 (N_7824,N_7735,N_7725);
and U7825 (N_7825,N_7603,N_7586);
and U7826 (N_7826,N_7502,N_7622);
xor U7827 (N_7827,N_7723,N_7679);
xnor U7828 (N_7828,N_7670,N_7658);
and U7829 (N_7829,N_7583,N_7599);
nand U7830 (N_7830,N_7566,N_7523);
nor U7831 (N_7831,N_7677,N_7538);
and U7832 (N_7832,N_7709,N_7625);
xor U7833 (N_7833,N_7619,N_7598);
nor U7834 (N_7834,N_7667,N_7585);
xnor U7835 (N_7835,N_7635,N_7558);
nand U7836 (N_7836,N_7637,N_7701);
or U7837 (N_7837,N_7687,N_7681);
nor U7838 (N_7838,N_7703,N_7680);
or U7839 (N_7839,N_7715,N_7514);
and U7840 (N_7840,N_7689,N_7676);
xnor U7841 (N_7841,N_7624,N_7642);
nand U7842 (N_7842,N_7584,N_7665);
nor U7843 (N_7843,N_7633,N_7612);
or U7844 (N_7844,N_7731,N_7690);
and U7845 (N_7845,N_7547,N_7659);
nor U7846 (N_7846,N_7593,N_7542);
nand U7847 (N_7847,N_7611,N_7577);
and U7848 (N_7848,N_7537,N_7530);
or U7849 (N_7849,N_7513,N_7548);
nor U7850 (N_7850,N_7700,N_7673);
xor U7851 (N_7851,N_7519,N_7527);
or U7852 (N_7852,N_7686,N_7614);
or U7853 (N_7853,N_7738,N_7564);
nor U7854 (N_7854,N_7610,N_7720);
nor U7855 (N_7855,N_7650,N_7729);
or U7856 (N_7856,N_7682,N_7613);
or U7857 (N_7857,N_7521,N_7571);
or U7858 (N_7858,N_7727,N_7707);
and U7859 (N_7859,N_7510,N_7522);
and U7860 (N_7860,N_7698,N_7570);
xnor U7861 (N_7861,N_7602,N_7572);
xnor U7862 (N_7862,N_7644,N_7728);
or U7863 (N_7863,N_7578,N_7685);
nand U7864 (N_7864,N_7630,N_7716);
nand U7865 (N_7865,N_7712,N_7569);
nand U7866 (N_7866,N_7617,N_7649);
nand U7867 (N_7867,N_7555,N_7643);
or U7868 (N_7868,N_7556,N_7640);
xnor U7869 (N_7869,N_7702,N_7674);
xor U7870 (N_7870,N_7600,N_7631);
nand U7871 (N_7871,N_7565,N_7638);
xnor U7872 (N_7872,N_7739,N_7609);
or U7873 (N_7873,N_7621,N_7629);
nor U7874 (N_7874,N_7741,N_7574);
nand U7875 (N_7875,N_7733,N_7532);
and U7876 (N_7876,N_7547,N_7539);
xor U7877 (N_7877,N_7743,N_7645);
nor U7878 (N_7878,N_7508,N_7580);
or U7879 (N_7879,N_7506,N_7562);
nand U7880 (N_7880,N_7708,N_7655);
xnor U7881 (N_7881,N_7605,N_7619);
and U7882 (N_7882,N_7571,N_7699);
and U7883 (N_7883,N_7749,N_7699);
and U7884 (N_7884,N_7664,N_7725);
or U7885 (N_7885,N_7615,N_7731);
or U7886 (N_7886,N_7637,N_7658);
and U7887 (N_7887,N_7706,N_7687);
or U7888 (N_7888,N_7715,N_7634);
nor U7889 (N_7889,N_7597,N_7725);
nor U7890 (N_7890,N_7662,N_7615);
nand U7891 (N_7891,N_7545,N_7673);
and U7892 (N_7892,N_7736,N_7606);
nand U7893 (N_7893,N_7711,N_7588);
nor U7894 (N_7894,N_7601,N_7642);
nor U7895 (N_7895,N_7579,N_7528);
nand U7896 (N_7896,N_7603,N_7684);
or U7897 (N_7897,N_7550,N_7659);
and U7898 (N_7898,N_7742,N_7566);
nand U7899 (N_7899,N_7524,N_7635);
and U7900 (N_7900,N_7597,N_7546);
and U7901 (N_7901,N_7707,N_7717);
nand U7902 (N_7902,N_7599,N_7624);
nor U7903 (N_7903,N_7559,N_7571);
nand U7904 (N_7904,N_7702,N_7668);
nand U7905 (N_7905,N_7691,N_7653);
or U7906 (N_7906,N_7501,N_7612);
or U7907 (N_7907,N_7554,N_7639);
xor U7908 (N_7908,N_7680,N_7577);
or U7909 (N_7909,N_7538,N_7660);
or U7910 (N_7910,N_7746,N_7646);
or U7911 (N_7911,N_7667,N_7560);
xnor U7912 (N_7912,N_7718,N_7656);
and U7913 (N_7913,N_7532,N_7546);
and U7914 (N_7914,N_7652,N_7709);
nor U7915 (N_7915,N_7592,N_7608);
or U7916 (N_7916,N_7576,N_7736);
nand U7917 (N_7917,N_7747,N_7676);
and U7918 (N_7918,N_7652,N_7668);
xor U7919 (N_7919,N_7736,N_7687);
and U7920 (N_7920,N_7737,N_7501);
and U7921 (N_7921,N_7741,N_7583);
or U7922 (N_7922,N_7647,N_7695);
and U7923 (N_7923,N_7658,N_7676);
or U7924 (N_7924,N_7515,N_7683);
nor U7925 (N_7925,N_7501,N_7728);
nand U7926 (N_7926,N_7607,N_7721);
xor U7927 (N_7927,N_7627,N_7551);
nand U7928 (N_7928,N_7522,N_7584);
and U7929 (N_7929,N_7506,N_7719);
and U7930 (N_7930,N_7698,N_7715);
nand U7931 (N_7931,N_7645,N_7700);
or U7932 (N_7932,N_7668,N_7547);
or U7933 (N_7933,N_7589,N_7675);
nor U7934 (N_7934,N_7717,N_7742);
xnor U7935 (N_7935,N_7655,N_7566);
or U7936 (N_7936,N_7654,N_7662);
or U7937 (N_7937,N_7741,N_7558);
or U7938 (N_7938,N_7684,N_7506);
nor U7939 (N_7939,N_7559,N_7619);
and U7940 (N_7940,N_7672,N_7593);
nand U7941 (N_7941,N_7638,N_7513);
or U7942 (N_7942,N_7697,N_7695);
nand U7943 (N_7943,N_7681,N_7551);
nor U7944 (N_7944,N_7679,N_7741);
and U7945 (N_7945,N_7731,N_7522);
xor U7946 (N_7946,N_7554,N_7685);
and U7947 (N_7947,N_7578,N_7629);
xnor U7948 (N_7948,N_7626,N_7694);
or U7949 (N_7949,N_7512,N_7625);
nor U7950 (N_7950,N_7718,N_7501);
xor U7951 (N_7951,N_7662,N_7653);
nand U7952 (N_7952,N_7505,N_7715);
nor U7953 (N_7953,N_7681,N_7619);
nand U7954 (N_7954,N_7552,N_7697);
xor U7955 (N_7955,N_7747,N_7589);
nor U7956 (N_7956,N_7580,N_7677);
or U7957 (N_7957,N_7728,N_7566);
and U7958 (N_7958,N_7653,N_7698);
nor U7959 (N_7959,N_7513,N_7645);
nor U7960 (N_7960,N_7709,N_7514);
xnor U7961 (N_7961,N_7728,N_7726);
nand U7962 (N_7962,N_7579,N_7611);
xor U7963 (N_7963,N_7601,N_7549);
and U7964 (N_7964,N_7732,N_7605);
xnor U7965 (N_7965,N_7563,N_7578);
nand U7966 (N_7966,N_7582,N_7633);
xnor U7967 (N_7967,N_7537,N_7703);
and U7968 (N_7968,N_7681,N_7719);
nand U7969 (N_7969,N_7715,N_7648);
and U7970 (N_7970,N_7666,N_7714);
and U7971 (N_7971,N_7713,N_7664);
nand U7972 (N_7972,N_7644,N_7632);
and U7973 (N_7973,N_7605,N_7567);
xor U7974 (N_7974,N_7552,N_7533);
nor U7975 (N_7975,N_7656,N_7686);
nor U7976 (N_7976,N_7638,N_7739);
nor U7977 (N_7977,N_7732,N_7518);
or U7978 (N_7978,N_7630,N_7574);
nor U7979 (N_7979,N_7721,N_7675);
and U7980 (N_7980,N_7587,N_7550);
or U7981 (N_7981,N_7652,N_7679);
or U7982 (N_7982,N_7512,N_7583);
xor U7983 (N_7983,N_7654,N_7699);
nor U7984 (N_7984,N_7560,N_7634);
xnor U7985 (N_7985,N_7669,N_7732);
xor U7986 (N_7986,N_7662,N_7506);
nand U7987 (N_7987,N_7527,N_7630);
or U7988 (N_7988,N_7701,N_7715);
and U7989 (N_7989,N_7501,N_7747);
or U7990 (N_7990,N_7614,N_7729);
and U7991 (N_7991,N_7532,N_7564);
nand U7992 (N_7992,N_7623,N_7590);
xnor U7993 (N_7993,N_7698,N_7747);
xnor U7994 (N_7994,N_7557,N_7541);
nand U7995 (N_7995,N_7653,N_7724);
or U7996 (N_7996,N_7682,N_7524);
or U7997 (N_7997,N_7588,N_7604);
and U7998 (N_7998,N_7569,N_7621);
nor U7999 (N_7999,N_7723,N_7580);
nand U8000 (N_8000,N_7770,N_7850);
or U8001 (N_8001,N_7824,N_7844);
nor U8002 (N_8002,N_7835,N_7771);
nand U8003 (N_8003,N_7934,N_7952);
nor U8004 (N_8004,N_7906,N_7759);
and U8005 (N_8005,N_7888,N_7860);
nor U8006 (N_8006,N_7983,N_7796);
nor U8007 (N_8007,N_7892,N_7955);
or U8008 (N_8008,N_7830,N_7876);
and U8009 (N_8009,N_7994,N_7772);
xnor U8010 (N_8010,N_7811,N_7899);
nor U8011 (N_8011,N_7935,N_7886);
nand U8012 (N_8012,N_7942,N_7808);
xor U8013 (N_8013,N_7853,N_7848);
nand U8014 (N_8014,N_7962,N_7982);
nor U8015 (N_8015,N_7863,N_7800);
nand U8016 (N_8016,N_7907,N_7946);
or U8017 (N_8017,N_7857,N_7929);
xor U8018 (N_8018,N_7949,N_7838);
xnor U8019 (N_8019,N_7924,N_7862);
xnor U8020 (N_8020,N_7781,N_7993);
nor U8021 (N_8021,N_7939,N_7856);
nand U8022 (N_8022,N_7768,N_7883);
and U8023 (N_8023,N_7938,N_7865);
or U8024 (N_8024,N_7911,N_7843);
xor U8025 (N_8025,N_7918,N_7902);
nand U8026 (N_8026,N_7915,N_7933);
and U8027 (N_8027,N_7976,N_7973);
or U8028 (N_8028,N_7867,N_7917);
nor U8029 (N_8029,N_7943,N_7782);
nor U8030 (N_8030,N_7926,N_7836);
xnor U8031 (N_8031,N_7941,N_7971);
nand U8032 (N_8032,N_7990,N_7810);
nor U8033 (N_8033,N_7769,N_7931);
nor U8034 (N_8034,N_7947,N_7777);
nand U8035 (N_8035,N_7855,N_7871);
xor U8036 (N_8036,N_7995,N_7847);
xor U8037 (N_8037,N_7859,N_7984);
and U8038 (N_8038,N_7783,N_7903);
nor U8039 (N_8039,N_7758,N_7951);
xnor U8040 (N_8040,N_7764,N_7980);
xnor U8041 (N_8041,N_7922,N_7798);
or U8042 (N_8042,N_7760,N_7870);
and U8043 (N_8043,N_7750,N_7755);
and U8044 (N_8044,N_7972,N_7937);
xnor U8045 (N_8045,N_7891,N_7818);
nor U8046 (N_8046,N_7936,N_7900);
nand U8047 (N_8047,N_7928,N_7839);
nand U8048 (N_8048,N_7961,N_7894);
nand U8049 (N_8049,N_7914,N_7958);
nand U8050 (N_8050,N_7767,N_7794);
xor U8051 (N_8051,N_7812,N_7889);
nand U8052 (N_8052,N_7877,N_7775);
nand U8053 (N_8053,N_7806,N_7979);
or U8054 (N_8054,N_7908,N_7967);
nand U8055 (N_8055,N_7997,N_7815);
xor U8056 (N_8056,N_7920,N_7807);
nand U8057 (N_8057,N_7968,N_7765);
xor U8058 (N_8058,N_7895,N_7991);
nand U8059 (N_8059,N_7868,N_7791);
nor U8060 (N_8060,N_7978,N_7981);
nor U8061 (N_8061,N_7773,N_7956);
xnor U8062 (N_8062,N_7778,N_7814);
and U8063 (N_8063,N_7905,N_7989);
or U8064 (N_8064,N_7802,N_7963);
or U8065 (N_8065,N_7837,N_7885);
or U8066 (N_8066,N_7826,N_7756);
nand U8067 (N_8067,N_7959,N_7854);
nand U8068 (N_8068,N_7784,N_7998);
nand U8069 (N_8069,N_7884,N_7825);
nor U8070 (N_8070,N_7817,N_7823);
and U8071 (N_8071,N_7785,N_7801);
nor U8072 (N_8072,N_7923,N_7790);
nand U8073 (N_8073,N_7864,N_7831);
xor U8074 (N_8074,N_7833,N_7988);
nor U8075 (N_8075,N_7845,N_7879);
xnor U8076 (N_8076,N_7927,N_7913);
nand U8077 (N_8077,N_7851,N_7992);
and U8078 (N_8078,N_7819,N_7919);
nor U8079 (N_8079,N_7893,N_7799);
nor U8080 (N_8080,N_7762,N_7809);
and U8081 (N_8081,N_7820,N_7897);
and U8082 (N_8082,N_7869,N_7986);
xnor U8083 (N_8083,N_7950,N_7852);
xnor U8084 (N_8084,N_7912,N_7930);
or U8085 (N_8085,N_7803,N_7829);
and U8086 (N_8086,N_7880,N_7987);
and U8087 (N_8087,N_7896,N_7975);
or U8088 (N_8088,N_7948,N_7954);
nor U8089 (N_8089,N_7858,N_7916);
or U8090 (N_8090,N_7828,N_7834);
nor U8091 (N_8091,N_7925,N_7813);
nand U8092 (N_8092,N_7763,N_7872);
nor U8093 (N_8093,N_7953,N_7754);
nor U8094 (N_8094,N_7985,N_7804);
nor U8095 (N_8095,N_7932,N_7827);
xor U8096 (N_8096,N_7887,N_7786);
nor U8097 (N_8097,N_7840,N_7874);
nand U8098 (N_8098,N_7761,N_7873);
and U8099 (N_8099,N_7752,N_7832);
and U8100 (N_8100,N_7977,N_7849);
nor U8101 (N_8101,N_7766,N_7910);
nand U8102 (N_8102,N_7821,N_7996);
and U8103 (N_8103,N_7898,N_7751);
nand U8104 (N_8104,N_7966,N_7957);
nor U8105 (N_8105,N_7793,N_7960);
or U8106 (N_8106,N_7964,N_7999);
xor U8107 (N_8107,N_7816,N_7805);
and U8108 (N_8108,N_7878,N_7970);
nor U8109 (N_8109,N_7945,N_7757);
nor U8110 (N_8110,N_7822,N_7944);
nand U8111 (N_8111,N_7901,N_7787);
or U8112 (N_8112,N_7776,N_7792);
and U8113 (N_8113,N_7890,N_7753);
nor U8114 (N_8114,N_7921,N_7789);
nor U8115 (N_8115,N_7881,N_7861);
or U8116 (N_8116,N_7904,N_7774);
xor U8117 (N_8117,N_7779,N_7797);
xor U8118 (N_8118,N_7969,N_7909);
nor U8119 (N_8119,N_7965,N_7866);
or U8120 (N_8120,N_7882,N_7795);
or U8121 (N_8121,N_7788,N_7841);
xnor U8122 (N_8122,N_7846,N_7974);
or U8123 (N_8123,N_7842,N_7780);
xnor U8124 (N_8124,N_7875,N_7940);
and U8125 (N_8125,N_7927,N_7807);
nand U8126 (N_8126,N_7939,N_7868);
xor U8127 (N_8127,N_7903,N_7855);
or U8128 (N_8128,N_7904,N_7997);
or U8129 (N_8129,N_7937,N_7769);
and U8130 (N_8130,N_7897,N_7917);
nor U8131 (N_8131,N_7898,N_7947);
nor U8132 (N_8132,N_7963,N_7911);
nor U8133 (N_8133,N_7970,N_7949);
or U8134 (N_8134,N_7755,N_7811);
and U8135 (N_8135,N_7876,N_7887);
nand U8136 (N_8136,N_7879,N_7938);
nand U8137 (N_8137,N_7821,N_7797);
nor U8138 (N_8138,N_7875,N_7997);
and U8139 (N_8139,N_7962,N_7904);
nand U8140 (N_8140,N_7813,N_7894);
nand U8141 (N_8141,N_7848,N_7927);
xnor U8142 (N_8142,N_7974,N_7932);
nor U8143 (N_8143,N_7782,N_7975);
or U8144 (N_8144,N_7991,N_7859);
or U8145 (N_8145,N_7821,N_7872);
nor U8146 (N_8146,N_7942,N_7890);
or U8147 (N_8147,N_7915,N_7780);
xnor U8148 (N_8148,N_7807,N_7952);
and U8149 (N_8149,N_7912,N_7842);
and U8150 (N_8150,N_7955,N_7804);
or U8151 (N_8151,N_7964,N_7769);
nor U8152 (N_8152,N_7937,N_7875);
or U8153 (N_8153,N_7960,N_7771);
nand U8154 (N_8154,N_7829,N_7820);
nand U8155 (N_8155,N_7775,N_7994);
nand U8156 (N_8156,N_7792,N_7775);
and U8157 (N_8157,N_7805,N_7965);
or U8158 (N_8158,N_7847,N_7891);
nand U8159 (N_8159,N_7879,N_7794);
xor U8160 (N_8160,N_7898,N_7771);
nand U8161 (N_8161,N_7914,N_7842);
nand U8162 (N_8162,N_7783,N_7952);
or U8163 (N_8163,N_7995,N_7998);
nand U8164 (N_8164,N_7830,N_7805);
or U8165 (N_8165,N_7843,N_7808);
xnor U8166 (N_8166,N_7751,N_7994);
xor U8167 (N_8167,N_7869,N_7961);
nor U8168 (N_8168,N_7761,N_7837);
nand U8169 (N_8169,N_7854,N_7803);
nor U8170 (N_8170,N_7821,N_7896);
nor U8171 (N_8171,N_7993,N_7924);
xor U8172 (N_8172,N_7919,N_7836);
nor U8173 (N_8173,N_7956,N_7797);
or U8174 (N_8174,N_7826,N_7812);
nor U8175 (N_8175,N_7884,N_7912);
nor U8176 (N_8176,N_7831,N_7951);
xnor U8177 (N_8177,N_7835,N_7892);
nand U8178 (N_8178,N_7949,N_7984);
or U8179 (N_8179,N_7761,N_7801);
xor U8180 (N_8180,N_7768,N_7787);
nand U8181 (N_8181,N_7998,N_7935);
and U8182 (N_8182,N_7942,N_7889);
nor U8183 (N_8183,N_7822,N_7838);
nand U8184 (N_8184,N_7926,N_7959);
xor U8185 (N_8185,N_7767,N_7847);
or U8186 (N_8186,N_7903,N_7993);
xor U8187 (N_8187,N_7955,N_7861);
and U8188 (N_8188,N_7867,N_7861);
and U8189 (N_8189,N_7964,N_7761);
nor U8190 (N_8190,N_7853,N_7970);
or U8191 (N_8191,N_7871,N_7952);
nand U8192 (N_8192,N_7862,N_7766);
and U8193 (N_8193,N_7820,N_7863);
and U8194 (N_8194,N_7933,N_7819);
xnor U8195 (N_8195,N_7859,N_7751);
and U8196 (N_8196,N_7812,N_7902);
and U8197 (N_8197,N_7841,N_7935);
xnor U8198 (N_8198,N_7752,N_7925);
xnor U8199 (N_8199,N_7870,N_7765);
xor U8200 (N_8200,N_7883,N_7867);
xnor U8201 (N_8201,N_7831,N_7910);
xnor U8202 (N_8202,N_7976,N_7991);
nand U8203 (N_8203,N_7974,N_7761);
and U8204 (N_8204,N_7953,N_7945);
and U8205 (N_8205,N_7770,N_7767);
and U8206 (N_8206,N_7944,N_7829);
or U8207 (N_8207,N_7835,N_7972);
xor U8208 (N_8208,N_7758,N_7752);
or U8209 (N_8209,N_7950,N_7936);
nand U8210 (N_8210,N_7762,N_7900);
xnor U8211 (N_8211,N_7823,N_7824);
or U8212 (N_8212,N_7841,N_7942);
or U8213 (N_8213,N_7879,N_7842);
xnor U8214 (N_8214,N_7905,N_7779);
nor U8215 (N_8215,N_7864,N_7792);
and U8216 (N_8216,N_7809,N_7967);
nor U8217 (N_8217,N_7823,N_7797);
and U8218 (N_8218,N_7943,N_7871);
xor U8219 (N_8219,N_7857,N_7760);
xor U8220 (N_8220,N_7916,N_7991);
and U8221 (N_8221,N_7966,N_7750);
nand U8222 (N_8222,N_7932,N_7893);
or U8223 (N_8223,N_7781,N_7928);
or U8224 (N_8224,N_7830,N_7774);
nor U8225 (N_8225,N_7779,N_7834);
nand U8226 (N_8226,N_7846,N_7833);
or U8227 (N_8227,N_7836,N_7902);
xor U8228 (N_8228,N_7789,N_7821);
xnor U8229 (N_8229,N_7937,N_7773);
nor U8230 (N_8230,N_7777,N_7910);
or U8231 (N_8231,N_7934,N_7800);
nand U8232 (N_8232,N_7845,N_7901);
nand U8233 (N_8233,N_7865,N_7880);
or U8234 (N_8234,N_7901,N_7910);
xor U8235 (N_8235,N_7893,N_7865);
nor U8236 (N_8236,N_7972,N_7903);
nor U8237 (N_8237,N_7794,N_7915);
nand U8238 (N_8238,N_7879,N_7937);
and U8239 (N_8239,N_7802,N_7911);
and U8240 (N_8240,N_7914,N_7841);
or U8241 (N_8241,N_7815,N_7883);
nor U8242 (N_8242,N_7924,N_7932);
or U8243 (N_8243,N_7996,N_7857);
xor U8244 (N_8244,N_7983,N_7929);
or U8245 (N_8245,N_7885,N_7810);
nand U8246 (N_8246,N_7877,N_7821);
or U8247 (N_8247,N_7891,N_7828);
and U8248 (N_8248,N_7988,N_7959);
nor U8249 (N_8249,N_7957,N_7834);
nor U8250 (N_8250,N_8036,N_8022);
nor U8251 (N_8251,N_8236,N_8003);
or U8252 (N_8252,N_8084,N_8006);
nand U8253 (N_8253,N_8123,N_8212);
or U8254 (N_8254,N_8023,N_8217);
nor U8255 (N_8255,N_8100,N_8037);
and U8256 (N_8256,N_8031,N_8027);
nand U8257 (N_8257,N_8173,N_8240);
xnor U8258 (N_8258,N_8140,N_8149);
nand U8259 (N_8259,N_8075,N_8159);
nor U8260 (N_8260,N_8184,N_8202);
nor U8261 (N_8261,N_8118,N_8034);
or U8262 (N_8262,N_8231,N_8205);
xor U8263 (N_8263,N_8158,N_8201);
or U8264 (N_8264,N_8210,N_8168);
and U8265 (N_8265,N_8093,N_8204);
nand U8266 (N_8266,N_8119,N_8108);
or U8267 (N_8267,N_8090,N_8230);
and U8268 (N_8268,N_8152,N_8129);
nor U8269 (N_8269,N_8109,N_8166);
xor U8270 (N_8270,N_8033,N_8193);
xor U8271 (N_8271,N_8150,N_8076);
nand U8272 (N_8272,N_8190,N_8067);
xor U8273 (N_8273,N_8025,N_8001);
nand U8274 (N_8274,N_8163,N_8048);
and U8275 (N_8275,N_8046,N_8183);
nand U8276 (N_8276,N_8091,N_8207);
nand U8277 (N_8277,N_8079,N_8132);
nand U8278 (N_8278,N_8131,N_8174);
xor U8279 (N_8279,N_8224,N_8078);
or U8280 (N_8280,N_8229,N_8156);
nand U8281 (N_8281,N_8213,N_8115);
xor U8282 (N_8282,N_8007,N_8248);
xor U8283 (N_8283,N_8055,N_8060);
nor U8284 (N_8284,N_8170,N_8239);
or U8285 (N_8285,N_8234,N_8215);
xnor U8286 (N_8286,N_8203,N_8062);
nor U8287 (N_8287,N_8222,N_8134);
nor U8288 (N_8288,N_8186,N_8110);
or U8289 (N_8289,N_8216,N_8113);
nor U8290 (N_8290,N_8112,N_8087);
xor U8291 (N_8291,N_8018,N_8228);
nand U8292 (N_8292,N_8194,N_8104);
and U8293 (N_8293,N_8105,N_8219);
nor U8294 (N_8294,N_8160,N_8126);
or U8295 (N_8295,N_8179,N_8107);
xnor U8296 (N_8296,N_8148,N_8211);
xnor U8297 (N_8297,N_8214,N_8041);
xor U8298 (N_8298,N_8220,N_8139);
and U8299 (N_8299,N_8012,N_8232);
nor U8300 (N_8300,N_8083,N_8095);
nor U8301 (N_8301,N_8127,N_8245);
nand U8302 (N_8302,N_8049,N_8032);
nand U8303 (N_8303,N_8061,N_8035);
or U8304 (N_8304,N_8082,N_8077);
xor U8305 (N_8305,N_8181,N_8209);
or U8306 (N_8306,N_8121,N_8050);
and U8307 (N_8307,N_8208,N_8144);
nor U8308 (N_8308,N_8045,N_8120);
and U8309 (N_8309,N_8014,N_8017);
or U8310 (N_8310,N_8019,N_8068);
nand U8311 (N_8311,N_8070,N_8157);
xor U8312 (N_8312,N_8238,N_8058);
nor U8313 (N_8313,N_8071,N_8124);
xnor U8314 (N_8314,N_8028,N_8011);
xor U8315 (N_8315,N_8000,N_8054);
nand U8316 (N_8316,N_8151,N_8111);
and U8317 (N_8317,N_8089,N_8218);
nand U8318 (N_8318,N_8180,N_8226);
and U8319 (N_8319,N_8147,N_8069);
and U8320 (N_8320,N_8191,N_8165);
and U8321 (N_8321,N_8088,N_8164);
nor U8322 (N_8322,N_8010,N_8233);
nand U8323 (N_8323,N_8169,N_8161);
or U8324 (N_8324,N_8008,N_8167);
and U8325 (N_8325,N_8044,N_8221);
and U8326 (N_8326,N_8247,N_8146);
nand U8327 (N_8327,N_8242,N_8094);
nor U8328 (N_8328,N_8080,N_8063);
nand U8329 (N_8329,N_8013,N_8065);
xor U8330 (N_8330,N_8106,N_8133);
nand U8331 (N_8331,N_8128,N_8135);
xor U8332 (N_8332,N_8145,N_8197);
xnor U8333 (N_8333,N_8086,N_8030);
and U8334 (N_8334,N_8200,N_8235);
xor U8335 (N_8335,N_8243,N_8199);
or U8336 (N_8336,N_8096,N_8249);
nand U8337 (N_8337,N_8122,N_8114);
or U8338 (N_8338,N_8066,N_8020);
and U8339 (N_8339,N_8040,N_8039);
or U8340 (N_8340,N_8103,N_8241);
or U8341 (N_8341,N_8136,N_8162);
and U8342 (N_8342,N_8246,N_8099);
nand U8343 (N_8343,N_8198,N_8097);
and U8344 (N_8344,N_8098,N_8237);
nand U8345 (N_8345,N_8155,N_8004);
nand U8346 (N_8346,N_8051,N_8130);
nor U8347 (N_8347,N_8142,N_8052);
nor U8348 (N_8348,N_8015,N_8223);
or U8349 (N_8349,N_8189,N_8138);
xnor U8350 (N_8350,N_8137,N_8227);
and U8351 (N_8351,N_8154,N_8016);
or U8352 (N_8352,N_8196,N_8225);
or U8353 (N_8353,N_8182,N_8064);
and U8354 (N_8354,N_8042,N_8143);
and U8355 (N_8355,N_8206,N_8029);
xor U8356 (N_8356,N_8175,N_8057);
or U8357 (N_8357,N_8085,N_8009);
nor U8358 (N_8358,N_8005,N_8047);
and U8359 (N_8359,N_8172,N_8177);
xor U8360 (N_8360,N_8059,N_8056);
nor U8361 (N_8361,N_8026,N_8053);
nand U8362 (N_8362,N_8074,N_8125);
xor U8363 (N_8363,N_8092,N_8038);
nand U8364 (N_8364,N_8153,N_8188);
xor U8365 (N_8365,N_8178,N_8021);
nor U8366 (N_8366,N_8024,N_8002);
nor U8367 (N_8367,N_8185,N_8187);
nor U8368 (N_8368,N_8072,N_8101);
xor U8369 (N_8369,N_8195,N_8073);
nand U8370 (N_8370,N_8171,N_8102);
and U8371 (N_8371,N_8043,N_8141);
or U8372 (N_8372,N_8081,N_8116);
xor U8373 (N_8373,N_8117,N_8176);
and U8374 (N_8374,N_8244,N_8192);
nand U8375 (N_8375,N_8179,N_8123);
xnor U8376 (N_8376,N_8052,N_8013);
and U8377 (N_8377,N_8222,N_8049);
nand U8378 (N_8378,N_8007,N_8040);
nor U8379 (N_8379,N_8248,N_8076);
nand U8380 (N_8380,N_8080,N_8081);
nor U8381 (N_8381,N_8097,N_8236);
nor U8382 (N_8382,N_8117,N_8131);
or U8383 (N_8383,N_8167,N_8003);
and U8384 (N_8384,N_8061,N_8137);
nand U8385 (N_8385,N_8184,N_8182);
nor U8386 (N_8386,N_8134,N_8180);
or U8387 (N_8387,N_8100,N_8128);
or U8388 (N_8388,N_8230,N_8186);
xnor U8389 (N_8389,N_8044,N_8097);
nand U8390 (N_8390,N_8218,N_8009);
xor U8391 (N_8391,N_8212,N_8199);
or U8392 (N_8392,N_8127,N_8030);
nor U8393 (N_8393,N_8158,N_8108);
and U8394 (N_8394,N_8191,N_8086);
and U8395 (N_8395,N_8249,N_8034);
nor U8396 (N_8396,N_8225,N_8113);
or U8397 (N_8397,N_8078,N_8023);
nand U8398 (N_8398,N_8157,N_8002);
xnor U8399 (N_8399,N_8129,N_8193);
or U8400 (N_8400,N_8232,N_8241);
nor U8401 (N_8401,N_8167,N_8057);
nor U8402 (N_8402,N_8210,N_8091);
or U8403 (N_8403,N_8211,N_8041);
or U8404 (N_8404,N_8045,N_8099);
nor U8405 (N_8405,N_8214,N_8211);
or U8406 (N_8406,N_8230,N_8122);
and U8407 (N_8407,N_8163,N_8244);
xnor U8408 (N_8408,N_8224,N_8191);
nor U8409 (N_8409,N_8156,N_8052);
nor U8410 (N_8410,N_8203,N_8176);
nor U8411 (N_8411,N_8186,N_8145);
or U8412 (N_8412,N_8104,N_8161);
xnor U8413 (N_8413,N_8200,N_8157);
xnor U8414 (N_8414,N_8142,N_8128);
and U8415 (N_8415,N_8159,N_8225);
nor U8416 (N_8416,N_8126,N_8061);
nor U8417 (N_8417,N_8133,N_8032);
nand U8418 (N_8418,N_8062,N_8038);
and U8419 (N_8419,N_8198,N_8138);
xor U8420 (N_8420,N_8204,N_8158);
and U8421 (N_8421,N_8128,N_8058);
xor U8422 (N_8422,N_8117,N_8170);
or U8423 (N_8423,N_8174,N_8219);
nor U8424 (N_8424,N_8100,N_8066);
xor U8425 (N_8425,N_8246,N_8230);
nand U8426 (N_8426,N_8102,N_8013);
xor U8427 (N_8427,N_8019,N_8045);
xor U8428 (N_8428,N_8049,N_8058);
and U8429 (N_8429,N_8193,N_8189);
nand U8430 (N_8430,N_8173,N_8106);
nor U8431 (N_8431,N_8103,N_8150);
nand U8432 (N_8432,N_8147,N_8218);
nand U8433 (N_8433,N_8032,N_8029);
and U8434 (N_8434,N_8249,N_8105);
and U8435 (N_8435,N_8212,N_8044);
nor U8436 (N_8436,N_8185,N_8154);
nor U8437 (N_8437,N_8228,N_8030);
or U8438 (N_8438,N_8200,N_8142);
nand U8439 (N_8439,N_8070,N_8184);
or U8440 (N_8440,N_8149,N_8014);
xnor U8441 (N_8441,N_8117,N_8112);
nor U8442 (N_8442,N_8070,N_8061);
xor U8443 (N_8443,N_8175,N_8129);
xor U8444 (N_8444,N_8061,N_8243);
xnor U8445 (N_8445,N_8215,N_8036);
nor U8446 (N_8446,N_8013,N_8240);
nand U8447 (N_8447,N_8057,N_8081);
nand U8448 (N_8448,N_8170,N_8187);
or U8449 (N_8449,N_8090,N_8038);
nand U8450 (N_8450,N_8094,N_8028);
nor U8451 (N_8451,N_8094,N_8116);
nor U8452 (N_8452,N_8164,N_8120);
or U8453 (N_8453,N_8096,N_8237);
or U8454 (N_8454,N_8062,N_8182);
or U8455 (N_8455,N_8139,N_8019);
or U8456 (N_8456,N_8115,N_8049);
nand U8457 (N_8457,N_8013,N_8183);
xor U8458 (N_8458,N_8111,N_8246);
or U8459 (N_8459,N_8187,N_8034);
xor U8460 (N_8460,N_8071,N_8173);
nor U8461 (N_8461,N_8168,N_8073);
and U8462 (N_8462,N_8078,N_8070);
or U8463 (N_8463,N_8122,N_8181);
xor U8464 (N_8464,N_8191,N_8119);
nand U8465 (N_8465,N_8148,N_8171);
nor U8466 (N_8466,N_8071,N_8046);
nor U8467 (N_8467,N_8132,N_8150);
xor U8468 (N_8468,N_8141,N_8076);
xor U8469 (N_8469,N_8238,N_8048);
or U8470 (N_8470,N_8056,N_8048);
nor U8471 (N_8471,N_8070,N_8150);
and U8472 (N_8472,N_8206,N_8192);
nand U8473 (N_8473,N_8104,N_8215);
nand U8474 (N_8474,N_8026,N_8191);
nand U8475 (N_8475,N_8030,N_8224);
and U8476 (N_8476,N_8078,N_8066);
or U8477 (N_8477,N_8000,N_8133);
or U8478 (N_8478,N_8107,N_8211);
and U8479 (N_8479,N_8232,N_8023);
or U8480 (N_8480,N_8126,N_8145);
nand U8481 (N_8481,N_8138,N_8144);
and U8482 (N_8482,N_8176,N_8056);
nor U8483 (N_8483,N_8048,N_8179);
xnor U8484 (N_8484,N_8161,N_8158);
nor U8485 (N_8485,N_8004,N_8222);
xor U8486 (N_8486,N_8132,N_8082);
and U8487 (N_8487,N_8125,N_8043);
or U8488 (N_8488,N_8048,N_8015);
nor U8489 (N_8489,N_8159,N_8037);
nor U8490 (N_8490,N_8201,N_8108);
and U8491 (N_8491,N_8203,N_8029);
nor U8492 (N_8492,N_8132,N_8221);
nor U8493 (N_8493,N_8175,N_8220);
and U8494 (N_8494,N_8154,N_8007);
xor U8495 (N_8495,N_8149,N_8087);
nor U8496 (N_8496,N_8229,N_8042);
and U8497 (N_8497,N_8125,N_8084);
and U8498 (N_8498,N_8121,N_8084);
nor U8499 (N_8499,N_8169,N_8028);
xor U8500 (N_8500,N_8487,N_8284);
xnor U8501 (N_8501,N_8485,N_8326);
nand U8502 (N_8502,N_8424,N_8266);
nor U8503 (N_8503,N_8365,N_8455);
xnor U8504 (N_8504,N_8389,N_8464);
xor U8505 (N_8505,N_8440,N_8277);
nand U8506 (N_8506,N_8263,N_8355);
nor U8507 (N_8507,N_8437,N_8443);
xnor U8508 (N_8508,N_8406,N_8411);
and U8509 (N_8509,N_8279,N_8462);
nor U8510 (N_8510,N_8410,N_8470);
and U8511 (N_8511,N_8373,N_8461);
nor U8512 (N_8512,N_8404,N_8472);
and U8513 (N_8513,N_8376,N_8403);
xnor U8514 (N_8514,N_8271,N_8377);
xor U8515 (N_8515,N_8489,N_8301);
or U8516 (N_8516,N_8310,N_8275);
and U8517 (N_8517,N_8401,N_8451);
nand U8518 (N_8518,N_8330,N_8346);
and U8519 (N_8519,N_8315,N_8388);
nor U8520 (N_8520,N_8251,N_8436);
nand U8521 (N_8521,N_8299,N_8328);
xnor U8522 (N_8522,N_8285,N_8446);
nor U8523 (N_8523,N_8349,N_8296);
nor U8524 (N_8524,N_8405,N_8370);
or U8525 (N_8525,N_8253,N_8313);
nand U8526 (N_8526,N_8260,N_8293);
nor U8527 (N_8527,N_8413,N_8382);
nand U8528 (N_8528,N_8474,N_8289);
or U8529 (N_8529,N_8281,N_8269);
or U8530 (N_8530,N_8323,N_8320);
and U8531 (N_8531,N_8454,N_8264);
nand U8532 (N_8532,N_8426,N_8308);
or U8533 (N_8533,N_8300,N_8316);
or U8534 (N_8534,N_8286,N_8449);
xnor U8535 (N_8535,N_8429,N_8475);
nand U8536 (N_8536,N_8407,N_8351);
nor U8537 (N_8537,N_8386,N_8331);
or U8538 (N_8538,N_8456,N_8460);
or U8539 (N_8539,N_8458,N_8379);
nor U8540 (N_8540,N_8337,N_8262);
nand U8541 (N_8541,N_8473,N_8398);
xor U8542 (N_8542,N_8329,N_8479);
nor U8543 (N_8543,N_8309,N_8481);
and U8544 (N_8544,N_8254,N_8419);
nor U8545 (N_8545,N_8468,N_8422);
and U8546 (N_8546,N_8255,N_8327);
and U8547 (N_8547,N_8493,N_8412);
nor U8548 (N_8548,N_8304,N_8463);
nor U8549 (N_8549,N_8268,N_8290);
and U8550 (N_8550,N_8369,N_8273);
nand U8551 (N_8551,N_8321,N_8274);
or U8552 (N_8552,N_8391,N_8342);
xnor U8553 (N_8553,N_8343,N_8291);
nand U8554 (N_8554,N_8261,N_8257);
nor U8555 (N_8555,N_8392,N_8420);
nor U8556 (N_8556,N_8394,N_8427);
nand U8557 (N_8557,N_8423,N_8417);
or U8558 (N_8558,N_8267,N_8256);
nor U8559 (N_8559,N_8364,N_8444);
and U8560 (N_8560,N_8498,N_8356);
xor U8561 (N_8561,N_8402,N_8488);
nand U8562 (N_8562,N_8288,N_8335);
or U8563 (N_8563,N_8385,N_8495);
xnor U8564 (N_8564,N_8397,N_8367);
and U8565 (N_8565,N_8457,N_8390);
nor U8566 (N_8566,N_8490,N_8372);
nand U8567 (N_8567,N_8368,N_8425);
and U8568 (N_8568,N_8438,N_8396);
nand U8569 (N_8569,N_8361,N_8441);
or U8570 (N_8570,N_8465,N_8312);
and U8571 (N_8571,N_8354,N_8278);
nor U8572 (N_8572,N_8374,N_8276);
nor U8573 (N_8573,N_8341,N_8258);
nor U8574 (N_8574,N_8452,N_8294);
xor U8575 (N_8575,N_8430,N_8305);
xnor U8576 (N_8576,N_8387,N_8471);
nor U8577 (N_8577,N_8434,N_8395);
nor U8578 (N_8578,N_8408,N_8332);
nor U8579 (N_8579,N_8371,N_8380);
and U8580 (N_8580,N_8287,N_8435);
and U8581 (N_8581,N_8283,N_8339);
and U8582 (N_8582,N_8482,N_8348);
nor U8583 (N_8583,N_8478,N_8322);
nand U8584 (N_8584,N_8466,N_8492);
or U8585 (N_8585,N_8298,N_8448);
xnor U8586 (N_8586,N_8303,N_8432);
nand U8587 (N_8587,N_8428,N_8483);
and U8588 (N_8588,N_8325,N_8494);
nand U8589 (N_8589,N_8250,N_8282);
and U8590 (N_8590,N_8334,N_8362);
nor U8591 (N_8591,N_8375,N_8306);
nand U8592 (N_8592,N_8307,N_8447);
nor U8593 (N_8593,N_8357,N_8295);
or U8594 (N_8594,N_8333,N_8352);
and U8595 (N_8595,N_8442,N_8344);
nor U8596 (N_8596,N_8358,N_8459);
xor U8597 (N_8597,N_8336,N_8499);
and U8598 (N_8598,N_8416,N_8311);
or U8599 (N_8599,N_8319,N_8353);
nand U8600 (N_8600,N_8252,N_8445);
or U8601 (N_8601,N_8384,N_8486);
or U8602 (N_8602,N_8476,N_8317);
and U8603 (N_8603,N_8409,N_8270);
xor U8604 (N_8604,N_8360,N_8347);
or U8605 (N_8605,N_8421,N_8340);
nor U8606 (N_8606,N_8366,N_8383);
or U8607 (N_8607,N_8318,N_8414);
xnor U8608 (N_8608,N_8477,N_8491);
nor U8609 (N_8609,N_8399,N_8302);
and U8610 (N_8610,N_8265,N_8338);
nand U8611 (N_8611,N_8467,N_8280);
nor U8612 (N_8612,N_8496,N_8480);
nor U8613 (N_8613,N_8297,N_8350);
nand U8614 (N_8614,N_8359,N_8381);
xnor U8615 (N_8615,N_8439,N_8484);
nor U8616 (N_8616,N_8415,N_8292);
xnor U8617 (N_8617,N_8450,N_8259);
or U8618 (N_8618,N_8324,N_8345);
xor U8619 (N_8619,N_8314,N_8378);
xor U8620 (N_8620,N_8363,N_8497);
xor U8621 (N_8621,N_8469,N_8418);
nand U8622 (N_8622,N_8393,N_8453);
nand U8623 (N_8623,N_8433,N_8400);
or U8624 (N_8624,N_8272,N_8431);
nor U8625 (N_8625,N_8417,N_8389);
nand U8626 (N_8626,N_8356,N_8255);
nor U8627 (N_8627,N_8465,N_8408);
nand U8628 (N_8628,N_8262,N_8347);
nand U8629 (N_8629,N_8401,N_8304);
nor U8630 (N_8630,N_8319,N_8337);
and U8631 (N_8631,N_8490,N_8451);
nand U8632 (N_8632,N_8464,N_8324);
xor U8633 (N_8633,N_8272,N_8459);
and U8634 (N_8634,N_8288,N_8305);
and U8635 (N_8635,N_8402,N_8476);
nand U8636 (N_8636,N_8264,N_8465);
nand U8637 (N_8637,N_8431,N_8353);
and U8638 (N_8638,N_8308,N_8450);
or U8639 (N_8639,N_8327,N_8442);
nand U8640 (N_8640,N_8288,N_8312);
nor U8641 (N_8641,N_8496,N_8279);
nand U8642 (N_8642,N_8340,N_8337);
nand U8643 (N_8643,N_8469,N_8327);
and U8644 (N_8644,N_8445,N_8417);
nor U8645 (N_8645,N_8496,N_8322);
or U8646 (N_8646,N_8478,N_8390);
nand U8647 (N_8647,N_8350,N_8296);
xor U8648 (N_8648,N_8381,N_8254);
nand U8649 (N_8649,N_8435,N_8252);
xor U8650 (N_8650,N_8265,N_8283);
and U8651 (N_8651,N_8296,N_8250);
nand U8652 (N_8652,N_8363,N_8293);
or U8653 (N_8653,N_8432,N_8333);
xor U8654 (N_8654,N_8315,N_8301);
xor U8655 (N_8655,N_8322,N_8449);
or U8656 (N_8656,N_8257,N_8262);
or U8657 (N_8657,N_8299,N_8367);
or U8658 (N_8658,N_8405,N_8477);
or U8659 (N_8659,N_8343,N_8378);
or U8660 (N_8660,N_8354,N_8273);
nand U8661 (N_8661,N_8480,N_8363);
or U8662 (N_8662,N_8350,N_8255);
xor U8663 (N_8663,N_8470,N_8269);
xnor U8664 (N_8664,N_8339,N_8342);
nor U8665 (N_8665,N_8277,N_8495);
or U8666 (N_8666,N_8373,N_8446);
or U8667 (N_8667,N_8442,N_8489);
nor U8668 (N_8668,N_8355,N_8315);
nor U8669 (N_8669,N_8368,N_8455);
nor U8670 (N_8670,N_8465,N_8479);
nor U8671 (N_8671,N_8423,N_8388);
or U8672 (N_8672,N_8378,N_8442);
nor U8673 (N_8673,N_8423,N_8480);
nand U8674 (N_8674,N_8405,N_8317);
and U8675 (N_8675,N_8416,N_8357);
nor U8676 (N_8676,N_8331,N_8299);
nand U8677 (N_8677,N_8265,N_8381);
nand U8678 (N_8678,N_8316,N_8401);
xor U8679 (N_8679,N_8391,N_8446);
nor U8680 (N_8680,N_8407,N_8476);
and U8681 (N_8681,N_8354,N_8498);
or U8682 (N_8682,N_8416,N_8355);
nor U8683 (N_8683,N_8369,N_8403);
or U8684 (N_8684,N_8310,N_8288);
nand U8685 (N_8685,N_8322,N_8381);
or U8686 (N_8686,N_8410,N_8351);
or U8687 (N_8687,N_8298,N_8276);
and U8688 (N_8688,N_8464,N_8431);
nand U8689 (N_8689,N_8330,N_8416);
and U8690 (N_8690,N_8375,N_8276);
nand U8691 (N_8691,N_8481,N_8324);
or U8692 (N_8692,N_8370,N_8372);
and U8693 (N_8693,N_8351,N_8485);
nor U8694 (N_8694,N_8490,N_8472);
nand U8695 (N_8695,N_8381,N_8287);
xnor U8696 (N_8696,N_8323,N_8251);
nor U8697 (N_8697,N_8372,N_8361);
nor U8698 (N_8698,N_8374,N_8417);
and U8699 (N_8699,N_8264,N_8309);
and U8700 (N_8700,N_8312,N_8280);
nor U8701 (N_8701,N_8474,N_8329);
and U8702 (N_8702,N_8429,N_8383);
nor U8703 (N_8703,N_8251,N_8488);
nor U8704 (N_8704,N_8393,N_8352);
nand U8705 (N_8705,N_8458,N_8487);
nand U8706 (N_8706,N_8462,N_8476);
xor U8707 (N_8707,N_8257,N_8382);
nor U8708 (N_8708,N_8283,N_8336);
nand U8709 (N_8709,N_8446,N_8321);
xnor U8710 (N_8710,N_8473,N_8357);
nor U8711 (N_8711,N_8332,N_8322);
nand U8712 (N_8712,N_8284,N_8296);
nand U8713 (N_8713,N_8439,N_8291);
nand U8714 (N_8714,N_8303,N_8295);
and U8715 (N_8715,N_8403,N_8436);
and U8716 (N_8716,N_8474,N_8437);
or U8717 (N_8717,N_8280,N_8362);
nand U8718 (N_8718,N_8375,N_8442);
or U8719 (N_8719,N_8439,N_8341);
nor U8720 (N_8720,N_8482,N_8464);
xnor U8721 (N_8721,N_8417,N_8454);
nor U8722 (N_8722,N_8496,N_8401);
xor U8723 (N_8723,N_8291,N_8305);
and U8724 (N_8724,N_8499,N_8256);
or U8725 (N_8725,N_8472,N_8434);
and U8726 (N_8726,N_8268,N_8441);
nor U8727 (N_8727,N_8351,N_8257);
or U8728 (N_8728,N_8313,N_8392);
or U8729 (N_8729,N_8498,N_8310);
nor U8730 (N_8730,N_8400,N_8319);
xor U8731 (N_8731,N_8462,N_8322);
and U8732 (N_8732,N_8471,N_8286);
xor U8733 (N_8733,N_8413,N_8312);
or U8734 (N_8734,N_8463,N_8380);
or U8735 (N_8735,N_8368,N_8317);
nor U8736 (N_8736,N_8484,N_8405);
nand U8737 (N_8737,N_8295,N_8334);
nor U8738 (N_8738,N_8427,N_8403);
or U8739 (N_8739,N_8428,N_8446);
xor U8740 (N_8740,N_8394,N_8397);
or U8741 (N_8741,N_8420,N_8325);
or U8742 (N_8742,N_8407,N_8491);
nor U8743 (N_8743,N_8289,N_8442);
nand U8744 (N_8744,N_8265,N_8359);
xnor U8745 (N_8745,N_8331,N_8393);
nand U8746 (N_8746,N_8311,N_8342);
and U8747 (N_8747,N_8470,N_8495);
nor U8748 (N_8748,N_8450,N_8497);
and U8749 (N_8749,N_8495,N_8354);
or U8750 (N_8750,N_8564,N_8515);
nand U8751 (N_8751,N_8700,N_8508);
and U8752 (N_8752,N_8736,N_8609);
nand U8753 (N_8753,N_8617,N_8559);
or U8754 (N_8754,N_8713,N_8527);
nor U8755 (N_8755,N_8732,N_8737);
and U8756 (N_8756,N_8656,N_8503);
nand U8757 (N_8757,N_8697,N_8516);
xor U8758 (N_8758,N_8744,N_8718);
nand U8759 (N_8759,N_8646,N_8593);
nand U8760 (N_8760,N_8526,N_8687);
or U8761 (N_8761,N_8678,N_8579);
nor U8762 (N_8762,N_8521,N_8641);
and U8763 (N_8763,N_8531,N_8691);
or U8764 (N_8764,N_8553,N_8556);
nor U8765 (N_8765,N_8557,N_8729);
nand U8766 (N_8766,N_8639,N_8525);
xnor U8767 (N_8767,N_8662,N_8710);
or U8768 (N_8768,N_8601,N_8623);
nor U8769 (N_8769,N_8549,N_8613);
and U8770 (N_8770,N_8707,N_8621);
and U8771 (N_8771,N_8524,N_8541);
nor U8772 (N_8772,N_8501,N_8620);
and U8773 (N_8773,N_8704,N_8546);
and U8774 (N_8774,N_8708,N_8666);
xor U8775 (N_8775,N_8683,N_8535);
nand U8776 (N_8776,N_8528,N_8518);
and U8777 (N_8777,N_8611,N_8667);
and U8778 (N_8778,N_8625,N_8569);
and U8779 (N_8779,N_8500,N_8676);
nor U8780 (N_8780,N_8709,N_8693);
nor U8781 (N_8781,N_8606,N_8536);
and U8782 (N_8782,N_8547,N_8634);
nor U8783 (N_8783,N_8624,N_8604);
and U8784 (N_8784,N_8738,N_8598);
or U8785 (N_8785,N_8520,N_8504);
xor U8786 (N_8786,N_8699,N_8726);
xor U8787 (N_8787,N_8689,N_8505);
and U8788 (N_8788,N_8533,N_8510);
xor U8789 (N_8789,N_8522,N_8651);
xnor U8790 (N_8790,N_8675,N_8565);
and U8791 (N_8791,N_8542,N_8669);
nand U8792 (N_8792,N_8637,N_8686);
nand U8793 (N_8793,N_8746,N_8595);
nor U8794 (N_8794,N_8748,N_8645);
and U8795 (N_8795,N_8714,N_8723);
nor U8796 (N_8796,N_8706,N_8673);
nor U8797 (N_8797,N_8696,N_8690);
nand U8798 (N_8798,N_8650,N_8674);
nand U8799 (N_8799,N_8592,N_8552);
or U8800 (N_8800,N_8562,N_8657);
nor U8801 (N_8801,N_8519,N_8749);
nand U8802 (N_8802,N_8733,N_8698);
nand U8803 (N_8803,N_8643,N_8597);
and U8804 (N_8804,N_8692,N_8717);
xor U8805 (N_8805,N_8603,N_8716);
nand U8806 (N_8806,N_8636,N_8685);
nand U8807 (N_8807,N_8586,N_8722);
nor U8808 (N_8808,N_8741,N_8551);
and U8809 (N_8809,N_8594,N_8665);
nor U8810 (N_8810,N_8555,N_8682);
or U8811 (N_8811,N_8640,N_8628);
nand U8812 (N_8812,N_8627,N_8633);
nand U8813 (N_8813,N_8728,N_8629);
nor U8814 (N_8814,N_8511,N_8560);
or U8815 (N_8815,N_8608,N_8548);
nand U8816 (N_8816,N_8544,N_8513);
xnor U8817 (N_8817,N_8602,N_8725);
and U8818 (N_8818,N_8581,N_8571);
and U8819 (N_8819,N_8638,N_8580);
xnor U8820 (N_8820,N_8661,N_8576);
and U8821 (N_8821,N_8721,N_8743);
or U8822 (N_8822,N_8745,N_8740);
and U8823 (N_8823,N_8703,N_8622);
or U8824 (N_8824,N_8618,N_8724);
or U8825 (N_8825,N_8507,N_8550);
xnor U8826 (N_8826,N_8605,N_8631);
nand U8827 (N_8827,N_8626,N_8652);
nor U8828 (N_8828,N_8660,N_8567);
nor U8829 (N_8829,N_8539,N_8590);
and U8830 (N_8830,N_8668,N_8715);
or U8831 (N_8831,N_8572,N_8719);
or U8832 (N_8832,N_8712,N_8701);
nor U8833 (N_8833,N_8577,N_8612);
nor U8834 (N_8834,N_8663,N_8570);
nand U8835 (N_8835,N_8514,N_8530);
and U8836 (N_8836,N_8596,N_8720);
and U8837 (N_8837,N_8670,N_8731);
nor U8838 (N_8838,N_8509,N_8658);
nand U8839 (N_8839,N_8563,N_8664);
nor U8840 (N_8840,N_8512,N_8735);
xnor U8841 (N_8841,N_8554,N_8659);
xor U8842 (N_8842,N_8705,N_8727);
or U8843 (N_8843,N_8589,N_8672);
or U8844 (N_8844,N_8647,N_8679);
or U8845 (N_8845,N_8642,N_8615);
xnor U8846 (N_8846,N_8694,N_8568);
nand U8847 (N_8847,N_8543,N_8730);
and U8848 (N_8848,N_8654,N_8600);
nor U8849 (N_8849,N_8632,N_8529);
and U8850 (N_8850,N_8739,N_8607);
nor U8851 (N_8851,N_8653,N_8574);
and U8852 (N_8852,N_8711,N_8558);
xor U8853 (N_8853,N_8583,N_8742);
xor U8854 (N_8854,N_8630,N_8695);
or U8855 (N_8855,N_8599,N_8648);
and U8856 (N_8856,N_8591,N_8561);
and U8857 (N_8857,N_8582,N_8502);
or U8858 (N_8858,N_8585,N_8747);
and U8859 (N_8859,N_8575,N_8688);
and U8860 (N_8860,N_8588,N_8677);
xor U8861 (N_8861,N_8532,N_8614);
or U8862 (N_8862,N_8540,N_8573);
and U8863 (N_8863,N_8534,N_8681);
or U8864 (N_8864,N_8584,N_8545);
xnor U8865 (N_8865,N_8523,N_8671);
or U8866 (N_8866,N_8655,N_8680);
xor U8867 (N_8867,N_8587,N_8610);
or U8868 (N_8868,N_8619,N_8538);
nor U8869 (N_8869,N_8649,N_8684);
or U8870 (N_8870,N_8702,N_8578);
xor U8871 (N_8871,N_8537,N_8506);
nor U8872 (N_8872,N_8566,N_8644);
and U8873 (N_8873,N_8616,N_8734);
and U8874 (N_8874,N_8635,N_8517);
nor U8875 (N_8875,N_8541,N_8584);
nand U8876 (N_8876,N_8626,N_8550);
xnor U8877 (N_8877,N_8626,N_8684);
and U8878 (N_8878,N_8593,N_8501);
nand U8879 (N_8879,N_8500,N_8580);
nor U8880 (N_8880,N_8664,N_8593);
and U8881 (N_8881,N_8616,N_8686);
nand U8882 (N_8882,N_8732,N_8689);
nor U8883 (N_8883,N_8534,N_8646);
nand U8884 (N_8884,N_8572,N_8623);
and U8885 (N_8885,N_8651,N_8610);
xnor U8886 (N_8886,N_8679,N_8584);
nand U8887 (N_8887,N_8523,N_8628);
nor U8888 (N_8888,N_8567,N_8503);
nor U8889 (N_8889,N_8689,N_8741);
nand U8890 (N_8890,N_8696,N_8557);
or U8891 (N_8891,N_8506,N_8689);
xnor U8892 (N_8892,N_8511,N_8671);
xnor U8893 (N_8893,N_8573,N_8724);
and U8894 (N_8894,N_8579,N_8611);
and U8895 (N_8895,N_8746,N_8606);
and U8896 (N_8896,N_8731,N_8581);
nand U8897 (N_8897,N_8591,N_8649);
or U8898 (N_8898,N_8609,N_8601);
and U8899 (N_8899,N_8647,N_8671);
or U8900 (N_8900,N_8670,N_8706);
and U8901 (N_8901,N_8562,N_8688);
and U8902 (N_8902,N_8618,N_8527);
or U8903 (N_8903,N_8546,N_8668);
xnor U8904 (N_8904,N_8698,N_8649);
xor U8905 (N_8905,N_8686,N_8702);
xnor U8906 (N_8906,N_8737,N_8510);
nor U8907 (N_8907,N_8624,N_8599);
xor U8908 (N_8908,N_8550,N_8650);
and U8909 (N_8909,N_8571,N_8741);
nand U8910 (N_8910,N_8703,N_8558);
nand U8911 (N_8911,N_8615,N_8525);
and U8912 (N_8912,N_8561,N_8734);
xnor U8913 (N_8913,N_8517,N_8607);
or U8914 (N_8914,N_8698,N_8622);
nand U8915 (N_8915,N_8506,N_8728);
or U8916 (N_8916,N_8534,N_8650);
or U8917 (N_8917,N_8525,N_8644);
nand U8918 (N_8918,N_8505,N_8591);
xor U8919 (N_8919,N_8683,N_8515);
xnor U8920 (N_8920,N_8560,N_8709);
xnor U8921 (N_8921,N_8577,N_8621);
nor U8922 (N_8922,N_8629,N_8522);
nor U8923 (N_8923,N_8607,N_8621);
nor U8924 (N_8924,N_8621,N_8625);
xnor U8925 (N_8925,N_8649,N_8556);
or U8926 (N_8926,N_8529,N_8726);
nand U8927 (N_8927,N_8597,N_8726);
or U8928 (N_8928,N_8571,N_8564);
or U8929 (N_8929,N_8603,N_8569);
nor U8930 (N_8930,N_8587,N_8529);
nor U8931 (N_8931,N_8531,N_8718);
nor U8932 (N_8932,N_8585,N_8686);
or U8933 (N_8933,N_8527,N_8710);
or U8934 (N_8934,N_8502,N_8545);
xnor U8935 (N_8935,N_8744,N_8711);
or U8936 (N_8936,N_8572,N_8747);
and U8937 (N_8937,N_8719,N_8567);
xnor U8938 (N_8938,N_8532,N_8595);
nand U8939 (N_8939,N_8516,N_8664);
and U8940 (N_8940,N_8653,N_8606);
or U8941 (N_8941,N_8728,N_8677);
xnor U8942 (N_8942,N_8734,N_8657);
nor U8943 (N_8943,N_8696,N_8518);
or U8944 (N_8944,N_8665,N_8529);
xnor U8945 (N_8945,N_8527,N_8600);
or U8946 (N_8946,N_8604,N_8563);
or U8947 (N_8947,N_8738,N_8583);
nor U8948 (N_8948,N_8617,N_8585);
or U8949 (N_8949,N_8706,N_8647);
or U8950 (N_8950,N_8695,N_8641);
xor U8951 (N_8951,N_8590,N_8688);
nand U8952 (N_8952,N_8594,N_8612);
nand U8953 (N_8953,N_8510,N_8742);
or U8954 (N_8954,N_8686,N_8667);
nor U8955 (N_8955,N_8584,N_8590);
xnor U8956 (N_8956,N_8661,N_8527);
nand U8957 (N_8957,N_8731,N_8502);
and U8958 (N_8958,N_8609,N_8657);
or U8959 (N_8959,N_8605,N_8619);
and U8960 (N_8960,N_8517,N_8648);
nor U8961 (N_8961,N_8710,N_8656);
xor U8962 (N_8962,N_8602,N_8511);
nor U8963 (N_8963,N_8665,N_8748);
nor U8964 (N_8964,N_8606,N_8544);
nand U8965 (N_8965,N_8743,N_8615);
nor U8966 (N_8966,N_8536,N_8512);
or U8967 (N_8967,N_8630,N_8539);
nand U8968 (N_8968,N_8725,N_8718);
or U8969 (N_8969,N_8728,N_8703);
xor U8970 (N_8970,N_8679,N_8736);
and U8971 (N_8971,N_8733,N_8646);
or U8972 (N_8972,N_8518,N_8722);
nand U8973 (N_8973,N_8571,N_8661);
nand U8974 (N_8974,N_8552,N_8542);
xor U8975 (N_8975,N_8698,N_8689);
or U8976 (N_8976,N_8514,N_8683);
xnor U8977 (N_8977,N_8543,N_8671);
and U8978 (N_8978,N_8569,N_8654);
xnor U8979 (N_8979,N_8703,N_8720);
xnor U8980 (N_8980,N_8509,N_8610);
or U8981 (N_8981,N_8616,N_8518);
nor U8982 (N_8982,N_8640,N_8698);
nand U8983 (N_8983,N_8696,N_8716);
xnor U8984 (N_8984,N_8703,N_8568);
nor U8985 (N_8985,N_8565,N_8511);
and U8986 (N_8986,N_8684,N_8616);
and U8987 (N_8987,N_8523,N_8728);
nor U8988 (N_8988,N_8636,N_8587);
and U8989 (N_8989,N_8657,N_8579);
nor U8990 (N_8990,N_8749,N_8727);
and U8991 (N_8991,N_8559,N_8568);
nor U8992 (N_8992,N_8687,N_8723);
or U8993 (N_8993,N_8650,N_8606);
or U8994 (N_8994,N_8722,N_8712);
nand U8995 (N_8995,N_8591,N_8567);
or U8996 (N_8996,N_8657,N_8701);
nor U8997 (N_8997,N_8705,N_8607);
nor U8998 (N_8998,N_8681,N_8612);
xnor U8999 (N_8999,N_8744,N_8738);
xor U9000 (N_9000,N_8895,N_8859);
nand U9001 (N_9001,N_8795,N_8943);
and U9002 (N_9002,N_8897,N_8957);
and U9003 (N_9003,N_8869,N_8761);
xnor U9004 (N_9004,N_8758,N_8992);
and U9005 (N_9005,N_8860,N_8796);
or U9006 (N_9006,N_8851,N_8790);
and U9007 (N_9007,N_8995,N_8912);
xnor U9008 (N_9008,N_8752,N_8827);
xor U9009 (N_9009,N_8838,N_8824);
or U9010 (N_9010,N_8867,N_8904);
xor U9011 (N_9011,N_8769,N_8978);
nor U9012 (N_9012,N_8926,N_8905);
xnor U9013 (N_9013,N_8817,N_8945);
xnor U9014 (N_9014,N_8839,N_8765);
or U9015 (N_9015,N_8892,N_8887);
nor U9016 (N_9016,N_8885,N_8993);
nor U9017 (N_9017,N_8914,N_8846);
nand U9018 (N_9018,N_8811,N_8850);
and U9019 (N_9019,N_8830,N_8880);
and U9020 (N_9020,N_8999,N_8858);
nor U9021 (N_9021,N_8944,N_8823);
and U9022 (N_9022,N_8847,N_8994);
xor U9023 (N_9023,N_8816,N_8854);
xor U9024 (N_9024,N_8930,N_8845);
xor U9025 (N_9025,N_8987,N_8813);
and U9026 (N_9026,N_8783,N_8770);
or U9027 (N_9027,N_8879,N_8865);
nor U9028 (N_9028,N_8797,N_8857);
nand U9029 (N_9029,N_8925,N_8900);
nor U9030 (N_9030,N_8810,N_8946);
nor U9031 (N_9031,N_8840,N_8950);
or U9032 (N_9032,N_8911,N_8753);
nor U9033 (N_9033,N_8990,N_8964);
or U9034 (N_9034,N_8763,N_8906);
nand U9035 (N_9035,N_8873,N_8982);
and U9036 (N_9036,N_8951,N_8980);
nor U9037 (N_9037,N_8807,N_8955);
xor U9038 (N_9038,N_8821,N_8938);
nor U9039 (N_9039,N_8862,N_8890);
nand U9040 (N_9040,N_8803,N_8874);
or U9041 (N_9041,N_8787,N_8836);
and U9042 (N_9042,N_8808,N_8908);
nor U9043 (N_9043,N_8798,N_8901);
nor U9044 (N_9044,N_8909,N_8806);
xnor U9045 (N_9045,N_8917,N_8876);
or U9046 (N_9046,N_8976,N_8921);
and U9047 (N_9047,N_8948,N_8775);
nand U9048 (N_9048,N_8963,N_8868);
xor U9049 (N_9049,N_8768,N_8893);
nand U9050 (N_9050,N_8910,N_8920);
and U9051 (N_9051,N_8861,N_8971);
xnor U9052 (N_9052,N_8849,N_8941);
or U9053 (N_9053,N_8961,N_8962);
nor U9054 (N_9054,N_8812,N_8800);
nor U9055 (N_9055,N_8779,N_8788);
nor U9056 (N_9056,N_8866,N_8888);
or U9057 (N_9057,N_8934,N_8872);
and U9058 (N_9058,N_8907,N_8924);
nor U9059 (N_9059,N_8988,N_8781);
nor U9060 (N_9060,N_8772,N_8767);
nand U9061 (N_9061,N_8815,N_8997);
nor U9062 (N_9062,N_8891,N_8991);
nand U9063 (N_9063,N_8764,N_8933);
or U9064 (N_9064,N_8931,N_8958);
or U9065 (N_9065,N_8985,N_8979);
nor U9066 (N_9066,N_8884,N_8972);
or U9067 (N_9067,N_8801,N_8947);
nor U9068 (N_9068,N_8762,N_8886);
xor U9069 (N_9069,N_8835,N_8927);
or U9070 (N_9070,N_8814,N_8833);
or U9071 (N_9071,N_8902,N_8932);
and U9072 (N_9072,N_8952,N_8818);
nor U9073 (N_9073,N_8953,N_8974);
xnor U9074 (N_9074,N_8989,N_8751);
or U9075 (N_9075,N_8949,N_8929);
nand U9076 (N_9076,N_8793,N_8954);
or U9077 (N_9077,N_8799,N_8848);
or U9078 (N_9078,N_8981,N_8754);
nand U9079 (N_9079,N_8883,N_8882);
or U9080 (N_9080,N_8969,N_8805);
xor U9081 (N_9081,N_8970,N_8960);
or U9082 (N_9082,N_8928,N_8896);
nand U9083 (N_9083,N_8864,N_8791);
xnor U9084 (N_9084,N_8828,N_8973);
or U9085 (N_9085,N_8771,N_8998);
nor U9086 (N_9086,N_8760,N_8842);
nor U9087 (N_9087,N_8756,N_8829);
xor U9088 (N_9088,N_8863,N_8878);
xor U9089 (N_9089,N_8777,N_8881);
and U9090 (N_9090,N_8871,N_8959);
or U9091 (N_9091,N_8913,N_8843);
xnor U9092 (N_9092,N_8841,N_8825);
nand U9093 (N_9093,N_8967,N_8837);
xnor U9094 (N_9094,N_8782,N_8870);
nand U9095 (N_9095,N_8919,N_8802);
nor U9096 (N_9096,N_8785,N_8822);
nand U9097 (N_9097,N_8986,N_8996);
nand U9098 (N_9098,N_8794,N_8832);
xor U9099 (N_9099,N_8834,N_8774);
xnor U9100 (N_9100,N_8977,N_8789);
nand U9101 (N_9101,N_8937,N_8903);
nor U9102 (N_9102,N_8918,N_8915);
nand U9103 (N_9103,N_8819,N_8975);
and U9104 (N_9104,N_8935,N_8826);
and U9105 (N_9105,N_8984,N_8898);
nor U9106 (N_9106,N_8809,N_8956);
xor U9107 (N_9107,N_8820,N_8922);
nor U9108 (N_9108,N_8877,N_8983);
or U9109 (N_9109,N_8776,N_8939);
xor U9110 (N_9110,N_8844,N_8852);
or U9111 (N_9111,N_8916,N_8855);
and U9112 (N_9112,N_8853,N_8780);
nor U9113 (N_9113,N_8784,N_8750);
and U9114 (N_9114,N_8778,N_8773);
and U9115 (N_9115,N_8966,N_8965);
or U9116 (N_9116,N_8792,N_8968);
nand U9117 (N_9117,N_8875,N_8766);
nand U9118 (N_9118,N_8889,N_8804);
nor U9119 (N_9119,N_8786,N_8757);
or U9120 (N_9120,N_8936,N_8831);
nor U9121 (N_9121,N_8759,N_8923);
xor U9122 (N_9122,N_8894,N_8899);
nand U9123 (N_9123,N_8755,N_8940);
and U9124 (N_9124,N_8856,N_8942);
xnor U9125 (N_9125,N_8867,N_8923);
or U9126 (N_9126,N_8835,N_8766);
xor U9127 (N_9127,N_8848,N_8802);
or U9128 (N_9128,N_8903,N_8893);
or U9129 (N_9129,N_8948,N_8851);
nor U9130 (N_9130,N_8936,N_8939);
or U9131 (N_9131,N_8952,N_8945);
xor U9132 (N_9132,N_8759,N_8953);
xnor U9133 (N_9133,N_8809,N_8829);
or U9134 (N_9134,N_8801,N_8965);
and U9135 (N_9135,N_8981,N_8926);
or U9136 (N_9136,N_8911,N_8842);
nand U9137 (N_9137,N_8907,N_8928);
nand U9138 (N_9138,N_8806,N_8980);
xor U9139 (N_9139,N_8919,N_8985);
or U9140 (N_9140,N_8764,N_8789);
nand U9141 (N_9141,N_8980,N_8968);
nand U9142 (N_9142,N_8872,N_8799);
nand U9143 (N_9143,N_8995,N_8831);
nand U9144 (N_9144,N_8989,N_8971);
nand U9145 (N_9145,N_8870,N_8761);
nor U9146 (N_9146,N_8989,N_8789);
xor U9147 (N_9147,N_8824,N_8881);
xor U9148 (N_9148,N_8819,N_8876);
xnor U9149 (N_9149,N_8775,N_8821);
xor U9150 (N_9150,N_8964,N_8974);
nor U9151 (N_9151,N_8928,N_8904);
or U9152 (N_9152,N_8816,N_8852);
nor U9153 (N_9153,N_8901,N_8767);
and U9154 (N_9154,N_8931,N_8833);
xor U9155 (N_9155,N_8966,N_8946);
nor U9156 (N_9156,N_8994,N_8978);
xnor U9157 (N_9157,N_8751,N_8902);
nor U9158 (N_9158,N_8806,N_8751);
or U9159 (N_9159,N_8818,N_8945);
nor U9160 (N_9160,N_8788,N_8885);
and U9161 (N_9161,N_8845,N_8792);
xor U9162 (N_9162,N_8895,N_8923);
nor U9163 (N_9163,N_8976,N_8919);
nand U9164 (N_9164,N_8758,N_8925);
nor U9165 (N_9165,N_8999,N_8996);
nand U9166 (N_9166,N_8810,N_8801);
nand U9167 (N_9167,N_8929,N_8786);
nor U9168 (N_9168,N_8765,N_8947);
or U9169 (N_9169,N_8833,N_8788);
nand U9170 (N_9170,N_8767,N_8782);
nor U9171 (N_9171,N_8969,N_8764);
or U9172 (N_9172,N_8990,N_8838);
nand U9173 (N_9173,N_8944,N_8901);
nand U9174 (N_9174,N_8971,N_8753);
xnor U9175 (N_9175,N_8936,N_8846);
xnor U9176 (N_9176,N_8850,N_8993);
nor U9177 (N_9177,N_8983,N_8963);
nand U9178 (N_9178,N_8999,N_8886);
or U9179 (N_9179,N_8896,N_8899);
xor U9180 (N_9180,N_8953,N_8872);
and U9181 (N_9181,N_8867,N_8864);
and U9182 (N_9182,N_8984,N_8972);
nand U9183 (N_9183,N_8827,N_8811);
and U9184 (N_9184,N_8778,N_8922);
nand U9185 (N_9185,N_8939,N_8958);
nand U9186 (N_9186,N_8770,N_8852);
xnor U9187 (N_9187,N_8846,N_8984);
or U9188 (N_9188,N_8816,N_8979);
and U9189 (N_9189,N_8860,N_8769);
nor U9190 (N_9190,N_8837,N_8929);
nand U9191 (N_9191,N_8983,N_8800);
nand U9192 (N_9192,N_8780,N_8934);
and U9193 (N_9193,N_8855,N_8932);
or U9194 (N_9194,N_8776,N_8839);
and U9195 (N_9195,N_8872,N_8892);
nand U9196 (N_9196,N_8925,N_8763);
nor U9197 (N_9197,N_8752,N_8974);
xor U9198 (N_9198,N_8792,N_8785);
xnor U9199 (N_9199,N_8846,N_8786);
xor U9200 (N_9200,N_8931,N_8968);
xnor U9201 (N_9201,N_8780,N_8982);
nand U9202 (N_9202,N_8869,N_8916);
nand U9203 (N_9203,N_8812,N_8798);
nor U9204 (N_9204,N_8797,N_8862);
xnor U9205 (N_9205,N_8791,N_8946);
or U9206 (N_9206,N_8998,N_8941);
xor U9207 (N_9207,N_8978,N_8872);
and U9208 (N_9208,N_8870,N_8774);
nand U9209 (N_9209,N_8848,N_8785);
nand U9210 (N_9210,N_8988,N_8836);
and U9211 (N_9211,N_8765,N_8960);
and U9212 (N_9212,N_8988,N_8785);
and U9213 (N_9213,N_8814,N_8932);
nor U9214 (N_9214,N_8985,N_8771);
and U9215 (N_9215,N_8763,N_8962);
nand U9216 (N_9216,N_8936,N_8959);
nand U9217 (N_9217,N_8807,N_8756);
nand U9218 (N_9218,N_8963,N_8819);
xor U9219 (N_9219,N_8986,N_8994);
nor U9220 (N_9220,N_8943,N_8799);
nor U9221 (N_9221,N_8797,N_8811);
and U9222 (N_9222,N_8910,N_8978);
or U9223 (N_9223,N_8928,N_8773);
xor U9224 (N_9224,N_8927,N_8886);
and U9225 (N_9225,N_8992,N_8838);
and U9226 (N_9226,N_8788,N_8916);
xor U9227 (N_9227,N_8793,N_8824);
or U9228 (N_9228,N_8758,N_8761);
xor U9229 (N_9229,N_8867,N_8974);
xnor U9230 (N_9230,N_8949,N_8870);
nand U9231 (N_9231,N_8851,N_8902);
xnor U9232 (N_9232,N_8879,N_8848);
nand U9233 (N_9233,N_8863,N_8908);
or U9234 (N_9234,N_8780,N_8786);
or U9235 (N_9235,N_8906,N_8836);
nor U9236 (N_9236,N_8880,N_8762);
or U9237 (N_9237,N_8851,N_8951);
nand U9238 (N_9238,N_8762,N_8942);
and U9239 (N_9239,N_8952,N_8886);
nor U9240 (N_9240,N_8764,N_8768);
xnor U9241 (N_9241,N_8996,N_8987);
and U9242 (N_9242,N_8932,N_8869);
xnor U9243 (N_9243,N_8969,N_8853);
or U9244 (N_9244,N_8997,N_8971);
xnor U9245 (N_9245,N_8827,N_8839);
nor U9246 (N_9246,N_8892,N_8778);
nand U9247 (N_9247,N_8894,N_8818);
nor U9248 (N_9248,N_8903,N_8857);
nor U9249 (N_9249,N_8895,N_8877);
xor U9250 (N_9250,N_9081,N_9085);
nand U9251 (N_9251,N_9118,N_9165);
nand U9252 (N_9252,N_9181,N_9088);
and U9253 (N_9253,N_9034,N_9220);
or U9254 (N_9254,N_9050,N_9046);
and U9255 (N_9255,N_9238,N_9035);
or U9256 (N_9256,N_9195,N_9073);
or U9257 (N_9257,N_9078,N_9037);
or U9258 (N_9258,N_9048,N_9199);
or U9259 (N_9259,N_9143,N_9194);
or U9260 (N_9260,N_9042,N_9201);
xnor U9261 (N_9261,N_9090,N_9124);
nor U9262 (N_9262,N_9086,N_9141);
nand U9263 (N_9263,N_9144,N_9249);
or U9264 (N_9264,N_9089,N_9028);
nand U9265 (N_9265,N_9160,N_9242);
nor U9266 (N_9266,N_9129,N_9147);
and U9267 (N_9267,N_9184,N_9043);
nor U9268 (N_9268,N_9064,N_9196);
nand U9269 (N_9269,N_9151,N_9159);
xor U9270 (N_9270,N_9113,N_9231);
nor U9271 (N_9271,N_9071,N_9172);
and U9272 (N_9272,N_9014,N_9218);
nand U9273 (N_9273,N_9183,N_9169);
and U9274 (N_9274,N_9222,N_9134);
and U9275 (N_9275,N_9191,N_9177);
and U9276 (N_9276,N_9011,N_9167);
or U9277 (N_9277,N_9152,N_9044);
xor U9278 (N_9278,N_9032,N_9163);
xor U9279 (N_9279,N_9108,N_9017);
nand U9280 (N_9280,N_9153,N_9036);
or U9281 (N_9281,N_9084,N_9119);
nor U9282 (N_9282,N_9182,N_9197);
xnor U9283 (N_9283,N_9004,N_9247);
nand U9284 (N_9284,N_9052,N_9135);
nor U9285 (N_9285,N_9217,N_9031);
nor U9286 (N_9286,N_9030,N_9038);
and U9287 (N_9287,N_9072,N_9007);
or U9288 (N_9288,N_9080,N_9010);
nand U9289 (N_9289,N_9100,N_9066);
and U9290 (N_9290,N_9161,N_9221);
nor U9291 (N_9291,N_9101,N_9154);
nand U9292 (N_9292,N_9106,N_9095);
nand U9293 (N_9293,N_9005,N_9003);
and U9294 (N_9294,N_9103,N_9128);
xor U9295 (N_9295,N_9123,N_9002);
or U9296 (N_9296,N_9168,N_9099);
nand U9297 (N_9297,N_9000,N_9051);
nand U9298 (N_9298,N_9130,N_9175);
and U9299 (N_9299,N_9202,N_9156);
nand U9300 (N_9300,N_9213,N_9212);
nand U9301 (N_9301,N_9176,N_9246);
nand U9302 (N_9302,N_9013,N_9021);
and U9303 (N_9303,N_9219,N_9243);
xnor U9304 (N_9304,N_9012,N_9192);
xnor U9305 (N_9305,N_9096,N_9069);
xor U9306 (N_9306,N_9205,N_9015);
xor U9307 (N_9307,N_9207,N_9233);
xor U9308 (N_9308,N_9245,N_9214);
xnor U9309 (N_9309,N_9076,N_9230);
nor U9310 (N_9310,N_9041,N_9077);
and U9311 (N_9311,N_9132,N_9056);
and U9312 (N_9312,N_9001,N_9166);
or U9313 (N_9313,N_9223,N_9225);
nand U9314 (N_9314,N_9067,N_9098);
nor U9315 (N_9315,N_9203,N_9186);
nor U9316 (N_9316,N_9114,N_9171);
xor U9317 (N_9317,N_9209,N_9226);
nor U9318 (N_9318,N_9107,N_9237);
or U9319 (N_9319,N_9137,N_9215);
nor U9320 (N_9320,N_9040,N_9060);
or U9321 (N_9321,N_9102,N_9127);
or U9322 (N_9322,N_9244,N_9227);
or U9323 (N_9323,N_9235,N_9150);
and U9324 (N_9324,N_9239,N_9248);
nand U9325 (N_9325,N_9131,N_9204);
or U9326 (N_9326,N_9087,N_9138);
or U9327 (N_9327,N_9234,N_9211);
nor U9328 (N_9328,N_9216,N_9068);
xor U9329 (N_9329,N_9029,N_9091);
nor U9330 (N_9330,N_9120,N_9190);
nand U9331 (N_9331,N_9241,N_9180);
xnor U9332 (N_9332,N_9025,N_9016);
xor U9333 (N_9333,N_9027,N_9039);
xnor U9334 (N_9334,N_9062,N_9094);
nand U9335 (N_9335,N_9047,N_9126);
nand U9336 (N_9336,N_9117,N_9173);
xnor U9337 (N_9337,N_9122,N_9045);
and U9338 (N_9338,N_9059,N_9210);
xnor U9339 (N_9339,N_9170,N_9193);
or U9340 (N_9340,N_9065,N_9092);
and U9341 (N_9341,N_9033,N_9155);
nor U9342 (N_9342,N_9208,N_9162);
or U9343 (N_9343,N_9061,N_9093);
xnor U9344 (N_9344,N_9139,N_9054);
nor U9345 (N_9345,N_9110,N_9149);
and U9346 (N_9346,N_9200,N_9185);
xor U9347 (N_9347,N_9228,N_9157);
or U9348 (N_9348,N_9049,N_9112);
or U9349 (N_9349,N_9079,N_9178);
and U9350 (N_9350,N_9024,N_9082);
nor U9351 (N_9351,N_9164,N_9136);
nor U9352 (N_9352,N_9097,N_9224);
and U9353 (N_9353,N_9009,N_9115);
xor U9354 (N_9354,N_9133,N_9020);
nor U9355 (N_9355,N_9109,N_9008);
nor U9356 (N_9356,N_9187,N_9019);
nor U9357 (N_9357,N_9158,N_9063);
nand U9358 (N_9358,N_9022,N_9074);
or U9359 (N_9359,N_9111,N_9232);
and U9360 (N_9360,N_9070,N_9148);
and U9361 (N_9361,N_9018,N_9075);
and U9362 (N_9362,N_9055,N_9188);
nor U9363 (N_9363,N_9142,N_9058);
nor U9364 (N_9364,N_9121,N_9140);
and U9365 (N_9365,N_9240,N_9198);
xnor U9366 (N_9366,N_9206,N_9146);
xor U9367 (N_9367,N_9189,N_9179);
xor U9368 (N_9368,N_9174,N_9229);
nor U9369 (N_9369,N_9083,N_9145);
or U9370 (N_9370,N_9236,N_9023);
or U9371 (N_9371,N_9026,N_9116);
nor U9372 (N_9372,N_9125,N_9105);
nor U9373 (N_9373,N_9006,N_9053);
nor U9374 (N_9374,N_9104,N_9057);
nor U9375 (N_9375,N_9225,N_9020);
nand U9376 (N_9376,N_9054,N_9121);
xor U9377 (N_9377,N_9124,N_9114);
nand U9378 (N_9378,N_9009,N_9078);
nor U9379 (N_9379,N_9230,N_9214);
nand U9380 (N_9380,N_9073,N_9107);
or U9381 (N_9381,N_9099,N_9102);
or U9382 (N_9382,N_9089,N_9151);
nor U9383 (N_9383,N_9235,N_9014);
xnor U9384 (N_9384,N_9125,N_9119);
nand U9385 (N_9385,N_9030,N_9181);
nand U9386 (N_9386,N_9113,N_9210);
nor U9387 (N_9387,N_9192,N_9200);
nand U9388 (N_9388,N_9013,N_9211);
xor U9389 (N_9389,N_9005,N_9099);
nor U9390 (N_9390,N_9121,N_9067);
xnor U9391 (N_9391,N_9079,N_9161);
nand U9392 (N_9392,N_9234,N_9186);
and U9393 (N_9393,N_9188,N_9201);
and U9394 (N_9394,N_9224,N_9014);
xnor U9395 (N_9395,N_9079,N_9113);
xor U9396 (N_9396,N_9177,N_9049);
and U9397 (N_9397,N_9019,N_9034);
nand U9398 (N_9398,N_9058,N_9086);
or U9399 (N_9399,N_9198,N_9008);
xnor U9400 (N_9400,N_9107,N_9214);
nor U9401 (N_9401,N_9212,N_9015);
xnor U9402 (N_9402,N_9053,N_9236);
or U9403 (N_9403,N_9227,N_9044);
or U9404 (N_9404,N_9113,N_9095);
and U9405 (N_9405,N_9179,N_9016);
xnor U9406 (N_9406,N_9092,N_9142);
nor U9407 (N_9407,N_9171,N_9035);
or U9408 (N_9408,N_9016,N_9050);
nor U9409 (N_9409,N_9044,N_9099);
nand U9410 (N_9410,N_9201,N_9034);
and U9411 (N_9411,N_9157,N_9032);
nand U9412 (N_9412,N_9149,N_9097);
nand U9413 (N_9413,N_9074,N_9238);
nor U9414 (N_9414,N_9233,N_9169);
nand U9415 (N_9415,N_9064,N_9157);
nand U9416 (N_9416,N_9247,N_9178);
nand U9417 (N_9417,N_9133,N_9240);
xnor U9418 (N_9418,N_9229,N_9002);
xor U9419 (N_9419,N_9156,N_9238);
nor U9420 (N_9420,N_9087,N_9003);
and U9421 (N_9421,N_9043,N_9190);
or U9422 (N_9422,N_9163,N_9017);
nor U9423 (N_9423,N_9097,N_9092);
xnor U9424 (N_9424,N_9018,N_9063);
and U9425 (N_9425,N_9116,N_9018);
nand U9426 (N_9426,N_9032,N_9119);
xor U9427 (N_9427,N_9082,N_9100);
or U9428 (N_9428,N_9141,N_9185);
xor U9429 (N_9429,N_9163,N_9145);
or U9430 (N_9430,N_9116,N_9025);
or U9431 (N_9431,N_9071,N_9197);
xor U9432 (N_9432,N_9173,N_9075);
xnor U9433 (N_9433,N_9182,N_9051);
and U9434 (N_9434,N_9126,N_9171);
or U9435 (N_9435,N_9051,N_9108);
nand U9436 (N_9436,N_9014,N_9178);
or U9437 (N_9437,N_9023,N_9134);
nand U9438 (N_9438,N_9179,N_9111);
nand U9439 (N_9439,N_9026,N_9091);
nand U9440 (N_9440,N_9089,N_9246);
xor U9441 (N_9441,N_9071,N_9101);
nor U9442 (N_9442,N_9236,N_9171);
nand U9443 (N_9443,N_9106,N_9195);
xnor U9444 (N_9444,N_9120,N_9048);
xnor U9445 (N_9445,N_9173,N_9047);
nor U9446 (N_9446,N_9089,N_9053);
nand U9447 (N_9447,N_9059,N_9074);
nor U9448 (N_9448,N_9097,N_9245);
and U9449 (N_9449,N_9137,N_9089);
nor U9450 (N_9450,N_9114,N_9217);
and U9451 (N_9451,N_9151,N_9058);
or U9452 (N_9452,N_9149,N_9162);
or U9453 (N_9453,N_9137,N_9176);
nor U9454 (N_9454,N_9093,N_9010);
xnor U9455 (N_9455,N_9040,N_9006);
or U9456 (N_9456,N_9188,N_9037);
xor U9457 (N_9457,N_9022,N_9075);
nand U9458 (N_9458,N_9087,N_9032);
and U9459 (N_9459,N_9102,N_9210);
nor U9460 (N_9460,N_9114,N_9128);
nor U9461 (N_9461,N_9122,N_9152);
nor U9462 (N_9462,N_9018,N_9228);
or U9463 (N_9463,N_9077,N_9237);
nor U9464 (N_9464,N_9078,N_9080);
nor U9465 (N_9465,N_9080,N_9149);
nand U9466 (N_9466,N_9148,N_9151);
xor U9467 (N_9467,N_9074,N_9164);
nor U9468 (N_9468,N_9146,N_9005);
xor U9469 (N_9469,N_9052,N_9076);
nor U9470 (N_9470,N_9072,N_9140);
nor U9471 (N_9471,N_9062,N_9034);
xor U9472 (N_9472,N_9063,N_9232);
and U9473 (N_9473,N_9078,N_9030);
and U9474 (N_9474,N_9171,N_9240);
or U9475 (N_9475,N_9127,N_9142);
xnor U9476 (N_9476,N_9140,N_9106);
xor U9477 (N_9477,N_9163,N_9135);
nand U9478 (N_9478,N_9020,N_9187);
nand U9479 (N_9479,N_9245,N_9220);
and U9480 (N_9480,N_9002,N_9098);
or U9481 (N_9481,N_9102,N_9151);
nor U9482 (N_9482,N_9103,N_9116);
or U9483 (N_9483,N_9140,N_9165);
or U9484 (N_9484,N_9094,N_9017);
or U9485 (N_9485,N_9054,N_9238);
nand U9486 (N_9486,N_9012,N_9191);
and U9487 (N_9487,N_9182,N_9240);
and U9488 (N_9488,N_9147,N_9123);
nand U9489 (N_9489,N_9176,N_9076);
nor U9490 (N_9490,N_9126,N_9177);
nand U9491 (N_9491,N_9150,N_9067);
or U9492 (N_9492,N_9019,N_9082);
xor U9493 (N_9493,N_9230,N_9101);
nor U9494 (N_9494,N_9238,N_9228);
xor U9495 (N_9495,N_9095,N_9003);
and U9496 (N_9496,N_9015,N_9065);
nor U9497 (N_9497,N_9215,N_9111);
nand U9498 (N_9498,N_9156,N_9060);
nand U9499 (N_9499,N_9222,N_9061);
and U9500 (N_9500,N_9487,N_9450);
nor U9501 (N_9501,N_9259,N_9439);
xor U9502 (N_9502,N_9492,N_9495);
nand U9503 (N_9503,N_9467,N_9386);
nor U9504 (N_9504,N_9436,N_9412);
nand U9505 (N_9505,N_9320,N_9445);
nor U9506 (N_9506,N_9483,N_9301);
or U9507 (N_9507,N_9423,N_9254);
xnor U9508 (N_9508,N_9388,N_9465);
nand U9509 (N_9509,N_9323,N_9340);
nor U9510 (N_9510,N_9250,N_9486);
nand U9511 (N_9511,N_9309,N_9394);
nand U9512 (N_9512,N_9258,N_9441);
xor U9513 (N_9513,N_9261,N_9269);
nor U9514 (N_9514,N_9270,N_9472);
nor U9515 (N_9515,N_9319,N_9331);
and U9516 (N_9516,N_9416,N_9325);
nor U9517 (N_9517,N_9390,N_9440);
xnor U9518 (N_9518,N_9494,N_9335);
nor U9519 (N_9519,N_9462,N_9350);
or U9520 (N_9520,N_9358,N_9449);
or U9521 (N_9521,N_9456,N_9410);
nor U9522 (N_9522,N_9489,N_9329);
or U9523 (N_9523,N_9364,N_9466);
nor U9524 (N_9524,N_9368,N_9404);
nor U9525 (N_9525,N_9266,N_9318);
nor U9526 (N_9526,N_9262,N_9382);
and U9527 (N_9527,N_9279,N_9479);
nand U9528 (N_9528,N_9473,N_9470);
and U9529 (N_9529,N_9268,N_9265);
and U9530 (N_9530,N_9286,N_9293);
and U9531 (N_9531,N_9316,N_9327);
xnor U9532 (N_9532,N_9347,N_9337);
nor U9533 (N_9533,N_9359,N_9498);
xor U9534 (N_9534,N_9446,N_9491);
and U9535 (N_9535,N_9384,N_9264);
nor U9536 (N_9536,N_9289,N_9344);
and U9537 (N_9537,N_9361,N_9338);
or U9538 (N_9538,N_9447,N_9274);
nor U9539 (N_9539,N_9408,N_9444);
nand U9540 (N_9540,N_9252,N_9306);
xor U9541 (N_9541,N_9413,N_9385);
xor U9542 (N_9542,N_9438,N_9474);
or U9543 (N_9543,N_9392,N_9477);
or U9544 (N_9544,N_9260,N_9488);
and U9545 (N_9545,N_9343,N_9435);
nor U9546 (N_9546,N_9377,N_9356);
or U9547 (N_9547,N_9428,N_9396);
nor U9548 (N_9548,N_9499,N_9280);
and U9549 (N_9549,N_9346,N_9395);
or U9550 (N_9550,N_9481,N_9371);
nor U9551 (N_9551,N_9271,N_9480);
nand U9552 (N_9552,N_9458,N_9399);
or U9553 (N_9553,N_9400,N_9354);
xnor U9554 (N_9554,N_9418,N_9313);
nor U9555 (N_9555,N_9314,N_9294);
nor U9556 (N_9556,N_9424,N_9490);
and U9557 (N_9557,N_9464,N_9454);
nand U9558 (N_9558,N_9496,N_9452);
and U9559 (N_9559,N_9457,N_9253);
nand U9560 (N_9560,N_9326,N_9349);
nand U9561 (N_9561,N_9433,N_9308);
and U9562 (N_9562,N_9283,N_9415);
nand U9563 (N_9563,N_9275,N_9332);
nor U9564 (N_9564,N_9453,N_9353);
or U9565 (N_9565,N_9409,N_9310);
xor U9566 (N_9566,N_9284,N_9379);
and U9567 (N_9567,N_9398,N_9305);
nand U9568 (N_9568,N_9317,N_9297);
nand U9569 (N_9569,N_9407,N_9485);
xnor U9570 (N_9570,N_9351,N_9478);
xor U9571 (N_9571,N_9366,N_9475);
nand U9572 (N_9572,N_9468,N_9391);
or U9573 (N_9573,N_9362,N_9461);
nor U9574 (N_9574,N_9282,N_9272);
or U9575 (N_9575,N_9311,N_9405);
or U9576 (N_9576,N_9370,N_9427);
or U9577 (N_9577,N_9321,N_9263);
xnor U9578 (N_9578,N_9425,N_9484);
xnor U9579 (N_9579,N_9304,N_9292);
nand U9580 (N_9580,N_9476,N_9328);
and U9581 (N_9581,N_9448,N_9345);
xor U9582 (N_9582,N_9469,N_9296);
nand U9583 (N_9583,N_9276,N_9429);
nand U9584 (N_9584,N_9442,N_9455);
nor U9585 (N_9585,N_9251,N_9267);
or U9586 (N_9586,N_9497,N_9380);
nand U9587 (N_9587,N_9322,N_9375);
nand U9588 (N_9588,N_9493,N_9312);
nor U9589 (N_9589,N_9426,N_9373);
nand U9590 (N_9590,N_9459,N_9393);
and U9591 (N_9591,N_9300,N_9403);
nand U9592 (N_9592,N_9376,N_9334);
nand U9593 (N_9593,N_9273,N_9299);
or U9594 (N_9594,N_9411,N_9401);
and U9595 (N_9595,N_9451,N_9421);
nor U9596 (N_9596,N_9430,N_9291);
nor U9597 (N_9597,N_9342,N_9372);
or U9598 (N_9598,N_9255,N_9257);
or U9599 (N_9599,N_9437,N_9295);
or U9600 (N_9600,N_9397,N_9363);
nand U9601 (N_9601,N_9369,N_9333);
or U9602 (N_9602,N_9288,N_9389);
xor U9603 (N_9603,N_9434,N_9281);
xor U9604 (N_9604,N_9277,N_9443);
nor U9605 (N_9605,N_9287,N_9460);
xor U9606 (N_9606,N_9463,N_9307);
nor U9607 (N_9607,N_9365,N_9414);
nor U9608 (N_9608,N_9278,N_9471);
and U9609 (N_9609,N_9303,N_9348);
nand U9610 (N_9610,N_9341,N_9315);
nor U9611 (N_9611,N_9378,N_9330);
nand U9612 (N_9612,N_9417,N_9360);
nor U9613 (N_9613,N_9339,N_9419);
nor U9614 (N_9614,N_9381,N_9432);
nand U9615 (N_9615,N_9406,N_9431);
nor U9616 (N_9616,N_9402,N_9302);
and U9617 (N_9617,N_9324,N_9352);
and U9618 (N_9618,N_9387,N_9357);
nor U9619 (N_9619,N_9290,N_9256);
nor U9620 (N_9620,N_9298,N_9367);
nor U9621 (N_9621,N_9420,N_9374);
nand U9622 (N_9622,N_9355,N_9336);
nand U9623 (N_9623,N_9422,N_9383);
and U9624 (N_9624,N_9482,N_9285);
and U9625 (N_9625,N_9485,N_9496);
nand U9626 (N_9626,N_9398,N_9360);
nor U9627 (N_9627,N_9463,N_9355);
nand U9628 (N_9628,N_9258,N_9342);
or U9629 (N_9629,N_9302,N_9497);
xor U9630 (N_9630,N_9348,N_9402);
nor U9631 (N_9631,N_9376,N_9457);
nand U9632 (N_9632,N_9378,N_9418);
or U9633 (N_9633,N_9392,N_9398);
nand U9634 (N_9634,N_9420,N_9435);
nand U9635 (N_9635,N_9474,N_9477);
or U9636 (N_9636,N_9332,N_9354);
and U9637 (N_9637,N_9278,N_9494);
nand U9638 (N_9638,N_9321,N_9310);
or U9639 (N_9639,N_9278,N_9318);
nor U9640 (N_9640,N_9252,N_9423);
nand U9641 (N_9641,N_9436,N_9346);
nor U9642 (N_9642,N_9277,N_9462);
xor U9643 (N_9643,N_9286,N_9354);
and U9644 (N_9644,N_9277,N_9409);
and U9645 (N_9645,N_9345,N_9273);
and U9646 (N_9646,N_9266,N_9362);
or U9647 (N_9647,N_9478,N_9254);
nand U9648 (N_9648,N_9370,N_9261);
or U9649 (N_9649,N_9366,N_9325);
or U9650 (N_9650,N_9355,N_9410);
nand U9651 (N_9651,N_9354,N_9394);
nor U9652 (N_9652,N_9397,N_9430);
xnor U9653 (N_9653,N_9353,N_9361);
xnor U9654 (N_9654,N_9435,N_9457);
and U9655 (N_9655,N_9274,N_9356);
or U9656 (N_9656,N_9284,N_9421);
nor U9657 (N_9657,N_9472,N_9329);
or U9658 (N_9658,N_9302,N_9458);
xnor U9659 (N_9659,N_9449,N_9280);
nand U9660 (N_9660,N_9459,N_9335);
and U9661 (N_9661,N_9428,N_9459);
or U9662 (N_9662,N_9470,N_9436);
and U9663 (N_9663,N_9486,N_9260);
or U9664 (N_9664,N_9469,N_9325);
and U9665 (N_9665,N_9403,N_9323);
nand U9666 (N_9666,N_9361,N_9419);
xor U9667 (N_9667,N_9255,N_9286);
xor U9668 (N_9668,N_9283,N_9387);
nor U9669 (N_9669,N_9405,N_9282);
or U9670 (N_9670,N_9386,N_9302);
nand U9671 (N_9671,N_9350,N_9496);
nor U9672 (N_9672,N_9422,N_9428);
nor U9673 (N_9673,N_9287,N_9253);
xnor U9674 (N_9674,N_9487,N_9262);
nor U9675 (N_9675,N_9486,N_9466);
xor U9676 (N_9676,N_9414,N_9299);
and U9677 (N_9677,N_9417,N_9445);
and U9678 (N_9678,N_9255,N_9372);
xnor U9679 (N_9679,N_9350,N_9376);
nand U9680 (N_9680,N_9305,N_9382);
nand U9681 (N_9681,N_9349,N_9384);
or U9682 (N_9682,N_9342,N_9323);
nand U9683 (N_9683,N_9259,N_9348);
nor U9684 (N_9684,N_9486,N_9406);
or U9685 (N_9685,N_9495,N_9310);
or U9686 (N_9686,N_9302,N_9387);
nand U9687 (N_9687,N_9269,N_9459);
and U9688 (N_9688,N_9468,N_9319);
nand U9689 (N_9689,N_9324,N_9347);
and U9690 (N_9690,N_9433,N_9342);
nand U9691 (N_9691,N_9421,N_9385);
or U9692 (N_9692,N_9419,N_9376);
xor U9693 (N_9693,N_9273,N_9458);
or U9694 (N_9694,N_9427,N_9316);
nand U9695 (N_9695,N_9353,N_9464);
or U9696 (N_9696,N_9421,N_9325);
nor U9697 (N_9697,N_9283,N_9258);
xor U9698 (N_9698,N_9274,N_9322);
nand U9699 (N_9699,N_9497,N_9277);
and U9700 (N_9700,N_9380,N_9392);
nor U9701 (N_9701,N_9320,N_9414);
and U9702 (N_9702,N_9477,N_9343);
xnor U9703 (N_9703,N_9388,N_9308);
or U9704 (N_9704,N_9301,N_9306);
nor U9705 (N_9705,N_9404,N_9489);
or U9706 (N_9706,N_9352,N_9404);
or U9707 (N_9707,N_9388,N_9394);
xnor U9708 (N_9708,N_9412,N_9408);
or U9709 (N_9709,N_9424,N_9355);
or U9710 (N_9710,N_9378,N_9362);
and U9711 (N_9711,N_9463,N_9264);
nor U9712 (N_9712,N_9455,N_9341);
xor U9713 (N_9713,N_9394,N_9469);
nor U9714 (N_9714,N_9368,N_9416);
nand U9715 (N_9715,N_9470,N_9480);
xor U9716 (N_9716,N_9269,N_9407);
and U9717 (N_9717,N_9487,N_9410);
nor U9718 (N_9718,N_9372,N_9389);
xor U9719 (N_9719,N_9295,N_9256);
or U9720 (N_9720,N_9474,N_9491);
nand U9721 (N_9721,N_9474,N_9375);
nand U9722 (N_9722,N_9406,N_9255);
or U9723 (N_9723,N_9457,N_9317);
and U9724 (N_9724,N_9468,N_9314);
or U9725 (N_9725,N_9349,N_9482);
xor U9726 (N_9726,N_9369,N_9388);
nor U9727 (N_9727,N_9459,N_9483);
or U9728 (N_9728,N_9487,N_9484);
and U9729 (N_9729,N_9278,N_9269);
nor U9730 (N_9730,N_9341,N_9340);
or U9731 (N_9731,N_9441,N_9288);
and U9732 (N_9732,N_9399,N_9454);
xnor U9733 (N_9733,N_9303,N_9451);
or U9734 (N_9734,N_9250,N_9493);
nor U9735 (N_9735,N_9482,N_9286);
nand U9736 (N_9736,N_9491,N_9311);
xor U9737 (N_9737,N_9407,N_9315);
nand U9738 (N_9738,N_9447,N_9448);
nand U9739 (N_9739,N_9403,N_9362);
and U9740 (N_9740,N_9418,N_9422);
nand U9741 (N_9741,N_9261,N_9332);
and U9742 (N_9742,N_9437,N_9257);
or U9743 (N_9743,N_9396,N_9392);
or U9744 (N_9744,N_9433,N_9413);
or U9745 (N_9745,N_9440,N_9351);
nor U9746 (N_9746,N_9436,N_9380);
or U9747 (N_9747,N_9440,N_9362);
xnor U9748 (N_9748,N_9254,N_9459);
and U9749 (N_9749,N_9438,N_9257);
nand U9750 (N_9750,N_9593,N_9529);
nand U9751 (N_9751,N_9614,N_9734);
nor U9752 (N_9752,N_9581,N_9696);
nand U9753 (N_9753,N_9578,N_9711);
nand U9754 (N_9754,N_9673,N_9690);
and U9755 (N_9755,N_9516,N_9528);
nand U9756 (N_9756,N_9553,N_9557);
or U9757 (N_9757,N_9710,N_9740);
xor U9758 (N_9758,N_9548,N_9527);
or U9759 (N_9759,N_9642,N_9598);
nor U9760 (N_9760,N_9520,N_9532);
or U9761 (N_9761,N_9742,N_9725);
nor U9762 (N_9762,N_9621,N_9603);
nor U9763 (N_9763,N_9706,N_9641);
xor U9764 (N_9764,N_9580,N_9712);
nor U9765 (N_9765,N_9629,N_9656);
xor U9766 (N_9766,N_9654,N_9661);
nor U9767 (N_9767,N_9558,N_9594);
or U9768 (N_9768,N_9583,N_9645);
nand U9769 (N_9769,N_9501,N_9615);
and U9770 (N_9770,N_9585,N_9588);
and U9771 (N_9771,N_9650,N_9522);
or U9772 (N_9772,N_9510,N_9688);
and U9773 (N_9773,N_9533,N_9617);
and U9774 (N_9774,N_9502,N_9749);
and U9775 (N_9775,N_9745,N_9554);
or U9776 (N_9776,N_9570,N_9653);
or U9777 (N_9777,N_9595,N_9640);
or U9778 (N_9778,N_9544,N_9525);
or U9779 (N_9779,N_9715,N_9552);
nand U9780 (N_9780,N_9589,N_9675);
nand U9781 (N_9781,N_9550,N_9722);
or U9782 (N_9782,N_9514,N_9545);
xor U9783 (N_9783,N_9733,N_9607);
nor U9784 (N_9784,N_9649,N_9700);
and U9785 (N_9785,N_9587,N_9647);
and U9786 (N_9786,N_9542,N_9663);
nand U9787 (N_9787,N_9644,N_9625);
xnor U9788 (N_9788,N_9618,N_9597);
and U9789 (N_9789,N_9718,N_9643);
nor U9790 (N_9790,N_9592,N_9569);
or U9791 (N_9791,N_9692,N_9600);
nor U9792 (N_9792,N_9687,N_9665);
or U9793 (N_9793,N_9508,N_9743);
or U9794 (N_9794,N_9674,N_9596);
or U9795 (N_9795,N_9556,N_9691);
xor U9796 (N_9796,N_9567,N_9561);
or U9797 (N_9797,N_9504,N_9681);
nor U9798 (N_9798,N_9739,N_9731);
nand U9799 (N_9799,N_9735,N_9748);
nor U9800 (N_9800,N_9565,N_9573);
xor U9801 (N_9801,N_9659,N_9500);
nor U9802 (N_9802,N_9684,N_9732);
and U9803 (N_9803,N_9666,N_9686);
and U9804 (N_9804,N_9543,N_9513);
xor U9805 (N_9805,N_9623,N_9697);
nor U9806 (N_9806,N_9729,N_9721);
xnor U9807 (N_9807,N_9536,N_9616);
xor U9808 (N_9808,N_9652,N_9677);
and U9809 (N_9809,N_9564,N_9579);
xor U9810 (N_9810,N_9628,N_9605);
nor U9811 (N_9811,N_9541,N_9609);
or U9812 (N_9812,N_9546,N_9519);
and U9813 (N_9813,N_9727,N_9699);
and U9814 (N_9814,N_9584,N_9606);
nor U9815 (N_9815,N_9555,N_9620);
nand U9816 (N_9816,N_9648,N_9512);
xnor U9817 (N_9817,N_9702,N_9651);
or U9818 (N_9818,N_9637,N_9575);
xnor U9819 (N_9819,N_9586,N_9549);
xor U9820 (N_9820,N_9540,N_9678);
xor U9821 (N_9821,N_9568,N_9622);
nand U9822 (N_9822,N_9746,N_9559);
nor U9823 (N_9823,N_9703,N_9517);
nor U9824 (N_9824,N_9741,N_9657);
nor U9825 (N_9825,N_9724,N_9682);
nand U9826 (N_9826,N_9719,N_9693);
nand U9827 (N_9827,N_9679,N_9547);
nand U9828 (N_9828,N_9574,N_9638);
and U9829 (N_9829,N_9515,N_9672);
nand U9830 (N_9830,N_9744,N_9627);
and U9831 (N_9831,N_9613,N_9671);
nand U9832 (N_9832,N_9599,N_9572);
nor U9833 (N_9833,N_9523,N_9660);
xor U9834 (N_9834,N_9576,N_9505);
nand U9835 (N_9835,N_9612,N_9658);
and U9836 (N_9836,N_9705,N_9503);
xnor U9837 (N_9837,N_9631,N_9602);
or U9838 (N_9838,N_9726,N_9611);
xnor U9839 (N_9839,N_9701,N_9716);
and U9840 (N_9840,N_9539,N_9591);
and U9841 (N_9841,N_9608,N_9689);
nand U9842 (N_9842,N_9680,N_9582);
nand U9843 (N_9843,N_9619,N_9624);
nand U9844 (N_9844,N_9590,N_9626);
or U9845 (N_9845,N_9737,N_9521);
xnor U9846 (N_9846,N_9634,N_9566);
xnor U9847 (N_9847,N_9538,N_9695);
xor U9848 (N_9848,N_9662,N_9537);
nor U9849 (N_9849,N_9670,N_9562);
nor U9850 (N_9850,N_9604,N_9630);
nand U9851 (N_9851,N_9563,N_9531);
nand U9852 (N_9852,N_9669,N_9571);
nand U9853 (N_9853,N_9655,N_9635);
xor U9854 (N_9854,N_9511,N_9676);
nor U9855 (N_9855,N_9723,N_9713);
xor U9856 (N_9856,N_9714,N_9560);
xnor U9857 (N_9857,N_9534,N_9535);
or U9858 (N_9858,N_9524,N_9633);
or U9859 (N_9859,N_9506,N_9639);
xnor U9860 (N_9860,N_9728,N_9704);
nand U9861 (N_9861,N_9518,N_9601);
nor U9862 (N_9862,N_9632,N_9736);
xnor U9863 (N_9863,N_9526,N_9610);
and U9864 (N_9864,N_9683,N_9730);
and U9865 (N_9865,N_9530,N_9646);
or U9866 (N_9866,N_9507,N_9551);
and U9867 (N_9867,N_9709,N_9720);
nor U9868 (N_9868,N_9738,N_9694);
nand U9869 (N_9869,N_9664,N_9577);
and U9870 (N_9870,N_9667,N_9708);
nor U9871 (N_9871,N_9685,N_9717);
or U9872 (N_9872,N_9668,N_9636);
and U9873 (N_9873,N_9698,N_9747);
or U9874 (N_9874,N_9509,N_9707);
or U9875 (N_9875,N_9566,N_9578);
xor U9876 (N_9876,N_9687,N_9677);
nor U9877 (N_9877,N_9600,N_9732);
and U9878 (N_9878,N_9676,N_9687);
nand U9879 (N_9879,N_9500,N_9570);
nand U9880 (N_9880,N_9547,N_9731);
xor U9881 (N_9881,N_9594,N_9569);
or U9882 (N_9882,N_9734,N_9517);
or U9883 (N_9883,N_9709,N_9644);
and U9884 (N_9884,N_9724,N_9717);
nand U9885 (N_9885,N_9694,N_9661);
nor U9886 (N_9886,N_9628,N_9551);
xor U9887 (N_9887,N_9524,N_9646);
or U9888 (N_9888,N_9690,N_9728);
nand U9889 (N_9889,N_9694,N_9698);
xnor U9890 (N_9890,N_9655,N_9587);
nor U9891 (N_9891,N_9728,N_9738);
and U9892 (N_9892,N_9513,N_9590);
xnor U9893 (N_9893,N_9518,N_9565);
or U9894 (N_9894,N_9670,N_9516);
nor U9895 (N_9895,N_9719,N_9514);
or U9896 (N_9896,N_9657,N_9565);
nand U9897 (N_9897,N_9727,N_9593);
or U9898 (N_9898,N_9600,N_9654);
or U9899 (N_9899,N_9663,N_9659);
or U9900 (N_9900,N_9736,N_9619);
or U9901 (N_9901,N_9741,N_9556);
or U9902 (N_9902,N_9719,N_9731);
or U9903 (N_9903,N_9748,N_9653);
nor U9904 (N_9904,N_9607,N_9745);
xor U9905 (N_9905,N_9579,N_9537);
or U9906 (N_9906,N_9678,N_9749);
and U9907 (N_9907,N_9629,N_9642);
and U9908 (N_9908,N_9695,N_9592);
and U9909 (N_9909,N_9580,N_9645);
nor U9910 (N_9910,N_9550,N_9658);
nor U9911 (N_9911,N_9667,N_9678);
xnor U9912 (N_9912,N_9635,N_9529);
or U9913 (N_9913,N_9550,N_9642);
xnor U9914 (N_9914,N_9543,N_9587);
nor U9915 (N_9915,N_9554,N_9672);
xnor U9916 (N_9916,N_9677,N_9538);
xor U9917 (N_9917,N_9591,N_9677);
nand U9918 (N_9918,N_9514,N_9519);
nand U9919 (N_9919,N_9627,N_9696);
nand U9920 (N_9920,N_9692,N_9696);
xor U9921 (N_9921,N_9729,N_9636);
nor U9922 (N_9922,N_9607,N_9579);
nor U9923 (N_9923,N_9526,N_9669);
xnor U9924 (N_9924,N_9537,N_9655);
nand U9925 (N_9925,N_9523,N_9687);
xor U9926 (N_9926,N_9700,N_9549);
or U9927 (N_9927,N_9645,N_9628);
nand U9928 (N_9928,N_9631,N_9515);
xnor U9929 (N_9929,N_9664,N_9667);
nand U9930 (N_9930,N_9679,N_9625);
and U9931 (N_9931,N_9556,N_9661);
and U9932 (N_9932,N_9667,N_9675);
and U9933 (N_9933,N_9511,N_9566);
xnor U9934 (N_9934,N_9531,N_9590);
nor U9935 (N_9935,N_9533,N_9616);
and U9936 (N_9936,N_9650,N_9693);
and U9937 (N_9937,N_9590,N_9504);
nand U9938 (N_9938,N_9672,N_9503);
and U9939 (N_9939,N_9512,N_9577);
nand U9940 (N_9940,N_9710,N_9598);
nor U9941 (N_9941,N_9638,N_9594);
nand U9942 (N_9942,N_9677,N_9528);
or U9943 (N_9943,N_9635,N_9692);
nand U9944 (N_9944,N_9521,N_9695);
xnor U9945 (N_9945,N_9543,N_9644);
xor U9946 (N_9946,N_9591,N_9664);
and U9947 (N_9947,N_9691,N_9593);
xnor U9948 (N_9948,N_9530,N_9558);
xnor U9949 (N_9949,N_9617,N_9530);
and U9950 (N_9950,N_9532,N_9583);
or U9951 (N_9951,N_9541,N_9514);
or U9952 (N_9952,N_9695,N_9616);
or U9953 (N_9953,N_9647,N_9634);
and U9954 (N_9954,N_9730,N_9635);
xnor U9955 (N_9955,N_9543,N_9746);
xor U9956 (N_9956,N_9512,N_9550);
nand U9957 (N_9957,N_9508,N_9635);
nor U9958 (N_9958,N_9716,N_9630);
nor U9959 (N_9959,N_9724,N_9660);
and U9960 (N_9960,N_9637,N_9684);
xor U9961 (N_9961,N_9592,N_9553);
nand U9962 (N_9962,N_9722,N_9524);
or U9963 (N_9963,N_9700,N_9568);
nand U9964 (N_9964,N_9618,N_9525);
xor U9965 (N_9965,N_9684,N_9602);
nor U9966 (N_9966,N_9572,N_9595);
xor U9967 (N_9967,N_9642,N_9638);
and U9968 (N_9968,N_9704,N_9646);
and U9969 (N_9969,N_9716,N_9549);
xnor U9970 (N_9970,N_9583,N_9621);
nand U9971 (N_9971,N_9637,N_9577);
nor U9972 (N_9972,N_9602,N_9667);
and U9973 (N_9973,N_9697,N_9635);
nand U9974 (N_9974,N_9696,N_9511);
nor U9975 (N_9975,N_9686,N_9639);
and U9976 (N_9976,N_9742,N_9654);
and U9977 (N_9977,N_9537,N_9555);
and U9978 (N_9978,N_9604,N_9635);
nand U9979 (N_9979,N_9641,N_9536);
xnor U9980 (N_9980,N_9642,N_9608);
and U9981 (N_9981,N_9703,N_9580);
nor U9982 (N_9982,N_9546,N_9645);
nand U9983 (N_9983,N_9651,N_9539);
and U9984 (N_9984,N_9664,N_9594);
and U9985 (N_9985,N_9702,N_9626);
or U9986 (N_9986,N_9567,N_9658);
nor U9987 (N_9987,N_9733,N_9586);
xor U9988 (N_9988,N_9667,N_9534);
nor U9989 (N_9989,N_9713,N_9615);
and U9990 (N_9990,N_9706,N_9652);
xnor U9991 (N_9991,N_9650,N_9611);
nand U9992 (N_9992,N_9653,N_9596);
or U9993 (N_9993,N_9622,N_9728);
xnor U9994 (N_9994,N_9632,N_9693);
and U9995 (N_9995,N_9740,N_9525);
xor U9996 (N_9996,N_9612,N_9692);
nor U9997 (N_9997,N_9626,N_9567);
and U9998 (N_9998,N_9657,N_9595);
nand U9999 (N_9999,N_9515,N_9742);
nand U10000 (N_10000,N_9767,N_9863);
xnor U10001 (N_10001,N_9795,N_9770);
xnor U10002 (N_10002,N_9983,N_9978);
and U10003 (N_10003,N_9921,N_9977);
and U10004 (N_10004,N_9836,N_9968);
nor U10005 (N_10005,N_9932,N_9781);
and U10006 (N_10006,N_9786,N_9934);
xnor U10007 (N_10007,N_9779,N_9828);
nor U10008 (N_10008,N_9778,N_9876);
or U10009 (N_10009,N_9787,N_9850);
or U10010 (N_10010,N_9973,N_9829);
xor U10011 (N_10011,N_9844,N_9764);
xnor U10012 (N_10012,N_9999,N_9814);
or U10013 (N_10013,N_9939,N_9959);
or U10014 (N_10014,N_9990,N_9841);
and U10015 (N_10015,N_9963,N_9857);
nand U10016 (N_10016,N_9759,N_9957);
xnor U10017 (N_10017,N_9879,N_9794);
and U10018 (N_10018,N_9886,N_9905);
nand U10019 (N_10019,N_9773,N_9981);
and U10020 (N_10020,N_9871,N_9769);
nand U10021 (N_10021,N_9907,N_9910);
xnor U10022 (N_10022,N_9766,N_9761);
xnor U10023 (N_10023,N_9837,N_9803);
xor U10024 (N_10024,N_9908,N_9797);
and U10025 (N_10025,N_9793,N_9920);
and U10026 (N_10026,N_9943,N_9987);
or U10027 (N_10027,N_9972,N_9895);
nor U10028 (N_10028,N_9897,N_9866);
nor U10029 (N_10029,N_9979,N_9812);
xnor U10030 (N_10030,N_9833,N_9783);
xor U10031 (N_10031,N_9865,N_9958);
nor U10032 (N_10032,N_9901,N_9950);
nor U10033 (N_10033,N_9845,N_9894);
nand U10034 (N_10034,N_9855,N_9808);
xnor U10035 (N_10035,N_9846,N_9853);
nor U10036 (N_10036,N_9928,N_9782);
xnor U10037 (N_10037,N_9929,N_9776);
nor U10038 (N_10038,N_9838,N_9917);
and U10039 (N_10039,N_9948,N_9811);
and U10040 (N_10040,N_9935,N_9964);
and U10041 (N_10041,N_9751,N_9996);
or U10042 (N_10042,N_9989,N_9951);
and U10043 (N_10043,N_9896,N_9768);
nor U10044 (N_10044,N_9997,N_9818);
nand U10045 (N_10045,N_9822,N_9898);
or U10046 (N_10046,N_9835,N_9757);
and U10047 (N_10047,N_9780,N_9752);
or U10048 (N_10048,N_9946,N_9777);
or U10049 (N_10049,N_9931,N_9792);
nand U10050 (N_10050,N_9930,N_9810);
xor U10051 (N_10051,N_9848,N_9960);
xor U10052 (N_10052,N_9949,N_9824);
xor U10053 (N_10053,N_9861,N_9914);
xor U10054 (N_10054,N_9750,N_9937);
or U10055 (N_10055,N_9839,N_9944);
xnor U10056 (N_10056,N_9980,N_9851);
nor U10057 (N_10057,N_9970,N_9969);
or U10058 (N_10058,N_9756,N_9762);
xnor U10059 (N_10059,N_9878,N_9801);
nand U10060 (N_10060,N_9986,N_9900);
or U10061 (N_10061,N_9933,N_9947);
and U10062 (N_10062,N_9892,N_9916);
nor U10063 (N_10063,N_9860,N_9988);
or U10064 (N_10064,N_9925,N_9985);
or U10065 (N_10065,N_9758,N_9961);
nand U10066 (N_10066,N_9971,N_9984);
xor U10067 (N_10067,N_9965,N_9877);
and U10068 (N_10068,N_9912,N_9952);
nand U10069 (N_10069,N_9940,N_9854);
xnor U10070 (N_10070,N_9904,N_9753);
nand U10071 (N_10071,N_9809,N_9923);
xor U10072 (N_10072,N_9800,N_9856);
or U10073 (N_10073,N_9956,N_9823);
nand U10074 (N_10074,N_9870,N_9843);
or U10075 (N_10075,N_9785,N_9874);
or U10076 (N_10076,N_9941,N_9906);
nand U10077 (N_10077,N_9884,N_9899);
and U10078 (N_10078,N_9890,N_9991);
nor U10079 (N_10079,N_9755,N_9831);
nand U10080 (N_10080,N_9887,N_9953);
xnor U10081 (N_10081,N_9967,N_9820);
xnor U10082 (N_10082,N_9775,N_9966);
nand U10083 (N_10083,N_9821,N_9858);
and U10084 (N_10084,N_9789,N_9784);
nor U10085 (N_10085,N_9926,N_9883);
and U10086 (N_10086,N_9765,N_9903);
nor U10087 (N_10087,N_9873,N_9847);
xnor U10088 (N_10088,N_9815,N_9992);
nor U10089 (N_10089,N_9927,N_9882);
nor U10090 (N_10090,N_9771,N_9813);
or U10091 (N_10091,N_9954,N_9834);
or U10092 (N_10092,N_9888,N_9826);
and U10093 (N_10093,N_9942,N_9945);
or U10094 (N_10094,N_9852,N_9902);
xor U10095 (N_10095,N_9788,N_9763);
xnor U10096 (N_10096,N_9976,N_9993);
xor U10097 (N_10097,N_9868,N_9772);
or U10098 (N_10098,N_9938,N_9842);
nand U10099 (N_10099,N_9840,N_9982);
and U10100 (N_10100,N_9881,N_9754);
nor U10101 (N_10101,N_9790,N_9832);
nand U10102 (N_10102,N_9875,N_9805);
nand U10103 (N_10103,N_9859,N_9798);
or U10104 (N_10104,N_9799,N_9911);
nand U10105 (N_10105,N_9975,N_9915);
and U10106 (N_10106,N_9849,N_9867);
or U10107 (N_10107,N_9955,N_9807);
and U10108 (N_10108,N_9919,N_9994);
nand U10109 (N_10109,N_9774,N_9885);
nor U10110 (N_10110,N_9802,N_9936);
xor U10111 (N_10111,N_9825,N_9827);
nor U10112 (N_10112,N_9891,N_9889);
nor U10113 (N_10113,N_9962,N_9816);
nand U10114 (N_10114,N_9872,N_9974);
or U10115 (N_10115,N_9869,N_9880);
and U10116 (N_10116,N_9819,N_9830);
or U10117 (N_10117,N_9893,N_9760);
nand U10118 (N_10118,N_9862,N_9804);
and U10119 (N_10119,N_9924,N_9913);
and U10120 (N_10120,N_9998,N_9806);
and U10121 (N_10121,N_9995,N_9918);
nor U10122 (N_10122,N_9817,N_9796);
and U10123 (N_10123,N_9909,N_9922);
xor U10124 (N_10124,N_9791,N_9864);
or U10125 (N_10125,N_9819,N_9829);
nand U10126 (N_10126,N_9861,N_9957);
nor U10127 (N_10127,N_9816,N_9998);
nor U10128 (N_10128,N_9909,N_9962);
nand U10129 (N_10129,N_9927,N_9837);
xnor U10130 (N_10130,N_9870,N_9836);
nand U10131 (N_10131,N_9984,N_9988);
and U10132 (N_10132,N_9973,N_9992);
and U10133 (N_10133,N_9894,N_9963);
and U10134 (N_10134,N_9774,N_9781);
xor U10135 (N_10135,N_9884,N_9754);
nor U10136 (N_10136,N_9868,N_9943);
nand U10137 (N_10137,N_9977,N_9949);
xnor U10138 (N_10138,N_9822,N_9880);
or U10139 (N_10139,N_9793,N_9886);
xnor U10140 (N_10140,N_9760,N_9787);
nand U10141 (N_10141,N_9948,N_9801);
and U10142 (N_10142,N_9905,N_9772);
or U10143 (N_10143,N_9800,N_9787);
xor U10144 (N_10144,N_9795,N_9988);
and U10145 (N_10145,N_9989,N_9830);
and U10146 (N_10146,N_9780,N_9895);
and U10147 (N_10147,N_9780,N_9936);
nor U10148 (N_10148,N_9876,N_9806);
and U10149 (N_10149,N_9957,N_9947);
or U10150 (N_10150,N_9881,N_9850);
or U10151 (N_10151,N_9999,N_9977);
nor U10152 (N_10152,N_9943,N_9873);
xnor U10153 (N_10153,N_9766,N_9842);
nand U10154 (N_10154,N_9881,N_9902);
or U10155 (N_10155,N_9977,N_9764);
nor U10156 (N_10156,N_9962,N_9770);
or U10157 (N_10157,N_9996,N_9843);
and U10158 (N_10158,N_9944,N_9767);
or U10159 (N_10159,N_9795,N_9832);
xor U10160 (N_10160,N_9886,N_9871);
or U10161 (N_10161,N_9909,N_9872);
or U10162 (N_10162,N_9904,N_9981);
or U10163 (N_10163,N_9964,N_9886);
or U10164 (N_10164,N_9880,N_9885);
or U10165 (N_10165,N_9893,N_9842);
nand U10166 (N_10166,N_9785,N_9821);
xnor U10167 (N_10167,N_9970,N_9829);
nor U10168 (N_10168,N_9834,N_9765);
xor U10169 (N_10169,N_9933,N_9994);
xor U10170 (N_10170,N_9936,N_9949);
nand U10171 (N_10171,N_9932,N_9953);
or U10172 (N_10172,N_9916,N_9987);
nand U10173 (N_10173,N_9751,N_9844);
and U10174 (N_10174,N_9856,N_9950);
xnor U10175 (N_10175,N_9806,N_9837);
nor U10176 (N_10176,N_9974,N_9858);
and U10177 (N_10177,N_9842,N_9964);
and U10178 (N_10178,N_9837,N_9916);
nand U10179 (N_10179,N_9927,N_9851);
and U10180 (N_10180,N_9891,N_9864);
or U10181 (N_10181,N_9893,N_9915);
or U10182 (N_10182,N_9910,N_9911);
xnor U10183 (N_10183,N_9839,N_9917);
xor U10184 (N_10184,N_9756,N_9979);
and U10185 (N_10185,N_9785,N_9987);
nand U10186 (N_10186,N_9766,N_9851);
and U10187 (N_10187,N_9851,N_9865);
or U10188 (N_10188,N_9895,N_9919);
or U10189 (N_10189,N_9796,N_9990);
or U10190 (N_10190,N_9851,N_9883);
and U10191 (N_10191,N_9883,N_9751);
and U10192 (N_10192,N_9763,N_9902);
nor U10193 (N_10193,N_9772,N_9823);
or U10194 (N_10194,N_9832,N_9893);
or U10195 (N_10195,N_9963,N_9785);
nor U10196 (N_10196,N_9809,N_9826);
or U10197 (N_10197,N_9957,N_9799);
nor U10198 (N_10198,N_9920,N_9855);
nand U10199 (N_10199,N_9771,N_9950);
and U10200 (N_10200,N_9919,N_9978);
xnor U10201 (N_10201,N_9856,N_9972);
or U10202 (N_10202,N_9812,N_9831);
nand U10203 (N_10203,N_9957,N_9830);
nand U10204 (N_10204,N_9764,N_9867);
nor U10205 (N_10205,N_9973,N_9902);
nor U10206 (N_10206,N_9871,N_9971);
and U10207 (N_10207,N_9932,N_9867);
nand U10208 (N_10208,N_9817,N_9779);
nand U10209 (N_10209,N_9756,N_9890);
nand U10210 (N_10210,N_9830,N_9766);
nand U10211 (N_10211,N_9783,N_9845);
xor U10212 (N_10212,N_9793,N_9820);
nor U10213 (N_10213,N_9991,N_9854);
nor U10214 (N_10214,N_9924,N_9931);
xor U10215 (N_10215,N_9833,N_9990);
xor U10216 (N_10216,N_9952,N_9841);
or U10217 (N_10217,N_9900,N_9962);
nand U10218 (N_10218,N_9921,N_9910);
nor U10219 (N_10219,N_9836,N_9817);
nor U10220 (N_10220,N_9874,N_9836);
nand U10221 (N_10221,N_9857,N_9990);
or U10222 (N_10222,N_9859,N_9825);
nand U10223 (N_10223,N_9877,N_9828);
nand U10224 (N_10224,N_9818,N_9988);
nor U10225 (N_10225,N_9799,N_9932);
or U10226 (N_10226,N_9921,N_9999);
xor U10227 (N_10227,N_9912,N_9866);
nand U10228 (N_10228,N_9831,N_9759);
xor U10229 (N_10229,N_9911,N_9899);
nand U10230 (N_10230,N_9949,N_9755);
nand U10231 (N_10231,N_9988,N_9947);
nand U10232 (N_10232,N_9792,N_9922);
xor U10233 (N_10233,N_9887,N_9756);
or U10234 (N_10234,N_9759,N_9878);
or U10235 (N_10235,N_9868,N_9823);
and U10236 (N_10236,N_9939,N_9862);
nand U10237 (N_10237,N_9866,N_9874);
nand U10238 (N_10238,N_9878,N_9876);
xor U10239 (N_10239,N_9763,N_9899);
or U10240 (N_10240,N_9766,N_9970);
or U10241 (N_10241,N_9872,N_9915);
xnor U10242 (N_10242,N_9849,N_9788);
nor U10243 (N_10243,N_9955,N_9859);
and U10244 (N_10244,N_9973,N_9830);
or U10245 (N_10245,N_9853,N_9776);
nor U10246 (N_10246,N_9806,N_9898);
nand U10247 (N_10247,N_9750,N_9763);
xor U10248 (N_10248,N_9875,N_9904);
nor U10249 (N_10249,N_9991,N_9907);
xnor U10250 (N_10250,N_10135,N_10205);
or U10251 (N_10251,N_10060,N_10078);
nor U10252 (N_10252,N_10087,N_10005);
nand U10253 (N_10253,N_10222,N_10168);
xnor U10254 (N_10254,N_10185,N_10088);
nor U10255 (N_10255,N_10158,N_10100);
or U10256 (N_10256,N_10031,N_10022);
and U10257 (N_10257,N_10121,N_10244);
and U10258 (N_10258,N_10011,N_10091);
or U10259 (N_10259,N_10124,N_10196);
nand U10260 (N_10260,N_10190,N_10199);
xnor U10261 (N_10261,N_10177,N_10148);
nor U10262 (N_10262,N_10044,N_10113);
and U10263 (N_10263,N_10117,N_10136);
nand U10264 (N_10264,N_10049,N_10055);
or U10265 (N_10265,N_10075,N_10242);
nand U10266 (N_10266,N_10125,N_10238);
nor U10267 (N_10267,N_10167,N_10192);
and U10268 (N_10268,N_10206,N_10154);
xnor U10269 (N_10269,N_10162,N_10059);
nor U10270 (N_10270,N_10133,N_10226);
xor U10271 (N_10271,N_10051,N_10095);
and U10272 (N_10272,N_10183,N_10076);
xor U10273 (N_10273,N_10042,N_10062);
xor U10274 (N_10274,N_10093,N_10215);
nand U10275 (N_10275,N_10094,N_10203);
nand U10276 (N_10276,N_10026,N_10126);
xor U10277 (N_10277,N_10046,N_10036);
and U10278 (N_10278,N_10157,N_10116);
nor U10279 (N_10279,N_10020,N_10072);
nand U10280 (N_10280,N_10163,N_10037);
nand U10281 (N_10281,N_10227,N_10128);
xnor U10282 (N_10282,N_10082,N_10077);
nor U10283 (N_10283,N_10234,N_10114);
nor U10284 (N_10284,N_10147,N_10195);
nor U10285 (N_10285,N_10096,N_10006);
or U10286 (N_10286,N_10212,N_10249);
xnor U10287 (N_10287,N_10170,N_10000);
and U10288 (N_10288,N_10235,N_10086);
and U10289 (N_10289,N_10040,N_10023);
and U10290 (N_10290,N_10034,N_10092);
and U10291 (N_10291,N_10200,N_10204);
nand U10292 (N_10292,N_10104,N_10225);
and U10293 (N_10293,N_10240,N_10065);
xor U10294 (N_10294,N_10236,N_10134);
or U10295 (N_10295,N_10129,N_10013);
nand U10296 (N_10296,N_10138,N_10211);
nor U10297 (N_10297,N_10045,N_10039);
nor U10298 (N_10298,N_10053,N_10202);
xor U10299 (N_10299,N_10233,N_10010);
or U10300 (N_10300,N_10207,N_10122);
or U10301 (N_10301,N_10214,N_10180);
nand U10302 (N_10302,N_10109,N_10153);
and U10303 (N_10303,N_10107,N_10182);
and U10304 (N_10304,N_10108,N_10213);
and U10305 (N_10305,N_10230,N_10181);
or U10306 (N_10306,N_10223,N_10210);
or U10307 (N_10307,N_10015,N_10101);
xnor U10308 (N_10308,N_10152,N_10239);
and U10309 (N_10309,N_10145,N_10245);
nand U10310 (N_10310,N_10047,N_10007);
xnor U10311 (N_10311,N_10074,N_10057);
or U10312 (N_10312,N_10019,N_10130);
or U10313 (N_10313,N_10208,N_10149);
nand U10314 (N_10314,N_10179,N_10186);
nor U10315 (N_10315,N_10220,N_10142);
nor U10316 (N_10316,N_10219,N_10194);
and U10317 (N_10317,N_10118,N_10068);
or U10318 (N_10318,N_10127,N_10028);
and U10319 (N_10319,N_10012,N_10171);
nand U10320 (N_10320,N_10033,N_10050);
nor U10321 (N_10321,N_10106,N_10029);
or U10322 (N_10322,N_10178,N_10120);
or U10323 (N_10323,N_10132,N_10216);
xor U10324 (N_10324,N_10054,N_10073);
nand U10325 (N_10325,N_10246,N_10081);
nor U10326 (N_10326,N_10035,N_10080);
and U10327 (N_10327,N_10024,N_10069);
or U10328 (N_10328,N_10009,N_10191);
nor U10329 (N_10329,N_10189,N_10061);
or U10330 (N_10330,N_10218,N_10144);
nor U10331 (N_10331,N_10159,N_10248);
or U10332 (N_10332,N_10139,N_10166);
nor U10333 (N_10333,N_10017,N_10198);
xnor U10334 (N_10334,N_10008,N_10111);
nand U10335 (N_10335,N_10103,N_10030);
nor U10336 (N_10336,N_10197,N_10001);
xnor U10337 (N_10337,N_10105,N_10066);
nor U10338 (N_10338,N_10174,N_10164);
xor U10339 (N_10339,N_10193,N_10131);
and U10340 (N_10340,N_10071,N_10175);
nand U10341 (N_10341,N_10165,N_10064);
nand U10342 (N_10342,N_10123,N_10027);
or U10343 (N_10343,N_10079,N_10089);
nand U10344 (N_10344,N_10228,N_10003);
nand U10345 (N_10345,N_10224,N_10097);
and U10346 (N_10346,N_10004,N_10021);
nor U10347 (N_10347,N_10090,N_10099);
nor U10348 (N_10348,N_10025,N_10188);
and U10349 (N_10349,N_10155,N_10176);
xor U10350 (N_10350,N_10112,N_10085);
or U10351 (N_10351,N_10169,N_10229);
or U10352 (N_10352,N_10115,N_10187);
nand U10353 (N_10353,N_10083,N_10067);
xor U10354 (N_10354,N_10098,N_10070);
nor U10355 (N_10355,N_10151,N_10237);
nor U10356 (N_10356,N_10110,N_10014);
or U10357 (N_10357,N_10063,N_10141);
and U10358 (N_10358,N_10140,N_10143);
xor U10359 (N_10359,N_10146,N_10217);
xnor U10360 (N_10360,N_10043,N_10160);
nor U10361 (N_10361,N_10209,N_10231);
and U10362 (N_10362,N_10156,N_10241);
nor U10363 (N_10363,N_10201,N_10102);
xnor U10364 (N_10364,N_10056,N_10137);
nor U10365 (N_10365,N_10041,N_10243);
and U10366 (N_10366,N_10084,N_10119);
xor U10367 (N_10367,N_10150,N_10232);
nand U10368 (N_10368,N_10172,N_10058);
and U10369 (N_10369,N_10173,N_10048);
xnor U10370 (N_10370,N_10018,N_10052);
or U10371 (N_10371,N_10032,N_10002);
xnor U10372 (N_10372,N_10016,N_10038);
xor U10373 (N_10373,N_10184,N_10161);
and U10374 (N_10374,N_10247,N_10221);
xnor U10375 (N_10375,N_10198,N_10105);
nand U10376 (N_10376,N_10043,N_10197);
xor U10377 (N_10377,N_10032,N_10101);
and U10378 (N_10378,N_10117,N_10081);
or U10379 (N_10379,N_10201,N_10117);
and U10380 (N_10380,N_10041,N_10065);
or U10381 (N_10381,N_10059,N_10083);
nor U10382 (N_10382,N_10134,N_10135);
or U10383 (N_10383,N_10203,N_10035);
or U10384 (N_10384,N_10137,N_10212);
or U10385 (N_10385,N_10142,N_10240);
nor U10386 (N_10386,N_10024,N_10014);
nand U10387 (N_10387,N_10202,N_10174);
nand U10388 (N_10388,N_10211,N_10027);
nor U10389 (N_10389,N_10070,N_10074);
nand U10390 (N_10390,N_10199,N_10125);
and U10391 (N_10391,N_10032,N_10124);
nand U10392 (N_10392,N_10123,N_10031);
and U10393 (N_10393,N_10230,N_10163);
and U10394 (N_10394,N_10068,N_10077);
xor U10395 (N_10395,N_10110,N_10192);
xor U10396 (N_10396,N_10194,N_10119);
nand U10397 (N_10397,N_10177,N_10109);
xor U10398 (N_10398,N_10023,N_10221);
xor U10399 (N_10399,N_10090,N_10237);
nand U10400 (N_10400,N_10166,N_10005);
nor U10401 (N_10401,N_10232,N_10061);
xnor U10402 (N_10402,N_10014,N_10015);
nor U10403 (N_10403,N_10109,N_10035);
and U10404 (N_10404,N_10056,N_10134);
and U10405 (N_10405,N_10174,N_10230);
and U10406 (N_10406,N_10100,N_10000);
and U10407 (N_10407,N_10112,N_10237);
nand U10408 (N_10408,N_10088,N_10072);
xor U10409 (N_10409,N_10209,N_10137);
or U10410 (N_10410,N_10000,N_10035);
xnor U10411 (N_10411,N_10096,N_10066);
xor U10412 (N_10412,N_10106,N_10164);
and U10413 (N_10413,N_10087,N_10200);
xor U10414 (N_10414,N_10238,N_10047);
nand U10415 (N_10415,N_10079,N_10077);
or U10416 (N_10416,N_10191,N_10108);
nor U10417 (N_10417,N_10095,N_10064);
nand U10418 (N_10418,N_10064,N_10086);
and U10419 (N_10419,N_10114,N_10133);
xor U10420 (N_10420,N_10225,N_10164);
xor U10421 (N_10421,N_10045,N_10194);
xnor U10422 (N_10422,N_10012,N_10004);
or U10423 (N_10423,N_10041,N_10058);
and U10424 (N_10424,N_10069,N_10197);
or U10425 (N_10425,N_10101,N_10081);
nand U10426 (N_10426,N_10154,N_10002);
nor U10427 (N_10427,N_10116,N_10235);
nand U10428 (N_10428,N_10230,N_10015);
nand U10429 (N_10429,N_10224,N_10013);
and U10430 (N_10430,N_10019,N_10238);
and U10431 (N_10431,N_10027,N_10157);
nor U10432 (N_10432,N_10107,N_10207);
and U10433 (N_10433,N_10119,N_10104);
nand U10434 (N_10434,N_10133,N_10094);
nand U10435 (N_10435,N_10044,N_10101);
nor U10436 (N_10436,N_10193,N_10010);
nand U10437 (N_10437,N_10198,N_10180);
nand U10438 (N_10438,N_10007,N_10044);
nor U10439 (N_10439,N_10113,N_10245);
nor U10440 (N_10440,N_10245,N_10058);
nand U10441 (N_10441,N_10208,N_10037);
nor U10442 (N_10442,N_10068,N_10231);
or U10443 (N_10443,N_10059,N_10193);
or U10444 (N_10444,N_10111,N_10168);
and U10445 (N_10445,N_10045,N_10243);
or U10446 (N_10446,N_10191,N_10214);
or U10447 (N_10447,N_10175,N_10083);
and U10448 (N_10448,N_10240,N_10187);
or U10449 (N_10449,N_10229,N_10221);
nand U10450 (N_10450,N_10225,N_10098);
nand U10451 (N_10451,N_10072,N_10141);
nor U10452 (N_10452,N_10157,N_10052);
nor U10453 (N_10453,N_10096,N_10248);
nand U10454 (N_10454,N_10167,N_10031);
and U10455 (N_10455,N_10208,N_10024);
or U10456 (N_10456,N_10140,N_10228);
or U10457 (N_10457,N_10121,N_10041);
and U10458 (N_10458,N_10065,N_10201);
nor U10459 (N_10459,N_10189,N_10032);
nand U10460 (N_10460,N_10069,N_10201);
nand U10461 (N_10461,N_10026,N_10234);
nand U10462 (N_10462,N_10048,N_10123);
and U10463 (N_10463,N_10244,N_10063);
or U10464 (N_10464,N_10150,N_10007);
nor U10465 (N_10465,N_10196,N_10022);
nand U10466 (N_10466,N_10024,N_10129);
nor U10467 (N_10467,N_10115,N_10147);
nor U10468 (N_10468,N_10247,N_10213);
and U10469 (N_10469,N_10012,N_10005);
nand U10470 (N_10470,N_10117,N_10166);
xnor U10471 (N_10471,N_10110,N_10126);
xnor U10472 (N_10472,N_10073,N_10088);
and U10473 (N_10473,N_10226,N_10189);
xor U10474 (N_10474,N_10103,N_10142);
or U10475 (N_10475,N_10121,N_10004);
or U10476 (N_10476,N_10178,N_10103);
nand U10477 (N_10477,N_10039,N_10161);
xor U10478 (N_10478,N_10071,N_10065);
nand U10479 (N_10479,N_10138,N_10034);
or U10480 (N_10480,N_10022,N_10237);
and U10481 (N_10481,N_10026,N_10165);
or U10482 (N_10482,N_10029,N_10163);
nor U10483 (N_10483,N_10207,N_10137);
and U10484 (N_10484,N_10046,N_10220);
or U10485 (N_10485,N_10073,N_10209);
nand U10486 (N_10486,N_10071,N_10111);
and U10487 (N_10487,N_10055,N_10133);
or U10488 (N_10488,N_10068,N_10119);
nor U10489 (N_10489,N_10215,N_10018);
and U10490 (N_10490,N_10172,N_10046);
or U10491 (N_10491,N_10099,N_10119);
nand U10492 (N_10492,N_10214,N_10005);
and U10493 (N_10493,N_10119,N_10233);
nor U10494 (N_10494,N_10111,N_10093);
nor U10495 (N_10495,N_10035,N_10185);
and U10496 (N_10496,N_10147,N_10164);
nor U10497 (N_10497,N_10037,N_10164);
nand U10498 (N_10498,N_10029,N_10098);
nor U10499 (N_10499,N_10048,N_10177);
nand U10500 (N_10500,N_10402,N_10251);
or U10501 (N_10501,N_10433,N_10374);
or U10502 (N_10502,N_10396,N_10491);
nor U10503 (N_10503,N_10260,N_10441);
nor U10504 (N_10504,N_10343,N_10315);
nor U10505 (N_10505,N_10366,N_10274);
nor U10506 (N_10506,N_10280,N_10253);
nor U10507 (N_10507,N_10304,N_10470);
nor U10508 (N_10508,N_10313,N_10482);
nand U10509 (N_10509,N_10365,N_10461);
or U10510 (N_10510,N_10383,N_10310);
xnor U10511 (N_10511,N_10475,N_10279);
nor U10512 (N_10512,N_10400,N_10312);
nand U10513 (N_10513,N_10484,N_10275);
or U10514 (N_10514,N_10476,N_10339);
xnor U10515 (N_10515,N_10474,N_10259);
xor U10516 (N_10516,N_10273,N_10330);
xor U10517 (N_10517,N_10466,N_10277);
nor U10518 (N_10518,N_10369,N_10447);
xor U10519 (N_10519,N_10497,N_10303);
nand U10520 (N_10520,N_10490,N_10286);
nor U10521 (N_10521,N_10377,N_10450);
xor U10522 (N_10522,N_10337,N_10326);
nand U10523 (N_10523,N_10266,N_10299);
nand U10524 (N_10524,N_10291,N_10472);
xnor U10525 (N_10525,N_10479,N_10332);
or U10526 (N_10526,N_10424,N_10406);
nor U10527 (N_10527,N_10449,N_10348);
xnor U10528 (N_10528,N_10354,N_10270);
and U10529 (N_10529,N_10397,N_10434);
and U10530 (N_10530,N_10480,N_10483);
or U10531 (N_10531,N_10283,N_10296);
and U10532 (N_10532,N_10281,N_10361);
and U10533 (N_10533,N_10351,N_10294);
nor U10534 (N_10534,N_10499,N_10265);
or U10535 (N_10535,N_10298,N_10427);
and U10536 (N_10536,N_10327,N_10272);
nand U10537 (N_10537,N_10276,N_10368);
and U10538 (N_10538,N_10385,N_10469);
and U10539 (N_10539,N_10496,N_10269);
and U10540 (N_10540,N_10459,N_10321);
or U10541 (N_10541,N_10429,N_10495);
nand U10542 (N_10542,N_10297,N_10443);
nand U10543 (N_10543,N_10408,N_10422);
and U10544 (N_10544,N_10306,N_10454);
nand U10545 (N_10545,N_10381,N_10481);
nor U10546 (N_10546,N_10324,N_10371);
or U10547 (N_10547,N_10372,N_10393);
nand U10548 (N_10548,N_10311,N_10442);
or U10549 (N_10549,N_10421,N_10420);
nand U10550 (N_10550,N_10413,N_10319);
and U10551 (N_10551,N_10473,N_10318);
and U10552 (N_10552,N_10370,N_10367);
nor U10553 (N_10553,N_10460,N_10417);
or U10554 (N_10554,N_10452,N_10255);
or U10555 (N_10555,N_10412,N_10347);
nor U10556 (N_10556,N_10399,N_10358);
xor U10557 (N_10557,N_10320,N_10308);
and U10558 (N_10558,N_10316,N_10256);
nor U10559 (N_10559,N_10389,N_10287);
or U10560 (N_10560,N_10446,N_10468);
nand U10561 (N_10561,N_10426,N_10355);
nand U10562 (N_10562,N_10431,N_10419);
or U10563 (N_10563,N_10464,N_10444);
nand U10564 (N_10564,N_10488,N_10250);
nor U10565 (N_10565,N_10388,N_10493);
and U10566 (N_10566,N_10252,N_10439);
nand U10567 (N_10567,N_10409,N_10489);
nor U10568 (N_10568,N_10329,N_10263);
or U10569 (N_10569,N_10403,N_10349);
xnor U10570 (N_10570,N_10357,N_10317);
xnor U10571 (N_10571,N_10457,N_10325);
xor U10572 (N_10572,N_10432,N_10344);
nor U10573 (N_10573,N_10435,N_10392);
and U10574 (N_10574,N_10328,N_10462);
nand U10575 (N_10575,N_10451,N_10302);
or U10576 (N_10576,N_10382,N_10305);
nor U10577 (N_10577,N_10363,N_10458);
nor U10578 (N_10578,N_10423,N_10282);
or U10579 (N_10579,N_10341,N_10254);
and U10580 (N_10580,N_10331,N_10336);
nor U10581 (N_10581,N_10453,N_10428);
nor U10582 (N_10582,N_10307,N_10338);
xor U10583 (N_10583,N_10465,N_10437);
nor U10584 (N_10584,N_10295,N_10445);
nor U10585 (N_10585,N_10333,N_10362);
or U10586 (N_10586,N_10404,N_10373);
nand U10587 (N_10587,N_10456,N_10498);
and U10588 (N_10588,N_10414,N_10467);
and U10589 (N_10589,N_10418,N_10322);
nand U10590 (N_10590,N_10384,N_10309);
nor U10591 (N_10591,N_10261,N_10395);
or U10592 (N_10592,N_10264,N_10364);
xnor U10593 (N_10593,N_10440,N_10352);
xor U10594 (N_10594,N_10375,N_10268);
nor U10595 (N_10595,N_10293,N_10285);
or U10596 (N_10596,N_10284,N_10314);
nor U10597 (N_10597,N_10415,N_10401);
nor U10598 (N_10598,N_10323,N_10300);
nor U10599 (N_10599,N_10345,N_10463);
nor U10600 (N_10600,N_10492,N_10391);
or U10601 (N_10601,N_10455,N_10376);
and U10602 (N_10602,N_10478,N_10289);
xor U10603 (N_10603,N_10487,N_10335);
or U10604 (N_10604,N_10271,N_10471);
or U10605 (N_10605,N_10438,N_10290);
xor U10606 (N_10606,N_10448,N_10257);
and U10607 (N_10607,N_10436,N_10411);
or U10608 (N_10608,N_10378,N_10346);
xor U10609 (N_10609,N_10379,N_10342);
and U10610 (N_10610,N_10477,N_10334);
xnor U10611 (N_10611,N_10410,N_10380);
xnor U10612 (N_10612,N_10416,N_10267);
nand U10613 (N_10613,N_10425,N_10356);
nor U10614 (N_10614,N_10390,N_10394);
and U10615 (N_10615,N_10288,N_10262);
or U10616 (N_10616,N_10386,N_10405);
xnor U10617 (N_10617,N_10485,N_10292);
nand U10618 (N_10618,N_10340,N_10494);
nor U10619 (N_10619,N_10430,N_10387);
and U10620 (N_10620,N_10359,N_10258);
or U10621 (N_10621,N_10353,N_10301);
or U10622 (N_10622,N_10350,N_10486);
nand U10623 (N_10623,N_10407,N_10360);
xor U10624 (N_10624,N_10278,N_10398);
or U10625 (N_10625,N_10452,N_10444);
and U10626 (N_10626,N_10422,N_10392);
nand U10627 (N_10627,N_10321,N_10326);
nand U10628 (N_10628,N_10426,N_10288);
and U10629 (N_10629,N_10398,N_10476);
nor U10630 (N_10630,N_10323,N_10251);
and U10631 (N_10631,N_10366,N_10350);
xnor U10632 (N_10632,N_10254,N_10494);
nand U10633 (N_10633,N_10280,N_10452);
nand U10634 (N_10634,N_10269,N_10292);
or U10635 (N_10635,N_10310,N_10288);
nor U10636 (N_10636,N_10252,N_10390);
xor U10637 (N_10637,N_10266,N_10339);
xnor U10638 (N_10638,N_10251,N_10417);
xor U10639 (N_10639,N_10304,N_10393);
and U10640 (N_10640,N_10328,N_10361);
and U10641 (N_10641,N_10262,N_10447);
nand U10642 (N_10642,N_10468,N_10253);
and U10643 (N_10643,N_10493,N_10348);
nand U10644 (N_10644,N_10283,N_10399);
nand U10645 (N_10645,N_10481,N_10307);
nor U10646 (N_10646,N_10307,N_10409);
nand U10647 (N_10647,N_10353,N_10484);
or U10648 (N_10648,N_10491,N_10251);
nor U10649 (N_10649,N_10277,N_10479);
nand U10650 (N_10650,N_10353,N_10362);
nand U10651 (N_10651,N_10416,N_10343);
xor U10652 (N_10652,N_10279,N_10337);
and U10653 (N_10653,N_10277,N_10278);
nand U10654 (N_10654,N_10380,N_10479);
nand U10655 (N_10655,N_10300,N_10311);
and U10656 (N_10656,N_10361,N_10292);
and U10657 (N_10657,N_10325,N_10492);
xnor U10658 (N_10658,N_10498,N_10267);
nand U10659 (N_10659,N_10435,N_10386);
nor U10660 (N_10660,N_10412,N_10390);
or U10661 (N_10661,N_10324,N_10365);
and U10662 (N_10662,N_10280,N_10431);
and U10663 (N_10663,N_10399,N_10490);
nand U10664 (N_10664,N_10261,N_10373);
and U10665 (N_10665,N_10402,N_10406);
nand U10666 (N_10666,N_10303,N_10408);
nand U10667 (N_10667,N_10413,N_10345);
xnor U10668 (N_10668,N_10402,N_10291);
nand U10669 (N_10669,N_10294,N_10364);
or U10670 (N_10670,N_10405,N_10351);
nand U10671 (N_10671,N_10287,N_10474);
nor U10672 (N_10672,N_10452,N_10309);
or U10673 (N_10673,N_10489,N_10280);
xnor U10674 (N_10674,N_10374,N_10291);
xnor U10675 (N_10675,N_10455,N_10476);
nor U10676 (N_10676,N_10422,N_10272);
or U10677 (N_10677,N_10273,N_10309);
and U10678 (N_10678,N_10445,N_10339);
nand U10679 (N_10679,N_10352,N_10391);
or U10680 (N_10680,N_10343,N_10462);
nand U10681 (N_10681,N_10268,N_10252);
xnor U10682 (N_10682,N_10429,N_10289);
and U10683 (N_10683,N_10410,N_10306);
and U10684 (N_10684,N_10497,N_10374);
or U10685 (N_10685,N_10253,N_10306);
nor U10686 (N_10686,N_10256,N_10377);
nor U10687 (N_10687,N_10452,N_10450);
or U10688 (N_10688,N_10313,N_10403);
nor U10689 (N_10689,N_10287,N_10424);
xor U10690 (N_10690,N_10367,N_10296);
nor U10691 (N_10691,N_10293,N_10343);
nand U10692 (N_10692,N_10460,N_10272);
nor U10693 (N_10693,N_10476,N_10466);
and U10694 (N_10694,N_10453,N_10319);
nand U10695 (N_10695,N_10358,N_10454);
or U10696 (N_10696,N_10293,N_10289);
and U10697 (N_10697,N_10317,N_10325);
nand U10698 (N_10698,N_10319,N_10411);
and U10699 (N_10699,N_10264,N_10355);
or U10700 (N_10700,N_10372,N_10294);
or U10701 (N_10701,N_10273,N_10267);
or U10702 (N_10702,N_10250,N_10432);
nand U10703 (N_10703,N_10497,N_10458);
and U10704 (N_10704,N_10312,N_10361);
xnor U10705 (N_10705,N_10486,N_10489);
or U10706 (N_10706,N_10421,N_10364);
or U10707 (N_10707,N_10454,N_10443);
nor U10708 (N_10708,N_10354,N_10432);
xor U10709 (N_10709,N_10453,N_10347);
nor U10710 (N_10710,N_10420,N_10317);
or U10711 (N_10711,N_10405,N_10253);
or U10712 (N_10712,N_10330,N_10366);
and U10713 (N_10713,N_10308,N_10259);
nor U10714 (N_10714,N_10393,N_10324);
or U10715 (N_10715,N_10423,N_10317);
nor U10716 (N_10716,N_10264,N_10423);
or U10717 (N_10717,N_10334,N_10298);
xor U10718 (N_10718,N_10332,N_10329);
xnor U10719 (N_10719,N_10285,N_10457);
or U10720 (N_10720,N_10485,N_10336);
xnor U10721 (N_10721,N_10343,N_10460);
or U10722 (N_10722,N_10359,N_10481);
xnor U10723 (N_10723,N_10394,N_10393);
and U10724 (N_10724,N_10405,N_10371);
xnor U10725 (N_10725,N_10415,N_10277);
or U10726 (N_10726,N_10409,N_10306);
or U10727 (N_10727,N_10346,N_10254);
and U10728 (N_10728,N_10365,N_10416);
nor U10729 (N_10729,N_10355,N_10499);
nand U10730 (N_10730,N_10280,N_10442);
or U10731 (N_10731,N_10371,N_10285);
nand U10732 (N_10732,N_10288,N_10420);
xor U10733 (N_10733,N_10334,N_10399);
nand U10734 (N_10734,N_10492,N_10385);
nand U10735 (N_10735,N_10294,N_10394);
xnor U10736 (N_10736,N_10412,N_10407);
nor U10737 (N_10737,N_10492,N_10329);
and U10738 (N_10738,N_10477,N_10263);
xnor U10739 (N_10739,N_10323,N_10363);
xor U10740 (N_10740,N_10376,N_10491);
or U10741 (N_10741,N_10369,N_10407);
and U10742 (N_10742,N_10300,N_10414);
and U10743 (N_10743,N_10449,N_10409);
nand U10744 (N_10744,N_10323,N_10418);
or U10745 (N_10745,N_10272,N_10405);
or U10746 (N_10746,N_10453,N_10366);
and U10747 (N_10747,N_10277,N_10307);
and U10748 (N_10748,N_10357,N_10261);
nor U10749 (N_10749,N_10325,N_10403);
nor U10750 (N_10750,N_10748,N_10631);
xnor U10751 (N_10751,N_10566,N_10561);
nor U10752 (N_10752,N_10592,N_10694);
nand U10753 (N_10753,N_10547,N_10524);
or U10754 (N_10754,N_10539,N_10659);
nand U10755 (N_10755,N_10721,N_10649);
or U10756 (N_10756,N_10571,N_10552);
or U10757 (N_10757,N_10706,N_10682);
nor U10758 (N_10758,N_10641,N_10651);
nand U10759 (N_10759,N_10620,N_10719);
nor U10760 (N_10760,N_10577,N_10500);
or U10761 (N_10761,N_10621,N_10633);
nor U10762 (N_10762,N_10570,N_10676);
xor U10763 (N_10763,N_10588,N_10532);
nor U10764 (N_10764,N_10734,N_10579);
or U10765 (N_10765,N_10614,N_10715);
and U10766 (N_10766,N_10675,N_10622);
nand U10767 (N_10767,N_10521,N_10737);
and U10768 (N_10768,N_10663,N_10615);
nor U10769 (N_10769,N_10697,N_10696);
nor U10770 (N_10770,N_10701,N_10745);
xnor U10771 (N_10771,N_10596,N_10687);
nand U10772 (N_10772,N_10530,N_10638);
and U10773 (N_10773,N_10546,N_10616);
or U10774 (N_10774,N_10670,N_10681);
xnor U10775 (N_10775,N_10514,N_10541);
or U10776 (N_10776,N_10587,N_10518);
and U10777 (N_10777,N_10535,N_10599);
or U10778 (N_10778,N_10644,N_10613);
xor U10779 (N_10779,N_10655,N_10728);
and U10780 (N_10780,N_10685,N_10590);
and U10781 (N_10781,N_10538,N_10511);
and U10782 (N_10782,N_10628,N_10502);
xor U10783 (N_10783,N_10686,N_10553);
xnor U10784 (N_10784,N_10597,N_10700);
nand U10785 (N_10785,N_10662,N_10679);
or U10786 (N_10786,N_10568,N_10704);
nand U10787 (N_10787,N_10680,N_10550);
nor U10788 (N_10788,N_10658,N_10718);
xnor U10789 (N_10789,N_10742,N_10705);
or U10790 (N_10790,N_10564,N_10639);
and U10791 (N_10791,N_10531,N_10747);
and U10792 (N_10792,N_10605,N_10740);
xor U10793 (N_10793,N_10690,N_10643);
xnor U10794 (N_10794,N_10657,N_10743);
xnor U10795 (N_10795,N_10674,N_10708);
and U10796 (N_10796,N_10572,N_10732);
and U10797 (N_10797,N_10668,N_10723);
or U10798 (N_10798,N_10640,N_10736);
xor U10799 (N_10799,N_10600,N_10543);
nand U10800 (N_10800,N_10529,N_10664);
nor U10801 (N_10801,N_10666,N_10602);
nor U10802 (N_10802,N_10729,N_10556);
or U10803 (N_10803,N_10523,N_10671);
xnor U10804 (N_10804,N_10584,N_10519);
or U10805 (N_10805,N_10522,N_10578);
xnor U10806 (N_10806,N_10510,N_10576);
or U10807 (N_10807,N_10717,N_10710);
and U10808 (N_10808,N_10626,N_10610);
xor U10809 (N_10809,N_10595,N_10582);
xor U10810 (N_10810,N_10581,N_10515);
nand U10811 (N_10811,N_10637,N_10669);
nand U10812 (N_10812,N_10738,N_10630);
nor U10813 (N_10813,N_10544,N_10563);
or U10814 (N_10814,N_10709,N_10665);
and U10815 (N_10815,N_10567,N_10629);
xor U10816 (N_10816,N_10560,N_10730);
nor U10817 (N_10817,N_10635,N_10648);
nand U10818 (N_10818,N_10517,N_10672);
nand U10819 (N_10819,N_10661,N_10702);
and U10820 (N_10820,N_10632,N_10739);
xnor U10821 (N_10821,N_10727,N_10591);
xor U10822 (N_10822,N_10619,N_10609);
nor U10823 (N_10823,N_10562,N_10735);
and U10824 (N_10824,N_10548,N_10513);
xor U10825 (N_10825,N_10545,N_10692);
nor U10826 (N_10826,N_10501,N_10520);
or U10827 (N_10827,N_10527,N_10693);
and U10828 (N_10828,N_10627,N_10575);
nand U10829 (N_10829,N_10646,N_10713);
nand U10830 (N_10830,N_10683,N_10606);
and U10831 (N_10831,N_10589,N_10583);
and U10832 (N_10832,N_10585,N_10634);
nand U10833 (N_10833,N_10722,N_10650);
xnor U10834 (N_10834,N_10534,N_10569);
xor U10835 (N_10835,N_10586,N_10625);
nor U10836 (N_10836,N_10645,N_10716);
xor U10837 (N_10837,N_10660,N_10617);
nor U10838 (N_10838,N_10607,N_10654);
nor U10839 (N_10839,N_10604,N_10652);
or U10840 (N_10840,N_10557,N_10698);
and U10841 (N_10841,N_10512,N_10549);
nor U10842 (N_10842,N_10526,N_10509);
xor U10843 (N_10843,N_10733,N_10720);
xor U10844 (N_10844,N_10554,N_10678);
nor U10845 (N_10845,N_10555,N_10691);
or U10846 (N_10846,N_10695,N_10508);
xor U10847 (N_10847,N_10558,N_10624);
xnor U10848 (N_10848,N_10725,N_10598);
nand U10849 (N_10849,N_10507,N_10749);
nand U10850 (N_10850,N_10593,N_10603);
nand U10851 (N_10851,N_10594,N_10537);
xor U10852 (N_10852,N_10689,N_10699);
xnor U10853 (N_10853,N_10505,N_10703);
xnor U10854 (N_10854,N_10623,N_10653);
and U10855 (N_10855,N_10528,N_10525);
nand U10856 (N_10856,N_10506,N_10580);
or U10857 (N_10857,N_10667,N_10551);
nor U10858 (N_10858,N_10608,N_10542);
or U10859 (N_10859,N_10533,N_10642);
xnor U10860 (N_10860,N_10559,N_10540);
and U10861 (N_10861,N_10746,N_10636);
and U10862 (N_10862,N_10724,N_10707);
and U10863 (N_10863,N_10503,N_10731);
nor U10864 (N_10864,N_10611,N_10618);
and U10865 (N_10865,N_10504,N_10516);
nand U10866 (N_10866,N_10565,N_10677);
nor U10867 (N_10867,N_10536,N_10744);
or U10868 (N_10868,N_10656,N_10647);
and U10869 (N_10869,N_10601,N_10673);
and U10870 (N_10870,N_10688,N_10612);
and U10871 (N_10871,N_10714,N_10684);
nor U10872 (N_10872,N_10741,N_10711);
nand U10873 (N_10873,N_10574,N_10726);
nand U10874 (N_10874,N_10712,N_10573);
and U10875 (N_10875,N_10655,N_10581);
xnor U10876 (N_10876,N_10622,N_10652);
xnor U10877 (N_10877,N_10689,N_10598);
nor U10878 (N_10878,N_10658,N_10695);
or U10879 (N_10879,N_10589,N_10563);
xnor U10880 (N_10880,N_10541,N_10506);
nand U10881 (N_10881,N_10707,N_10668);
nor U10882 (N_10882,N_10570,N_10510);
or U10883 (N_10883,N_10598,N_10526);
xnor U10884 (N_10884,N_10739,N_10738);
and U10885 (N_10885,N_10748,N_10583);
or U10886 (N_10886,N_10742,N_10623);
nand U10887 (N_10887,N_10606,N_10559);
and U10888 (N_10888,N_10679,N_10656);
xor U10889 (N_10889,N_10548,N_10568);
nor U10890 (N_10890,N_10601,N_10506);
or U10891 (N_10891,N_10723,N_10521);
or U10892 (N_10892,N_10617,N_10719);
nor U10893 (N_10893,N_10657,N_10737);
nand U10894 (N_10894,N_10691,N_10507);
xor U10895 (N_10895,N_10641,N_10602);
and U10896 (N_10896,N_10534,N_10525);
xor U10897 (N_10897,N_10604,N_10640);
and U10898 (N_10898,N_10618,N_10605);
nor U10899 (N_10899,N_10701,N_10741);
xnor U10900 (N_10900,N_10521,N_10621);
xor U10901 (N_10901,N_10546,N_10605);
nor U10902 (N_10902,N_10698,N_10541);
xor U10903 (N_10903,N_10608,N_10509);
and U10904 (N_10904,N_10734,N_10593);
xor U10905 (N_10905,N_10657,N_10679);
xnor U10906 (N_10906,N_10714,N_10632);
nand U10907 (N_10907,N_10557,N_10631);
or U10908 (N_10908,N_10627,N_10711);
nor U10909 (N_10909,N_10684,N_10620);
nand U10910 (N_10910,N_10746,N_10634);
xnor U10911 (N_10911,N_10551,N_10627);
or U10912 (N_10912,N_10582,N_10557);
xnor U10913 (N_10913,N_10597,N_10633);
and U10914 (N_10914,N_10582,N_10507);
or U10915 (N_10915,N_10583,N_10612);
nand U10916 (N_10916,N_10534,N_10602);
or U10917 (N_10917,N_10693,N_10678);
or U10918 (N_10918,N_10721,N_10681);
or U10919 (N_10919,N_10569,N_10536);
xor U10920 (N_10920,N_10574,N_10565);
or U10921 (N_10921,N_10625,N_10636);
or U10922 (N_10922,N_10536,N_10595);
nand U10923 (N_10923,N_10582,N_10545);
xnor U10924 (N_10924,N_10506,N_10632);
nand U10925 (N_10925,N_10741,N_10588);
nand U10926 (N_10926,N_10725,N_10729);
nor U10927 (N_10927,N_10617,N_10609);
xnor U10928 (N_10928,N_10526,N_10643);
nor U10929 (N_10929,N_10722,N_10615);
xor U10930 (N_10930,N_10674,N_10503);
nand U10931 (N_10931,N_10671,N_10635);
or U10932 (N_10932,N_10714,N_10642);
and U10933 (N_10933,N_10558,N_10525);
nand U10934 (N_10934,N_10558,N_10662);
or U10935 (N_10935,N_10505,N_10641);
nor U10936 (N_10936,N_10500,N_10727);
xor U10937 (N_10937,N_10718,N_10670);
and U10938 (N_10938,N_10608,N_10586);
nor U10939 (N_10939,N_10653,N_10723);
nor U10940 (N_10940,N_10526,N_10685);
nand U10941 (N_10941,N_10566,N_10678);
nand U10942 (N_10942,N_10560,N_10691);
or U10943 (N_10943,N_10715,N_10732);
nor U10944 (N_10944,N_10535,N_10553);
or U10945 (N_10945,N_10525,N_10586);
nor U10946 (N_10946,N_10707,N_10691);
or U10947 (N_10947,N_10695,N_10669);
xnor U10948 (N_10948,N_10573,N_10652);
nand U10949 (N_10949,N_10699,N_10623);
and U10950 (N_10950,N_10729,N_10695);
xor U10951 (N_10951,N_10575,N_10520);
xnor U10952 (N_10952,N_10683,N_10639);
xnor U10953 (N_10953,N_10646,N_10625);
or U10954 (N_10954,N_10670,N_10612);
or U10955 (N_10955,N_10596,N_10696);
nor U10956 (N_10956,N_10531,N_10628);
or U10957 (N_10957,N_10618,N_10519);
and U10958 (N_10958,N_10517,N_10647);
xnor U10959 (N_10959,N_10558,N_10649);
nand U10960 (N_10960,N_10569,N_10682);
xor U10961 (N_10961,N_10710,N_10695);
and U10962 (N_10962,N_10736,N_10598);
nor U10963 (N_10963,N_10695,N_10666);
nor U10964 (N_10964,N_10646,N_10577);
and U10965 (N_10965,N_10561,N_10632);
nor U10966 (N_10966,N_10579,N_10558);
nor U10967 (N_10967,N_10701,N_10677);
nand U10968 (N_10968,N_10664,N_10616);
xor U10969 (N_10969,N_10707,N_10713);
and U10970 (N_10970,N_10573,N_10738);
nand U10971 (N_10971,N_10707,N_10591);
and U10972 (N_10972,N_10597,N_10680);
nor U10973 (N_10973,N_10554,N_10556);
nor U10974 (N_10974,N_10691,N_10548);
xor U10975 (N_10975,N_10634,N_10609);
and U10976 (N_10976,N_10727,N_10529);
or U10977 (N_10977,N_10641,N_10545);
nand U10978 (N_10978,N_10526,N_10620);
nand U10979 (N_10979,N_10555,N_10720);
nand U10980 (N_10980,N_10584,N_10619);
nor U10981 (N_10981,N_10706,N_10672);
and U10982 (N_10982,N_10506,N_10739);
and U10983 (N_10983,N_10500,N_10572);
and U10984 (N_10984,N_10716,N_10524);
nand U10985 (N_10985,N_10608,N_10697);
nand U10986 (N_10986,N_10738,N_10569);
nor U10987 (N_10987,N_10544,N_10655);
or U10988 (N_10988,N_10721,N_10701);
or U10989 (N_10989,N_10584,N_10541);
nand U10990 (N_10990,N_10722,N_10543);
and U10991 (N_10991,N_10729,N_10582);
nor U10992 (N_10992,N_10597,N_10523);
xor U10993 (N_10993,N_10748,N_10668);
nor U10994 (N_10994,N_10576,N_10671);
or U10995 (N_10995,N_10554,N_10576);
nor U10996 (N_10996,N_10726,N_10666);
xnor U10997 (N_10997,N_10501,N_10636);
nor U10998 (N_10998,N_10677,N_10516);
or U10999 (N_10999,N_10663,N_10535);
nand U11000 (N_11000,N_10864,N_10997);
and U11001 (N_11001,N_10959,N_10951);
xor U11002 (N_11002,N_10834,N_10767);
and U11003 (N_11003,N_10833,N_10880);
nor U11004 (N_11004,N_10875,N_10946);
and U11005 (N_11005,N_10927,N_10799);
nor U11006 (N_11006,N_10846,N_10999);
nor U11007 (N_11007,N_10934,N_10964);
nand U11008 (N_11008,N_10801,N_10994);
and U11009 (N_11009,N_10942,N_10992);
xnor U11010 (N_11010,N_10973,N_10769);
and U11011 (N_11011,N_10970,N_10904);
or U11012 (N_11012,N_10775,N_10868);
nor U11013 (N_11013,N_10911,N_10975);
nand U11014 (N_11014,N_10863,N_10930);
and U11015 (N_11015,N_10874,N_10764);
nor U11016 (N_11016,N_10807,N_10836);
nand U11017 (N_11017,N_10832,N_10779);
or U11018 (N_11018,N_10956,N_10826);
xnor U11019 (N_11019,N_10884,N_10870);
xnor U11020 (N_11020,N_10815,N_10757);
nand U11021 (N_11021,N_10952,N_10941);
or U11022 (N_11022,N_10995,N_10782);
or U11023 (N_11023,N_10899,N_10928);
nor U11024 (N_11024,N_10900,N_10982);
and U11025 (N_11025,N_10953,N_10990);
nand U11026 (N_11026,N_10753,N_10981);
xnor U11027 (N_11027,N_10831,N_10871);
and U11028 (N_11028,N_10802,N_10845);
nor U11029 (N_11029,N_10985,N_10803);
and U11030 (N_11030,N_10897,N_10931);
nor U11031 (N_11031,N_10867,N_10783);
xnor U11032 (N_11032,N_10784,N_10908);
nor U11033 (N_11033,N_10816,N_10776);
and U11034 (N_11034,N_10772,N_10835);
xnor U11035 (N_11035,N_10854,N_10910);
nand U11036 (N_11036,N_10977,N_10983);
or U11037 (N_11037,N_10881,N_10932);
and U11038 (N_11038,N_10991,N_10887);
nor U11039 (N_11039,N_10998,N_10967);
nand U11040 (N_11040,N_10786,N_10762);
and U11041 (N_11041,N_10770,N_10976);
xor U11042 (N_11042,N_10936,N_10787);
nor U11043 (N_11043,N_10929,N_10894);
nor U11044 (N_11044,N_10751,N_10958);
nand U11045 (N_11045,N_10890,N_10792);
xor U11046 (N_11046,N_10750,N_10918);
or U11047 (N_11047,N_10872,N_10765);
nand U11048 (N_11048,N_10912,N_10771);
nor U11049 (N_11049,N_10780,N_10889);
xnor U11050 (N_11050,N_10778,N_10773);
nand U11051 (N_11051,N_10923,N_10922);
and U11052 (N_11052,N_10789,N_10858);
nor U11053 (N_11053,N_10980,N_10841);
or U11054 (N_11054,N_10913,N_10901);
or U11055 (N_11055,N_10837,N_10969);
nor U11056 (N_11056,N_10804,N_10903);
or U11057 (N_11057,N_10921,N_10896);
and U11058 (N_11058,N_10905,N_10791);
nand U11059 (N_11059,N_10949,N_10862);
nor U11060 (N_11060,N_10938,N_10813);
nor U11061 (N_11061,N_10948,N_10971);
xnor U11062 (N_11062,N_10883,N_10935);
and U11063 (N_11063,N_10754,N_10796);
nor U11064 (N_11064,N_10962,N_10760);
or U11065 (N_11065,N_10957,N_10756);
xor U11066 (N_11066,N_10893,N_10853);
xnor U11067 (N_11067,N_10926,N_10752);
nor U11068 (N_11068,N_10916,N_10869);
xnor U11069 (N_11069,N_10861,N_10924);
xor U11070 (N_11070,N_10989,N_10965);
and U11071 (N_11071,N_10808,N_10960);
or U11072 (N_11072,N_10920,N_10848);
and U11073 (N_11073,N_10843,N_10943);
xnor U11074 (N_11074,N_10827,N_10895);
nor U11075 (N_11075,N_10891,N_10825);
nor U11076 (N_11076,N_10915,N_10909);
nand U11077 (N_11077,N_10755,N_10996);
nor U11078 (N_11078,N_10842,N_10954);
nand U11079 (N_11079,N_10945,N_10968);
xor U11080 (N_11080,N_10947,N_10800);
and U11081 (N_11081,N_10849,N_10774);
nor U11082 (N_11082,N_10852,N_10993);
xnor U11083 (N_11083,N_10972,N_10902);
or U11084 (N_11084,N_10763,N_10781);
nand U11085 (N_11085,N_10919,N_10797);
and U11086 (N_11086,N_10823,N_10876);
xor U11087 (N_11087,N_10820,N_10859);
and U11088 (N_11088,N_10839,N_10788);
and U11089 (N_11089,N_10814,N_10933);
or U11090 (N_11090,N_10855,N_10822);
nor U11091 (N_11091,N_10877,N_10955);
and U11092 (N_11092,N_10811,N_10925);
xor U11093 (N_11093,N_10950,N_10795);
nand U11094 (N_11094,N_10939,N_10873);
nand U11095 (N_11095,N_10898,N_10847);
xor U11096 (N_11096,N_10865,N_10860);
nor U11097 (N_11097,N_10790,N_10857);
or U11098 (N_11098,N_10963,N_10809);
or U11099 (N_11099,N_10761,N_10892);
or U11100 (N_11100,N_10866,N_10819);
nor U11101 (N_11101,N_10829,N_10777);
nand U11102 (N_11102,N_10879,N_10850);
xnor U11103 (N_11103,N_10907,N_10830);
or U11104 (N_11104,N_10914,N_10785);
and U11105 (N_11105,N_10979,N_10917);
or U11106 (N_11106,N_10974,N_10768);
and U11107 (N_11107,N_10844,N_10885);
nor U11108 (N_11108,N_10987,N_10759);
nor U11109 (N_11109,N_10888,N_10986);
nand U11110 (N_11110,N_10851,N_10810);
nor U11111 (N_11111,N_10961,N_10882);
xnor U11112 (N_11112,N_10984,N_10794);
nand U11113 (N_11113,N_10824,N_10812);
nor U11114 (N_11114,N_10856,N_10793);
xor U11115 (N_11115,N_10940,N_10878);
nand U11116 (N_11116,N_10838,N_10937);
nand U11117 (N_11117,N_10821,N_10906);
nor U11118 (N_11118,N_10818,N_10966);
xor U11119 (N_11119,N_10805,N_10988);
nor U11120 (N_11120,N_10840,N_10944);
and U11121 (N_11121,N_10886,N_10798);
xor U11122 (N_11122,N_10978,N_10806);
xor U11123 (N_11123,N_10758,N_10817);
xor U11124 (N_11124,N_10828,N_10766);
nor U11125 (N_11125,N_10865,N_10840);
nand U11126 (N_11126,N_10813,N_10941);
nor U11127 (N_11127,N_10788,N_10854);
nor U11128 (N_11128,N_10780,N_10930);
and U11129 (N_11129,N_10842,N_10765);
or U11130 (N_11130,N_10947,N_10924);
xnor U11131 (N_11131,N_10951,N_10863);
or U11132 (N_11132,N_10750,N_10776);
xnor U11133 (N_11133,N_10852,N_10914);
nand U11134 (N_11134,N_10946,N_10994);
or U11135 (N_11135,N_10841,N_10826);
and U11136 (N_11136,N_10977,N_10905);
or U11137 (N_11137,N_10772,N_10938);
or U11138 (N_11138,N_10982,N_10794);
or U11139 (N_11139,N_10828,N_10936);
and U11140 (N_11140,N_10957,N_10789);
nand U11141 (N_11141,N_10787,N_10938);
nand U11142 (N_11142,N_10773,N_10946);
nor U11143 (N_11143,N_10956,N_10936);
nand U11144 (N_11144,N_10846,N_10826);
xor U11145 (N_11145,N_10906,N_10772);
xnor U11146 (N_11146,N_10952,N_10906);
nor U11147 (N_11147,N_10927,N_10776);
nand U11148 (N_11148,N_10852,N_10958);
xnor U11149 (N_11149,N_10825,N_10901);
and U11150 (N_11150,N_10792,N_10899);
or U11151 (N_11151,N_10952,N_10935);
xnor U11152 (N_11152,N_10782,N_10855);
nor U11153 (N_11153,N_10833,N_10831);
or U11154 (N_11154,N_10815,N_10885);
and U11155 (N_11155,N_10861,N_10918);
xor U11156 (N_11156,N_10977,N_10753);
xor U11157 (N_11157,N_10885,N_10857);
nor U11158 (N_11158,N_10961,N_10939);
or U11159 (N_11159,N_10967,N_10819);
xnor U11160 (N_11160,N_10759,N_10850);
xnor U11161 (N_11161,N_10818,N_10795);
nand U11162 (N_11162,N_10901,N_10846);
xor U11163 (N_11163,N_10826,N_10932);
xor U11164 (N_11164,N_10797,N_10827);
nand U11165 (N_11165,N_10968,N_10950);
nor U11166 (N_11166,N_10978,N_10993);
nand U11167 (N_11167,N_10788,N_10885);
and U11168 (N_11168,N_10968,N_10801);
nor U11169 (N_11169,N_10771,N_10999);
xnor U11170 (N_11170,N_10783,N_10997);
nor U11171 (N_11171,N_10975,N_10848);
or U11172 (N_11172,N_10856,N_10902);
nor U11173 (N_11173,N_10781,N_10799);
and U11174 (N_11174,N_10920,N_10927);
nor U11175 (N_11175,N_10907,N_10762);
xnor U11176 (N_11176,N_10953,N_10940);
nor U11177 (N_11177,N_10997,N_10921);
or U11178 (N_11178,N_10932,N_10929);
nor U11179 (N_11179,N_10903,N_10840);
xnor U11180 (N_11180,N_10957,N_10925);
xor U11181 (N_11181,N_10764,N_10843);
nor U11182 (N_11182,N_10877,N_10886);
or U11183 (N_11183,N_10796,N_10772);
and U11184 (N_11184,N_10926,N_10788);
xnor U11185 (N_11185,N_10909,N_10948);
xor U11186 (N_11186,N_10957,N_10859);
and U11187 (N_11187,N_10783,N_10767);
xor U11188 (N_11188,N_10924,N_10978);
nand U11189 (N_11189,N_10875,N_10816);
xnor U11190 (N_11190,N_10986,N_10870);
nor U11191 (N_11191,N_10928,N_10824);
and U11192 (N_11192,N_10757,N_10837);
nor U11193 (N_11193,N_10970,N_10911);
nand U11194 (N_11194,N_10804,N_10915);
nand U11195 (N_11195,N_10787,N_10977);
nand U11196 (N_11196,N_10888,N_10830);
and U11197 (N_11197,N_10939,N_10807);
nand U11198 (N_11198,N_10785,N_10874);
or U11199 (N_11199,N_10896,N_10962);
nand U11200 (N_11200,N_10994,N_10964);
or U11201 (N_11201,N_10800,N_10994);
and U11202 (N_11202,N_10834,N_10881);
or U11203 (N_11203,N_10821,N_10972);
or U11204 (N_11204,N_10872,N_10949);
nor U11205 (N_11205,N_10855,N_10985);
nand U11206 (N_11206,N_10836,N_10928);
and U11207 (N_11207,N_10981,N_10781);
xor U11208 (N_11208,N_10908,N_10879);
nor U11209 (N_11209,N_10869,N_10881);
nand U11210 (N_11210,N_10925,N_10991);
xor U11211 (N_11211,N_10994,N_10871);
or U11212 (N_11212,N_10911,N_10893);
and U11213 (N_11213,N_10785,N_10985);
xnor U11214 (N_11214,N_10939,N_10819);
or U11215 (N_11215,N_10967,N_10791);
or U11216 (N_11216,N_10912,N_10898);
xor U11217 (N_11217,N_10838,N_10783);
nor U11218 (N_11218,N_10926,N_10777);
nand U11219 (N_11219,N_10825,N_10999);
or U11220 (N_11220,N_10872,N_10999);
and U11221 (N_11221,N_10825,N_10763);
nand U11222 (N_11222,N_10752,N_10994);
or U11223 (N_11223,N_10811,N_10906);
or U11224 (N_11224,N_10929,N_10805);
and U11225 (N_11225,N_10910,N_10859);
and U11226 (N_11226,N_10965,N_10912);
xor U11227 (N_11227,N_10822,N_10887);
nor U11228 (N_11228,N_10916,N_10970);
xor U11229 (N_11229,N_10999,N_10996);
or U11230 (N_11230,N_10934,N_10920);
xnor U11231 (N_11231,N_10927,N_10793);
xor U11232 (N_11232,N_10830,N_10948);
xor U11233 (N_11233,N_10933,N_10909);
or U11234 (N_11234,N_10902,N_10913);
or U11235 (N_11235,N_10934,N_10875);
nor U11236 (N_11236,N_10972,N_10998);
or U11237 (N_11237,N_10903,N_10861);
and U11238 (N_11238,N_10810,N_10960);
and U11239 (N_11239,N_10872,N_10893);
xor U11240 (N_11240,N_10900,N_10995);
and U11241 (N_11241,N_10838,N_10919);
xnor U11242 (N_11242,N_10897,N_10895);
nor U11243 (N_11243,N_10851,N_10894);
or U11244 (N_11244,N_10986,N_10928);
nor U11245 (N_11245,N_10915,N_10901);
and U11246 (N_11246,N_10798,N_10991);
nor U11247 (N_11247,N_10967,N_10910);
nand U11248 (N_11248,N_10906,N_10833);
and U11249 (N_11249,N_10930,N_10924);
or U11250 (N_11250,N_11031,N_11204);
and U11251 (N_11251,N_11115,N_11103);
xnor U11252 (N_11252,N_11214,N_11181);
xnor U11253 (N_11253,N_11047,N_11163);
or U11254 (N_11254,N_11043,N_11046);
xor U11255 (N_11255,N_11127,N_11039);
and U11256 (N_11256,N_11035,N_11036);
xor U11257 (N_11257,N_11034,N_11002);
nand U11258 (N_11258,N_11062,N_11219);
or U11259 (N_11259,N_11227,N_11205);
and U11260 (N_11260,N_11107,N_11105);
xnor U11261 (N_11261,N_11144,N_11230);
nand U11262 (N_11262,N_11086,N_11179);
and U11263 (N_11263,N_11173,N_11059);
or U11264 (N_11264,N_11054,N_11048);
and U11265 (N_11265,N_11057,N_11114);
and U11266 (N_11266,N_11042,N_11037);
nor U11267 (N_11267,N_11167,N_11072);
or U11268 (N_11268,N_11212,N_11033);
nor U11269 (N_11269,N_11003,N_11011);
or U11270 (N_11270,N_11170,N_11073);
nand U11271 (N_11271,N_11207,N_11118);
nand U11272 (N_11272,N_11005,N_11156);
xor U11273 (N_11273,N_11010,N_11069);
or U11274 (N_11274,N_11040,N_11116);
or U11275 (N_11275,N_11178,N_11218);
xor U11276 (N_11276,N_11094,N_11247);
or U11277 (N_11277,N_11134,N_11159);
and U11278 (N_11278,N_11143,N_11229);
nor U11279 (N_11279,N_11238,N_11097);
or U11280 (N_11280,N_11199,N_11180);
nand U11281 (N_11281,N_11175,N_11133);
or U11282 (N_11282,N_11130,N_11157);
nand U11283 (N_11283,N_11213,N_11067);
xor U11284 (N_11284,N_11209,N_11102);
nand U11285 (N_11285,N_11095,N_11222);
xor U11286 (N_11286,N_11112,N_11078);
nand U11287 (N_11287,N_11138,N_11171);
and U11288 (N_11288,N_11136,N_11210);
or U11289 (N_11289,N_11142,N_11166);
xnor U11290 (N_11290,N_11197,N_11091);
nor U11291 (N_11291,N_11109,N_11004);
nand U11292 (N_11292,N_11188,N_11125);
nand U11293 (N_11293,N_11221,N_11060);
nor U11294 (N_11294,N_11027,N_11141);
or U11295 (N_11295,N_11187,N_11017);
and U11296 (N_11296,N_11122,N_11055);
nand U11297 (N_11297,N_11101,N_11201);
nand U11298 (N_11298,N_11018,N_11110);
xor U11299 (N_11299,N_11019,N_11202);
nand U11300 (N_11300,N_11131,N_11032);
and U11301 (N_11301,N_11126,N_11085);
xor U11302 (N_11302,N_11020,N_11198);
nand U11303 (N_11303,N_11243,N_11029);
or U11304 (N_11304,N_11172,N_11082);
xnor U11305 (N_11305,N_11071,N_11211);
and U11306 (N_11306,N_11161,N_11015);
xor U11307 (N_11307,N_11242,N_11239);
xnor U11308 (N_11308,N_11012,N_11000);
nand U11309 (N_11309,N_11006,N_11160);
xnor U11310 (N_11310,N_11149,N_11226);
and U11311 (N_11311,N_11026,N_11132);
and U11312 (N_11312,N_11164,N_11056);
nor U11313 (N_11313,N_11120,N_11215);
nor U11314 (N_11314,N_11025,N_11185);
and U11315 (N_11315,N_11203,N_11089);
or U11316 (N_11316,N_11236,N_11129);
nand U11317 (N_11317,N_11088,N_11066);
nand U11318 (N_11318,N_11053,N_11087);
nor U11319 (N_11319,N_11194,N_11246);
nand U11320 (N_11320,N_11140,N_11068);
xnor U11321 (N_11321,N_11177,N_11190);
and U11322 (N_11322,N_11145,N_11220);
nand U11323 (N_11323,N_11135,N_11223);
and U11324 (N_11324,N_11007,N_11021);
xor U11325 (N_11325,N_11045,N_11041);
and U11326 (N_11326,N_11113,N_11061);
or U11327 (N_11327,N_11234,N_11154);
and U11328 (N_11328,N_11150,N_11165);
nand U11329 (N_11329,N_11058,N_11249);
nand U11330 (N_11330,N_11158,N_11146);
nor U11331 (N_11331,N_11030,N_11099);
xnor U11332 (N_11332,N_11092,N_11241);
nor U11333 (N_11333,N_11208,N_11080);
or U11334 (N_11334,N_11162,N_11193);
nand U11335 (N_11335,N_11051,N_11106);
nor U11336 (N_11336,N_11075,N_11216);
nand U11337 (N_11337,N_11152,N_11237);
or U11338 (N_11338,N_11076,N_11148);
xor U11339 (N_11339,N_11083,N_11153);
and U11340 (N_11340,N_11038,N_11128);
xnor U11341 (N_11341,N_11217,N_11123);
and U11342 (N_11342,N_11151,N_11195);
xnor U11343 (N_11343,N_11024,N_11233);
xnor U11344 (N_11344,N_11155,N_11119);
or U11345 (N_11345,N_11196,N_11182);
nand U11346 (N_11346,N_11189,N_11248);
and U11347 (N_11347,N_11064,N_11001);
nor U11348 (N_11348,N_11014,N_11232);
nand U11349 (N_11349,N_11023,N_11231);
nand U11350 (N_11350,N_11235,N_11184);
and U11351 (N_11351,N_11065,N_11147);
and U11352 (N_11352,N_11050,N_11174);
or U11353 (N_11353,N_11240,N_11108);
nand U11354 (N_11354,N_11186,N_11100);
nand U11355 (N_11355,N_11224,N_11009);
or U11356 (N_11356,N_11139,N_11191);
or U11357 (N_11357,N_11016,N_11070);
nor U11358 (N_11358,N_11063,N_11090);
or U11359 (N_11359,N_11096,N_11200);
nor U11360 (N_11360,N_11124,N_11052);
nand U11361 (N_11361,N_11013,N_11206);
or U11362 (N_11362,N_11044,N_11245);
and U11363 (N_11363,N_11104,N_11228);
nor U11364 (N_11364,N_11225,N_11168);
or U11365 (N_11365,N_11049,N_11183);
nor U11366 (N_11366,N_11022,N_11192);
or U11367 (N_11367,N_11111,N_11074);
nor U11368 (N_11368,N_11084,N_11008);
or U11369 (N_11369,N_11244,N_11117);
xor U11370 (N_11370,N_11093,N_11081);
xnor U11371 (N_11371,N_11028,N_11077);
or U11372 (N_11372,N_11079,N_11169);
nor U11373 (N_11373,N_11098,N_11121);
xor U11374 (N_11374,N_11176,N_11137);
and U11375 (N_11375,N_11089,N_11163);
or U11376 (N_11376,N_11100,N_11143);
nor U11377 (N_11377,N_11177,N_11231);
or U11378 (N_11378,N_11117,N_11056);
and U11379 (N_11379,N_11218,N_11119);
and U11380 (N_11380,N_11192,N_11150);
xnor U11381 (N_11381,N_11009,N_11187);
nand U11382 (N_11382,N_11014,N_11233);
and U11383 (N_11383,N_11045,N_11035);
xor U11384 (N_11384,N_11034,N_11122);
and U11385 (N_11385,N_11118,N_11163);
xor U11386 (N_11386,N_11177,N_11034);
or U11387 (N_11387,N_11230,N_11161);
xor U11388 (N_11388,N_11148,N_11061);
and U11389 (N_11389,N_11001,N_11078);
xnor U11390 (N_11390,N_11177,N_11054);
xnor U11391 (N_11391,N_11146,N_11163);
nor U11392 (N_11392,N_11084,N_11156);
xor U11393 (N_11393,N_11001,N_11034);
and U11394 (N_11394,N_11071,N_11145);
and U11395 (N_11395,N_11207,N_11007);
nand U11396 (N_11396,N_11140,N_11058);
or U11397 (N_11397,N_11247,N_11149);
nand U11398 (N_11398,N_11161,N_11114);
and U11399 (N_11399,N_11117,N_11079);
and U11400 (N_11400,N_11216,N_11245);
nor U11401 (N_11401,N_11148,N_11002);
or U11402 (N_11402,N_11246,N_11071);
xor U11403 (N_11403,N_11054,N_11058);
and U11404 (N_11404,N_11048,N_11146);
nor U11405 (N_11405,N_11239,N_11174);
and U11406 (N_11406,N_11074,N_11045);
nand U11407 (N_11407,N_11153,N_11032);
xnor U11408 (N_11408,N_11211,N_11086);
or U11409 (N_11409,N_11145,N_11002);
xnor U11410 (N_11410,N_11014,N_11194);
and U11411 (N_11411,N_11207,N_11159);
xnor U11412 (N_11412,N_11005,N_11240);
nand U11413 (N_11413,N_11229,N_11209);
xor U11414 (N_11414,N_11103,N_11062);
and U11415 (N_11415,N_11042,N_11145);
xnor U11416 (N_11416,N_11018,N_11118);
nand U11417 (N_11417,N_11248,N_11097);
nor U11418 (N_11418,N_11221,N_11037);
xor U11419 (N_11419,N_11117,N_11071);
nand U11420 (N_11420,N_11213,N_11162);
nand U11421 (N_11421,N_11187,N_11240);
and U11422 (N_11422,N_11025,N_11222);
or U11423 (N_11423,N_11150,N_11139);
xor U11424 (N_11424,N_11234,N_11245);
or U11425 (N_11425,N_11156,N_11225);
xor U11426 (N_11426,N_11200,N_11135);
and U11427 (N_11427,N_11136,N_11242);
and U11428 (N_11428,N_11198,N_11005);
nor U11429 (N_11429,N_11016,N_11085);
nand U11430 (N_11430,N_11009,N_11248);
and U11431 (N_11431,N_11043,N_11193);
or U11432 (N_11432,N_11185,N_11182);
nor U11433 (N_11433,N_11084,N_11113);
nor U11434 (N_11434,N_11141,N_11249);
nand U11435 (N_11435,N_11023,N_11192);
or U11436 (N_11436,N_11008,N_11171);
nand U11437 (N_11437,N_11071,N_11079);
and U11438 (N_11438,N_11024,N_11030);
or U11439 (N_11439,N_11217,N_11132);
and U11440 (N_11440,N_11096,N_11103);
or U11441 (N_11441,N_11170,N_11024);
xnor U11442 (N_11442,N_11054,N_11204);
or U11443 (N_11443,N_11168,N_11244);
xnor U11444 (N_11444,N_11231,N_11159);
or U11445 (N_11445,N_11245,N_11219);
or U11446 (N_11446,N_11081,N_11064);
nor U11447 (N_11447,N_11236,N_11014);
nand U11448 (N_11448,N_11173,N_11092);
nor U11449 (N_11449,N_11110,N_11049);
nor U11450 (N_11450,N_11123,N_11130);
and U11451 (N_11451,N_11248,N_11191);
xor U11452 (N_11452,N_11199,N_11225);
nor U11453 (N_11453,N_11029,N_11156);
nor U11454 (N_11454,N_11174,N_11079);
xor U11455 (N_11455,N_11228,N_11244);
or U11456 (N_11456,N_11188,N_11078);
nand U11457 (N_11457,N_11188,N_11072);
or U11458 (N_11458,N_11156,N_11210);
xnor U11459 (N_11459,N_11213,N_11072);
nor U11460 (N_11460,N_11044,N_11125);
nand U11461 (N_11461,N_11064,N_11169);
and U11462 (N_11462,N_11121,N_11027);
nor U11463 (N_11463,N_11244,N_11150);
or U11464 (N_11464,N_11000,N_11183);
nor U11465 (N_11465,N_11019,N_11013);
or U11466 (N_11466,N_11223,N_11195);
nand U11467 (N_11467,N_11066,N_11156);
and U11468 (N_11468,N_11053,N_11029);
nor U11469 (N_11469,N_11215,N_11003);
nand U11470 (N_11470,N_11243,N_11139);
nor U11471 (N_11471,N_11169,N_11060);
nand U11472 (N_11472,N_11145,N_11119);
or U11473 (N_11473,N_11086,N_11133);
nor U11474 (N_11474,N_11172,N_11131);
xor U11475 (N_11475,N_11138,N_11195);
nor U11476 (N_11476,N_11114,N_11059);
xnor U11477 (N_11477,N_11169,N_11222);
nor U11478 (N_11478,N_11049,N_11046);
nand U11479 (N_11479,N_11129,N_11227);
nor U11480 (N_11480,N_11036,N_11103);
or U11481 (N_11481,N_11240,N_11055);
nor U11482 (N_11482,N_11140,N_11014);
nand U11483 (N_11483,N_11220,N_11041);
nand U11484 (N_11484,N_11229,N_11072);
nand U11485 (N_11485,N_11094,N_11142);
or U11486 (N_11486,N_11118,N_11129);
or U11487 (N_11487,N_11041,N_11193);
nor U11488 (N_11488,N_11177,N_11056);
or U11489 (N_11489,N_11023,N_11193);
xnor U11490 (N_11490,N_11064,N_11062);
xnor U11491 (N_11491,N_11062,N_11138);
nor U11492 (N_11492,N_11032,N_11157);
and U11493 (N_11493,N_11052,N_11101);
or U11494 (N_11494,N_11062,N_11020);
or U11495 (N_11495,N_11109,N_11043);
xnor U11496 (N_11496,N_11000,N_11153);
nand U11497 (N_11497,N_11161,N_11094);
or U11498 (N_11498,N_11073,N_11121);
and U11499 (N_11499,N_11037,N_11046);
nor U11500 (N_11500,N_11323,N_11321);
nor U11501 (N_11501,N_11422,N_11478);
or U11502 (N_11502,N_11455,N_11493);
and U11503 (N_11503,N_11452,N_11479);
and U11504 (N_11504,N_11324,N_11477);
nand U11505 (N_11505,N_11473,N_11379);
or U11506 (N_11506,N_11263,N_11398);
or U11507 (N_11507,N_11347,N_11318);
nand U11508 (N_11508,N_11485,N_11410);
nor U11509 (N_11509,N_11377,N_11295);
nor U11510 (N_11510,N_11349,N_11360);
and U11511 (N_11511,N_11399,N_11285);
xor U11512 (N_11512,N_11405,N_11425);
nand U11513 (N_11513,N_11258,N_11339);
xnor U11514 (N_11514,N_11395,N_11294);
xor U11515 (N_11515,N_11494,N_11465);
or U11516 (N_11516,N_11299,N_11463);
and U11517 (N_11517,N_11256,N_11322);
xor U11518 (N_11518,N_11257,N_11404);
nor U11519 (N_11519,N_11328,N_11315);
xor U11520 (N_11520,N_11301,N_11305);
and U11521 (N_11521,N_11302,N_11427);
and U11522 (N_11522,N_11312,N_11391);
and U11523 (N_11523,N_11464,N_11453);
xnor U11524 (N_11524,N_11412,N_11325);
or U11525 (N_11525,N_11401,N_11262);
nand U11526 (N_11526,N_11260,N_11409);
or U11527 (N_11527,N_11486,N_11259);
nand U11528 (N_11528,N_11434,N_11298);
or U11529 (N_11529,N_11431,N_11397);
or U11530 (N_11530,N_11288,N_11439);
xnor U11531 (N_11531,N_11444,N_11253);
nor U11532 (N_11532,N_11419,N_11363);
and U11533 (N_11533,N_11413,N_11394);
nor U11534 (N_11534,N_11320,N_11313);
xnor U11535 (N_11535,N_11447,N_11343);
or U11536 (N_11536,N_11255,N_11383);
and U11537 (N_11537,N_11375,N_11384);
nor U11538 (N_11538,N_11454,N_11458);
xnor U11539 (N_11539,N_11346,N_11378);
nand U11540 (N_11540,N_11462,N_11286);
nor U11541 (N_11541,N_11406,N_11438);
or U11542 (N_11542,N_11317,N_11496);
or U11543 (N_11543,N_11270,N_11371);
and U11544 (N_11544,N_11393,N_11332);
nor U11545 (N_11545,N_11426,N_11304);
nand U11546 (N_11546,N_11326,N_11475);
xor U11547 (N_11547,N_11386,N_11306);
nand U11548 (N_11548,N_11316,N_11442);
nor U11549 (N_11549,N_11250,N_11390);
nand U11550 (N_11550,N_11293,N_11277);
xor U11551 (N_11551,N_11381,N_11373);
or U11552 (N_11552,N_11296,N_11376);
xor U11553 (N_11553,N_11490,N_11411);
xnor U11554 (N_11554,N_11300,N_11388);
or U11555 (N_11555,N_11267,N_11430);
nor U11556 (N_11556,N_11408,N_11433);
and U11557 (N_11557,N_11344,N_11336);
nor U11558 (N_11558,N_11290,N_11443);
xnor U11559 (N_11559,N_11483,N_11348);
and U11560 (N_11560,N_11457,N_11366);
xnor U11561 (N_11561,N_11415,N_11416);
or U11562 (N_11562,N_11351,N_11310);
xnor U11563 (N_11563,N_11273,N_11382);
and U11564 (N_11564,N_11329,N_11327);
and U11565 (N_11565,N_11499,N_11340);
and U11566 (N_11566,N_11470,N_11265);
or U11567 (N_11567,N_11414,N_11400);
nand U11568 (N_11568,N_11402,N_11441);
or U11569 (N_11569,N_11283,N_11380);
or U11570 (N_11570,N_11354,N_11303);
xor U11571 (N_11571,N_11274,N_11264);
and U11572 (N_11572,N_11392,N_11484);
nand U11573 (N_11573,N_11334,N_11284);
xnor U11574 (N_11574,N_11374,N_11424);
and U11575 (N_11575,N_11418,N_11492);
xnor U11576 (N_11576,N_11331,N_11387);
xnor U11577 (N_11577,N_11271,N_11450);
or U11578 (N_11578,N_11461,N_11309);
nand U11579 (N_11579,N_11367,N_11417);
or U11580 (N_11580,N_11252,N_11289);
or U11581 (N_11581,N_11440,N_11342);
nor U11582 (N_11582,N_11498,N_11488);
nand U11583 (N_11583,N_11369,N_11368);
nand U11584 (N_11584,N_11269,N_11272);
or U11585 (N_11585,N_11308,N_11278);
nor U11586 (N_11586,N_11389,N_11370);
nand U11587 (N_11587,N_11468,N_11338);
and U11588 (N_11588,N_11497,N_11420);
xor U11589 (N_11589,N_11495,N_11423);
xor U11590 (N_11590,N_11362,N_11385);
xor U11591 (N_11591,N_11435,N_11482);
and U11592 (N_11592,N_11432,N_11449);
and U11593 (N_11593,N_11357,N_11345);
and U11594 (N_11594,N_11279,N_11451);
nor U11595 (N_11595,N_11335,N_11407);
and U11596 (N_11596,N_11469,N_11352);
or U11597 (N_11597,N_11436,N_11281);
xor U11598 (N_11598,N_11311,N_11314);
and U11599 (N_11599,N_11456,N_11421);
nand U11600 (N_11600,N_11429,N_11489);
nor U11601 (N_11601,N_11356,N_11372);
nand U11602 (N_11602,N_11353,N_11291);
nand U11603 (N_11603,N_11282,N_11476);
and U11604 (N_11604,N_11365,N_11459);
nor U11605 (N_11605,N_11359,N_11471);
and U11606 (N_11606,N_11330,N_11337);
and U11607 (N_11607,N_11251,N_11446);
and U11608 (N_11608,N_11261,N_11355);
nor U11609 (N_11609,N_11297,N_11254);
and U11610 (N_11610,N_11276,N_11466);
xnor U11611 (N_11611,N_11467,N_11364);
or U11612 (N_11612,N_11307,N_11445);
nor U11613 (N_11613,N_11472,N_11319);
xor U11614 (N_11614,N_11358,N_11287);
and U11615 (N_11615,N_11481,N_11292);
or U11616 (N_11616,N_11275,N_11480);
nand U11617 (N_11617,N_11460,N_11428);
and U11618 (N_11618,N_11266,N_11474);
and U11619 (N_11619,N_11268,N_11333);
xor U11620 (N_11620,N_11491,N_11350);
xnor U11621 (N_11621,N_11403,N_11280);
xor U11622 (N_11622,N_11487,N_11437);
and U11623 (N_11623,N_11361,N_11396);
nand U11624 (N_11624,N_11448,N_11341);
nor U11625 (N_11625,N_11491,N_11441);
or U11626 (N_11626,N_11450,N_11488);
nand U11627 (N_11627,N_11479,N_11383);
and U11628 (N_11628,N_11435,N_11328);
xnor U11629 (N_11629,N_11462,N_11452);
and U11630 (N_11630,N_11337,N_11452);
nand U11631 (N_11631,N_11451,N_11382);
nor U11632 (N_11632,N_11424,N_11342);
nand U11633 (N_11633,N_11394,N_11469);
nand U11634 (N_11634,N_11343,N_11498);
or U11635 (N_11635,N_11269,N_11453);
xor U11636 (N_11636,N_11375,N_11443);
nor U11637 (N_11637,N_11391,N_11478);
or U11638 (N_11638,N_11408,N_11412);
nor U11639 (N_11639,N_11445,N_11368);
nor U11640 (N_11640,N_11309,N_11433);
and U11641 (N_11641,N_11467,N_11386);
nor U11642 (N_11642,N_11480,N_11259);
xor U11643 (N_11643,N_11351,N_11380);
xnor U11644 (N_11644,N_11405,N_11422);
nand U11645 (N_11645,N_11461,N_11429);
or U11646 (N_11646,N_11339,N_11352);
and U11647 (N_11647,N_11370,N_11299);
nand U11648 (N_11648,N_11412,N_11405);
or U11649 (N_11649,N_11321,N_11263);
xor U11650 (N_11650,N_11457,N_11310);
xnor U11651 (N_11651,N_11429,N_11446);
nand U11652 (N_11652,N_11292,N_11441);
and U11653 (N_11653,N_11411,N_11267);
or U11654 (N_11654,N_11456,N_11358);
and U11655 (N_11655,N_11489,N_11317);
and U11656 (N_11656,N_11365,N_11334);
nor U11657 (N_11657,N_11465,N_11346);
and U11658 (N_11658,N_11417,N_11447);
nand U11659 (N_11659,N_11424,N_11422);
or U11660 (N_11660,N_11322,N_11399);
nand U11661 (N_11661,N_11455,N_11250);
and U11662 (N_11662,N_11327,N_11358);
or U11663 (N_11663,N_11396,N_11474);
or U11664 (N_11664,N_11401,N_11340);
or U11665 (N_11665,N_11433,N_11304);
xor U11666 (N_11666,N_11495,N_11287);
or U11667 (N_11667,N_11471,N_11295);
or U11668 (N_11668,N_11403,N_11376);
xnor U11669 (N_11669,N_11363,N_11438);
or U11670 (N_11670,N_11347,N_11293);
and U11671 (N_11671,N_11475,N_11348);
xor U11672 (N_11672,N_11470,N_11283);
xnor U11673 (N_11673,N_11310,N_11452);
and U11674 (N_11674,N_11473,N_11491);
nand U11675 (N_11675,N_11297,N_11498);
nand U11676 (N_11676,N_11390,N_11352);
xnor U11677 (N_11677,N_11340,N_11489);
nand U11678 (N_11678,N_11363,N_11441);
xnor U11679 (N_11679,N_11389,N_11258);
nand U11680 (N_11680,N_11293,N_11256);
nand U11681 (N_11681,N_11345,N_11463);
nand U11682 (N_11682,N_11321,N_11252);
nor U11683 (N_11683,N_11255,N_11378);
or U11684 (N_11684,N_11287,N_11444);
and U11685 (N_11685,N_11466,N_11315);
nand U11686 (N_11686,N_11250,N_11274);
or U11687 (N_11687,N_11349,N_11286);
and U11688 (N_11688,N_11454,N_11448);
nor U11689 (N_11689,N_11478,N_11273);
or U11690 (N_11690,N_11443,N_11461);
and U11691 (N_11691,N_11442,N_11444);
nand U11692 (N_11692,N_11415,N_11309);
xor U11693 (N_11693,N_11385,N_11276);
and U11694 (N_11694,N_11473,N_11269);
and U11695 (N_11695,N_11375,N_11496);
or U11696 (N_11696,N_11463,N_11411);
xor U11697 (N_11697,N_11324,N_11303);
nor U11698 (N_11698,N_11288,N_11397);
or U11699 (N_11699,N_11393,N_11483);
or U11700 (N_11700,N_11400,N_11256);
nand U11701 (N_11701,N_11384,N_11439);
and U11702 (N_11702,N_11334,N_11256);
or U11703 (N_11703,N_11315,N_11499);
xnor U11704 (N_11704,N_11369,N_11357);
nor U11705 (N_11705,N_11419,N_11454);
or U11706 (N_11706,N_11309,N_11322);
nor U11707 (N_11707,N_11415,N_11458);
nor U11708 (N_11708,N_11314,N_11495);
xor U11709 (N_11709,N_11395,N_11375);
nor U11710 (N_11710,N_11434,N_11344);
or U11711 (N_11711,N_11465,N_11257);
and U11712 (N_11712,N_11288,N_11420);
nor U11713 (N_11713,N_11445,N_11432);
or U11714 (N_11714,N_11329,N_11322);
xor U11715 (N_11715,N_11357,N_11443);
or U11716 (N_11716,N_11264,N_11275);
xnor U11717 (N_11717,N_11272,N_11456);
nor U11718 (N_11718,N_11462,N_11272);
xor U11719 (N_11719,N_11272,N_11476);
or U11720 (N_11720,N_11430,N_11335);
xor U11721 (N_11721,N_11269,N_11404);
and U11722 (N_11722,N_11309,N_11486);
or U11723 (N_11723,N_11291,N_11415);
nand U11724 (N_11724,N_11299,N_11250);
or U11725 (N_11725,N_11420,N_11298);
and U11726 (N_11726,N_11347,N_11371);
nor U11727 (N_11727,N_11268,N_11361);
xor U11728 (N_11728,N_11337,N_11361);
nand U11729 (N_11729,N_11338,N_11473);
nor U11730 (N_11730,N_11492,N_11499);
nor U11731 (N_11731,N_11430,N_11388);
and U11732 (N_11732,N_11433,N_11335);
xnor U11733 (N_11733,N_11480,N_11318);
nor U11734 (N_11734,N_11325,N_11257);
xor U11735 (N_11735,N_11469,N_11278);
nand U11736 (N_11736,N_11413,N_11332);
nand U11737 (N_11737,N_11388,N_11370);
nand U11738 (N_11738,N_11472,N_11268);
nor U11739 (N_11739,N_11395,N_11462);
or U11740 (N_11740,N_11432,N_11420);
xor U11741 (N_11741,N_11452,N_11421);
nand U11742 (N_11742,N_11486,N_11446);
or U11743 (N_11743,N_11271,N_11490);
nand U11744 (N_11744,N_11392,N_11252);
nand U11745 (N_11745,N_11342,N_11263);
or U11746 (N_11746,N_11282,N_11463);
nand U11747 (N_11747,N_11341,N_11402);
nor U11748 (N_11748,N_11380,N_11355);
or U11749 (N_11749,N_11352,N_11287);
xor U11750 (N_11750,N_11742,N_11624);
or U11751 (N_11751,N_11636,N_11599);
nand U11752 (N_11752,N_11530,N_11737);
nor U11753 (N_11753,N_11716,N_11645);
and U11754 (N_11754,N_11718,N_11560);
nand U11755 (N_11755,N_11655,N_11638);
nor U11756 (N_11756,N_11697,N_11672);
and U11757 (N_11757,N_11527,N_11605);
nor U11758 (N_11758,N_11677,N_11695);
nor U11759 (N_11759,N_11715,N_11734);
or U11760 (N_11760,N_11643,N_11710);
or U11761 (N_11761,N_11627,N_11646);
and U11762 (N_11762,N_11671,N_11708);
and U11763 (N_11763,N_11714,N_11520);
and U11764 (N_11764,N_11588,N_11691);
nor U11765 (N_11765,N_11614,N_11709);
nand U11766 (N_11766,N_11582,N_11681);
nor U11767 (N_11767,N_11705,N_11618);
nor U11768 (N_11768,N_11704,N_11522);
xnor U11769 (N_11769,N_11601,N_11583);
xnor U11770 (N_11770,N_11569,N_11620);
or U11771 (N_11771,N_11541,N_11699);
nor U11772 (N_11772,N_11612,N_11741);
and U11773 (N_11773,N_11647,N_11679);
xor U11774 (N_11774,N_11509,N_11553);
or U11775 (N_11775,N_11639,N_11552);
and U11776 (N_11776,N_11564,N_11698);
or U11777 (N_11777,N_11577,N_11634);
or U11778 (N_11778,N_11503,N_11533);
and U11779 (N_11779,N_11657,N_11508);
nor U11780 (N_11780,N_11661,N_11515);
or U11781 (N_11781,N_11502,N_11743);
nand U11782 (N_11782,N_11619,N_11732);
or U11783 (N_11783,N_11514,N_11543);
or U11784 (N_11784,N_11728,N_11525);
nor U11785 (N_11785,N_11607,N_11633);
or U11786 (N_11786,N_11635,N_11632);
and U11787 (N_11787,N_11551,N_11547);
and U11788 (N_11788,N_11740,N_11707);
xnor U11789 (N_11789,N_11680,N_11623);
or U11790 (N_11790,N_11631,N_11596);
nor U11791 (N_11791,N_11600,N_11526);
nor U11792 (N_11792,N_11745,N_11559);
and U11793 (N_11793,N_11687,N_11589);
and U11794 (N_11794,N_11669,N_11688);
and U11795 (N_11795,N_11719,N_11660);
nand U11796 (N_11796,N_11720,N_11587);
or U11797 (N_11797,N_11717,N_11706);
nor U11798 (N_11798,N_11575,N_11640);
xnor U11799 (N_11799,N_11505,N_11531);
or U11800 (N_11800,N_11593,N_11517);
or U11801 (N_11801,N_11629,N_11696);
xor U11802 (N_11802,N_11590,N_11524);
or U11803 (N_11803,N_11665,N_11521);
nor U11804 (N_11804,N_11692,N_11573);
nor U11805 (N_11805,N_11504,N_11610);
nand U11806 (N_11806,N_11676,N_11506);
xnor U11807 (N_11807,N_11744,N_11650);
xnor U11808 (N_11808,N_11544,N_11659);
xor U11809 (N_11809,N_11511,N_11586);
nand U11810 (N_11810,N_11644,N_11637);
xnor U11811 (N_11811,N_11673,N_11642);
or U11812 (N_11812,N_11554,N_11733);
or U11813 (N_11813,N_11566,N_11611);
nand U11814 (N_11814,N_11548,N_11653);
xnor U11815 (N_11815,N_11556,N_11726);
xor U11816 (N_11816,N_11529,N_11641);
or U11817 (N_11817,N_11562,N_11536);
nor U11818 (N_11818,N_11594,N_11723);
or U11819 (N_11819,N_11736,N_11739);
or U11820 (N_11820,N_11724,N_11722);
xnor U11821 (N_11821,N_11546,N_11658);
or U11822 (N_11822,N_11670,N_11565);
xor U11823 (N_11823,N_11702,N_11689);
or U11824 (N_11824,N_11545,N_11703);
nand U11825 (N_11825,N_11735,N_11535);
or U11826 (N_11826,N_11602,N_11628);
nor U11827 (N_11827,N_11685,N_11609);
nand U11828 (N_11828,N_11523,N_11507);
or U11829 (N_11829,N_11570,N_11510);
nand U11830 (N_11830,N_11550,N_11501);
or U11831 (N_11831,N_11667,N_11557);
or U11832 (N_11832,N_11630,N_11662);
nor U11833 (N_11833,N_11598,N_11749);
xnor U11834 (N_11834,N_11581,N_11578);
nor U11835 (N_11835,N_11542,N_11652);
nand U11836 (N_11836,N_11537,N_11686);
and U11837 (N_11837,N_11608,N_11549);
nor U11838 (N_11838,N_11592,N_11712);
or U11839 (N_11839,N_11567,N_11555);
and U11840 (N_11840,N_11580,N_11538);
and U11841 (N_11841,N_11666,N_11597);
xor U11842 (N_11842,N_11654,N_11664);
or U11843 (N_11843,N_11591,N_11738);
nand U11844 (N_11844,N_11615,N_11617);
nand U11845 (N_11845,N_11613,N_11516);
or U11846 (N_11846,N_11729,N_11579);
nand U11847 (N_11847,N_11700,N_11725);
xor U11848 (N_11848,N_11721,N_11713);
and U11849 (N_11849,N_11684,N_11678);
nor U11850 (N_11850,N_11595,N_11621);
nand U11851 (N_11851,N_11585,N_11656);
nor U11852 (N_11852,N_11747,N_11682);
and U11853 (N_11853,N_11576,N_11574);
and U11854 (N_11854,N_11694,N_11540);
xnor U11855 (N_11855,N_11518,N_11606);
nor U11856 (N_11856,N_11663,N_11563);
xnor U11857 (N_11857,N_11727,N_11748);
and U11858 (N_11858,N_11648,N_11603);
nand U11859 (N_11859,N_11571,N_11622);
or U11860 (N_11860,N_11539,N_11701);
and U11861 (N_11861,N_11512,N_11690);
nor U11862 (N_11862,N_11731,N_11558);
xor U11863 (N_11863,N_11568,N_11674);
or U11864 (N_11864,N_11534,N_11649);
or U11865 (N_11865,N_11532,N_11616);
nand U11866 (N_11866,N_11513,N_11561);
nand U11867 (N_11867,N_11693,N_11626);
nand U11868 (N_11868,N_11584,N_11730);
nor U11869 (N_11869,N_11668,N_11683);
or U11870 (N_11870,N_11572,N_11711);
nand U11871 (N_11871,N_11746,N_11519);
or U11872 (N_11872,N_11625,N_11528);
nor U11873 (N_11873,N_11500,N_11651);
nand U11874 (N_11874,N_11604,N_11675);
nor U11875 (N_11875,N_11604,N_11700);
xor U11876 (N_11876,N_11597,N_11537);
nand U11877 (N_11877,N_11740,N_11639);
xor U11878 (N_11878,N_11697,N_11623);
xor U11879 (N_11879,N_11739,N_11529);
nor U11880 (N_11880,N_11694,N_11557);
nor U11881 (N_11881,N_11569,N_11673);
nor U11882 (N_11882,N_11507,N_11670);
nand U11883 (N_11883,N_11734,N_11546);
xnor U11884 (N_11884,N_11574,N_11693);
xor U11885 (N_11885,N_11538,N_11532);
or U11886 (N_11886,N_11698,N_11691);
nor U11887 (N_11887,N_11511,N_11527);
nand U11888 (N_11888,N_11711,N_11590);
nor U11889 (N_11889,N_11524,N_11667);
nor U11890 (N_11890,N_11668,N_11667);
nand U11891 (N_11891,N_11736,N_11545);
or U11892 (N_11892,N_11551,N_11660);
or U11893 (N_11893,N_11730,N_11679);
or U11894 (N_11894,N_11643,N_11747);
nand U11895 (N_11895,N_11501,N_11553);
xnor U11896 (N_11896,N_11739,N_11611);
or U11897 (N_11897,N_11584,N_11622);
or U11898 (N_11898,N_11512,N_11698);
nor U11899 (N_11899,N_11518,N_11727);
and U11900 (N_11900,N_11518,N_11643);
and U11901 (N_11901,N_11697,N_11636);
and U11902 (N_11902,N_11642,N_11630);
and U11903 (N_11903,N_11552,N_11702);
or U11904 (N_11904,N_11690,N_11612);
and U11905 (N_11905,N_11574,N_11738);
nor U11906 (N_11906,N_11714,N_11659);
xor U11907 (N_11907,N_11674,N_11632);
and U11908 (N_11908,N_11744,N_11729);
xor U11909 (N_11909,N_11723,N_11609);
and U11910 (N_11910,N_11668,N_11538);
nor U11911 (N_11911,N_11569,N_11635);
and U11912 (N_11912,N_11719,N_11662);
or U11913 (N_11913,N_11687,N_11598);
xnor U11914 (N_11914,N_11613,N_11727);
or U11915 (N_11915,N_11707,N_11656);
nand U11916 (N_11916,N_11654,N_11628);
nand U11917 (N_11917,N_11684,N_11699);
or U11918 (N_11918,N_11747,N_11629);
and U11919 (N_11919,N_11531,N_11618);
or U11920 (N_11920,N_11603,N_11591);
nand U11921 (N_11921,N_11718,N_11567);
or U11922 (N_11922,N_11608,N_11644);
nor U11923 (N_11923,N_11568,N_11708);
and U11924 (N_11924,N_11693,N_11513);
nand U11925 (N_11925,N_11518,N_11676);
and U11926 (N_11926,N_11705,N_11634);
or U11927 (N_11927,N_11626,N_11605);
nor U11928 (N_11928,N_11593,N_11530);
xor U11929 (N_11929,N_11637,N_11721);
nor U11930 (N_11930,N_11692,N_11733);
and U11931 (N_11931,N_11569,N_11743);
xor U11932 (N_11932,N_11620,N_11700);
nand U11933 (N_11933,N_11713,N_11672);
nand U11934 (N_11934,N_11689,N_11657);
xor U11935 (N_11935,N_11703,N_11702);
xor U11936 (N_11936,N_11591,N_11723);
or U11937 (N_11937,N_11529,N_11631);
xnor U11938 (N_11938,N_11513,N_11657);
and U11939 (N_11939,N_11721,N_11644);
nor U11940 (N_11940,N_11645,N_11616);
nor U11941 (N_11941,N_11726,N_11737);
nor U11942 (N_11942,N_11559,N_11691);
or U11943 (N_11943,N_11563,N_11617);
nor U11944 (N_11944,N_11632,N_11669);
or U11945 (N_11945,N_11704,N_11564);
nor U11946 (N_11946,N_11539,N_11666);
and U11947 (N_11947,N_11559,N_11551);
or U11948 (N_11948,N_11716,N_11555);
xor U11949 (N_11949,N_11746,N_11714);
nor U11950 (N_11950,N_11639,N_11670);
nand U11951 (N_11951,N_11688,N_11504);
or U11952 (N_11952,N_11689,N_11512);
or U11953 (N_11953,N_11652,N_11679);
or U11954 (N_11954,N_11640,N_11594);
nand U11955 (N_11955,N_11725,N_11563);
nor U11956 (N_11956,N_11517,N_11505);
nand U11957 (N_11957,N_11527,N_11555);
xnor U11958 (N_11958,N_11565,N_11530);
or U11959 (N_11959,N_11700,N_11625);
or U11960 (N_11960,N_11644,N_11749);
or U11961 (N_11961,N_11601,N_11679);
nand U11962 (N_11962,N_11709,N_11581);
xor U11963 (N_11963,N_11540,N_11646);
xor U11964 (N_11964,N_11579,N_11565);
xor U11965 (N_11965,N_11620,N_11639);
or U11966 (N_11966,N_11721,N_11571);
nor U11967 (N_11967,N_11500,N_11733);
xnor U11968 (N_11968,N_11536,N_11666);
nor U11969 (N_11969,N_11629,N_11562);
nand U11970 (N_11970,N_11514,N_11541);
nand U11971 (N_11971,N_11528,N_11506);
or U11972 (N_11972,N_11747,N_11571);
and U11973 (N_11973,N_11677,N_11601);
xor U11974 (N_11974,N_11517,N_11558);
nand U11975 (N_11975,N_11717,N_11648);
xor U11976 (N_11976,N_11583,N_11706);
or U11977 (N_11977,N_11722,N_11521);
and U11978 (N_11978,N_11538,N_11503);
or U11979 (N_11979,N_11504,N_11654);
xnor U11980 (N_11980,N_11530,N_11532);
nor U11981 (N_11981,N_11681,N_11715);
nor U11982 (N_11982,N_11646,N_11527);
xor U11983 (N_11983,N_11637,N_11748);
xnor U11984 (N_11984,N_11653,N_11534);
or U11985 (N_11985,N_11666,N_11642);
or U11986 (N_11986,N_11715,N_11678);
or U11987 (N_11987,N_11501,N_11715);
or U11988 (N_11988,N_11678,N_11601);
nor U11989 (N_11989,N_11679,N_11586);
nand U11990 (N_11990,N_11629,N_11716);
xnor U11991 (N_11991,N_11641,N_11739);
or U11992 (N_11992,N_11604,N_11520);
nor U11993 (N_11993,N_11709,N_11714);
and U11994 (N_11994,N_11737,N_11613);
xnor U11995 (N_11995,N_11624,N_11684);
nand U11996 (N_11996,N_11576,N_11718);
nor U11997 (N_11997,N_11585,N_11556);
nand U11998 (N_11998,N_11691,N_11533);
or U11999 (N_11999,N_11641,N_11690);
nand U12000 (N_12000,N_11957,N_11865);
and U12001 (N_12001,N_11831,N_11984);
xor U12002 (N_12002,N_11869,N_11890);
nand U12003 (N_12003,N_11927,N_11794);
nor U12004 (N_12004,N_11968,N_11939);
xnor U12005 (N_12005,N_11854,N_11889);
xnor U12006 (N_12006,N_11789,N_11929);
xor U12007 (N_12007,N_11975,N_11818);
xnor U12008 (N_12008,N_11809,N_11881);
and U12009 (N_12009,N_11944,N_11763);
nor U12010 (N_12010,N_11837,N_11756);
nand U12011 (N_12011,N_11878,N_11933);
nor U12012 (N_12012,N_11788,N_11852);
nor U12013 (N_12013,N_11775,N_11985);
nand U12014 (N_12014,N_11851,N_11992);
nand U12015 (N_12015,N_11971,N_11772);
and U12016 (N_12016,N_11770,N_11955);
or U12017 (N_12017,N_11754,N_11844);
nor U12018 (N_12018,N_11974,N_11931);
or U12019 (N_12019,N_11947,N_11849);
nor U12020 (N_12020,N_11903,N_11839);
xor U12021 (N_12021,N_11857,N_11954);
xor U12022 (N_12022,N_11817,N_11990);
or U12023 (N_12023,N_11815,N_11853);
and U12024 (N_12024,N_11926,N_11988);
nand U12025 (N_12025,N_11995,N_11977);
xor U12026 (N_12026,N_11959,N_11879);
nand U12027 (N_12027,N_11783,N_11780);
nand U12028 (N_12028,N_11885,N_11829);
and U12029 (N_12029,N_11883,N_11846);
nand U12030 (N_12030,N_11886,N_11960);
or U12031 (N_12031,N_11916,N_11768);
nor U12032 (N_12032,N_11790,N_11871);
or U12033 (N_12033,N_11918,N_11950);
or U12034 (N_12034,N_11765,N_11972);
and U12035 (N_12035,N_11755,N_11764);
nand U12036 (N_12036,N_11895,N_11993);
xor U12037 (N_12037,N_11920,N_11751);
xor U12038 (N_12038,N_11937,N_11862);
or U12039 (N_12039,N_11820,N_11996);
nor U12040 (N_12040,N_11834,N_11843);
or U12041 (N_12041,N_11914,N_11795);
and U12042 (N_12042,N_11987,N_11847);
nor U12043 (N_12043,N_11860,N_11911);
xnor U12044 (N_12044,N_11900,N_11962);
and U12045 (N_12045,N_11896,N_11766);
nand U12046 (N_12046,N_11757,N_11932);
nand U12047 (N_12047,N_11796,N_11824);
or U12048 (N_12048,N_11936,N_11943);
or U12049 (N_12049,N_11951,N_11953);
nand U12050 (N_12050,N_11759,N_11876);
and U12051 (N_12051,N_11774,N_11841);
or U12052 (N_12052,N_11956,N_11980);
nand U12053 (N_12053,N_11905,N_11884);
xnor U12054 (N_12054,N_11803,N_11859);
nor U12055 (N_12055,N_11899,N_11840);
or U12056 (N_12056,N_11835,N_11942);
nand U12057 (N_12057,N_11752,N_11753);
xnor U12058 (N_12058,N_11806,N_11930);
and U12059 (N_12059,N_11825,N_11779);
xnor U12060 (N_12060,N_11867,N_11791);
and U12061 (N_12061,N_11750,N_11981);
and U12062 (N_12062,N_11946,N_11804);
xnor U12063 (N_12063,N_11925,N_11907);
and U12064 (N_12064,N_11868,N_11917);
xnor U12065 (N_12065,N_11976,N_11938);
or U12066 (N_12066,N_11855,N_11940);
nor U12067 (N_12067,N_11888,N_11861);
xor U12068 (N_12068,N_11912,N_11948);
xnor U12069 (N_12069,N_11773,N_11802);
nand U12070 (N_12070,N_11758,N_11991);
and U12071 (N_12071,N_11836,N_11863);
xnor U12072 (N_12072,N_11893,N_11810);
nor U12073 (N_12073,N_11866,N_11819);
nand U12074 (N_12074,N_11776,N_11811);
nor U12075 (N_12075,N_11761,N_11812);
and U12076 (N_12076,N_11833,N_11874);
xnor U12077 (N_12077,N_11807,N_11921);
and U12078 (N_12078,N_11923,N_11813);
nor U12079 (N_12079,N_11787,N_11842);
nand U12080 (N_12080,N_11964,N_11828);
or U12081 (N_12081,N_11848,N_11873);
nor U12082 (N_12082,N_11904,N_11919);
nand U12083 (N_12083,N_11799,N_11928);
and U12084 (N_12084,N_11994,N_11778);
or U12085 (N_12085,N_11798,N_11870);
and U12086 (N_12086,N_11941,N_11821);
xor U12087 (N_12087,N_11967,N_11762);
and U12088 (N_12088,N_11800,N_11897);
xor U12089 (N_12089,N_11808,N_11973);
nor U12090 (N_12090,N_11894,N_11767);
nor U12091 (N_12091,N_11983,N_11826);
nor U12092 (N_12092,N_11781,N_11830);
and U12093 (N_12093,N_11997,N_11797);
xor U12094 (N_12094,N_11958,N_11979);
and U12095 (N_12095,N_11908,N_11934);
or U12096 (N_12096,N_11965,N_11827);
and U12097 (N_12097,N_11963,N_11838);
nor U12098 (N_12098,N_11935,N_11793);
nand U12099 (N_12099,N_11880,N_11782);
nand U12100 (N_12100,N_11832,N_11961);
and U12101 (N_12101,N_11982,N_11882);
nor U12102 (N_12102,N_11922,N_11760);
and U12103 (N_12103,N_11945,N_11887);
xor U12104 (N_12104,N_11909,N_11875);
xor U12105 (N_12105,N_11816,N_11949);
nand U12106 (N_12106,N_11771,N_11902);
or U12107 (N_12107,N_11952,N_11915);
and U12108 (N_12108,N_11801,N_11856);
nor U12109 (N_12109,N_11784,N_11998);
and U12110 (N_12110,N_11913,N_11989);
or U12111 (N_12111,N_11924,N_11970);
or U12112 (N_12112,N_11858,N_11986);
xor U12113 (N_12113,N_11891,N_11966);
or U12114 (N_12114,N_11814,N_11777);
nor U12115 (N_12115,N_11786,N_11969);
and U12116 (N_12116,N_11999,N_11805);
or U12117 (N_12117,N_11877,N_11906);
nor U12118 (N_12118,N_11910,N_11872);
xnor U12119 (N_12119,N_11785,N_11845);
nand U12120 (N_12120,N_11901,N_11823);
xnor U12121 (N_12121,N_11792,N_11850);
and U12122 (N_12122,N_11978,N_11892);
and U12123 (N_12123,N_11898,N_11822);
nor U12124 (N_12124,N_11864,N_11769);
and U12125 (N_12125,N_11968,N_11788);
or U12126 (N_12126,N_11879,N_11863);
and U12127 (N_12127,N_11916,N_11862);
nor U12128 (N_12128,N_11879,N_11878);
xor U12129 (N_12129,N_11901,N_11903);
xnor U12130 (N_12130,N_11911,N_11853);
nand U12131 (N_12131,N_11974,N_11873);
and U12132 (N_12132,N_11883,N_11946);
nand U12133 (N_12133,N_11854,N_11782);
or U12134 (N_12134,N_11974,N_11959);
nor U12135 (N_12135,N_11818,N_11807);
xnor U12136 (N_12136,N_11942,N_11877);
and U12137 (N_12137,N_11788,N_11777);
nand U12138 (N_12138,N_11923,N_11946);
and U12139 (N_12139,N_11774,N_11850);
nor U12140 (N_12140,N_11780,N_11898);
and U12141 (N_12141,N_11792,N_11927);
or U12142 (N_12142,N_11763,N_11852);
or U12143 (N_12143,N_11757,N_11782);
or U12144 (N_12144,N_11960,N_11780);
nor U12145 (N_12145,N_11931,N_11845);
nand U12146 (N_12146,N_11856,N_11770);
or U12147 (N_12147,N_11767,N_11840);
or U12148 (N_12148,N_11936,N_11940);
or U12149 (N_12149,N_11760,N_11838);
nor U12150 (N_12150,N_11881,N_11966);
and U12151 (N_12151,N_11987,N_11784);
nand U12152 (N_12152,N_11770,N_11934);
nand U12153 (N_12153,N_11889,N_11937);
nor U12154 (N_12154,N_11967,N_11940);
or U12155 (N_12155,N_11857,N_11761);
and U12156 (N_12156,N_11948,N_11790);
nor U12157 (N_12157,N_11772,N_11855);
xor U12158 (N_12158,N_11910,N_11944);
xor U12159 (N_12159,N_11940,N_11919);
and U12160 (N_12160,N_11965,N_11761);
nand U12161 (N_12161,N_11916,N_11866);
nand U12162 (N_12162,N_11773,N_11928);
xnor U12163 (N_12163,N_11751,N_11865);
xor U12164 (N_12164,N_11839,N_11958);
and U12165 (N_12165,N_11859,N_11989);
nand U12166 (N_12166,N_11878,N_11906);
xnor U12167 (N_12167,N_11932,N_11765);
and U12168 (N_12168,N_11890,N_11855);
xor U12169 (N_12169,N_11900,N_11968);
and U12170 (N_12170,N_11865,N_11895);
or U12171 (N_12171,N_11923,N_11773);
or U12172 (N_12172,N_11792,N_11799);
or U12173 (N_12173,N_11770,N_11760);
or U12174 (N_12174,N_11767,N_11750);
and U12175 (N_12175,N_11836,N_11890);
xnor U12176 (N_12176,N_11826,N_11915);
xor U12177 (N_12177,N_11787,N_11914);
or U12178 (N_12178,N_11833,N_11967);
and U12179 (N_12179,N_11984,N_11824);
nor U12180 (N_12180,N_11969,N_11862);
nand U12181 (N_12181,N_11763,N_11853);
or U12182 (N_12182,N_11774,N_11933);
or U12183 (N_12183,N_11867,N_11866);
or U12184 (N_12184,N_11873,N_11794);
or U12185 (N_12185,N_11835,N_11843);
or U12186 (N_12186,N_11891,N_11984);
xnor U12187 (N_12187,N_11831,N_11940);
nor U12188 (N_12188,N_11791,N_11900);
and U12189 (N_12189,N_11972,N_11901);
nand U12190 (N_12190,N_11955,N_11919);
nand U12191 (N_12191,N_11956,N_11799);
or U12192 (N_12192,N_11982,N_11926);
nor U12193 (N_12193,N_11894,N_11772);
nor U12194 (N_12194,N_11911,N_11878);
nand U12195 (N_12195,N_11759,N_11928);
nor U12196 (N_12196,N_11942,N_11804);
nand U12197 (N_12197,N_11979,N_11774);
and U12198 (N_12198,N_11924,N_11959);
nor U12199 (N_12199,N_11846,N_11968);
or U12200 (N_12200,N_11751,N_11814);
and U12201 (N_12201,N_11876,N_11766);
nor U12202 (N_12202,N_11804,N_11878);
nor U12203 (N_12203,N_11756,N_11854);
nand U12204 (N_12204,N_11769,N_11784);
and U12205 (N_12205,N_11910,N_11997);
nand U12206 (N_12206,N_11959,N_11900);
or U12207 (N_12207,N_11879,N_11992);
xnor U12208 (N_12208,N_11946,N_11771);
nor U12209 (N_12209,N_11932,N_11847);
nor U12210 (N_12210,N_11926,N_11946);
and U12211 (N_12211,N_11862,N_11855);
nor U12212 (N_12212,N_11852,N_11751);
nand U12213 (N_12213,N_11788,N_11994);
nand U12214 (N_12214,N_11761,N_11816);
xor U12215 (N_12215,N_11860,N_11864);
or U12216 (N_12216,N_11857,N_11942);
nand U12217 (N_12217,N_11797,N_11786);
or U12218 (N_12218,N_11857,N_11895);
xor U12219 (N_12219,N_11755,N_11989);
or U12220 (N_12220,N_11829,N_11854);
or U12221 (N_12221,N_11776,N_11938);
xor U12222 (N_12222,N_11994,N_11897);
and U12223 (N_12223,N_11839,N_11995);
nand U12224 (N_12224,N_11773,N_11976);
or U12225 (N_12225,N_11801,N_11844);
nor U12226 (N_12226,N_11771,N_11981);
nor U12227 (N_12227,N_11988,N_11783);
and U12228 (N_12228,N_11960,N_11785);
and U12229 (N_12229,N_11780,N_11766);
or U12230 (N_12230,N_11836,N_11907);
nand U12231 (N_12231,N_11962,N_11996);
or U12232 (N_12232,N_11897,N_11762);
and U12233 (N_12233,N_11995,N_11974);
xor U12234 (N_12234,N_11938,N_11771);
nand U12235 (N_12235,N_11865,N_11775);
and U12236 (N_12236,N_11904,N_11848);
or U12237 (N_12237,N_11809,N_11859);
or U12238 (N_12238,N_11973,N_11835);
and U12239 (N_12239,N_11952,N_11764);
nor U12240 (N_12240,N_11832,N_11982);
and U12241 (N_12241,N_11811,N_11999);
and U12242 (N_12242,N_11862,N_11830);
and U12243 (N_12243,N_11771,N_11810);
and U12244 (N_12244,N_11815,N_11812);
nand U12245 (N_12245,N_11825,N_11753);
xnor U12246 (N_12246,N_11803,N_11798);
nor U12247 (N_12247,N_11968,N_11787);
nand U12248 (N_12248,N_11801,N_11933);
xor U12249 (N_12249,N_11904,N_11927);
xnor U12250 (N_12250,N_12182,N_12026);
nand U12251 (N_12251,N_12232,N_12191);
nand U12252 (N_12252,N_12062,N_12096);
nand U12253 (N_12253,N_12067,N_12201);
nand U12254 (N_12254,N_12030,N_12152);
or U12255 (N_12255,N_12170,N_12010);
or U12256 (N_12256,N_12113,N_12205);
and U12257 (N_12257,N_12072,N_12145);
xnor U12258 (N_12258,N_12206,N_12217);
and U12259 (N_12259,N_12155,N_12039);
xor U12260 (N_12260,N_12186,N_12209);
xor U12261 (N_12261,N_12169,N_12154);
nand U12262 (N_12262,N_12123,N_12080);
and U12263 (N_12263,N_12228,N_12004);
nor U12264 (N_12264,N_12198,N_12220);
nor U12265 (N_12265,N_12031,N_12181);
and U12266 (N_12266,N_12188,N_12167);
nor U12267 (N_12267,N_12204,N_12027);
nand U12268 (N_12268,N_12242,N_12024);
nor U12269 (N_12269,N_12107,N_12015);
nor U12270 (N_12270,N_12137,N_12227);
and U12271 (N_12271,N_12138,N_12184);
or U12272 (N_12272,N_12032,N_12022);
and U12273 (N_12273,N_12116,N_12019);
nor U12274 (N_12274,N_12165,N_12020);
or U12275 (N_12275,N_12049,N_12078);
xor U12276 (N_12276,N_12118,N_12238);
and U12277 (N_12277,N_12136,N_12061);
and U12278 (N_12278,N_12075,N_12210);
nor U12279 (N_12279,N_12091,N_12108);
and U12280 (N_12280,N_12065,N_12168);
nand U12281 (N_12281,N_12193,N_12213);
and U12282 (N_12282,N_12237,N_12239);
or U12283 (N_12283,N_12106,N_12208);
and U12284 (N_12284,N_12122,N_12175);
or U12285 (N_12285,N_12249,N_12161);
nor U12286 (N_12286,N_12203,N_12140);
nor U12287 (N_12287,N_12174,N_12009);
and U12288 (N_12288,N_12215,N_12159);
nand U12289 (N_12289,N_12218,N_12007);
nand U12290 (N_12290,N_12016,N_12094);
xor U12291 (N_12291,N_12124,N_12156);
xor U12292 (N_12292,N_12120,N_12003);
nand U12293 (N_12293,N_12105,N_12035);
xnor U12294 (N_12294,N_12157,N_12050);
nor U12295 (N_12295,N_12176,N_12102);
and U12296 (N_12296,N_12025,N_12223);
xor U12297 (N_12297,N_12090,N_12064);
xor U12298 (N_12298,N_12070,N_12044);
nand U12299 (N_12299,N_12112,N_12079);
nor U12300 (N_12300,N_12224,N_12097);
and U12301 (N_12301,N_12087,N_12162);
and U12302 (N_12302,N_12059,N_12054);
nand U12303 (N_12303,N_12246,N_12229);
and U12304 (N_12304,N_12014,N_12126);
xor U12305 (N_12305,N_12110,N_12041);
and U12306 (N_12306,N_12195,N_12178);
or U12307 (N_12307,N_12129,N_12052);
or U12308 (N_12308,N_12055,N_12194);
or U12309 (N_12309,N_12017,N_12074);
and U12310 (N_12310,N_12231,N_12190);
xor U12311 (N_12311,N_12244,N_12083);
or U12312 (N_12312,N_12021,N_12151);
nand U12313 (N_12313,N_12125,N_12199);
nand U12314 (N_12314,N_12144,N_12115);
and U12315 (N_12315,N_12164,N_12098);
nand U12316 (N_12316,N_12139,N_12141);
and U12317 (N_12317,N_12221,N_12212);
nor U12318 (N_12318,N_12095,N_12002);
nand U12319 (N_12319,N_12093,N_12158);
nand U12320 (N_12320,N_12234,N_12033);
or U12321 (N_12321,N_12233,N_12214);
xnor U12322 (N_12322,N_12187,N_12076);
nand U12323 (N_12323,N_12202,N_12149);
nor U12324 (N_12324,N_12185,N_12100);
xnor U12325 (N_12325,N_12127,N_12040);
xnor U12326 (N_12326,N_12018,N_12111);
xor U12327 (N_12327,N_12058,N_12063);
nand U12328 (N_12328,N_12046,N_12008);
xnor U12329 (N_12329,N_12177,N_12036);
nand U12330 (N_12330,N_12146,N_12057);
xor U12331 (N_12331,N_12099,N_12069);
or U12332 (N_12332,N_12131,N_12060);
nand U12333 (N_12333,N_12114,N_12092);
nor U12334 (N_12334,N_12183,N_12132);
nor U12335 (N_12335,N_12142,N_12005);
nor U12336 (N_12336,N_12082,N_12088);
or U12337 (N_12337,N_12066,N_12147);
and U12338 (N_12338,N_12029,N_12071);
and U12339 (N_12339,N_12230,N_12073);
nor U12340 (N_12340,N_12117,N_12163);
nor U12341 (N_12341,N_12068,N_12084);
and U12342 (N_12342,N_12056,N_12133);
nand U12343 (N_12343,N_12104,N_12130);
or U12344 (N_12344,N_12245,N_12171);
xor U12345 (N_12345,N_12189,N_12219);
nor U12346 (N_12346,N_12222,N_12081);
nor U12347 (N_12347,N_12011,N_12134);
nor U12348 (N_12348,N_12197,N_12172);
nand U12349 (N_12349,N_12034,N_12028);
or U12350 (N_12350,N_12143,N_12216);
nand U12351 (N_12351,N_12166,N_12045);
or U12352 (N_12352,N_12023,N_12135);
xor U12353 (N_12353,N_12089,N_12173);
nor U12354 (N_12354,N_12153,N_12051);
xnor U12355 (N_12355,N_12128,N_12006);
xor U12356 (N_12356,N_12119,N_12148);
nand U12357 (N_12357,N_12192,N_12048);
and U12358 (N_12358,N_12012,N_12103);
xor U12359 (N_12359,N_12037,N_12200);
nor U12360 (N_12360,N_12101,N_12179);
nor U12361 (N_12361,N_12150,N_12248);
xnor U12362 (N_12362,N_12000,N_12247);
nor U12363 (N_12363,N_12013,N_12196);
nand U12364 (N_12364,N_12180,N_12085);
and U12365 (N_12365,N_12047,N_12086);
or U12366 (N_12366,N_12038,N_12053);
and U12367 (N_12367,N_12001,N_12121);
or U12368 (N_12368,N_12207,N_12225);
nand U12369 (N_12369,N_12109,N_12235);
nand U12370 (N_12370,N_12160,N_12211);
nor U12371 (N_12371,N_12241,N_12043);
or U12372 (N_12372,N_12243,N_12042);
and U12373 (N_12373,N_12226,N_12077);
nor U12374 (N_12374,N_12240,N_12236);
or U12375 (N_12375,N_12199,N_12115);
nand U12376 (N_12376,N_12025,N_12041);
or U12377 (N_12377,N_12111,N_12165);
xnor U12378 (N_12378,N_12244,N_12039);
nor U12379 (N_12379,N_12153,N_12209);
nand U12380 (N_12380,N_12245,N_12174);
and U12381 (N_12381,N_12133,N_12089);
nor U12382 (N_12382,N_12188,N_12220);
and U12383 (N_12383,N_12211,N_12135);
and U12384 (N_12384,N_12026,N_12023);
xnor U12385 (N_12385,N_12028,N_12170);
or U12386 (N_12386,N_12077,N_12185);
xor U12387 (N_12387,N_12007,N_12024);
and U12388 (N_12388,N_12039,N_12165);
or U12389 (N_12389,N_12241,N_12179);
xor U12390 (N_12390,N_12137,N_12121);
and U12391 (N_12391,N_12016,N_12237);
nand U12392 (N_12392,N_12132,N_12073);
nor U12393 (N_12393,N_12048,N_12195);
and U12394 (N_12394,N_12114,N_12223);
and U12395 (N_12395,N_12096,N_12105);
nand U12396 (N_12396,N_12126,N_12211);
and U12397 (N_12397,N_12150,N_12087);
nand U12398 (N_12398,N_12209,N_12238);
nand U12399 (N_12399,N_12168,N_12221);
nor U12400 (N_12400,N_12023,N_12009);
or U12401 (N_12401,N_12123,N_12130);
nor U12402 (N_12402,N_12070,N_12199);
and U12403 (N_12403,N_12003,N_12055);
or U12404 (N_12404,N_12095,N_12223);
nand U12405 (N_12405,N_12076,N_12058);
or U12406 (N_12406,N_12152,N_12028);
xnor U12407 (N_12407,N_12079,N_12004);
or U12408 (N_12408,N_12144,N_12011);
and U12409 (N_12409,N_12047,N_12203);
nand U12410 (N_12410,N_12129,N_12033);
or U12411 (N_12411,N_12096,N_12170);
nor U12412 (N_12412,N_12040,N_12125);
and U12413 (N_12413,N_12130,N_12107);
nor U12414 (N_12414,N_12226,N_12123);
and U12415 (N_12415,N_12156,N_12077);
or U12416 (N_12416,N_12108,N_12219);
nor U12417 (N_12417,N_12151,N_12108);
nor U12418 (N_12418,N_12204,N_12235);
nor U12419 (N_12419,N_12237,N_12235);
xor U12420 (N_12420,N_12245,N_12225);
or U12421 (N_12421,N_12137,N_12194);
or U12422 (N_12422,N_12190,N_12215);
nor U12423 (N_12423,N_12185,N_12052);
xor U12424 (N_12424,N_12210,N_12244);
nor U12425 (N_12425,N_12030,N_12072);
nand U12426 (N_12426,N_12194,N_12154);
or U12427 (N_12427,N_12078,N_12176);
or U12428 (N_12428,N_12002,N_12156);
xnor U12429 (N_12429,N_12081,N_12124);
nor U12430 (N_12430,N_12105,N_12137);
xnor U12431 (N_12431,N_12032,N_12137);
nand U12432 (N_12432,N_12110,N_12240);
nand U12433 (N_12433,N_12249,N_12107);
and U12434 (N_12434,N_12082,N_12098);
nand U12435 (N_12435,N_12216,N_12196);
nand U12436 (N_12436,N_12202,N_12222);
nor U12437 (N_12437,N_12107,N_12165);
or U12438 (N_12438,N_12090,N_12011);
nor U12439 (N_12439,N_12001,N_12235);
nand U12440 (N_12440,N_12077,N_12154);
nand U12441 (N_12441,N_12093,N_12068);
nand U12442 (N_12442,N_12070,N_12164);
and U12443 (N_12443,N_12071,N_12096);
and U12444 (N_12444,N_12156,N_12000);
or U12445 (N_12445,N_12043,N_12066);
xor U12446 (N_12446,N_12170,N_12164);
or U12447 (N_12447,N_12131,N_12169);
nand U12448 (N_12448,N_12078,N_12140);
nand U12449 (N_12449,N_12215,N_12175);
xnor U12450 (N_12450,N_12064,N_12069);
or U12451 (N_12451,N_12200,N_12212);
or U12452 (N_12452,N_12221,N_12007);
xor U12453 (N_12453,N_12225,N_12187);
and U12454 (N_12454,N_12057,N_12138);
nor U12455 (N_12455,N_12110,N_12089);
and U12456 (N_12456,N_12089,N_12210);
nor U12457 (N_12457,N_12146,N_12038);
nand U12458 (N_12458,N_12230,N_12235);
xor U12459 (N_12459,N_12212,N_12178);
nand U12460 (N_12460,N_12144,N_12223);
nand U12461 (N_12461,N_12000,N_12184);
and U12462 (N_12462,N_12242,N_12152);
nor U12463 (N_12463,N_12066,N_12131);
xnor U12464 (N_12464,N_12052,N_12055);
xnor U12465 (N_12465,N_12114,N_12166);
and U12466 (N_12466,N_12043,N_12203);
nand U12467 (N_12467,N_12149,N_12084);
xnor U12468 (N_12468,N_12141,N_12102);
nand U12469 (N_12469,N_12122,N_12102);
nand U12470 (N_12470,N_12079,N_12194);
nand U12471 (N_12471,N_12242,N_12081);
and U12472 (N_12472,N_12189,N_12140);
nor U12473 (N_12473,N_12109,N_12199);
xnor U12474 (N_12474,N_12190,N_12104);
nand U12475 (N_12475,N_12064,N_12053);
xor U12476 (N_12476,N_12190,N_12102);
xnor U12477 (N_12477,N_12127,N_12107);
and U12478 (N_12478,N_12138,N_12073);
or U12479 (N_12479,N_12152,N_12175);
nand U12480 (N_12480,N_12226,N_12122);
nand U12481 (N_12481,N_12228,N_12159);
and U12482 (N_12482,N_12187,N_12095);
or U12483 (N_12483,N_12247,N_12028);
nor U12484 (N_12484,N_12160,N_12079);
and U12485 (N_12485,N_12134,N_12029);
nor U12486 (N_12486,N_12167,N_12020);
and U12487 (N_12487,N_12024,N_12042);
xnor U12488 (N_12488,N_12170,N_12197);
or U12489 (N_12489,N_12174,N_12033);
nand U12490 (N_12490,N_12123,N_12089);
nor U12491 (N_12491,N_12179,N_12034);
or U12492 (N_12492,N_12035,N_12156);
or U12493 (N_12493,N_12201,N_12112);
nor U12494 (N_12494,N_12032,N_12077);
nor U12495 (N_12495,N_12166,N_12126);
xnor U12496 (N_12496,N_12077,N_12130);
or U12497 (N_12497,N_12240,N_12014);
or U12498 (N_12498,N_12053,N_12080);
xor U12499 (N_12499,N_12049,N_12223);
nor U12500 (N_12500,N_12429,N_12445);
and U12501 (N_12501,N_12495,N_12402);
nand U12502 (N_12502,N_12266,N_12324);
nand U12503 (N_12503,N_12479,N_12449);
xor U12504 (N_12504,N_12262,N_12306);
xnor U12505 (N_12505,N_12448,N_12440);
nand U12506 (N_12506,N_12434,N_12451);
nand U12507 (N_12507,N_12388,N_12494);
nand U12508 (N_12508,N_12310,N_12299);
and U12509 (N_12509,N_12374,N_12257);
or U12510 (N_12510,N_12436,N_12423);
and U12511 (N_12511,N_12364,N_12304);
or U12512 (N_12512,N_12354,N_12256);
xor U12513 (N_12513,N_12400,N_12279);
nand U12514 (N_12514,N_12492,N_12255);
or U12515 (N_12515,N_12416,N_12444);
nand U12516 (N_12516,N_12293,N_12333);
nand U12517 (N_12517,N_12417,N_12322);
or U12518 (N_12518,N_12398,N_12365);
and U12519 (N_12519,N_12291,N_12483);
nor U12520 (N_12520,N_12358,N_12489);
or U12521 (N_12521,N_12287,N_12372);
and U12522 (N_12522,N_12419,N_12428);
or U12523 (N_12523,N_12356,N_12309);
or U12524 (N_12524,N_12447,N_12278);
nand U12525 (N_12525,N_12455,N_12397);
nand U12526 (N_12526,N_12410,N_12341);
xnor U12527 (N_12527,N_12264,N_12373);
xor U12528 (N_12528,N_12357,N_12361);
xnor U12529 (N_12529,N_12286,N_12270);
and U12530 (N_12530,N_12377,N_12290);
or U12531 (N_12531,N_12362,N_12457);
or U12532 (N_12532,N_12325,N_12426);
and U12533 (N_12533,N_12301,N_12389);
nand U12534 (N_12534,N_12353,N_12381);
and U12535 (N_12535,N_12369,N_12348);
or U12536 (N_12536,N_12273,N_12438);
xnor U12537 (N_12537,N_12418,N_12359);
or U12538 (N_12538,N_12307,N_12472);
nand U12539 (N_12539,N_12328,N_12387);
and U12540 (N_12540,N_12288,N_12459);
or U12541 (N_12541,N_12276,N_12330);
nor U12542 (N_12542,N_12297,N_12285);
nand U12543 (N_12543,N_12390,N_12496);
nand U12544 (N_12544,N_12269,N_12403);
nand U12545 (N_12545,N_12268,N_12280);
or U12546 (N_12546,N_12452,N_12326);
or U12547 (N_12547,N_12331,N_12318);
or U12548 (N_12548,N_12317,N_12401);
and U12549 (N_12549,N_12473,N_12383);
and U12550 (N_12550,N_12303,N_12250);
nor U12551 (N_12551,N_12407,N_12474);
and U12552 (N_12552,N_12493,N_12395);
nand U12553 (N_12553,N_12338,N_12368);
xnor U12554 (N_12554,N_12352,N_12355);
nand U12555 (N_12555,N_12454,N_12380);
xnor U12556 (N_12556,N_12392,N_12414);
nand U12557 (N_12557,N_12409,N_12430);
nor U12558 (N_12558,N_12378,N_12334);
xor U12559 (N_12559,N_12298,N_12295);
nand U12560 (N_12560,N_12439,N_12431);
nor U12561 (N_12561,N_12463,N_12350);
nand U12562 (N_12562,N_12399,N_12320);
nor U12563 (N_12563,N_12366,N_12453);
nor U12564 (N_12564,N_12487,N_12469);
and U12565 (N_12565,N_12261,N_12462);
xnor U12566 (N_12566,N_12284,N_12458);
xor U12567 (N_12567,N_12484,N_12482);
and U12568 (N_12568,N_12468,N_12498);
nand U12569 (N_12569,N_12442,N_12465);
nor U12570 (N_12570,N_12274,N_12277);
nor U12571 (N_12571,N_12421,N_12302);
xnor U12572 (N_12572,N_12323,N_12259);
nand U12573 (N_12573,N_12382,N_12425);
and U12574 (N_12574,N_12433,N_12321);
and U12575 (N_12575,N_12476,N_12258);
xnor U12576 (N_12576,N_12437,N_12342);
or U12577 (N_12577,N_12480,N_12490);
and U12578 (N_12578,N_12422,N_12396);
and U12579 (N_12579,N_12435,N_12450);
and U12580 (N_12580,N_12415,N_12360);
and U12581 (N_12581,N_12497,N_12376);
or U12582 (N_12582,N_12265,N_12367);
xnor U12583 (N_12583,N_12340,N_12427);
xor U12584 (N_12584,N_12394,N_12471);
nor U12585 (N_12585,N_12384,N_12443);
or U12586 (N_12586,N_12466,N_12281);
xor U12587 (N_12587,N_12253,N_12339);
or U12588 (N_12588,N_12470,N_12478);
xor U12589 (N_12589,N_12456,N_12485);
and U12590 (N_12590,N_12319,N_12336);
xor U12591 (N_12591,N_12337,N_12363);
nor U12592 (N_12592,N_12347,N_12271);
nor U12593 (N_12593,N_12263,N_12345);
nor U12594 (N_12594,N_12499,N_12349);
and U12595 (N_12595,N_12311,N_12344);
or U12596 (N_12596,N_12313,N_12477);
or U12597 (N_12597,N_12386,N_12289);
nor U12598 (N_12598,N_12267,N_12413);
and U12599 (N_12599,N_12486,N_12300);
and U12600 (N_12600,N_12346,N_12294);
nand U12601 (N_12601,N_12460,N_12308);
xnor U12602 (N_12602,N_12329,N_12464);
nand U12603 (N_12603,N_12379,N_12393);
nand U12604 (N_12604,N_12488,N_12316);
nor U12605 (N_12605,N_12404,N_12292);
or U12606 (N_12606,N_12312,N_12343);
xor U12607 (N_12607,N_12412,N_12252);
or U12608 (N_12608,N_12441,N_12408);
nand U12609 (N_12609,N_12475,N_12467);
or U12610 (N_12610,N_12424,N_12405);
or U12611 (N_12611,N_12305,N_12420);
nand U12612 (N_12612,N_12296,N_12491);
nand U12613 (N_12613,N_12327,N_12461);
nor U12614 (N_12614,N_12335,N_12481);
nor U12615 (N_12615,N_12283,N_12391);
nor U12616 (N_12616,N_12385,N_12275);
nor U12617 (N_12617,N_12272,N_12282);
or U12618 (N_12618,N_12371,N_12411);
xor U12619 (N_12619,N_12406,N_12332);
xnor U12620 (N_12620,N_12251,N_12432);
or U12621 (N_12621,N_12370,N_12351);
xnor U12622 (N_12622,N_12314,N_12315);
nor U12623 (N_12623,N_12254,N_12375);
nand U12624 (N_12624,N_12446,N_12260);
nand U12625 (N_12625,N_12277,N_12332);
nor U12626 (N_12626,N_12418,N_12413);
and U12627 (N_12627,N_12361,N_12373);
xor U12628 (N_12628,N_12437,N_12383);
nand U12629 (N_12629,N_12447,N_12381);
and U12630 (N_12630,N_12252,N_12377);
xor U12631 (N_12631,N_12277,N_12446);
and U12632 (N_12632,N_12285,N_12272);
or U12633 (N_12633,N_12475,N_12462);
or U12634 (N_12634,N_12254,N_12342);
xor U12635 (N_12635,N_12302,N_12290);
or U12636 (N_12636,N_12358,N_12404);
nand U12637 (N_12637,N_12396,N_12443);
nor U12638 (N_12638,N_12341,N_12481);
nor U12639 (N_12639,N_12356,N_12339);
and U12640 (N_12640,N_12408,N_12493);
nand U12641 (N_12641,N_12427,N_12417);
xor U12642 (N_12642,N_12326,N_12434);
and U12643 (N_12643,N_12465,N_12348);
nor U12644 (N_12644,N_12378,N_12382);
or U12645 (N_12645,N_12428,N_12432);
nor U12646 (N_12646,N_12392,N_12330);
xor U12647 (N_12647,N_12375,N_12351);
xnor U12648 (N_12648,N_12417,N_12476);
and U12649 (N_12649,N_12397,N_12374);
xnor U12650 (N_12650,N_12434,N_12308);
nor U12651 (N_12651,N_12329,N_12276);
and U12652 (N_12652,N_12441,N_12325);
xnor U12653 (N_12653,N_12455,N_12406);
nor U12654 (N_12654,N_12368,N_12451);
xnor U12655 (N_12655,N_12305,N_12322);
xor U12656 (N_12656,N_12453,N_12356);
xnor U12657 (N_12657,N_12464,N_12438);
and U12658 (N_12658,N_12363,N_12318);
nor U12659 (N_12659,N_12340,N_12462);
xor U12660 (N_12660,N_12486,N_12467);
nor U12661 (N_12661,N_12399,N_12317);
xnor U12662 (N_12662,N_12356,N_12264);
or U12663 (N_12663,N_12259,N_12482);
nor U12664 (N_12664,N_12284,N_12377);
and U12665 (N_12665,N_12493,N_12417);
or U12666 (N_12666,N_12357,N_12380);
and U12667 (N_12667,N_12418,N_12287);
and U12668 (N_12668,N_12307,N_12451);
or U12669 (N_12669,N_12470,N_12419);
or U12670 (N_12670,N_12311,N_12268);
nand U12671 (N_12671,N_12425,N_12464);
xnor U12672 (N_12672,N_12441,N_12261);
or U12673 (N_12673,N_12312,N_12472);
nor U12674 (N_12674,N_12366,N_12265);
or U12675 (N_12675,N_12489,N_12345);
nand U12676 (N_12676,N_12310,N_12473);
nor U12677 (N_12677,N_12499,N_12456);
nand U12678 (N_12678,N_12435,N_12342);
xor U12679 (N_12679,N_12340,N_12455);
xor U12680 (N_12680,N_12384,N_12360);
and U12681 (N_12681,N_12274,N_12266);
nor U12682 (N_12682,N_12306,N_12342);
or U12683 (N_12683,N_12404,N_12291);
or U12684 (N_12684,N_12392,N_12301);
or U12685 (N_12685,N_12400,N_12481);
or U12686 (N_12686,N_12276,N_12337);
xnor U12687 (N_12687,N_12347,N_12436);
nor U12688 (N_12688,N_12393,N_12271);
or U12689 (N_12689,N_12336,N_12467);
xor U12690 (N_12690,N_12442,N_12468);
or U12691 (N_12691,N_12408,N_12329);
xnor U12692 (N_12692,N_12383,N_12483);
and U12693 (N_12693,N_12316,N_12447);
or U12694 (N_12694,N_12469,N_12363);
and U12695 (N_12695,N_12433,N_12329);
and U12696 (N_12696,N_12458,N_12300);
xor U12697 (N_12697,N_12321,N_12330);
nor U12698 (N_12698,N_12455,N_12479);
xor U12699 (N_12699,N_12454,N_12292);
nor U12700 (N_12700,N_12295,N_12395);
nor U12701 (N_12701,N_12368,N_12494);
nor U12702 (N_12702,N_12406,N_12325);
nor U12703 (N_12703,N_12423,N_12460);
and U12704 (N_12704,N_12265,N_12494);
nor U12705 (N_12705,N_12479,N_12474);
and U12706 (N_12706,N_12300,N_12442);
nor U12707 (N_12707,N_12302,N_12480);
nand U12708 (N_12708,N_12289,N_12264);
or U12709 (N_12709,N_12455,N_12263);
xnor U12710 (N_12710,N_12393,N_12317);
or U12711 (N_12711,N_12467,N_12372);
xnor U12712 (N_12712,N_12258,N_12402);
or U12713 (N_12713,N_12423,N_12332);
nand U12714 (N_12714,N_12426,N_12308);
xor U12715 (N_12715,N_12253,N_12470);
or U12716 (N_12716,N_12412,N_12437);
nor U12717 (N_12717,N_12293,N_12448);
and U12718 (N_12718,N_12399,N_12430);
nand U12719 (N_12719,N_12371,N_12428);
nand U12720 (N_12720,N_12334,N_12382);
nor U12721 (N_12721,N_12435,N_12261);
nor U12722 (N_12722,N_12340,N_12387);
nor U12723 (N_12723,N_12443,N_12439);
xor U12724 (N_12724,N_12304,N_12303);
xor U12725 (N_12725,N_12252,N_12382);
or U12726 (N_12726,N_12291,N_12282);
nand U12727 (N_12727,N_12490,N_12345);
nand U12728 (N_12728,N_12494,N_12480);
nor U12729 (N_12729,N_12286,N_12306);
nand U12730 (N_12730,N_12484,N_12355);
and U12731 (N_12731,N_12255,N_12365);
or U12732 (N_12732,N_12432,N_12414);
or U12733 (N_12733,N_12265,N_12499);
nor U12734 (N_12734,N_12293,N_12284);
nand U12735 (N_12735,N_12429,N_12465);
nand U12736 (N_12736,N_12316,N_12340);
nor U12737 (N_12737,N_12278,N_12393);
and U12738 (N_12738,N_12304,N_12350);
and U12739 (N_12739,N_12283,N_12448);
or U12740 (N_12740,N_12476,N_12356);
and U12741 (N_12741,N_12365,N_12490);
xor U12742 (N_12742,N_12393,N_12339);
xor U12743 (N_12743,N_12353,N_12393);
nand U12744 (N_12744,N_12448,N_12354);
xor U12745 (N_12745,N_12370,N_12452);
nand U12746 (N_12746,N_12383,N_12311);
or U12747 (N_12747,N_12409,N_12369);
and U12748 (N_12748,N_12284,N_12279);
xor U12749 (N_12749,N_12386,N_12385);
or U12750 (N_12750,N_12663,N_12658);
xor U12751 (N_12751,N_12570,N_12548);
or U12752 (N_12752,N_12505,N_12659);
nand U12753 (N_12753,N_12699,N_12585);
and U12754 (N_12754,N_12673,N_12580);
nor U12755 (N_12755,N_12604,N_12613);
xor U12756 (N_12756,N_12631,N_12626);
or U12757 (N_12757,N_12589,N_12726);
nor U12758 (N_12758,N_12675,N_12743);
xnor U12759 (N_12759,N_12618,N_12724);
and U12760 (N_12760,N_12594,N_12596);
or U12761 (N_12761,N_12562,N_12552);
nand U12762 (N_12762,N_12534,N_12697);
nand U12763 (N_12763,N_12667,N_12744);
xnor U12764 (N_12764,N_12651,N_12561);
xor U12765 (N_12765,N_12539,N_12623);
nand U12766 (N_12766,N_12669,N_12737);
and U12767 (N_12767,N_12565,N_12664);
nand U12768 (N_12768,N_12621,N_12614);
xor U12769 (N_12769,N_12646,N_12642);
nand U12770 (N_12770,N_12502,N_12706);
nand U12771 (N_12771,N_12575,N_12602);
nor U12772 (N_12772,N_12571,N_12685);
nor U12773 (N_12773,N_12730,N_12718);
nor U12774 (N_12774,N_12683,N_12656);
xnor U12775 (N_12775,N_12703,N_12601);
nand U12776 (N_12776,N_12644,N_12680);
and U12777 (N_12777,N_12637,N_12603);
or U12778 (N_12778,N_12716,N_12510);
nor U12779 (N_12779,N_12694,N_12582);
or U12780 (N_12780,N_12628,N_12696);
nand U12781 (N_12781,N_12630,N_12723);
nor U12782 (N_12782,N_12678,N_12599);
nand U12783 (N_12783,N_12729,N_12660);
nand U12784 (N_12784,N_12702,N_12681);
nor U12785 (N_12785,N_12563,N_12523);
or U12786 (N_12786,N_12707,N_12600);
nand U12787 (N_12787,N_12544,N_12657);
xor U12788 (N_12788,N_12701,N_12624);
or U12789 (N_12789,N_12555,N_12513);
or U12790 (N_12790,N_12731,N_12719);
xnor U12791 (N_12791,N_12520,N_12521);
nand U12792 (N_12792,N_12512,N_12581);
nor U12793 (N_12793,N_12501,N_12738);
nand U12794 (N_12794,N_12745,N_12536);
nor U12795 (N_12795,N_12535,N_12721);
and U12796 (N_12796,N_12611,N_12591);
and U12797 (N_12797,N_12735,N_12511);
and U12798 (N_12798,N_12698,N_12676);
xnor U12799 (N_12799,N_12636,N_12748);
or U12800 (N_12800,N_12634,N_12610);
or U12801 (N_12801,N_12672,N_12720);
or U12802 (N_12802,N_12684,N_12715);
and U12803 (N_12803,N_12597,N_12717);
and U12804 (N_12804,N_12524,N_12627);
or U12805 (N_12805,N_12622,N_12527);
nand U12806 (N_12806,N_12519,N_12515);
nor U12807 (N_12807,N_12540,N_12643);
nand U12808 (N_12808,N_12617,N_12700);
or U12809 (N_12809,N_12648,N_12587);
xnor U12810 (N_12810,N_12528,N_12616);
and U12811 (N_12811,N_12525,N_12705);
or U12812 (N_12812,N_12689,N_12677);
nand U12813 (N_12813,N_12506,N_12674);
nand U12814 (N_12814,N_12560,N_12574);
nor U12815 (N_12815,N_12509,N_12736);
nor U12816 (N_12816,N_12584,N_12567);
nor U12817 (N_12817,N_12541,N_12526);
nand U12818 (N_12818,N_12522,N_12733);
and U12819 (N_12819,N_12609,N_12693);
or U12820 (N_12820,N_12714,N_12551);
xor U12821 (N_12821,N_12531,N_12692);
nor U12822 (N_12822,N_12655,N_12557);
xor U12823 (N_12823,N_12686,N_12529);
or U12824 (N_12824,N_12533,N_12641);
and U12825 (N_12825,N_12569,N_12554);
and U12826 (N_12826,N_12690,N_12516);
nor U12827 (N_12827,N_12568,N_12741);
nand U12828 (N_12828,N_12638,N_12620);
xor U12829 (N_12829,N_12605,N_12593);
or U12830 (N_12830,N_12632,N_12727);
nor U12831 (N_12831,N_12579,N_12635);
or U12832 (N_12832,N_12640,N_12661);
xnor U12833 (N_12833,N_12608,N_12665);
nand U12834 (N_12834,N_12566,N_12606);
xor U12835 (N_12835,N_12653,N_12691);
and U12836 (N_12836,N_12556,N_12629);
nor U12837 (N_12837,N_12532,N_12546);
nor U12838 (N_12838,N_12749,N_12530);
and U12839 (N_12839,N_12507,N_12722);
and U12840 (N_12840,N_12543,N_12670);
or U12841 (N_12841,N_12739,N_12654);
nor U12842 (N_12842,N_12711,N_12588);
xor U12843 (N_12843,N_12695,N_12709);
nand U12844 (N_12844,N_12558,N_12577);
nand U12845 (N_12845,N_12732,N_12572);
and U12846 (N_12846,N_12650,N_12559);
xor U12847 (N_12847,N_12514,N_12545);
and U12848 (N_12848,N_12537,N_12652);
or U12849 (N_12849,N_12712,N_12586);
nor U12850 (N_12850,N_12517,N_12740);
xor U12851 (N_12851,N_12679,N_12564);
nand U12852 (N_12852,N_12742,N_12747);
nand U12853 (N_12853,N_12538,N_12518);
xor U12854 (N_12854,N_12547,N_12595);
and U12855 (N_12855,N_12578,N_12573);
nand U12856 (N_12856,N_12542,N_12583);
or U12857 (N_12857,N_12612,N_12645);
or U12858 (N_12858,N_12590,N_12619);
xnor U12859 (N_12859,N_12734,N_12662);
nand U12860 (N_12860,N_12508,N_12671);
nor U12861 (N_12861,N_12666,N_12647);
nand U12862 (N_12862,N_12649,N_12728);
nor U12863 (N_12863,N_12687,N_12504);
and U12864 (N_12864,N_12639,N_12633);
nand U12865 (N_12865,N_12500,N_12704);
nand U12866 (N_12866,N_12688,N_12550);
or U12867 (N_12867,N_12549,N_12625);
nor U12868 (N_12868,N_12710,N_12713);
xnor U12869 (N_12869,N_12592,N_12553);
nor U12870 (N_12870,N_12576,N_12708);
xnor U12871 (N_12871,N_12668,N_12607);
nand U12872 (N_12872,N_12503,N_12746);
nand U12873 (N_12873,N_12725,N_12615);
nand U12874 (N_12874,N_12682,N_12598);
nand U12875 (N_12875,N_12741,N_12661);
nand U12876 (N_12876,N_12500,N_12718);
or U12877 (N_12877,N_12640,N_12546);
or U12878 (N_12878,N_12749,N_12720);
nand U12879 (N_12879,N_12638,N_12700);
xor U12880 (N_12880,N_12544,N_12677);
and U12881 (N_12881,N_12662,N_12614);
xnor U12882 (N_12882,N_12731,N_12741);
and U12883 (N_12883,N_12591,N_12676);
nand U12884 (N_12884,N_12691,N_12656);
nor U12885 (N_12885,N_12696,N_12713);
nand U12886 (N_12886,N_12663,N_12545);
nand U12887 (N_12887,N_12535,N_12727);
or U12888 (N_12888,N_12627,N_12587);
xnor U12889 (N_12889,N_12560,N_12661);
nor U12890 (N_12890,N_12726,N_12505);
nor U12891 (N_12891,N_12722,N_12745);
and U12892 (N_12892,N_12731,N_12713);
or U12893 (N_12893,N_12742,N_12529);
nand U12894 (N_12894,N_12629,N_12611);
and U12895 (N_12895,N_12695,N_12726);
nand U12896 (N_12896,N_12665,N_12684);
xnor U12897 (N_12897,N_12700,N_12531);
nor U12898 (N_12898,N_12527,N_12512);
xor U12899 (N_12899,N_12696,N_12637);
or U12900 (N_12900,N_12649,N_12648);
and U12901 (N_12901,N_12688,N_12571);
nor U12902 (N_12902,N_12582,N_12710);
and U12903 (N_12903,N_12714,N_12559);
xor U12904 (N_12904,N_12705,N_12555);
nand U12905 (N_12905,N_12712,N_12552);
nor U12906 (N_12906,N_12566,N_12733);
and U12907 (N_12907,N_12674,N_12583);
nor U12908 (N_12908,N_12747,N_12746);
xor U12909 (N_12909,N_12702,N_12549);
nand U12910 (N_12910,N_12513,N_12634);
nor U12911 (N_12911,N_12569,N_12564);
nor U12912 (N_12912,N_12714,N_12546);
xor U12913 (N_12913,N_12604,N_12695);
and U12914 (N_12914,N_12598,N_12590);
nand U12915 (N_12915,N_12603,N_12728);
nor U12916 (N_12916,N_12661,N_12687);
nor U12917 (N_12917,N_12562,N_12673);
xor U12918 (N_12918,N_12504,N_12654);
or U12919 (N_12919,N_12737,N_12668);
nor U12920 (N_12920,N_12727,N_12551);
and U12921 (N_12921,N_12744,N_12543);
nand U12922 (N_12922,N_12548,N_12721);
and U12923 (N_12923,N_12611,N_12718);
nand U12924 (N_12924,N_12684,N_12554);
or U12925 (N_12925,N_12633,N_12655);
or U12926 (N_12926,N_12566,N_12543);
nand U12927 (N_12927,N_12634,N_12501);
nand U12928 (N_12928,N_12687,N_12699);
or U12929 (N_12929,N_12600,N_12724);
or U12930 (N_12930,N_12662,N_12562);
xnor U12931 (N_12931,N_12544,N_12513);
and U12932 (N_12932,N_12697,N_12628);
or U12933 (N_12933,N_12518,N_12535);
nand U12934 (N_12934,N_12738,N_12519);
nand U12935 (N_12935,N_12595,N_12573);
and U12936 (N_12936,N_12671,N_12650);
nand U12937 (N_12937,N_12576,N_12624);
nand U12938 (N_12938,N_12699,N_12635);
nor U12939 (N_12939,N_12521,N_12574);
xor U12940 (N_12940,N_12724,N_12652);
xor U12941 (N_12941,N_12740,N_12626);
and U12942 (N_12942,N_12607,N_12714);
nand U12943 (N_12943,N_12575,N_12504);
or U12944 (N_12944,N_12571,N_12739);
xnor U12945 (N_12945,N_12613,N_12715);
and U12946 (N_12946,N_12638,N_12563);
xor U12947 (N_12947,N_12635,N_12538);
and U12948 (N_12948,N_12526,N_12720);
or U12949 (N_12949,N_12625,N_12729);
nor U12950 (N_12950,N_12728,N_12699);
or U12951 (N_12951,N_12529,N_12569);
or U12952 (N_12952,N_12541,N_12717);
nand U12953 (N_12953,N_12643,N_12726);
and U12954 (N_12954,N_12695,N_12743);
nor U12955 (N_12955,N_12645,N_12620);
nand U12956 (N_12956,N_12744,N_12736);
nand U12957 (N_12957,N_12680,N_12571);
nand U12958 (N_12958,N_12616,N_12539);
xnor U12959 (N_12959,N_12596,N_12724);
or U12960 (N_12960,N_12556,N_12709);
nor U12961 (N_12961,N_12586,N_12725);
or U12962 (N_12962,N_12665,N_12540);
nand U12963 (N_12963,N_12632,N_12719);
and U12964 (N_12964,N_12609,N_12741);
nand U12965 (N_12965,N_12597,N_12700);
nand U12966 (N_12966,N_12568,N_12529);
nor U12967 (N_12967,N_12694,N_12512);
and U12968 (N_12968,N_12740,N_12710);
nor U12969 (N_12969,N_12671,N_12648);
nand U12970 (N_12970,N_12625,N_12512);
xor U12971 (N_12971,N_12684,N_12545);
nor U12972 (N_12972,N_12683,N_12645);
nand U12973 (N_12973,N_12598,N_12734);
or U12974 (N_12974,N_12737,N_12562);
nand U12975 (N_12975,N_12596,N_12697);
and U12976 (N_12976,N_12727,N_12593);
nor U12977 (N_12977,N_12658,N_12726);
and U12978 (N_12978,N_12740,N_12658);
nand U12979 (N_12979,N_12695,N_12694);
and U12980 (N_12980,N_12702,N_12692);
xor U12981 (N_12981,N_12673,N_12629);
nand U12982 (N_12982,N_12511,N_12676);
nor U12983 (N_12983,N_12542,N_12731);
nand U12984 (N_12984,N_12597,N_12741);
and U12985 (N_12985,N_12503,N_12552);
or U12986 (N_12986,N_12558,N_12585);
xor U12987 (N_12987,N_12738,N_12518);
xnor U12988 (N_12988,N_12728,N_12723);
nand U12989 (N_12989,N_12745,N_12583);
nor U12990 (N_12990,N_12660,N_12606);
xnor U12991 (N_12991,N_12746,N_12678);
nand U12992 (N_12992,N_12519,N_12733);
nand U12993 (N_12993,N_12692,N_12512);
or U12994 (N_12994,N_12646,N_12525);
nor U12995 (N_12995,N_12517,N_12501);
xor U12996 (N_12996,N_12691,N_12522);
or U12997 (N_12997,N_12665,N_12661);
or U12998 (N_12998,N_12719,N_12578);
and U12999 (N_12999,N_12728,N_12563);
nor U13000 (N_13000,N_12815,N_12944);
xnor U13001 (N_13001,N_12978,N_12901);
nand U13002 (N_13002,N_12794,N_12832);
xnor U13003 (N_13003,N_12825,N_12782);
nor U13004 (N_13004,N_12792,N_12781);
xor U13005 (N_13005,N_12958,N_12925);
and U13006 (N_13006,N_12874,N_12882);
and U13007 (N_13007,N_12966,N_12904);
nand U13008 (N_13008,N_12865,N_12791);
or U13009 (N_13009,N_12891,N_12807);
and U13010 (N_13010,N_12780,N_12755);
and U13011 (N_13011,N_12992,N_12989);
or U13012 (N_13012,N_12840,N_12934);
and U13013 (N_13013,N_12753,N_12942);
or U13014 (N_13014,N_12758,N_12824);
nand U13015 (N_13015,N_12774,N_12864);
xnor U13016 (N_13016,N_12763,N_12835);
or U13017 (N_13017,N_12955,N_12796);
xnor U13018 (N_13018,N_12846,N_12750);
nand U13019 (N_13019,N_12998,N_12754);
nor U13020 (N_13020,N_12827,N_12823);
and U13021 (N_13021,N_12946,N_12893);
xor U13022 (N_13022,N_12980,N_12918);
xnor U13023 (N_13023,N_12974,N_12854);
nor U13024 (N_13024,N_12756,N_12964);
or U13025 (N_13025,N_12797,N_12852);
nand U13026 (N_13026,N_12994,N_12931);
and U13027 (N_13027,N_12784,N_12833);
nand U13028 (N_13028,N_12762,N_12943);
and U13029 (N_13029,N_12940,N_12887);
nor U13030 (N_13030,N_12976,N_12805);
and U13031 (N_13031,N_12801,N_12811);
nor U13032 (N_13032,N_12834,N_12919);
and U13033 (N_13033,N_12871,N_12902);
nor U13034 (N_13034,N_12808,N_12929);
or U13035 (N_13035,N_12802,N_12973);
xnor U13036 (N_13036,N_12937,N_12981);
and U13037 (N_13037,N_12848,N_12914);
nor U13038 (N_13038,N_12951,N_12959);
or U13039 (N_13039,N_12899,N_12799);
nand U13040 (N_13040,N_12972,N_12788);
or U13041 (N_13041,N_12819,N_12957);
xor U13042 (N_13042,N_12786,N_12770);
nor U13043 (N_13043,N_12868,N_12941);
and U13044 (N_13044,N_12869,N_12793);
and U13045 (N_13045,N_12847,N_12988);
nor U13046 (N_13046,N_12809,N_12987);
xor U13047 (N_13047,N_12836,N_12983);
xor U13048 (N_13048,N_12971,N_12773);
nand U13049 (N_13049,N_12890,N_12843);
nand U13050 (N_13050,N_12804,N_12867);
nand U13051 (N_13051,N_12900,N_12818);
nor U13052 (N_13052,N_12772,N_12768);
nand U13053 (N_13053,N_12814,N_12766);
nor U13054 (N_13054,N_12909,N_12845);
nor U13055 (N_13055,N_12894,N_12828);
xor U13056 (N_13056,N_12870,N_12928);
nor U13057 (N_13057,N_12922,N_12751);
and U13058 (N_13058,N_12884,N_12916);
nor U13059 (N_13059,N_12965,N_12990);
xor U13060 (N_13060,N_12985,N_12886);
nor U13061 (N_13061,N_12897,N_12935);
xnor U13062 (N_13062,N_12789,N_12875);
nand U13063 (N_13063,N_12949,N_12895);
nor U13064 (N_13064,N_12945,N_12950);
and U13065 (N_13065,N_12798,N_12986);
and U13066 (N_13066,N_12999,N_12997);
xnor U13067 (N_13067,N_12926,N_12851);
nand U13068 (N_13068,N_12936,N_12883);
nand U13069 (N_13069,N_12878,N_12858);
xnor U13070 (N_13070,N_12862,N_12906);
and U13071 (N_13071,N_12881,N_12830);
xor U13072 (N_13072,N_12927,N_12776);
xnor U13073 (N_13073,N_12790,N_12938);
and U13074 (N_13074,N_12775,N_12779);
and U13075 (N_13075,N_12841,N_12982);
or U13076 (N_13076,N_12996,N_12863);
nand U13077 (N_13077,N_12816,N_12948);
nand U13078 (N_13078,N_12889,N_12960);
nor U13079 (N_13079,N_12866,N_12961);
xor U13080 (N_13080,N_12760,N_12783);
nor U13081 (N_13081,N_12861,N_12910);
nand U13082 (N_13082,N_12759,N_12880);
xor U13083 (N_13083,N_12829,N_12903);
nand U13084 (N_13084,N_12907,N_12842);
or U13085 (N_13085,N_12810,N_12820);
xnor U13086 (N_13086,N_12991,N_12839);
or U13087 (N_13087,N_12806,N_12908);
nor U13088 (N_13088,N_12932,N_12920);
xor U13089 (N_13089,N_12822,N_12954);
xor U13090 (N_13090,N_12984,N_12837);
and U13091 (N_13091,N_12963,N_12913);
xor U13092 (N_13092,N_12764,N_12947);
nand U13093 (N_13093,N_12977,N_12892);
nor U13094 (N_13094,N_12821,N_12877);
or U13095 (N_13095,N_12787,N_12771);
nor U13096 (N_13096,N_12888,N_12898);
and U13097 (N_13097,N_12975,N_12857);
xor U13098 (N_13098,N_12915,N_12970);
or U13099 (N_13099,N_12924,N_12850);
nor U13100 (N_13100,N_12930,N_12879);
or U13101 (N_13101,N_12885,N_12933);
nand U13102 (N_13102,N_12859,N_12765);
or U13103 (N_13103,N_12856,N_12962);
nor U13104 (N_13104,N_12778,N_12817);
and U13105 (N_13105,N_12761,N_12911);
nand U13106 (N_13106,N_12838,N_12917);
xnor U13107 (N_13107,N_12873,N_12993);
nor U13108 (N_13108,N_12969,N_12967);
and U13109 (N_13109,N_12905,N_12872);
and U13110 (N_13110,N_12912,N_12800);
and U13111 (N_13111,N_12849,N_12785);
xor U13112 (N_13112,N_12812,N_12769);
or U13113 (N_13113,N_12979,N_12777);
xor U13114 (N_13114,N_12939,N_12995);
nor U13115 (N_13115,N_12767,N_12956);
nor U13116 (N_13116,N_12826,N_12860);
nand U13117 (N_13117,N_12813,N_12876);
and U13118 (N_13118,N_12896,N_12803);
and U13119 (N_13119,N_12921,N_12853);
nand U13120 (N_13120,N_12831,N_12844);
or U13121 (N_13121,N_12752,N_12952);
and U13122 (N_13122,N_12923,N_12757);
or U13123 (N_13123,N_12953,N_12795);
or U13124 (N_13124,N_12968,N_12855);
xor U13125 (N_13125,N_12981,N_12802);
and U13126 (N_13126,N_12881,N_12805);
or U13127 (N_13127,N_12795,N_12854);
nor U13128 (N_13128,N_12926,N_12922);
xor U13129 (N_13129,N_12754,N_12919);
nor U13130 (N_13130,N_12897,N_12954);
nand U13131 (N_13131,N_12770,N_12869);
nand U13132 (N_13132,N_12762,N_12869);
and U13133 (N_13133,N_12932,N_12934);
or U13134 (N_13134,N_12908,N_12865);
nor U13135 (N_13135,N_12760,N_12945);
xnor U13136 (N_13136,N_12980,N_12776);
and U13137 (N_13137,N_12928,N_12977);
nor U13138 (N_13138,N_12850,N_12837);
nor U13139 (N_13139,N_12938,N_12981);
xor U13140 (N_13140,N_12961,N_12951);
nor U13141 (N_13141,N_12965,N_12799);
nor U13142 (N_13142,N_12845,N_12921);
and U13143 (N_13143,N_12835,N_12965);
and U13144 (N_13144,N_12920,N_12847);
nand U13145 (N_13145,N_12789,N_12998);
nor U13146 (N_13146,N_12826,N_12865);
nand U13147 (N_13147,N_12851,N_12953);
xor U13148 (N_13148,N_12853,N_12897);
or U13149 (N_13149,N_12792,N_12820);
and U13150 (N_13150,N_12857,N_12831);
nor U13151 (N_13151,N_12979,N_12828);
nor U13152 (N_13152,N_12819,N_12848);
or U13153 (N_13153,N_12998,N_12965);
and U13154 (N_13154,N_12868,N_12986);
xnor U13155 (N_13155,N_12939,N_12842);
and U13156 (N_13156,N_12963,N_12933);
nand U13157 (N_13157,N_12844,N_12847);
and U13158 (N_13158,N_12916,N_12823);
and U13159 (N_13159,N_12955,N_12832);
nand U13160 (N_13160,N_12936,N_12960);
and U13161 (N_13161,N_12978,N_12861);
nand U13162 (N_13162,N_12829,N_12801);
xor U13163 (N_13163,N_12790,N_12985);
or U13164 (N_13164,N_12830,N_12892);
or U13165 (N_13165,N_12818,N_12889);
and U13166 (N_13166,N_12939,N_12941);
or U13167 (N_13167,N_12924,N_12832);
and U13168 (N_13168,N_12750,N_12876);
nor U13169 (N_13169,N_12810,N_12755);
or U13170 (N_13170,N_12779,N_12832);
or U13171 (N_13171,N_12798,N_12811);
and U13172 (N_13172,N_12992,N_12830);
xor U13173 (N_13173,N_12850,N_12814);
xnor U13174 (N_13174,N_12784,N_12763);
nand U13175 (N_13175,N_12935,N_12772);
xor U13176 (N_13176,N_12931,N_12872);
xnor U13177 (N_13177,N_12945,N_12858);
nor U13178 (N_13178,N_12834,N_12798);
nand U13179 (N_13179,N_12906,N_12841);
and U13180 (N_13180,N_12890,N_12905);
xor U13181 (N_13181,N_12979,N_12865);
or U13182 (N_13182,N_12770,N_12851);
and U13183 (N_13183,N_12942,N_12819);
and U13184 (N_13184,N_12854,N_12764);
nor U13185 (N_13185,N_12838,N_12789);
or U13186 (N_13186,N_12918,N_12997);
nand U13187 (N_13187,N_12899,N_12955);
nor U13188 (N_13188,N_12904,N_12786);
or U13189 (N_13189,N_12981,N_12758);
xnor U13190 (N_13190,N_12958,N_12831);
xor U13191 (N_13191,N_12812,N_12775);
nor U13192 (N_13192,N_12958,N_12965);
or U13193 (N_13193,N_12884,N_12897);
and U13194 (N_13194,N_12849,N_12884);
xnor U13195 (N_13195,N_12893,N_12883);
xnor U13196 (N_13196,N_12977,N_12936);
xor U13197 (N_13197,N_12875,N_12915);
or U13198 (N_13198,N_12973,N_12807);
nand U13199 (N_13199,N_12868,N_12882);
nand U13200 (N_13200,N_12901,N_12840);
nand U13201 (N_13201,N_12867,N_12918);
xnor U13202 (N_13202,N_12984,N_12891);
or U13203 (N_13203,N_12979,N_12846);
nand U13204 (N_13204,N_12999,N_12862);
nand U13205 (N_13205,N_12894,N_12821);
or U13206 (N_13206,N_12931,N_12976);
or U13207 (N_13207,N_12822,N_12864);
nand U13208 (N_13208,N_12881,N_12926);
or U13209 (N_13209,N_12916,N_12811);
or U13210 (N_13210,N_12872,N_12761);
nor U13211 (N_13211,N_12875,N_12828);
or U13212 (N_13212,N_12761,N_12813);
xnor U13213 (N_13213,N_12869,N_12758);
or U13214 (N_13214,N_12894,N_12856);
and U13215 (N_13215,N_12847,N_12793);
or U13216 (N_13216,N_12954,N_12858);
xnor U13217 (N_13217,N_12923,N_12761);
or U13218 (N_13218,N_12857,N_12999);
or U13219 (N_13219,N_12771,N_12823);
nand U13220 (N_13220,N_12867,N_12967);
xnor U13221 (N_13221,N_12767,N_12859);
nor U13222 (N_13222,N_12785,N_12806);
nor U13223 (N_13223,N_12987,N_12818);
nand U13224 (N_13224,N_12840,N_12807);
nor U13225 (N_13225,N_12758,N_12791);
and U13226 (N_13226,N_12867,N_12815);
nand U13227 (N_13227,N_12828,N_12951);
or U13228 (N_13228,N_12776,N_12863);
nand U13229 (N_13229,N_12773,N_12974);
and U13230 (N_13230,N_12763,N_12864);
nand U13231 (N_13231,N_12992,N_12845);
and U13232 (N_13232,N_12846,N_12890);
or U13233 (N_13233,N_12762,N_12952);
nor U13234 (N_13234,N_12980,N_12933);
nor U13235 (N_13235,N_12921,N_12969);
nand U13236 (N_13236,N_12801,N_12880);
nand U13237 (N_13237,N_12976,N_12893);
nand U13238 (N_13238,N_12950,N_12985);
nand U13239 (N_13239,N_12833,N_12752);
and U13240 (N_13240,N_12880,N_12998);
xor U13241 (N_13241,N_12973,N_12901);
nand U13242 (N_13242,N_12838,N_12903);
and U13243 (N_13243,N_12966,N_12874);
or U13244 (N_13244,N_12918,N_12961);
nand U13245 (N_13245,N_12959,N_12799);
and U13246 (N_13246,N_12931,N_12988);
and U13247 (N_13247,N_12833,N_12848);
nor U13248 (N_13248,N_12995,N_12912);
nor U13249 (N_13249,N_12778,N_12925);
and U13250 (N_13250,N_13185,N_13151);
nand U13251 (N_13251,N_13072,N_13237);
nand U13252 (N_13252,N_13187,N_13091);
nor U13253 (N_13253,N_13196,N_13041);
nand U13254 (N_13254,N_13108,N_13028);
nand U13255 (N_13255,N_13201,N_13023);
nor U13256 (N_13256,N_13199,N_13060);
nand U13257 (N_13257,N_13197,N_13010);
nand U13258 (N_13258,N_13156,N_13180);
and U13259 (N_13259,N_13068,N_13173);
nand U13260 (N_13260,N_13018,N_13070);
or U13261 (N_13261,N_13065,N_13188);
or U13262 (N_13262,N_13193,N_13054);
xor U13263 (N_13263,N_13118,N_13026);
and U13264 (N_13264,N_13110,N_13131);
or U13265 (N_13265,N_13117,N_13106);
xor U13266 (N_13266,N_13067,N_13172);
nor U13267 (N_13267,N_13008,N_13229);
nand U13268 (N_13268,N_13139,N_13051);
and U13269 (N_13269,N_13214,N_13094);
nand U13270 (N_13270,N_13063,N_13205);
and U13271 (N_13271,N_13169,N_13002);
nand U13272 (N_13272,N_13085,N_13078);
xnor U13273 (N_13273,N_13114,N_13092);
or U13274 (N_13274,N_13046,N_13116);
xor U13275 (N_13275,N_13003,N_13007);
nor U13276 (N_13276,N_13155,N_13195);
nor U13277 (N_13277,N_13079,N_13243);
and U13278 (N_13278,N_13074,N_13042);
or U13279 (N_13279,N_13038,N_13175);
nand U13280 (N_13280,N_13152,N_13133);
xor U13281 (N_13281,N_13025,N_13192);
or U13282 (N_13282,N_13064,N_13107);
xnor U13283 (N_13283,N_13202,N_13102);
or U13284 (N_13284,N_13045,N_13093);
or U13285 (N_13285,N_13037,N_13066);
and U13286 (N_13286,N_13032,N_13212);
nand U13287 (N_13287,N_13226,N_13061);
xor U13288 (N_13288,N_13055,N_13142);
or U13289 (N_13289,N_13194,N_13016);
nor U13290 (N_13290,N_13238,N_13020);
nand U13291 (N_13291,N_13005,N_13178);
nor U13292 (N_13292,N_13179,N_13167);
xnor U13293 (N_13293,N_13132,N_13150);
and U13294 (N_13294,N_13204,N_13119);
nand U13295 (N_13295,N_13144,N_13121);
nor U13296 (N_13296,N_13058,N_13249);
and U13297 (N_13297,N_13245,N_13113);
nand U13298 (N_13298,N_13052,N_13153);
nor U13299 (N_13299,N_13069,N_13022);
and U13300 (N_13300,N_13176,N_13228);
xor U13301 (N_13301,N_13220,N_13209);
xor U13302 (N_13302,N_13130,N_13240);
nand U13303 (N_13303,N_13103,N_13100);
nand U13304 (N_13304,N_13112,N_13182);
xor U13305 (N_13305,N_13084,N_13077);
nand U13306 (N_13306,N_13241,N_13216);
nand U13307 (N_13307,N_13081,N_13062);
xor U13308 (N_13308,N_13124,N_13009);
nor U13309 (N_13309,N_13036,N_13128);
xnor U13310 (N_13310,N_13236,N_13105);
xor U13311 (N_13311,N_13136,N_13098);
or U13312 (N_13312,N_13000,N_13125);
xnor U13313 (N_13313,N_13019,N_13076);
xnor U13314 (N_13314,N_13148,N_13244);
nand U13315 (N_13315,N_13021,N_13165);
or U13316 (N_13316,N_13191,N_13215);
xnor U13317 (N_13317,N_13177,N_13115);
xor U13318 (N_13318,N_13040,N_13053);
or U13319 (N_13319,N_13088,N_13219);
nand U13320 (N_13320,N_13223,N_13247);
nor U13321 (N_13321,N_13073,N_13101);
xnor U13322 (N_13322,N_13013,N_13159);
nor U13323 (N_13323,N_13186,N_13164);
or U13324 (N_13324,N_13127,N_13011);
or U13325 (N_13325,N_13122,N_13146);
nor U13326 (N_13326,N_13048,N_13012);
and U13327 (N_13327,N_13232,N_13047);
nor U13328 (N_13328,N_13154,N_13184);
and U13329 (N_13329,N_13057,N_13157);
and U13330 (N_13330,N_13083,N_13217);
nor U13331 (N_13331,N_13166,N_13143);
nor U13332 (N_13332,N_13031,N_13120);
and U13333 (N_13333,N_13160,N_13024);
nor U13334 (N_13334,N_13015,N_13233);
nor U13335 (N_13335,N_13129,N_13086);
nor U13336 (N_13336,N_13218,N_13001);
xnor U13337 (N_13337,N_13095,N_13044);
nor U13338 (N_13338,N_13030,N_13017);
nor U13339 (N_13339,N_13242,N_13089);
or U13340 (N_13340,N_13059,N_13227);
and U13341 (N_13341,N_13210,N_13162);
xor U13342 (N_13342,N_13140,N_13149);
and U13343 (N_13343,N_13246,N_13206);
or U13344 (N_13344,N_13207,N_13090);
or U13345 (N_13345,N_13004,N_13170);
nand U13346 (N_13346,N_13056,N_13145);
xnor U13347 (N_13347,N_13050,N_13181);
nand U13348 (N_13348,N_13161,N_13174);
nand U13349 (N_13349,N_13183,N_13158);
xor U13350 (N_13350,N_13006,N_13082);
nor U13351 (N_13351,N_13027,N_13141);
xnor U13352 (N_13352,N_13211,N_13034);
xor U13353 (N_13353,N_13235,N_13033);
xnor U13354 (N_13354,N_13080,N_13035);
nand U13355 (N_13355,N_13075,N_13111);
and U13356 (N_13356,N_13137,N_13147);
and U13357 (N_13357,N_13099,N_13029);
or U13358 (N_13358,N_13248,N_13134);
nor U13359 (N_13359,N_13087,N_13198);
and U13360 (N_13360,N_13097,N_13071);
and U13361 (N_13361,N_13203,N_13014);
nor U13362 (N_13362,N_13096,N_13135);
and U13363 (N_13363,N_13225,N_13231);
xnor U13364 (N_13364,N_13239,N_13168);
nor U13365 (N_13365,N_13234,N_13104);
nor U13366 (N_13366,N_13190,N_13043);
or U13367 (N_13367,N_13213,N_13171);
and U13368 (N_13368,N_13163,N_13049);
and U13369 (N_13369,N_13138,N_13221);
xnor U13370 (N_13370,N_13224,N_13123);
and U13371 (N_13371,N_13230,N_13109);
nand U13372 (N_13372,N_13208,N_13200);
xor U13373 (N_13373,N_13039,N_13126);
nand U13374 (N_13374,N_13222,N_13189);
nor U13375 (N_13375,N_13042,N_13073);
nor U13376 (N_13376,N_13024,N_13113);
xor U13377 (N_13377,N_13165,N_13218);
or U13378 (N_13378,N_13249,N_13155);
nor U13379 (N_13379,N_13065,N_13185);
xor U13380 (N_13380,N_13102,N_13192);
xor U13381 (N_13381,N_13122,N_13000);
nor U13382 (N_13382,N_13111,N_13235);
or U13383 (N_13383,N_13204,N_13148);
nand U13384 (N_13384,N_13084,N_13065);
xor U13385 (N_13385,N_13022,N_13238);
xor U13386 (N_13386,N_13159,N_13116);
xor U13387 (N_13387,N_13212,N_13100);
and U13388 (N_13388,N_13042,N_13244);
xor U13389 (N_13389,N_13173,N_13051);
nor U13390 (N_13390,N_13110,N_13050);
xor U13391 (N_13391,N_13224,N_13018);
xnor U13392 (N_13392,N_13191,N_13069);
nand U13393 (N_13393,N_13229,N_13017);
nor U13394 (N_13394,N_13168,N_13009);
or U13395 (N_13395,N_13194,N_13008);
nand U13396 (N_13396,N_13167,N_13232);
and U13397 (N_13397,N_13086,N_13218);
and U13398 (N_13398,N_13234,N_13230);
or U13399 (N_13399,N_13081,N_13232);
xor U13400 (N_13400,N_13206,N_13020);
nor U13401 (N_13401,N_13192,N_13137);
nor U13402 (N_13402,N_13225,N_13107);
and U13403 (N_13403,N_13015,N_13216);
or U13404 (N_13404,N_13087,N_13024);
or U13405 (N_13405,N_13060,N_13184);
and U13406 (N_13406,N_13214,N_13042);
nor U13407 (N_13407,N_13065,N_13027);
and U13408 (N_13408,N_13005,N_13199);
nor U13409 (N_13409,N_13247,N_13157);
or U13410 (N_13410,N_13075,N_13187);
and U13411 (N_13411,N_13193,N_13229);
nor U13412 (N_13412,N_13080,N_13064);
and U13413 (N_13413,N_13129,N_13228);
nand U13414 (N_13414,N_13187,N_13105);
or U13415 (N_13415,N_13204,N_13032);
xor U13416 (N_13416,N_13180,N_13029);
xor U13417 (N_13417,N_13131,N_13185);
nand U13418 (N_13418,N_13104,N_13197);
nand U13419 (N_13419,N_13090,N_13246);
nor U13420 (N_13420,N_13057,N_13037);
nand U13421 (N_13421,N_13157,N_13215);
and U13422 (N_13422,N_13084,N_13099);
nor U13423 (N_13423,N_13106,N_13104);
nor U13424 (N_13424,N_13117,N_13154);
nor U13425 (N_13425,N_13133,N_13020);
xnor U13426 (N_13426,N_13172,N_13077);
nand U13427 (N_13427,N_13018,N_13184);
nand U13428 (N_13428,N_13159,N_13047);
or U13429 (N_13429,N_13047,N_13161);
xnor U13430 (N_13430,N_13208,N_13085);
xor U13431 (N_13431,N_13146,N_13191);
or U13432 (N_13432,N_13063,N_13021);
nand U13433 (N_13433,N_13064,N_13109);
or U13434 (N_13434,N_13035,N_13028);
and U13435 (N_13435,N_13152,N_13093);
xor U13436 (N_13436,N_13028,N_13122);
or U13437 (N_13437,N_13037,N_13237);
and U13438 (N_13438,N_13187,N_13208);
or U13439 (N_13439,N_13025,N_13062);
nand U13440 (N_13440,N_13172,N_13236);
nor U13441 (N_13441,N_13099,N_13123);
and U13442 (N_13442,N_13235,N_13095);
xor U13443 (N_13443,N_13110,N_13066);
nor U13444 (N_13444,N_13189,N_13162);
or U13445 (N_13445,N_13157,N_13199);
nor U13446 (N_13446,N_13001,N_13152);
nor U13447 (N_13447,N_13230,N_13189);
and U13448 (N_13448,N_13235,N_13037);
and U13449 (N_13449,N_13166,N_13217);
or U13450 (N_13450,N_13136,N_13016);
nand U13451 (N_13451,N_13010,N_13120);
xor U13452 (N_13452,N_13058,N_13088);
nand U13453 (N_13453,N_13202,N_13134);
or U13454 (N_13454,N_13176,N_13099);
xnor U13455 (N_13455,N_13089,N_13066);
or U13456 (N_13456,N_13085,N_13193);
and U13457 (N_13457,N_13023,N_13184);
nand U13458 (N_13458,N_13222,N_13023);
nor U13459 (N_13459,N_13152,N_13145);
xor U13460 (N_13460,N_13054,N_13029);
and U13461 (N_13461,N_13083,N_13039);
nand U13462 (N_13462,N_13078,N_13006);
nor U13463 (N_13463,N_13000,N_13133);
or U13464 (N_13464,N_13014,N_13170);
xor U13465 (N_13465,N_13078,N_13205);
xor U13466 (N_13466,N_13208,N_13091);
and U13467 (N_13467,N_13106,N_13166);
or U13468 (N_13468,N_13154,N_13217);
and U13469 (N_13469,N_13198,N_13084);
nand U13470 (N_13470,N_13087,N_13166);
nor U13471 (N_13471,N_13140,N_13191);
and U13472 (N_13472,N_13152,N_13026);
xnor U13473 (N_13473,N_13125,N_13108);
and U13474 (N_13474,N_13095,N_13051);
or U13475 (N_13475,N_13177,N_13051);
nand U13476 (N_13476,N_13130,N_13157);
nand U13477 (N_13477,N_13134,N_13074);
or U13478 (N_13478,N_13223,N_13210);
xnor U13479 (N_13479,N_13056,N_13165);
nor U13480 (N_13480,N_13059,N_13198);
or U13481 (N_13481,N_13154,N_13240);
and U13482 (N_13482,N_13071,N_13062);
nand U13483 (N_13483,N_13210,N_13095);
nor U13484 (N_13484,N_13075,N_13041);
nand U13485 (N_13485,N_13093,N_13060);
nor U13486 (N_13486,N_13013,N_13025);
nand U13487 (N_13487,N_13222,N_13109);
xor U13488 (N_13488,N_13197,N_13000);
nor U13489 (N_13489,N_13036,N_13068);
nand U13490 (N_13490,N_13141,N_13244);
nand U13491 (N_13491,N_13015,N_13158);
nand U13492 (N_13492,N_13113,N_13109);
nor U13493 (N_13493,N_13236,N_13131);
or U13494 (N_13494,N_13079,N_13127);
xor U13495 (N_13495,N_13235,N_13164);
or U13496 (N_13496,N_13041,N_13089);
and U13497 (N_13497,N_13086,N_13094);
xnor U13498 (N_13498,N_13121,N_13190);
nor U13499 (N_13499,N_13194,N_13156);
nand U13500 (N_13500,N_13293,N_13367);
and U13501 (N_13501,N_13457,N_13345);
and U13502 (N_13502,N_13438,N_13442);
xor U13503 (N_13503,N_13302,N_13404);
nor U13504 (N_13504,N_13489,N_13405);
nand U13505 (N_13505,N_13390,N_13465);
nor U13506 (N_13506,N_13322,N_13412);
nand U13507 (N_13507,N_13466,N_13347);
and U13508 (N_13508,N_13298,N_13328);
or U13509 (N_13509,N_13313,N_13495);
or U13510 (N_13510,N_13349,N_13431);
xor U13511 (N_13511,N_13427,N_13401);
nor U13512 (N_13512,N_13352,N_13470);
xor U13513 (N_13513,N_13284,N_13496);
nand U13514 (N_13514,N_13464,N_13290);
nand U13515 (N_13515,N_13472,N_13282);
and U13516 (N_13516,N_13312,N_13388);
or U13517 (N_13517,N_13460,N_13294);
and U13518 (N_13518,N_13350,N_13392);
nor U13519 (N_13519,N_13451,N_13297);
xor U13520 (N_13520,N_13306,N_13428);
nand U13521 (N_13521,N_13452,N_13426);
xnor U13522 (N_13522,N_13276,N_13416);
nand U13523 (N_13523,N_13425,N_13351);
or U13524 (N_13524,N_13436,N_13320);
and U13525 (N_13525,N_13448,N_13286);
nand U13526 (N_13526,N_13391,N_13346);
or U13527 (N_13527,N_13471,N_13461);
nor U13528 (N_13528,N_13424,N_13359);
xor U13529 (N_13529,N_13422,N_13334);
and U13530 (N_13530,N_13371,N_13373);
and U13531 (N_13531,N_13273,N_13361);
and U13532 (N_13532,N_13274,N_13467);
nand U13533 (N_13533,N_13443,N_13376);
nor U13534 (N_13534,N_13270,N_13266);
or U13535 (N_13535,N_13354,N_13258);
nor U13536 (N_13536,N_13365,N_13263);
nor U13537 (N_13537,N_13333,N_13341);
nor U13538 (N_13538,N_13379,N_13413);
nand U13539 (N_13539,N_13393,N_13441);
nor U13540 (N_13540,N_13492,N_13387);
nand U13541 (N_13541,N_13479,N_13410);
xor U13542 (N_13542,N_13497,N_13317);
nor U13543 (N_13543,N_13364,N_13366);
nand U13544 (N_13544,N_13477,N_13475);
and U13545 (N_13545,N_13355,N_13321);
and U13546 (N_13546,N_13447,N_13295);
or U13547 (N_13547,N_13372,N_13303);
and U13548 (N_13548,N_13289,N_13307);
and U13549 (N_13549,N_13415,N_13257);
or U13550 (N_13550,N_13326,N_13279);
nor U13551 (N_13551,N_13421,N_13300);
and U13552 (N_13552,N_13325,N_13383);
nor U13553 (N_13553,N_13437,N_13285);
or U13554 (N_13554,N_13380,N_13480);
and U13555 (N_13555,N_13308,N_13356);
nand U13556 (N_13556,N_13456,N_13382);
and U13557 (N_13557,N_13264,N_13268);
or U13558 (N_13558,N_13414,N_13358);
nor U13559 (N_13559,N_13332,N_13408);
nor U13560 (N_13560,N_13260,N_13481);
nor U13561 (N_13561,N_13291,N_13487);
or U13562 (N_13562,N_13374,N_13450);
xnor U13563 (N_13563,N_13476,N_13433);
or U13564 (N_13564,N_13488,N_13250);
nand U13565 (N_13565,N_13329,N_13402);
xnor U13566 (N_13566,N_13339,N_13299);
nor U13567 (N_13567,N_13275,N_13251);
and U13568 (N_13568,N_13336,N_13344);
xnor U13569 (N_13569,N_13362,N_13269);
and U13570 (N_13570,N_13384,N_13440);
and U13571 (N_13571,N_13280,N_13324);
and U13572 (N_13572,N_13377,N_13357);
nand U13573 (N_13573,N_13439,N_13394);
nor U13574 (N_13574,N_13252,N_13493);
xor U13575 (N_13575,N_13309,N_13419);
xor U13576 (N_13576,N_13323,N_13490);
or U13577 (N_13577,N_13474,N_13429);
or U13578 (N_13578,N_13491,N_13473);
or U13579 (N_13579,N_13486,N_13417);
nor U13580 (N_13580,N_13259,N_13430);
xnor U13581 (N_13581,N_13316,N_13267);
and U13582 (N_13582,N_13305,N_13453);
or U13583 (N_13583,N_13288,N_13253);
nand U13584 (N_13584,N_13398,N_13482);
nand U13585 (N_13585,N_13484,N_13435);
nand U13586 (N_13586,N_13360,N_13272);
and U13587 (N_13587,N_13369,N_13459);
and U13588 (N_13588,N_13301,N_13330);
nand U13589 (N_13589,N_13319,N_13449);
xnor U13590 (N_13590,N_13418,N_13432);
or U13591 (N_13591,N_13283,N_13485);
and U13592 (N_13592,N_13375,N_13256);
nor U13593 (N_13593,N_13446,N_13277);
nor U13594 (N_13594,N_13254,N_13389);
xor U13595 (N_13595,N_13378,N_13311);
xor U13596 (N_13596,N_13385,N_13458);
and U13597 (N_13597,N_13411,N_13278);
nor U13598 (N_13598,N_13434,N_13370);
nor U13599 (N_13599,N_13400,N_13255);
xor U13600 (N_13600,N_13409,N_13338);
xnor U13601 (N_13601,N_13327,N_13469);
nand U13602 (N_13602,N_13494,N_13386);
nand U13603 (N_13603,N_13335,N_13315);
xnor U13604 (N_13604,N_13343,N_13397);
and U13605 (N_13605,N_13498,N_13478);
and U13606 (N_13606,N_13310,N_13281);
nor U13607 (N_13607,N_13271,N_13287);
nor U13608 (N_13608,N_13368,N_13261);
or U13609 (N_13609,N_13454,N_13331);
and U13610 (N_13610,N_13444,N_13262);
xnor U13611 (N_13611,N_13342,N_13483);
or U13612 (N_13612,N_13463,N_13407);
nor U13613 (N_13613,N_13381,N_13292);
nand U13614 (N_13614,N_13337,N_13423);
and U13615 (N_13615,N_13403,N_13499);
nand U13616 (N_13616,N_13340,N_13296);
and U13617 (N_13617,N_13420,N_13462);
or U13618 (N_13618,N_13314,N_13455);
or U13619 (N_13619,N_13445,N_13395);
nor U13620 (N_13620,N_13396,N_13318);
nor U13621 (N_13621,N_13265,N_13304);
nor U13622 (N_13622,N_13399,N_13406);
nor U13623 (N_13623,N_13468,N_13348);
and U13624 (N_13624,N_13353,N_13363);
or U13625 (N_13625,N_13364,N_13410);
and U13626 (N_13626,N_13359,N_13350);
or U13627 (N_13627,N_13266,N_13429);
nand U13628 (N_13628,N_13342,N_13303);
or U13629 (N_13629,N_13264,N_13435);
xnor U13630 (N_13630,N_13494,N_13316);
or U13631 (N_13631,N_13292,N_13433);
and U13632 (N_13632,N_13460,N_13431);
or U13633 (N_13633,N_13331,N_13295);
and U13634 (N_13634,N_13423,N_13495);
nor U13635 (N_13635,N_13464,N_13362);
and U13636 (N_13636,N_13353,N_13403);
nand U13637 (N_13637,N_13417,N_13343);
or U13638 (N_13638,N_13409,N_13407);
or U13639 (N_13639,N_13485,N_13269);
nand U13640 (N_13640,N_13372,N_13373);
xnor U13641 (N_13641,N_13255,N_13279);
nand U13642 (N_13642,N_13359,N_13409);
or U13643 (N_13643,N_13312,N_13460);
xor U13644 (N_13644,N_13449,N_13326);
nand U13645 (N_13645,N_13332,N_13324);
or U13646 (N_13646,N_13293,N_13432);
xnor U13647 (N_13647,N_13283,N_13296);
and U13648 (N_13648,N_13378,N_13297);
and U13649 (N_13649,N_13328,N_13309);
and U13650 (N_13650,N_13277,N_13407);
nand U13651 (N_13651,N_13457,N_13393);
nand U13652 (N_13652,N_13485,N_13496);
xor U13653 (N_13653,N_13339,N_13357);
xor U13654 (N_13654,N_13459,N_13368);
xor U13655 (N_13655,N_13317,N_13499);
nand U13656 (N_13656,N_13288,N_13418);
or U13657 (N_13657,N_13286,N_13435);
or U13658 (N_13658,N_13449,N_13367);
xor U13659 (N_13659,N_13433,N_13438);
nand U13660 (N_13660,N_13425,N_13428);
xor U13661 (N_13661,N_13379,N_13258);
nor U13662 (N_13662,N_13252,N_13255);
xor U13663 (N_13663,N_13259,N_13375);
nand U13664 (N_13664,N_13384,N_13483);
nand U13665 (N_13665,N_13258,N_13468);
xor U13666 (N_13666,N_13423,N_13427);
or U13667 (N_13667,N_13472,N_13311);
nor U13668 (N_13668,N_13317,N_13405);
nor U13669 (N_13669,N_13283,N_13332);
or U13670 (N_13670,N_13473,N_13309);
nand U13671 (N_13671,N_13384,N_13467);
xor U13672 (N_13672,N_13417,N_13306);
nand U13673 (N_13673,N_13317,N_13434);
nand U13674 (N_13674,N_13415,N_13456);
nand U13675 (N_13675,N_13381,N_13490);
nand U13676 (N_13676,N_13296,N_13250);
xor U13677 (N_13677,N_13315,N_13312);
nor U13678 (N_13678,N_13442,N_13276);
and U13679 (N_13679,N_13408,N_13393);
or U13680 (N_13680,N_13453,N_13279);
nor U13681 (N_13681,N_13428,N_13463);
nand U13682 (N_13682,N_13313,N_13494);
and U13683 (N_13683,N_13471,N_13283);
nand U13684 (N_13684,N_13403,N_13423);
nand U13685 (N_13685,N_13470,N_13463);
xor U13686 (N_13686,N_13428,N_13297);
and U13687 (N_13687,N_13400,N_13297);
or U13688 (N_13688,N_13447,N_13360);
nand U13689 (N_13689,N_13274,N_13342);
or U13690 (N_13690,N_13459,N_13305);
nand U13691 (N_13691,N_13371,N_13333);
nand U13692 (N_13692,N_13371,N_13351);
xor U13693 (N_13693,N_13459,N_13450);
or U13694 (N_13694,N_13489,N_13272);
nor U13695 (N_13695,N_13436,N_13321);
nand U13696 (N_13696,N_13373,N_13335);
nor U13697 (N_13697,N_13369,N_13283);
xor U13698 (N_13698,N_13268,N_13330);
nor U13699 (N_13699,N_13403,N_13380);
or U13700 (N_13700,N_13408,N_13339);
nand U13701 (N_13701,N_13290,N_13310);
or U13702 (N_13702,N_13322,N_13384);
or U13703 (N_13703,N_13310,N_13322);
nand U13704 (N_13704,N_13357,N_13305);
xnor U13705 (N_13705,N_13455,N_13272);
xnor U13706 (N_13706,N_13326,N_13456);
nand U13707 (N_13707,N_13253,N_13473);
nand U13708 (N_13708,N_13326,N_13352);
nand U13709 (N_13709,N_13406,N_13331);
nand U13710 (N_13710,N_13428,N_13394);
nor U13711 (N_13711,N_13314,N_13341);
xnor U13712 (N_13712,N_13396,N_13385);
nand U13713 (N_13713,N_13348,N_13317);
or U13714 (N_13714,N_13368,N_13404);
and U13715 (N_13715,N_13473,N_13405);
and U13716 (N_13716,N_13408,N_13465);
nor U13717 (N_13717,N_13271,N_13487);
xor U13718 (N_13718,N_13421,N_13382);
or U13719 (N_13719,N_13271,N_13428);
nor U13720 (N_13720,N_13472,N_13283);
nand U13721 (N_13721,N_13443,N_13470);
xnor U13722 (N_13722,N_13418,N_13390);
and U13723 (N_13723,N_13373,N_13385);
nand U13724 (N_13724,N_13314,N_13289);
nand U13725 (N_13725,N_13332,N_13256);
and U13726 (N_13726,N_13426,N_13388);
nor U13727 (N_13727,N_13384,N_13430);
nand U13728 (N_13728,N_13442,N_13480);
xnor U13729 (N_13729,N_13447,N_13258);
nor U13730 (N_13730,N_13323,N_13349);
nor U13731 (N_13731,N_13314,N_13278);
xor U13732 (N_13732,N_13442,N_13261);
nand U13733 (N_13733,N_13454,N_13467);
nand U13734 (N_13734,N_13315,N_13429);
and U13735 (N_13735,N_13365,N_13449);
or U13736 (N_13736,N_13326,N_13256);
or U13737 (N_13737,N_13497,N_13351);
nor U13738 (N_13738,N_13315,N_13441);
and U13739 (N_13739,N_13396,N_13435);
nor U13740 (N_13740,N_13270,N_13444);
nand U13741 (N_13741,N_13433,N_13260);
nand U13742 (N_13742,N_13266,N_13386);
nor U13743 (N_13743,N_13398,N_13270);
or U13744 (N_13744,N_13424,N_13437);
or U13745 (N_13745,N_13296,N_13407);
nand U13746 (N_13746,N_13367,N_13437);
xor U13747 (N_13747,N_13301,N_13319);
nand U13748 (N_13748,N_13265,N_13470);
nand U13749 (N_13749,N_13342,N_13250);
xor U13750 (N_13750,N_13687,N_13644);
and U13751 (N_13751,N_13618,N_13567);
nor U13752 (N_13752,N_13736,N_13616);
and U13753 (N_13753,N_13746,N_13628);
nand U13754 (N_13754,N_13528,N_13508);
and U13755 (N_13755,N_13617,N_13716);
nor U13756 (N_13756,N_13726,N_13586);
and U13757 (N_13757,N_13678,N_13589);
nand U13758 (N_13758,N_13661,N_13507);
nand U13759 (N_13759,N_13522,N_13540);
nand U13760 (N_13760,N_13509,N_13549);
xnor U13761 (N_13761,N_13636,N_13524);
or U13762 (N_13762,N_13610,N_13696);
nand U13763 (N_13763,N_13685,N_13526);
or U13764 (N_13764,N_13565,N_13557);
xnor U13765 (N_13765,N_13630,N_13662);
nor U13766 (N_13766,N_13633,N_13622);
nor U13767 (N_13767,N_13739,N_13733);
nor U13768 (N_13768,N_13723,N_13735);
nand U13769 (N_13769,N_13632,N_13655);
xnor U13770 (N_13770,N_13592,N_13527);
and U13771 (N_13771,N_13533,N_13569);
nor U13772 (N_13772,N_13690,N_13542);
nor U13773 (N_13773,N_13552,N_13707);
nor U13774 (N_13774,N_13715,N_13573);
nand U13775 (N_13775,N_13659,N_13672);
nor U13776 (N_13776,N_13681,N_13582);
xnor U13777 (N_13777,N_13580,N_13538);
or U13778 (N_13778,N_13682,N_13744);
or U13779 (N_13779,N_13611,N_13646);
xor U13780 (N_13780,N_13748,N_13559);
or U13781 (N_13781,N_13614,N_13639);
and U13782 (N_13782,N_13663,N_13667);
nand U13783 (N_13783,N_13654,N_13595);
and U13784 (N_13784,N_13749,N_13593);
or U13785 (N_13785,N_13642,N_13572);
nor U13786 (N_13786,N_13619,N_13574);
xor U13787 (N_13787,N_13698,N_13613);
nand U13788 (N_13788,N_13568,N_13673);
and U13789 (N_13789,N_13658,N_13608);
nor U13790 (N_13790,N_13517,N_13563);
and U13791 (N_13791,N_13712,N_13713);
nor U13792 (N_13792,N_13529,N_13692);
or U13793 (N_13793,N_13721,N_13742);
xnor U13794 (N_13794,N_13722,N_13547);
xor U13795 (N_13795,N_13640,N_13653);
and U13796 (N_13796,N_13703,N_13674);
nand U13797 (N_13797,N_13520,N_13629);
or U13798 (N_13798,N_13551,N_13679);
nand U13799 (N_13799,N_13506,N_13534);
or U13800 (N_13800,N_13603,N_13560);
nand U13801 (N_13801,N_13546,N_13695);
xor U13802 (N_13802,N_13558,N_13669);
or U13803 (N_13803,N_13544,N_13570);
and U13804 (N_13804,N_13596,N_13689);
and U13805 (N_13805,N_13605,N_13512);
and U13806 (N_13806,N_13743,N_13531);
or U13807 (N_13807,N_13624,N_13741);
nor U13808 (N_13808,N_13501,N_13647);
nor U13809 (N_13809,N_13649,N_13600);
or U13810 (N_13810,N_13519,N_13510);
xor U13811 (N_13811,N_13627,N_13700);
or U13812 (N_13812,N_13740,N_13583);
nand U13813 (N_13813,N_13747,N_13686);
nor U13814 (N_13814,N_13537,N_13541);
nor U13815 (N_13815,N_13631,N_13675);
or U13816 (N_13816,N_13651,N_13668);
xor U13817 (N_13817,N_13588,N_13607);
xnor U13818 (N_13818,N_13701,N_13677);
or U13819 (N_13819,N_13734,N_13585);
or U13820 (N_13820,N_13525,N_13590);
nor U13821 (N_13821,N_13575,N_13599);
nor U13822 (N_13822,N_13543,N_13587);
or U13823 (N_13823,N_13566,N_13718);
or U13824 (N_13824,N_13612,N_13516);
and U13825 (N_13825,N_13737,N_13719);
nor U13826 (N_13826,N_13708,N_13693);
nand U13827 (N_13827,N_13710,N_13556);
nand U13828 (N_13828,N_13641,N_13656);
xnor U13829 (N_13829,N_13523,N_13601);
xor U13830 (N_13830,N_13730,N_13694);
xor U13831 (N_13831,N_13635,N_13579);
nand U13832 (N_13832,N_13665,N_13697);
xor U13833 (N_13833,N_13513,N_13591);
nor U13834 (N_13834,N_13691,N_13732);
or U13835 (N_13835,N_13532,N_13514);
nand U13836 (N_13836,N_13604,N_13577);
or U13837 (N_13837,N_13745,N_13676);
and U13838 (N_13838,N_13626,N_13660);
xor U13839 (N_13839,N_13724,N_13666);
or U13840 (N_13840,N_13615,N_13578);
and U13841 (N_13841,N_13670,N_13539);
or U13842 (N_13842,N_13606,N_13511);
or U13843 (N_13843,N_13553,N_13720);
nand U13844 (N_13844,N_13683,N_13714);
nand U13845 (N_13845,N_13515,N_13684);
xor U13846 (N_13846,N_13706,N_13584);
and U13847 (N_13847,N_13688,N_13562);
and U13848 (N_13848,N_13671,N_13643);
nor U13849 (N_13849,N_13500,N_13727);
nand U13850 (N_13850,N_13609,N_13652);
and U13851 (N_13851,N_13576,N_13621);
or U13852 (N_13852,N_13650,N_13555);
or U13853 (N_13853,N_13709,N_13728);
or U13854 (N_13854,N_13680,N_13602);
or U13855 (N_13855,N_13504,N_13564);
xor U13856 (N_13856,N_13699,N_13657);
or U13857 (N_13857,N_13594,N_13637);
xnor U13858 (N_13858,N_13704,N_13535);
or U13859 (N_13859,N_13571,N_13518);
and U13860 (N_13860,N_13645,N_13554);
and U13861 (N_13861,N_13598,N_13545);
and U13862 (N_13862,N_13634,N_13521);
or U13863 (N_13863,N_13738,N_13548);
nand U13864 (N_13864,N_13729,N_13503);
xor U13865 (N_13865,N_13705,N_13717);
nand U13866 (N_13866,N_13550,N_13620);
and U13867 (N_13867,N_13502,N_13638);
nand U13868 (N_13868,N_13530,N_13597);
xor U13869 (N_13869,N_13536,N_13664);
and U13870 (N_13870,N_13625,N_13725);
or U13871 (N_13871,N_13505,N_13711);
xnor U13872 (N_13872,N_13702,N_13561);
and U13873 (N_13873,N_13731,N_13648);
nor U13874 (N_13874,N_13581,N_13623);
nand U13875 (N_13875,N_13741,N_13737);
and U13876 (N_13876,N_13644,N_13533);
xnor U13877 (N_13877,N_13541,N_13679);
nor U13878 (N_13878,N_13688,N_13749);
nand U13879 (N_13879,N_13557,N_13676);
and U13880 (N_13880,N_13699,N_13635);
nor U13881 (N_13881,N_13684,N_13567);
and U13882 (N_13882,N_13735,N_13706);
nor U13883 (N_13883,N_13697,N_13531);
or U13884 (N_13884,N_13720,N_13733);
nor U13885 (N_13885,N_13638,N_13676);
and U13886 (N_13886,N_13718,N_13743);
and U13887 (N_13887,N_13574,N_13618);
xnor U13888 (N_13888,N_13634,N_13660);
nand U13889 (N_13889,N_13632,N_13554);
xnor U13890 (N_13890,N_13623,N_13539);
or U13891 (N_13891,N_13525,N_13657);
xnor U13892 (N_13892,N_13535,N_13598);
or U13893 (N_13893,N_13613,N_13593);
xor U13894 (N_13894,N_13570,N_13716);
or U13895 (N_13895,N_13600,N_13573);
nor U13896 (N_13896,N_13591,N_13568);
and U13897 (N_13897,N_13585,N_13714);
nand U13898 (N_13898,N_13634,N_13598);
and U13899 (N_13899,N_13567,N_13745);
nor U13900 (N_13900,N_13520,N_13715);
and U13901 (N_13901,N_13541,N_13649);
or U13902 (N_13902,N_13511,N_13686);
or U13903 (N_13903,N_13644,N_13502);
nand U13904 (N_13904,N_13562,N_13516);
or U13905 (N_13905,N_13577,N_13629);
nor U13906 (N_13906,N_13636,N_13550);
or U13907 (N_13907,N_13543,N_13748);
nand U13908 (N_13908,N_13568,N_13561);
nor U13909 (N_13909,N_13550,N_13616);
nor U13910 (N_13910,N_13661,N_13706);
nand U13911 (N_13911,N_13554,N_13580);
or U13912 (N_13912,N_13514,N_13745);
and U13913 (N_13913,N_13684,N_13583);
xnor U13914 (N_13914,N_13507,N_13579);
and U13915 (N_13915,N_13731,N_13564);
xnor U13916 (N_13916,N_13742,N_13652);
xor U13917 (N_13917,N_13574,N_13725);
or U13918 (N_13918,N_13673,N_13672);
nor U13919 (N_13919,N_13669,N_13735);
nor U13920 (N_13920,N_13525,N_13512);
nor U13921 (N_13921,N_13708,N_13670);
or U13922 (N_13922,N_13599,N_13639);
or U13923 (N_13923,N_13566,N_13516);
or U13924 (N_13924,N_13531,N_13731);
and U13925 (N_13925,N_13661,N_13668);
nor U13926 (N_13926,N_13501,N_13533);
or U13927 (N_13927,N_13640,N_13578);
nor U13928 (N_13928,N_13513,N_13505);
nor U13929 (N_13929,N_13614,N_13734);
xor U13930 (N_13930,N_13641,N_13718);
nor U13931 (N_13931,N_13590,N_13744);
or U13932 (N_13932,N_13606,N_13739);
nor U13933 (N_13933,N_13625,N_13542);
nand U13934 (N_13934,N_13521,N_13633);
and U13935 (N_13935,N_13624,N_13501);
or U13936 (N_13936,N_13502,N_13696);
nand U13937 (N_13937,N_13560,N_13647);
nor U13938 (N_13938,N_13608,N_13626);
nor U13939 (N_13939,N_13587,N_13746);
xnor U13940 (N_13940,N_13642,N_13607);
or U13941 (N_13941,N_13567,N_13613);
xor U13942 (N_13942,N_13677,N_13558);
nor U13943 (N_13943,N_13511,N_13534);
xnor U13944 (N_13944,N_13579,N_13540);
or U13945 (N_13945,N_13506,N_13745);
xnor U13946 (N_13946,N_13734,N_13582);
and U13947 (N_13947,N_13624,N_13735);
nand U13948 (N_13948,N_13629,N_13613);
xor U13949 (N_13949,N_13655,N_13707);
xor U13950 (N_13950,N_13519,N_13731);
nand U13951 (N_13951,N_13636,N_13714);
and U13952 (N_13952,N_13706,N_13534);
or U13953 (N_13953,N_13528,N_13563);
and U13954 (N_13954,N_13640,N_13537);
nor U13955 (N_13955,N_13739,N_13678);
xor U13956 (N_13956,N_13604,N_13712);
xor U13957 (N_13957,N_13552,N_13590);
and U13958 (N_13958,N_13518,N_13592);
and U13959 (N_13959,N_13749,N_13507);
or U13960 (N_13960,N_13555,N_13552);
nand U13961 (N_13961,N_13570,N_13526);
or U13962 (N_13962,N_13587,N_13612);
or U13963 (N_13963,N_13612,N_13632);
or U13964 (N_13964,N_13701,N_13612);
nor U13965 (N_13965,N_13639,N_13604);
nor U13966 (N_13966,N_13729,N_13652);
and U13967 (N_13967,N_13522,N_13533);
and U13968 (N_13968,N_13643,N_13722);
nand U13969 (N_13969,N_13541,N_13579);
or U13970 (N_13970,N_13659,N_13584);
xnor U13971 (N_13971,N_13500,N_13568);
nand U13972 (N_13972,N_13739,N_13593);
nor U13973 (N_13973,N_13577,N_13573);
nand U13974 (N_13974,N_13606,N_13737);
nand U13975 (N_13975,N_13744,N_13739);
nor U13976 (N_13976,N_13726,N_13741);
nor U13977 (N_13977,N_13676,N_13694);
nor U13978 (N_13978,N_13511,N_13552);
xnor U13979 (N_13979,N_13541,N_13618);
nand U13980 (N_13980,N_13512,N_13724);
or U13981 (N_13981,N_13555,N_13721);
nor U13982 (N_13982,N_13598,N_13510);
and U13983 (N_13983,N_13584,N_13561);
and U13984 (N_13984,N_13739,N_13621);
nor U13985 (N_13985,N_13565,N_13594);
xor U13986 (N_13986,N_13748,N_13716);
xor U13987 (N_13987,N_13561,N_13746);
nand U13988 (N_13988,N_13681,N_13729);
xnor U13989 (N_13989,N_13529,N_13722);
or U13990 (N_13990,N_13598,N_13675);
nor U13991 (N_13991,N_13607,N_13522);
or U13992 (N_13992,N_13576,N_13709);
nor U13993 (N_13993,N_13559,N_13588);
xnor U13994 (N_13994,N_13630,N_13528);
xnor U13995 (N_13995,N_13712,N_13610);
or U13996 (N_13996,N_13601,N_13699);
and U13997 (N_13997,N_13641,N_13702);
xor U13998 (N_13998,N_13506,N_13588);
or U13999 (N_13999,N_13574,N_13549);
xor U14000 (N_14000,N_13797,N_13821);
xnor U14001 (N_14001,N_13896,N_13988);
nor U14002 (N_14002,N_13940,N_13930);
nand U14003 (N_14003,N_13751,N_13926);
nand U14004 (N_14004,N_13914,N_13997);
or U14005 (N_14005,N_13776,N_13928);
and U14006 (N_14006,N_13753,N_13848);
xor U14007 (N_14007,N_13841,N_13858);
xnor U14008 (N_14008,N_13781,N_13910);
xnor U14009 (N_14009,N_13990,N_13975);
xnor U14010 (N_14010,N_13810,N_13969);
xnor U14011 (N_14011,N_13767,N_13897);
or U14012 (N_14012,N_13917,N_13913);
xnor U14013 (N_14013,N_13970,N_13894);
and U14014 (N_14014,N_13980,N_13958);
nand U14015 (N_14015,N_13952,N_13992);
xor U14016 (N_14016,N_13864,N_13982);
xnor U14017 (N_14017,N_13840,N_13920);
and U14018 (N_14018,N_13770,N_13795);
xor U14019 (N_14019,N_13956,N_13921);
and U14020 (N_14020,N_13768,N_13993);
and U14021 (N_14021,N_13893,N_13777);
or U14022 (N_14022,N_13796,N_13812);
nand U14023 (N_14023,N_13785,N_13763);
nor U14024 (N_14024,N_13815,N_13862);
nand U14025 (N_14025,N_13750,N_13938);
nor U14026 (N_14026,N_13829,N_13919);
xor U14027 (N_14027,N_13847,N_13963);
nor U14028 (N_14028,N_13782,N_13927);
nand U14029 (N_14029,N_13849,N_13819);
xnor U14030 (N_14030,N_13998,N_13761);
nand U14031 (N_14031,N_13866,N_13895);
nand U14032 (N_14032,N_13948,N_13807);
nor U14033 (N_14033,N_13900,N_13892);
or U14034 (N_14034,N_13950,N_13861);
and U14035 (N_14035,N_13937,N_13856);
or U14036 (N_14036,N_13759,N_13813);
or U14037 (N_14037,N_13905,N_13916);
and U14038 (N_14038,N_13954,N_13853);
or U14039 (N_14039,N_13936,N_13838);
and U14040 (N_14040,N_13885,N_13825);
or U14041 (N_14041,N_13991,N_13964);
and U14042 (N_14042,N_13953,N_13774);
xor U14043 (N_14043,N_13822,N_13934);
or U14044 (N_14044,N_13945,N_13789);
and U14045 (N_14045,N_13806,N_13826);
and U14046 (N_14046,N_13933,N_13756);
nand U14047 (N_14047,N_13891,N_13762);
and U14048 (N_14048,N_13874,N_13901);
xor U14049 (N_14049,N_13983,N_13943);
and U14050 (N_14050,N_13788,N_13951);
nand U14051 (N_14051,N_13876,N_13863);
or U14052 (N_14052,N_13814,N_13946);
xor U14053 (N_14053,N_13965,N_13968);
or U14054 (N_14054,N_13771,N_13804);
xnor U14055 (N_14055,N_13974,N_13995);
nand U14056 (N_14056,N_13769,N_13909);
nor U14057 (N_14057,N_13820,N_13846);
nor U14058 (N_14058,N_13961,N_13899);
nor U14059 (N_14059,N_13884,N_13780);
or U14060 (N_14060,N_13879,N_13941);
xnor U14061 (N_14061,N_13903,N_13923);
nor U14062 (N_14062,N_13985,N_13857);
nand U14063 (N_14063,N_13989,N_13932);
and U14064 (N_14064,N_13787,N_13865);
and U14065 (N_14065,N_13845,N_13971);
xnor U14066 (N_14066,N_13764,N_13799);
nor U14067 (N_14067,N_13765,N_13783);
nor U14068 (N_14068,N_13830,N_13828);
xnor U14069 (N_14069,N_13859,N_13844);
and U14070 (N_14070,N_13809,N_13827);
xor U14071 (N_14071,N_13880,N_13877);
nand U14072 (N_14072,N_13868,N_13798);
xnor U14073 (N_14073,N_13855,N_13960);
and U14074 (N_14074,N_13922,N_13839);
nor U14075 (N_14075,N_13860,N_13870);
and U14076 (N_14076,N_13834,N_13888);
xnor U14077 (N_14077,N_13792,N_13786);
and U14078 (N_14078,N_13996,N_13925);
or U14079 (N_14079,N_13912,N_13955);
nor U14080 (N_14080,N_13784,N_13882);
nand U14081 (N_14081,N_13889,N_13779);
and U14082 (N_14082,N_13924,N_13754);
nor U14083 (N_14083,N_13816,N_13886);
nand U14084 (N_14084,N_13832,N_13793);
nor U14085 (N_14085,N_13871,N_13906);
nor U14086 (N_14086,N_13939,N_13875);
nand U14087 (N_14087,N_13851,N_13778);
nand U14088 (N_14088,N_13760,N_13872);
nor U14089 (N_14089,N_13775,N_13976);
and U14090 (N_14090,N_13805,N_13881);
nand U14091 (N_14091,N_13852,N_13907);
xnor U14092 (N_14092,N_13817,N_13766);
or U14093 (N_14093,N_13772,N_13883);
xor U14094 (N_14094,N_13842,N_13999);
xor U14095 (N_14095,N_13758,N_13869);
or U14096 (N_14096,N_13836,N_13947);
xor U14097 (N_14097,N_13801,N_13843);
and U14098 (N_14098,N_13935,N_13833);
or U14099 (N_14099,N_13929,N_13944);
xnor U14100 (N_14100,N_13898,N_13942);
nor U14101 (N_14101,N_13981,N_13915);
xor U14102 (N_14102,N_13949,N_13818);
xnor U14103 (N_14103,N_13931,N_13837);
and U14104 (N_14104,N_13831,N_13800);
nor U14105 (N_14105,N_13791,N_13904);
or U14106 (N_14106,N_13802,N_13823);
xor U14107 (N_14107,N_13873,N_13911);
xnor U14108 (N_14108,N_13986,N_13773);
and U14109 (N_14109,N_13978,N_13854);
or U14110 (N_14110,N_13824,N_13755);
and U14111 (N_14111,N_13811,N_13890);
nand U14112 (N_14112,N_13987,N_13757);
xnor U14113 (N_14113,N_13790,N_13803);
nor U14114 (N_14114,N_13887,N_13908);
or U14115 (N_14115,N_13977,N_13808);
and U14116 (N_14116,N_13979,N_13867);
or U14117 (N_14117,N_13902,N_13973);
or U14118 (N_14118,N_13966,N_13918);
nor U14119 (N_14119,N_13972,N_13959);
and U14120 (N_14120,N_13967,N_13962);
nand U14121 (N_14121,N_13994,N_13878);
nor U14122 (N_14122,N_13850,N_13957);
xnor U14123 (N_14123,N_13794,N_13752);
and U14124 (N_14124,N_13835,N_13984);
xor U14125 (N_14125,N_13923,N_13787);
xnor U14126 (N_14126,N_13893,N_13932);
and U14127 (N_14127,N_13962,N_13806);
nor U14128 (N_14128,N_13823,N_13806);
nor U14129 (N_14129,N_13894,N_13878);
and U14130 (N_14130,N_13809,N_13811);
or U14131 (N_14131,N_13789,N_13983);
or U14132 (N_14132,N_13937,N_13883);
xnor U14133 (N_14133,N_13795,N_13810);
xnor U14134 (N_14134,N_13813,N_13973);
nor U14135 (N_14135,N_13878,N_13753);
or U14136 (N_14136,N_13830,N_13871);
and U14137 (N_14137,N_13958,N_13766);
nor U14138 (N_14138,N_13762,N_13970);
or U14139 (N_14139,N_13983,N_13939);
nor U14140 (N_14140,N_13888,N_13833);
nor U14141 (N_14141,N_13862,N_13976);
xnor U14142 (N_14142,N_13877,N_13775);
nand U14143 (N_14143,N_13791,N_13933);
xnor U14144 (N_14144,N_13796,N_13867);
and U14145 (N_14145,N_13803,N_13946);
xor U14146 (N_14146,N_13796,N_13788);
xnor U14147 (N_14147,N_13781,N_13913);
nand U14148 (N_14148,N_13899,N_13783);
or U14149 (N_14149,N_13901,N_13900);
nor U14150 (N_14150,N_13866,N_13934);
nand U14151 (N_14151,N_13963,N_13783);
nor U14152 (N_14152,N_13917,N_13958);
or U14153 (N_14153,N_13939,N_13889);
or U14154 (N_14154,N_13832,N_13941);
and U14155 (N_14155,N_13757,N_13759);
or U14156 (N_14156,N_13823,N_13970);
xnor U14157 (N_14157,N_13781,N_13836);
xnor U14158 (N_14158,N_13955,N_13943);
nand U14159 (N_14159,N_13996,N_13875);
and U14160 (N_14160,N_13970,N_13843);
nand U14161 (N_14161,N_13835,N_13843);
xor U14162 (N_14162,N_13790,N_13946);
or U14163 (N_14163,N_13772,N_13803);
xor U14164 (N_14164,N_13824,N_13868);
nand U14165 (N_14165,N_13765,N_13966);
xnor U14166 (N_14166,N_13988,N_13925);
or U14167 (N_14167,N_13890,N_13782);
or U14168 (N_14168,N_13793,N_13820);
xor U14169 (N_14169,N_13868,N_13807);
xnor U14170 (N_14170,N_13863,N_13771);
nor U14171 (N_14171,N_13926,N_13816);
nor U14172 (N_14172,N_13795,N_13837);
and U14173 (N_14173,N_13845,N_13958);
and U14174 (N_14174,N_13990,N_13932);
xnor U14175 (N_14175,N_13795,N_13821);
nand U14176 (N_14176,N_13905,N_13784);
nor U14177 (N_14177,N_13990,N_13997);
xor U14178 (N_14178,N_13827,N_13780);
and U14179 (N_14179,N_13846,N_13891);
or U14180 (N_14180,N_13969,N_13852);
nand U14181 (N_14181,N_13880,N_13896);
or U14182 (N_14182,N_13980,N_13852);
nor U14183 (N_14183,N_13879,N_13942);
xor U14184 (N_14184,N_13945,N_13866);
nand U14185 (N_14185,N_13929,N_13787);
xnor U14186 (N_14186,N_13824,N_13968);
nand U14187 (N_14187,N_13784,N_13769);
nand U14188 (N_14188,N_13892,N_13760);
xnor U14189 (N_14189,N_13848,N_13961);
and U14190 (N_14190,N_13902,N_13846);
or U14191 (N_14191,N_13806,N_13885);
and U14192 (N_14192,N_13759,N_13936);
nand U14193 (N_14193,N_13856,N_13853);
nor U14194 (N_14194,N_13784,N_13853);
or U14195 (N_14195,N_13899,N_13886);
nand U14196 (N_14196,N_13760,N_13834);
and U14197 (N_14197,N_13754,N_13801);
and U14198 (N_14198,N_13945,N_13908);
nor U14199 (N_14199,N_13981,N_13766);
and U14200 (N_14200,N_13973,N_13796);
or U14201 (N_14201,N_13754,N_13887);
nand U14202 (N_14202,N_13922,N_13777);
xnor U14203 (N_14203,N_13904,N_13829);
nand U14204 (N_14204,N_13910,N_13771);
xnor U14205 (N_14205,N_13771,N_13879);
nor U14206 (N_14206,N_13864,N_13846);
or U14207 (N_14207,N_13841,N_13933);
or U14208 (N_14208,N_13799,N_13975);
and U14209 (N_14209,N_13909,N_13765);
or U14210 (N_14210,N_13878,N_13771);
nand U14211 (N_14211,N_13918,N_13818);
xor U14212 (N_14212,N_13999,N_13854);
xnor U14213 (N_14213,N_13865,N_13851);
nand U14214 (N_14214,N_13834,N_13830);
and U14215 (N_14215,N_13883,N_13836);
nand U14216 (N_14216,N_13815,N_13971);
and U14217 (N_14217,N_13894,N_13797);
and U14218 (N_14218,N_13825,N_13794);
or U14219 (N_14219,N_13919,N_13939);
nand U14220 (N_14220,N_13845,N_13997);
or U14221 (N_14221,N_13903,N_13768);
nand U14222 (N_14222,N_13756,N_13931);
and U14223 (N_14223,N_13931,N_13801);
or U14224 (N_14224,N_13995,N_13992);
nand U14225 (N_14225,N_13777,N_13765);
xnor U14226 (N_14226,N_13794,N_13780);
or U14227 (N_14227,N_13836,N_13937);
nor U14228 (N_14228,N_13883,N_13776);
nor U14229 (N_14229,N_13899,N_13862);
or U14230 (N_14230,N_13969,N_13948);
nand U14231 (N_14231,N_13975,N_13961);
xor U14232 (N_14232,N_13995,N_13861);
nor U14233 (N_14233,N_13882,N_13816);
xnor U14234 (N_14234,N_13812,N_13980);
and U14235 (N_14235,N_13837,N_13879);
nor U14236 (N_14236,N_13800,N_13897);
nor U14237 (N_14237,N_13820,N_13867);
or U14238 (N_14238,N_13923,N_13763);
nand U14239 (N_14239,N_13830,N_13935);
nor U14240 (N_14240,N_13910,N_13875);
nor U14241 (N_14241,N_13862,N_13842);
nand U14242 (N_14242,N_13975,N_13879);
or U14243 (N_14243,N_13875,N_13846);
nand U14244 (N_14244,N_13982,N_13935);
nor U14245 (N_14245,N_13975,N_13926);
nand U14246 (N_14246,N_13793,N_13812);
nand U14247 (N_14247,N_13901,N_13972);
xor U14248 (N_14248,N_13966,N_13962);
xnor U14249 (N_14249,N_13793,N_13854);
xnor U14250 (N_14250,N_14164,N_14158);
xnor U14251 (N_14251,N_14096,N_14049);
and U14252 (N_14252,N_14166,N_14013);
xnor U14253 (N_14253,N_14148,N_14167);
xor U14254 (N_14254,N_14106,N_14119);
xnor U14255 (N_14255,N_14007,N_14005);
nor U14256 (N_14256,N_14000,N_14059);
nor U14257 (N_14257,N_14047,N_14063);
or U14258 (N_14258,N_14198,N_14018);
nor U14259 (N_14259,N_14052,N_14051);
or U14260 (N_14260,N_14091,N_14233);
xor U14261 (N_14261,N_14110,N_14086);
nand U14262 (N_14262,N_14145,N_14033);
nor U14263 (N_14263,N_14090,N_14137);
or U14264 (N_14264,N_14234,N_14201);
nand U14265 (N_14265,N_14165,N_14154);
or U14266 (N_14266,N_14011,N_14131);
xor U14267 (N_14267,N_14141,N_14180);
nand U14268 (N_14268,N_14045,N_14153);
and U14269 (N_14269,N_14009,N_14043);
nor U14270 (N_14270,N_14161,N_14088);
or U14271 (N_14271,N_14179,N_14200);
nand U14272 (N_14272,N_14084,N_14210);
nor U14273 (N_14273,N_14229,N_14249);
or U14274 (N_14274,N_14177,N_14132);
and U14275 (N_14275,N_14117,N_14050);
xor U14276 (N_14276,N_14159,N_14127);
nand U14277 (N_14277,N_14103,N_14235);
and U14278 (N_14278,N_14204,N_14073);
nor U14279 (N_14279,N_14214,N_14072);
xor U14280 (N_14280,N_14243,N_14174);
or U14281 (N_14281,N_14218,N_14184);
or U14282 (N_14282,N_14195,N_14095);
nand U14283 (N_14283,N_14104,N_14207);
nand U14284 (N_14284,N_14206,N_14185);
nor U14285 (N_14285,N_14053,N_14240);
and U14286 (N_14286,N_14081,N_14055);
nor U14287 (N_14287,N_14160,N_14040);
nor U14288 (N_14288,N_14069,N_14037);
or U14289 (N_14289,N_14228,N_14039);
or U14290 (N_14290,N_14142,N_14056);
xor U14291 (N_14291,N_14006,N_14192);
or U14292 (N_14292,N_14169,N_14170);
xnor U14293 (N_14293,N_14028,N_14035);
nor U14294 (N_14294,N_14058,N_14173);
and U14295 (N_14295,N_14116,N_14187);
xnor U14296 (N_14296,N_14066,N_14038);
nand U14297 (N_14297,N_14019,N_14105);
nor U14298 (N_14298,N_14223,N_14188);
or U14299 (N_14299,N_14071,N_14034);
or U14300 (N_14300,N_14017,N_14060);
or U14301 (N_14301,N_14150,N_14093);
nand U14302 (N_14302,N_14026,N_14130);
or U14303 (N_14303,N_14118,N_14134);
or U14304 (N_14304,N_14189,N_14083);
nor U14305 (N_14305,N_14208,N_14212);
and U14306 (N_14306,N_14065,N_14002);
and U14307 (N_14307,N_14101,N_14178);
xnor U14308 (N_14308,N_14246,N_14054);
xnor U14309 (N_14309,N_14082,N_14021);
nand U14310 (N_14310,N_14183,N_14027);
or U14311 (N_14311,N_14205,N_14044);
nor U14312 (N_14312,N_14067,N_14216);
or U14313 (N_14313,N_14171,N_14176);
nor U14314 (N_14314,N_14213,N_14123);
or U14315 (N_14315,N_14016,N_14097);
nand U14316 (N_14316,N_14152,N_14114);
nor U14317 (N_14317,N_14068,N_14138);
and U14318 (N_14318,N_14133,N_14209);
or U14319 (N_14319,N_14237,N_14181);
nand U14320 (N_14320,N_14224,N_14041);
xor U14321 (N_14321,N_14100,N_14232);
or U14322 (N_14322,N_14139,N_14147);
or U14323 (N_14323,N_14194,N_14113);
nor U14324 (N_14324,N_14221,N_14230);
and U14325 (N_14325,N_14023,N_14182);
nand U14326 (N_14326,N_14220,N_14155);
xor U14327 (N_14327,N_14031,N_14140);
nor U14328 (N_14328,N_14241,N_14217);
nor U14329 (N_14329,N_14087,N_14135);
nand U14330 (N_14330,N_14239,N_14144);
or U14331 (N_14331,N_14227,N_14092);
nand U14332 (N_14332,N_14225,N_14226);
nand U14333 (N_14333,N_14245,N_14156);
or U14334 (N_14334,N_14057,N_14120);
nor U14335 (N_14335,N_14190,N_14036);
xor U14336 (N_14336,N_14129,N_14008);
and U14337 (N_14337,N_14115,N_14125);
nand U14338 (N_14338,N_14143,N_14111);
and U14339 (N_14339,N_14074,N_14247);
nor U14340 (N_14340,N_14076,N_14231);
or U14341 (N_14341,N_14048,N_14024);
and U14342 (N_14342,N_14203,N_14062);
or U14343 (N_14343,N_14077,N_14151);
xnor U14344 (N_14344,N_14149,N_14112);
nand U14345 (N_14345,N_14046,N_14197);
or U14346 (N_14346,N_14109,N_14196);
or U14347 (N_14347,N_14122,N_14128);
nor U14348 (N_14348,N_14121,N_14030);
nor U14349 (N_14349,N_14029,N_14136);
nand U14350 (N_14350,N_14064,N_14108);
or U14351 (N_14351,N_14102,N_14248);
xnor U14352 (N_14352,N_14079,N_14089);
and U14353 (N_14353,N_14211,N_14070);
nor U14354 (N_14354,N_14025,N_14078);
nand U14355 (N_14355,N_14015,N_14199);
and U14356 (N_14356,N_14193,N_14085);
and U14357 (N_14357,N_14061,N_14126);
nand U14358 (N_14358,N_14242,N_14146);
or U14359 (N_14359,N_14107,N_14162);
and U14360 (N_14360,N_14099,N_14191);
nor U14361 (N_14361,N_14098,N_14244);
nand U14362 (N_14362,N_14001,N_14003);
nand U14363 (N_14363,N_14215,N_14163);
nand U14364 (N_14364,N_14010,N_14222);
xor U14365 (N_14365,N_14004,N_14014);
or U14366 (N_14366,N_14012,N_14168);
nor U14367 (N_14367,N_14219,N_14094);
nand U14368 (N_14368,N_14238,N_14022);
and U14369 (N_14369,N_14080,N_14157);
or U14370 (N_14370,N_14236,N_14186);
nand U14371 (N_14371,N_14202,N_14124);
or U14372 (N_14372,N_14042,N_14172);
nor U14373 (N_14373,N_14175,N_14020);
nor U14374 (N_14374,N_14032,N_14075);
xnor U14375 (N_14375,N_14238,N_14208);
and U14376 (N_14376,N_14112,N_14168);
xnor U14377 (N_14377,N_14206,N_14073);
nor U14378 (N_14378,N_14079,N_14080);
and U14379 (N_14379,N_14160,N_14080);
xnor U14380 (N_14380,N_14085,N_14080);
and U14381 (N_14381,N_14062,N_14208);
or U14382 (N_14382,N_14213,N_14076);
nand U14383 (N_14383,N_14193,N_14240);
or U14384 (N_14384,N_14193,N_14044);
xnor U14385 (N_14385,N_14000,N_14138);
or U14386 (N_14386,N_14180,N_14167);
nor U14387 (N_14387,N_14055,N_14228);
nand U14388 (N_14388,N_14156,N_14011);
and U14389 (N_14389,N_14058,N_14003);
nor U14390 (N_14390,N_14241,N_14235);
xnor U14391 (N_14391,N_14220,N_14128);
or U14392 (N_14392,N_14170,N_14130);
and U14393 (N_14393,N_14182,N_14081);
xor U14394 (N_14394,N_14060,N_14006);
and U14395 (N_14395,N_14216,N_14110);
nand U14396 (N_14396,N_14065,N_14247);
xor U14397 (N_14397,N_14192,N_14219);
xnor U14398 (N_14398,N_14143,N_14060);
or U14399 (N_14399,N_14061,N_14085);
or U14400 (N_14400,N_14209,N_14082);
xnor U14401 (N_14401,N_14139,N_14148);
and U14402 (N_14402,N_14046,N_14069);
nor U14403 (N_14403,N_14025,N_14136);
nand U14404 (N_14404,N_14063,N_14091);
xnor U14405 (N_14405,N_14224,N_14245);
nor U14406 (N_14406,N_14006,N_14249);
nor U14407 (N_14407,N_14237,N_14224);
and U14408 (N_14408,N_14013,N_14202);
and U14409 (N_14409,N_14193,N_14088);
nor U14410 (N_14410,N_14057,N_14180);
nor U14411 (N_14411,N_14010,N_14042);
nand U14412 (N_14412,N_14095,N_14235);
nor U14413 (N_14413,N_14205,N_14103);
and U14414 (N_14414,N_14003,N_14047);
xnor U14415 (N_14415,N_14121,N_14202);
nor U14416 (N_14416,N_14184,N_14109);
nand U14417 (N_14417,N_14096,N_14241);
xor U14418 (N_14418,N_14211,N_14230);
nor U14419 (N_14419,N_14193,N_14076);
or U14420 (N_14420,N_14143,N_14119);
and U14421 (N_14421,N_14074,N_14219);
nand U14422 (N_14422,N_14233,N_14078);
and U14423 (N_14423,N_14050,N_14060);
or U14424 (N_14424,N_14194,N_14205);
and U14425 (N_14425,N_14070,N_14134);
or U14426 (N_14426,N_14057,N_14106);
and U14427 (N_14427,N_14041,N_14141);
or U14428 (N_14428,N_14200,N_14073);
nand U14429 (N_14429,N_14040,N_14029);
nor U14430 (N_14430,N_14223,N_14244);
nor U14431 (N_14431,N_14074,N_14021);
or U14432 (N_14432,N_14034,N_14142);
nand U14433 (N_14433,N_14224,N_14222);
and U14434 (N_14434,N_14168,N_14095);
nor U14435 (N_14435,N_14212,N_14042);
nor U14436 (N_14436,N_14233,N_14014);
or U14437 (N_14437,N_14135,N_14223);
or U14438 (N_14438,N_14128,N_14222);
and U14439 (N_14439,N_14128,N_14219);
nand U14440 (N_14440,N_14161,N_14081);
xor U14441 (N_14441,N_14057,N_14188);
and U14442 (N_14442,N_14025,N_14037);
and U14443 (N_14443,N_14117,N_14247);
nor U14444 (N_14444,N_14174,N_14124);
and U14445 (N_14445,N_14081,N_14197);
nor U14446 (N_14446,N_14194,N_14033);
and U14447 (N_14447,N_14220,N_14101);
xor U14448 (N_14448,N_14082,N_14064);
or U14449 (N_14449,N_14004,N_14180);
xor U14450 (N_14450,N_14210,N_14123);
xor U14451 (N_14451,N_14185,N_14032);
xor U14452 (N_14452,N_14070,N_14239);
xor U14453 (N_14453,N_14095,N_14017);
or U14454 (N_14454,N_14180,N_14220);
and U14455 (N_14455,N_14162,N_14080);
or U14456 (N_14456,N_14210,N_14038);
or U14457 (N_14457,N_14201,N_14082);
xor U14458 (N_14458,N_14240,N_14006);
and U14459 (N_14459,N_14184,N_14143);
xnor U14460 (N_14460,N_14034,N_14088);
nand U14461 (N_14461,N_14076,N_14012);
xnor U14462 (N_14462,N_14240,N_14072);
nand U14463 (N_14463,N_14235,N_14229);
xor U14464 (N_14464,N_14095,N_14090);
nand U14465 (N_14465,N_14203,N_14065);
nand U14466 (N_14466,N_14147,N_14074);
xnor U14467 (N_14467,N_14213,N_14209);
and U14468 (N_14468,N_14235,N_14002);
nor U14469 (N_14469,N_14249,N_14219);
or U14470 (N_14470,N_14054,N_14105);
xnor U14471 (N_14471,N_14194,N_14061);
and U14472 (N_14472,N_14002,N_14093);
nor U14473 (N_14473,N_14200,N_14097);
nor U14474 (N_14474,N_14046,N_14144);
nand U14475 (N_14475,N_14072,N_14025);
nor U14476 (N_14476,N_14195,N_14135);
xor U14477 (N_14477,N_14111,N_14177);
or U14478 (N_14478,N_14192,N_14204);
or U14479 (N_14479,N_14215,N_14232);
or U14480 (N_14480,N_14205,N_14002);
xor U14481 (N_14481,N_14097,N_14226);
or U14482 (N_14482,N_14151,N_14136);
or U14483 (N_14483,N_14165,N_14234);
and U14484 (N_14484,N_14165,N_14220);
and U14485 (N_14485,N_14061,N_14009);
and U14486 (N_14486,N_14004,N_14231);
or U14487 (N_14487,N_14180,N_14037);
nand U14488 (N_14488,N_14217,N_14222);
and U14489 (N_14489,N_14235,N_14075);
or U14490 (N_14490,N_14121,N_14113);
nand U14491 (N_14491,N_14085,N_14083);
xor U14492 (N_14492,N_14130,N_14057);
nor U14493 (N_14493,N_14112,N_14142);
xnor U14494 (N_14494,N_14055,N_14103);
nor U14495 (N_14495,N_14167,N_14237);
xnor U14496 (N_14496,N_14104,N_14105);
and U14497 (N_14497,N_14190,N_14196);
nand U14498 (N_14498,N_14004,N_14162);
and U14499 (N_14499,N_14195,N_14042);
xor U14500 (N_14500,N_14449,N_14450);
and U14501 (N_14501,N_14478,N_14255);
xor U14502 (N_14502,N_14258,N_14432);
and U14503 (N_14503,N_14490,N_14347);
xor U14504 (N_14504,N_14320,N_14497);
nor U14505 (N_14505,N_14305,N_14386);
nand U14506 (N_14506,N_14250,N_14302);
xor U14507 (N_14507,N_14273,N_14346);
or U14508 (N_14508,N_14408,N_14259);
xnor U14509 (N_14509,N_14392,N_14394);
nand U14510 (N_14510,N_14393,N_14485);
nor U14511 (N_14511,N_14266,N_14414);
nor U14512 (N_14512,N_14480,N_14253);
and U14513 (N_14513,N_14377,N_14365);
nand U14514 (N_14514,N_14401,N_14470);
xnor U14515 (N_14515,N_14256,N_14438);
xor U14516 (N_14516,N_14395,N_14337);
or U14517 (N_14517,N_14447,N_14477);
nor U14518 (N_14518,N_14442,N_14415);
xnor U14519 (N_14519,N_14344,N_14464);
xnor U14520 (N_14520,N_14328,N_14466);
and U14521 (N_14521,N_14371,N_14335);
or U14522 (N_14522,N_14251,N_14267);
nor U14523 (N_14523,N_14323,N_14360);
or U14524 (N_14524,N_14455,N_14318);
and U14525 (N_14525,N_14358,N_14304);
nor U14526 (N_14526,N_14364,N_14303);
nand U14527 (N_14527,N_14291,N_14434);
or U14528 (N_14528,N_14383,N_14276);
or U14529 (N_14529,N_14441,N_14451);
or U14530 (N_14530,N_14370,N_14325);
xnor U14531 (N_14531,N_14299,N_14496);
or U14532 (N_14532,N_14468,N_14287);
nor U14533 (N_14533,N_14473,N_14483);
nand U14534 (N_14534,N_14489,N_14257);
or U14535 (N_14535,N_14345,N_14396);
nand U14536 (N_14536,N_14301,N_14278);
xor U14537 (N_14537,N_14421,N_14437);
nand U14538 (N_14538,N_14382,N_14474);
nand U14539 (N_14539,N_14486,N_14352);
xor U14540 (N_14540,N_14491,N_14279);
nor U14541 (N_14541,N_14322,N_14402);
or U14542 (N_14542,N_14487,N_14356);
xor U14543 (N_14543,N_14385,N_14271);
or U14544 (N_14544,N_14330,N_14416);
and U14545 (N_14545,N_14495,N_14397);
or U14546 (N_14546,N_14380,N_14307);
or U14547 (N_14547,N_14390,N_14350);
nand U14548 (N_14548,N_14313,N_14265);
nor U14549 (N_14549,N_14406,N_14341);
nand U14550 (N_14550,N_14428,N_14332);
xor U14551 (N_14551,N_14445,N_14321);
nor U14552 (N_14552,N_14298,N_14420);
or U14553 (N_14553,N_14275,N_14462);
and U14554 (N_14554,N_14481,N_14423);
nand U14555 (N_14555,N_14270,N_14324);
and U14556 (N_14556,N_14425,N_14381);
nor U14557 (N_14557,N_14499,N_14319);
nor U14558 (N_14558,N_14262,N_14461);
or U14559 (N_14559,N_14430,N_14436);
xor U14560 (N_14560,N_14398,N_14351);
or U14561 (N_14561,N_14443,N_14424);
or U14562 (N_14562,N_14277,N_14280);
or U14563 (N_14563,N_14281,N_14479);
xnor U14564 (N_14564,N_14403,N_14407);
nor U14565 (N_14565,N_14329,N_14471);
xor U14566 (N_14566,N_14435,N_14254);
nor U14567 (N_14567,N_14463,N_14426);
nand U14568 (N_14568,N_14467,N_14340);
and U14569 (N_14569,N_14409,N_14327);
nand U14570 (N_14570,N_14376,N_14469);
or U14571 (N_14571,N_14348,N_14452);
xor U14572 (N_14572,N_14317,N_14284);
xor U14573 (N_14573,N_14498,N_14458);
and U14574 (N_14574,N_14404,N_14283);
nor U14575 (N_14575,N_14431,N_14412);
nor U14576 (N_14576,N_14448,N_14286);
nor U14577 (N_14577,N_14342,N_14482);
and U14578 (N_14578,N_14269,N_14295);
xnor U14579 (N_14579,N_14343,N_14354);
nand U14580 (N_14580,N_14369,N_14260);
nand U14581 (N_14581,N_14410,N_14338);
and U14582 (N_14582,N_14296,N_14353);
nor U14583 (N_14583,N_14336,N_14388);
nor U14584 (N_14584,N_14413,N_14440);
nor U14585 (N_14585,N_14312,N_14493);
nand U14586 (N_14586,N_14460,N_14368);
nor U14587 (N_14587,N_14268,N_14288);
nor U14588 (N_14588,N_14429,N_14306);
and U14589 (N_14589,N_14494,N_14282);
xor U14590 (N_14590,N_14405,N_14290);
nor U14591 (N_14591,N_14285,N_14422);
and U14592 (N_14592,N_14375,N_14439);
xor U14593 (N_14593,N_14293,N_14310);
nand U14594 (N_14594,N_14339,N_14387);
or U14595 (N_14595,N_14349,N_14309);
xor U14596 (N_14596,N_14400,N_14457);
nand U14597 (N_14597,N_14378,N_14361);
nand U14598 (N_14598,N_14316,N_14297);
nand U14599 (N_14599,N_14379,N_14488);
and U14600 (N_14600,N_14372,N_14472);
xor U14601 (N_14601,N_14331,N_14475);
nand U14602 (N_14602,N_14476,N_14465);
nand U14603 (N_14603,N_14384,N_14300);
nor U14604 (N_14604,N_14446,N_14334);
and U14605 (N_14605,N_14444,N_14459);
nand U14606 (N_14606,N_14374,N_14264);
nor U14607 (N_14607,N_14308,N_14355);
or U14608 (N_14608,N_14389,N_14492);
and U14609 (N_14609,N_14261,N_14453);
and U14610 (N_14610,N_14272,N_14289);
xor U14611 (N_14611,N_14411,N_14433);
and U14612 (N_14612,N_14357,N_14359);
and U14613 (N_14613,N_14427,N_14315);
xnor U14614 (N_14614,N_14417,N_14399);
xnor U14615 (N_14615,N_14252,N_14454);
and U14616 (N_14616,N_14484,N_14419);
and U14617 (N_14617,N_14292,N_14311);
xor U14618 (N_14618,N_14274,N_14363);
and U14619 (N_14619,N_14333,N_14456);
nand U14620 (N_14620,N_14362,N_14373);
xnor U14621 (N_14621,N_14391,N_14418);
xor U14622 (N_14622,N_14263,N_14366);
xor U14623 (N_14623,N_14326,N_14367);
nor U14624 (N_14624,N_14294,N_14314);
nand U14625 (N_14625,N_14486,N_14396);
nand U14626 (N_14626,N_14478,N_14289);
nor U14627 (N_14627,N_14474,N_14442);
or U14628 (N_14628,N_14364,N_14417);
xnor U14629 (N_14629,N_14459,N_14318);
or U14630 (N_14630,N_14382,N_14475);
and U14631 (N_14631,N_14389,N_14306);
or U14632 (N_14632,N_14383,N_14346);
nand U14633 (N_14633,N_14364,N_14429);
xor U14634 (N_14634,N_14299,N_14374);
nor U14635 (N_14635,N_14471,N_14395);
xnor U14636 (N_14636,N_14383,N_14426);
nand U14637 (N_14637,N_14296,N_14434);
or U14638 (N_14638,N_14263,N_14418);
or U14639 (N_14639,N_14450,N_14305);
nor U14640 (N_14640,N_14426,N_14297);
xor U14641 (N_14641,N_14434,N_14445);
and U14642 (N_14642,N_14414,N_14310);
and U14643 (N_14643,N_14385,N_14295);
xnor U14644 (N_14644,N_14341,N_14308);
and U14645 (N_14645,N_14281,N_14334);
xnor U14646 (N_14646,N_14294,N_14389);
nand U14647 (N_14647,N_14253,N_14289);
xnor U14648 (N_14648,N_14360,N_14479);
or U14649 (N_14649,N_14296,N_14469);
nor U14650 (N_14650,N_14298,N_14378);
nor U14651 (N_14651,N_14422,N_14278);
xor U14652 (N_14652,N_14404,N_14304);
and U14653 (N_14653,N_14478,N_14417);
xnor U14654 (N_14654,N_14324,N_14281);
or U14655 (N_14655,N_14406,N_14480);
nor U14656 (N_14656,N_14258,N_14479);
and U14657 (N_14657,N_14492,N_14254);
and U14658 (N_14658,N_14416,N_14353);
nand U14659 (N_14659,N_14376,N_14299);
nand U14660 (N_14660,N_14474,N_14310);
xnor U14661 (N_14661,N_14474,N_14390);
nor U14662 (N_14662,N_14271,N_14458);
xor U14663 (N_14663,N_14476,N_14357);
and U14664 (N_14664,N_14448,N_14427);
nand U14665 (N_14665,N_14431,N_14329);
xor U14666 (N_14666,N_14257,N_14431);
or U14667 (N_14667,N_14467,N_14464);
xnor U14668 (N_14668,N_14351,N_14438);
xnor U14669 (N_14669,N_14251,N_14335);
nor U14670 (N_14670,N_14396,N_14388);
or U14671 (N_14671,N_14479,N_14465);
xor U14672 (N_14672,N_14319,N_14431);
xnor U14673 (N_14673,N_14360,N_14325);
or U14674 (N_14674,N_14436,N_14317);
xnor U14675 (N_14675,N_14289,N_14420);
xor U14676 (N_14676,N_14424,N_14445);
and U14677 (N_14677,N_14277,N_14267);
nand U14678 (N_14678,N_14273,N_14481);
or U14679 (N_14679,N_14431,N_14327);
nor U14680 (N_14680,N_14416,N_14363);
nor U14681 (N_14681,N_14489,N_14425);
and U14682 (N_14682,N_14308,N_14325);
or U14683 (N_14683,N_14370,N_14465);
or U14684 (N_14684,N_14448,N_14260);
and U14685 (N_14685,N_14383,N_14385);
nand U14686 (N_14686,N_14438,N_14315);
or U14687 (N_14687,N_14361,N_14392);
nor U14688 (N_14688,N_14467,N_14292);
nor U14689 (N_14689,N_14491,N_14429);
or U14690 (N_14690,N_14355,N_14474);
nand U14691 (N_14691,N_14337,N_14261);
nand U14692 (N_14692,N_14256,N_14287);
xor U14693 (N_14693,N_14258,N_14273);
xor U14694 (N_14694,N_14426,N_14260);
nand U14695 (N_14695,N_14383,N_14387);
xor U14696 (N_14696,N_14454,N_14259);
or U14697 (N_14697,N_14402,N_14467);
or U14698 (N_14698,N_14499,N_14255);
nor U14699 (N_14699,N_14398,N_14328);
and U14700 (N_14700,N_14256,N_14384);
and U14701 (N_14701,N_14316,N_14398);
nor U14702 (N_14702,N_14386,N_14400);
xnor U14703 (N_14703,N_14370,N_14404);
or U14704 (N_14704,N_14252,N_14353);
or U14705 (N_14705,N_14326,N_14417);
nor U14706 (N_14706,N_14273,N_14447);
xor U14707 (N_14707,N_14348,N_14350);
nor U14708 (N_14708,N_14278,N_14465);
and U14709 (N_14709,N_14371,N_14394);
xor U14710 (N_14710,N_14341,N_14496);
nor U14711 (N_14711,N_14430,N_14251);
xor U14712 (N_14712,N_14409,N_14471);
nor U14713 (N_14713,N_14465,N_14380);
xnor U14714 (N_14714,N_14497,N_14308);
or U14715 (N_14715,N_14465,N_14301);
nand U14716 (N_14716,N_14462,N_14395);
and U14717 (N_14717,N_14384,N_14332);
nand U14718 (N_14718,N_14383,N_14484);
and U14719 (N_14719,N_14405,N_14426);
or U14720 (N_14720,N_14311,N_14369);
xor U14721 (N_14721,N_14353,N_14264);
or U14722 (N_14722,N_14386,N_14253);
nand U14723 (N_14723,N_14298,N_14387);
or U14724 (N_14724,N_14475,N_14371);
or U14725 (N_14725,N_14406,N_14440);
xor U14726 (N_14726,N_14369,N_14479);
xnor U14727 (N_14727,N_14461,N_14390);
or U14728 (N_14728,N_14293,N_14332);
and U14729 (N_14729,N_14467,N_14371);
nor U14730 (N_14730,N_14433,N_14379);
and U14731 (N_14731,N_14292,N_14273);
or U14732 (N_14732,N_14409,N_14312);
nor U14733 (N_14733,N_14272,N_14391);
or U14734 (N_14734,N_14336,N_14476);
nor U14735 (N_14735,N_14454,N_14446);
or U14736 (N_14736,N_14330,N_14479);
nor U14737 (N_14737,N_14333,N_14428);
and U14738 (N_14738,N_14428,N_14406);
nor U14739 (N_14739,N_14310,N_14326);
and U14740 (N_14740,N_14251,N_14498);
xor U14741 (N_14741,N_14381,N_14360);
xnor U14742 (N_14742,N_14430,N_14388);
nand U14743 (N_14743,N_14279,N_14314);
or U14744 (N_14744,N_14306,N_14367);
nor U14745 (N_14745,N_14433,N_14259);
or U14746 (N_14746,N_14330,N_14398);
xor U14747 (N_14747,N_14359,N_14429);
nand U14748 (N_14748,N_14416,N_14497);
xor U14749 (N_14749,N_14314,N_14432);
nor U14750 (N_14750,N_14627,N_14530);
xor U14751 (N_14751,N_14566,N_14719);
nand U14752 (N_14752,N_14541,N_14655);
nor U14753 (N_14753,N_14732,N_14722);
and U14754 (N_14754,N_14502,N_14569);
nand U14755 (N_14755,N_14677,N_14638);
nand U14756 (N_14756,N_14727,N_14728);
or U14757 (N_14757,N_14580,N_14549);
or U14758 (N_14758,N_14675,N_14529);
nand U14759 (N_14759,N_14747,N_14699);
and U14760 (N_14760,N_14698,N_14640);
or U14761 (N_14761,N_14508,N_14644);
nor U14762 (N_14762,N_14511,N_14577);
or U14763 (N_14763,N_14739,N_14731);
and U14764 (N_14764,N_14510,N_14573);
or U14765 (N_14765,N_14626,N_14715);
or U14766 (N_14766,N_14558,N_14632);
and U14767 (N_14767,N_14590,N_14745);
nor U14768 (N_14768,N_14528,N_14743);
nor U14769 (N_14769,N_14654,N_14714);
nor U14770 (N_14770,N_14726,N_14616);
or U14771 (N_14771,N_14648,N_14552);
and U14772 (N_14772,N_14553,N_14684);
nor U14773 (N_14773,N_14595,N_14519);
and U14774 (N_14774,N_14597,N_14668);
and U14775 (N_14775,N_14706,N_14562);
xnor U14776 (N_14776,N_14564,N_14701);
xor U14777 (N_14777,N_14544,N_14693);
and U14778 (N_14778,N_14666,N_14617);
or U14779 (N_14779,N_14734,N_14618);
or U14780 (N_14780,N_14650,N_14662);
or U14781 (N_14781,N_14665,N_14568);
xor U14782 (N_14782,N_14517,N_14691);
nor U14783 (N_14783,N_14619,N_14692);
xnor U14784 (N_14784,N_14651,N_14628);
nand U14785 (N_14785,N_14740,N_14574);
or U14786 (N_14786,N_14554,N_14524);
xor U14787 (N_14787,N_14697,N_14533);
nor U14788 (N_14788,N_14579,N_14563);
xnor U14789 (N_14789,N_14717,N_14676);
or U14790 (N_14790,N_14718,N_14713);
or U14791 (N_14791,N_14642,N_14503);
nor U14792 (N_14792,N_14601,N_14685);
nand U14793 (N_14793,N_14531,N_14730);
nand U14794 (N_14794,N_14622,N_14578);
xor U14795 (N_14795,N_14526,N_14672);
nand U14796 (N_14796,N_14705,N_14545);
nor U14797 (N_14797,N_14615,N_14603);
nand U14798 (N_14798,N_14532,N_14561);
nor U14799 (N_14799,N_14636,N_14741);
or U14800 (N_14800,N_14744,N_14604);
nand U14801 (N_14801,N_14647,N_14535);
or U14802 (N_14802,N_14605,N_14634);
nor U14803 (N_14803,N_14682,N_14559);
and U14804 (N_14804,N_14501,N_14625);
or U14805 (N_14805,N_14702,N_14661);
or U14806 (N_14806,N_14724,N_14704);
and U14807 (N_14807,N_14641,N_14639);
and U14808 (N_14808,N_14523,N_14610);
nand U14809 (N_14809,N_14594,N_14570);
and U14810 (N_14810,N_14703,N_14657);
and U14811 (N_14811,N_14635,N_14643);
or U14812 (N_14812,N_14613,N_14707);
nor U14813 (N_14813,N_14737,N_14509);
and U14814 (N_14814,N_14583,N_14671);
nand U14815 (N_14815,N_14630,N_14560);
nand U14816 (N_14816,N_14736,N_14599);
or U14817 (N_14817,N_14542,N_14735);
xor U14818 (N_14818,N_14556,N_14738);
and U14819 (N_14819,N_14712,N_14688);
or U14820 (N_14820,N_14695,N_14709);
nand U14821 (N_14821,N_14725,N_14637);
nand U14822 (N_14822,N_14652,N_14507);
xor U14823 (N_14823,N_14521,N_14557);
or U14824 (N_14824,N_14729,N_14572);
xor U14825 (N_14825,N_14538,N_14518);
or U14826 (N_14826,N_14674,N_14721);
nand U14827 (N_14827,N_14664,N_14505);
and U14828 (N_14828,N_14606,N_14582);
nand U14829 (N_14829,N_14525,N_14546);
or U14830 (N_14830,N_14659,N_14504);
xor U14831 (N_14831,N_14621,N_14588);
nor U14832 (N_14832,N_14587,N_14608);
or U14833 (N_14833,N_14686,N_14749);
or U14834 (N_14834,N_14711,N_14527);
xor U14835 (N_14835,N_14516,N_14536);
or U14836 (N_14836,N_14585,N_14584);
xor U14837 (N_14837,N_14681,N_14515);
nand U14838 (N_14838,N_14612,N_14689);
nand U14839 (N_14839,N_14567,N_14576);
nor U14840 (N_14840,N_14673,N_14540);
xor U14841 (N_14841,N_14512,N_14669);
xor U14842 (N_14842,N_14624,N_14522);
or U14843 (N_14843,N_14633,N_14680);
or U14844 (N_14844,N_14551,N_14649);
and U14845 (N_14845,N_14733,N_14539);
and U14846 (N_14846,N_14700,N_14710);
nand U14847 (N_14847,N_14645,N_14547);
nand U14848 (N_14848,N_14683,N_14629);
or U14849 (N_14849,N_14678,N_14581);
nor U14850 (N_14850,N_14742,N_14658);
and U14851 (N_14851,N_14550,N_14555);
nand U14852 (N_14852,N_14600,N_14506);
and U14853 (N_14853,N_14646,N_14667);
nand U14854 (N_14854,N_14598,N_14571);
or U14855 (N_14855,N_14609,N_14670);
xnor U14856 (N_14856,N_14602,N_14534);
nand U14857 (N_14857,N_14679,N_14514);
nand U14858 (N_14858,N_14513,N_14720);
nand U14859 (N_14859,N_14543,N_14591);
and U14860 (N_14860,N_14537,N_14589);
nor U14861 (N_14861,N_14656,N_14520);
and U14862 (N_14862,N_14620,N_14690);
and U14863 (N_14863,N_14592,N_14586);
and U14864 (N_14864,N_14623,N_14653);
nand U14865 (N_14865,N_14660,N_14548);
or U14866 (N_14866,N_14593,N_14716);
nor U14867 (N_14867,N_14575,N_14746);
nand U14868 (N_14868,N_14694,N_14687);
nand U14869 (N_14869,N_14611,N_14614);
nor U14870 (N_14870,N_14500,N_14565);
and U14871 (N_14871,N_14748,N_14696);
and U14872 (N_14872,N_14631,N_14663);
and U14873 (N_14873,N_14596,N_14607);
and U14874 (N_14874,N_14723,N_14708);
xor U14875 (N_14875,N_14550,N_14520);
nor U14876 (N_14876,N_14636,N_14562);
nor U14877 (N_14877,N_14660,N_14626);
xnor U14878 (N_14878,N_14545,N_14647);
and U14879 (N_14879,N_14524,N_14630);
or U14880 (N_14880,N_14679,N_14727);
xnor U14881 (N_14881,N_14547,N_14630);
or U14882 (N_14882,N_14513,N_14609);
or U14883 (N_14883,N_14506,N_14640);
nor U14884 (N_14884,N_14551,N_14662);
xor U14885 (N_14885,N_14599,N_14659);
xor U14886 (N_14886,N_14577,N_14571);
and U14887 (N_14887,N_14602,N_14682);
and U14888 (N_14888,N_14608,N_14511);
xnor U14889 (N_14889,N_14618,N_14624);
nand U14890 (N_14890,N_14607,N_14694);
nand U14891 (N_14891,N_14581,N_14698);
and U14892 (N_14892,N_14746,N_14576);
nand U14893 (N_14893,N_14743,N_14657);
xor U14894 (N_14894,N_14598,N_14520);
or U14895 (N_14895,N_14546,N_14520);
nor U14896 (N_14896,N_14560,N_14545);
or U14897 (N_14897,N_14583,N_14736);
nor U14898 (N_14898,N_14722,N_14746);
and U14899 (N_14899,N_14531,N_14549);
or U14900 (N_14900,N_14602,N_14729);
nand U14901 (N_14901,N_14610,N_14637);
nor U14902 (N_14902,N_14682,N_14614);
nor U14903 (N_14903,N_14725,N_14671);
and U14904 (N_14904,N_14576,N_14549);
xor U14905 (N_14905,N_14517,N_14613);
xnor U14906 (N_14906,N_14543,N_14660);
nor U14907 (N_14907,N_14504,N_14731);
or U14908 (N_14908,N_14663,N_14655);
nor U14909 (N_14909,N_14664,N_14590);
xor U14910 (N_14910,N_14667,N_14607);
xnor U14911 (N_14911,N_14539,N_14663);
nand U14912 (N_14912,N_14719,N_14523);
xnor U14913 (N_14913,N_14509,N_14603);
xor U14914 (N_14914,N_14525,N_14748);
and U14915 (N_14915,N_14671,N_14741);
nor U14916 (N_14916,N_14719,N_14571);
nand U14917 (N_14917,N_14730,N_14587);
nand U14918 (N_14918,N_14611,N_14612);
xnor U14919 (N_14919,N_14664,N_14719);
nor U14920 (N_14920,N_14575,N_14517);
xnor U14921 (N_14921,N_14542,N_14580);
nor U14922 (N_14922,N_14699,N_14711);
nand U14923 (N_14923,N_14636,N_14638);
nor U14924 (N_14924,N_14622,N_14539);
or U14925 (N_14925,N_14713,N_14740);
xor U14926 (N_14926,N_14617,N_14720);
nand U14927 (N_14927,N_14701,N_14561);
xnor U14928 (N_14928,N_14618,N_14738);
xnor U14929 (N_14929,N_14687,N_14743);
nor U14930 (N_14930,N_14520,N_14631);
nand U14931 (N_14931,N_14517,N_14726);
nor U14932 (N_14932,N_14503,N_14641);
and U14933 (N_14933,N_14651,N_14674);
or U14934 (N_14934,N_14617,N_14676);
nand U14935 (N_14935,N_14571,N_14521);
nor U14936 (N_14936,N_14567,N_14554);
nor U14937 (N_14937,N_14737,N_14522);
and U14938 (N_14938,N_14650,N_14694);
nor U14939 (N_14939,N_14617,N_14519);
nor U14940 (N_14940,N_14701,N_14601);
or U14941 (N_14941,N_14516,N_14570);
and U14942 (N_14942,N_14619,N_14588);
xor U14943 (N_14943,N_14501,N_14561);
xor U14944 (N_14944,N_14664,N_14730);
xor U14945 (N_14945,N_14700,N_14713);
xnor U14946 (N_14946,N_14584,N_14748);
or U14947 (N_14947,N_14671,N_14717);
and U14948 (N_14948,N_14565,N_14646);
and U14949 (N_14949,N_14700,N_14590);
nand U14950 (N_14950,N_14715,N_14644);
and U14951 (N_14951,N_14567,N_14701);
or U14952 (N_14952,N_14675,N_14650);
xor U14953 (N_14953,N_14576,N_14623);
and U14954 (N_14954,N_14724,N_14682);
nand U14955 (N_14955,N_14503,N_14724);
and U14956 (N_14956,N_14651,N_14659);
nand U14957 (N_14957,N_14734,N_14575);
xor U14958 (N_14958,N_14608,N_14747);
and U14959 (N_14959,N_14501,N_14516);
nor U14960 (N_14960,N_14636,N_14666);
nor U14961 (N_14961,N_14606,N_14621);
or U14962 (N_14962,N_14720,N_14645);
nand U14963 (N_14963,N_14520,N_14624);
or U14964 (N_14964,N_14689,N_14555);
xor U14965 (N_14965,N_14707,N_14654);
xnor U14966 (N_14966,N_14686,N_14502);
nor U14967 (N_14967,N_14643,N_14705);
nor U14968 (N_14968,N_14620,N_14665);
and U14969 (N_14969,N_14702,N_14743);
xnor U14970 (N_14970,N_14627,N_14616);
xnor U14971 (N_14971,N_14741,N_14720);
nor U14972 (N_14972,N_14732,N_14704);
and U14973 (N_14973,N_14696,N_14669);
xnor U14974 (N_14974,N_14560,N_14672);
xnor U14975 (N_14975,N_14587,N_14678);
and U14976 (N_14976,N_14554,N_14507);
or U14977 (N_14977,N_14672,N_14513);
or U14978 (N_14978,N_14719,N_14715);
or U14979 (N_14979,N_14685,N_14543);
xor U14980 (N_14980,N_14627,N_14658);
nor U14981 (N_14981,N_14728,N_14610);
nand U14982 (N_14982,N_14733,N_14681);
nor U14983 (N_14983,N_14564,N_14571);
xor U14984 (N_14984,N_14647,N_14724);
nand U14985 (N_14985,N_14644,N_14503);
and U14986 (N_14986,N_14527,N_14734);
and U14987 (N_14987,N_14560,N_14503);
or U14988 (N_14988,N_14582,N_14526);
nand U14989 (N_14989,N_14566,N_14744);
xnor U14990 (N_14990,N_14712,N_14617);
and U14991 (N_14991,N_14625,N_14525);
nor U14992 (N_14992,N_14730,N_14613);
nand U14993 (N_14993,N_14641,N_14584);
xor U14994 (N_14994,N_14500,N_14665);
and U14995 (N_14995,N_14638,N_14646);
or U14996 (N_14996,N_14527,N_14528);
and U14997 (N_14997,N_14679,N_14613);
or U14998 (N_14998,N_14651,N_14720);
xor U14999 (N_14999,N_14610,N_14709);
and U15000 (N_15000,N_14822,N_14756);
or U15001 (N_15001,N_14863,N_14800);
and U15002 (N_15002,N_14777,N_14834);
or U15003 (N_15003,N_14956,N_14793);
nor U15004 (N_15004,N_14960,N_14908);
nor U15005 (N_15005,N_14957,N_14818);
xnor U15006 (N_15006,N_14986,N_14928);
and U15007 (N_15007,N_14854,N_14764);
xor U15008 (N_15008,N_14811,N_14836);
and U15009 (N_15009,N_14761,N_14974);
nand U15010 (N_15010,N_14906,N_14867);
xnor U15011 (N_15011,N_14920,N_14897);
xnor U15012 (N_15012,N_14843,N_14758);
nor U15013 (N_15013,N_14815,N_14765);
xnor U15014 (N_15014,N_14855,N_14992);
nand U15015 (N_15015,N_14808,N_14766);
nand U15016 (N_15016,N_14926,N_14943);
or U15017 (N_15017,N_14880,N_14911);
or U15018 (N_15018,N_14768,N_14819);
nor U15019 (N_15019,N_14866,N_14796);
nand U15020 (N_15020,N_14752,N_14963);
or U15021 (N_15021,N_14892,N_14902);
xor U15022 (N_15022,N_14895,N_14791);
xnor U15023 (N_15023,N_14924,N_14944);
nand U15024 (N_15024,N_14996,N_14751);
and U15025 (N_15025,N_14998,N_14827);
nor U15026 (N_15026,N_14794,N_14910);
xor U15027 (N_15027,N_14885,N_14878);
nand U15028 (N_15028,N_14987,N_14909);
nor U15029 (N_15029,N_14929,N_14890);
and U15030 (N_15030,N_14889,N_14925);
nand U15031 (N_15031,N_14989,N_14813);
or U15032 (N_15032,N_14918,N_14784);
nor U15033 (N_15033,N_14828,N_14894);
and U15034 (N_15034,N_14806,N_14829);
and U15035 (N_15035,N_14973,N_14961);
or U15036 (N_15036,N_14759,N_14770);
xnor U15037 (N_15037,N_14869,N_14830);
nand U15038 (N_15038,N_14899,N_14883);
nor U15039 (N_15039,N_14955,N_14976);
nor U15040 (N_15040,N_14879,N_14984);
or U15041 (N_15041,N_14873,N_14862);
or U15042 (N_15042,N_14914,N_14875);
nand U15043 (N_15043,N_14958,N_14948);
nand U15044 (N_15044,N_14824,N_14864);
nand U15045 (N_15045,N_14763,N_14849);
or U15046 (N_15046,N_14913,N_14896);
xor U15047 (N_15047,N_14769,N_14851);
nor U15048 (N_15048,N_14951,N_14812);
nand U15049 (N_15049,N_14935,N_14970);
or U15050 (N_15050,N_14884,N_14847);
or U15051 (N_15051,N_14876,N_14850);
or U15052 (N_15052,N_14949,N_14816);
nor U15053 (N_15053,N_14952,N_14916);
nand U15054 (N_15054,N_14977,N_14945);
nor U15055 (N_15055,N_14831,N_14781);
or U15056 (N_15056,N_14814,N_14826);
nor U15057 (N_15057,N_14980,N_14904);
or U15058 (N_15058,N_14965,N_14807);
and U15059 (N_15059,N_14903,N_14979);
or U15060 (N_15060,N_14782,N_14792);
xor U15061 (N_15061,N_14757,N_14972);
xor U15062 (N_15062,N_14857,N_14861);
nand U15063 (N_15063,N_14941,N_14841);
and U15064 (N_15064,N_14981,N_14900);
or U15065 (N_15065,N_14832,N_14838);
nand U15066 (N_15066,N_14882,N_14860);
xor U15067 (N_15067,N_14785,N_14852);
nand U15068 (N_15068,N_14887,N_14778);
or U15069 (N_15069,N_14803,N_14772);
xor U15070 (N_15070,N_14898,N_14936);
and U15071 (N_15071,N_14959,N_14823);
nand U15072 (N_15072,N_14915,N_14912);
and U15073 (N_15073,N_14786,N_14966);
nor U15074 (N_15074,N_14870,N_14804);
nor U15075 (N_15075,N_14990,N_14801);
xor U15076 (N_15076,N_14946,N_14975);
and U15077 (N_15077,N_14771,N_14983);
nand U15078 (N_15078,N_14939,N_14930);
nor U15079 (N_15079,N_14940,N_14954);
nor U15080 (N_15080,N_14937,N_14856);
xor U15081 (N_15081,N_14934,N_14999);
nor U15082 (N_15082,N_14817,N_14888);
or U15083 (N_15083,N_14881,N_14877);
or U15084 (N_15084,N_14762,N_14947);
xor U15085 (N_15085,N_14886,N_14790);
xor U15086 (N_15086,N_14953,N_14893);
or U15087 (N_15087,N_14994,N_14971);
nor U15088 (N_15088,N_14802,N_14773);
nor U15089 (N_15089,N_14798,N_14988);
nor U15090 (N_15090,N_14969,N_14933);
nor U15091 (N_15091,N_14938,N_14907);
or U15092 (N_15092,N_14932,N_14874);
or U15093 (N_15093,N_14821,N_14997);
nor U15094 (N_15094,N_14922,N_14968);
nor U15095 (N_15095,N_14917,N_14775);
and U15096 (N_15096,N_14842,N_14787);
nand U15097 (N_15097,N_14844,N_14995);
nor U15098 (N_15098,N_14753,N_14846);
and U15099 (N_15099,N_14809,N_14927);
and U15100 (N_15100,N_14859,N_14825);
nor U15101 (N_15101,N_14891,N_14840);
xnor U15102 (N_15102,N_14776,N_14799);
nand U15103 (N_15103,N_14779,N_14872);
or U15104 (N_15104,N_14788,N_14978);
xor U15105 (N_15105,N_14962,N_14967);
xor U15106 (N_15106,N_14993,N_14868);
nand U15107 (N_15107,N_14871,N_14805);
or U15108 (N_15108,N_14901,N_14923);
or U15109 (N_15109,N_14905,N_14820);
nand U15110 (N_15110,N_14982,N_14865);
or U15111 (N_15111,N_14837,N_14964);
nor U15112 (N_15112,N_14835,N_14760);
and U15113 (N_15113,N_14797,N_14919);
nor U15114 (N_15114,N_14950,N_14810);
nor U15115 (N_15115,N_14795,N_14833);
nand U15116 (N_15116,N_14991,N_14750);
xnor U15117 (N_15117,N_14985,N_14789);
and U15118 (N_15118,N_14774,N_14942);
nor U15119 (N_15119,N_14853,N_14858);
xor U15120 (N_15120,N_14848,N_14931);
and U15121 (N_15121,N_14780,N_14783);
or U15122 (N_15122,N_14921,N_14839);
xor U15123 (N_15123,N_14845,N_14754);
nand U15124 (N_15124,N_14755,N_14767);
or U15125 (N_15125,N_14916,N_14822);
and U15126 (N_15126,N_14844,N_14903);
or U15127 (N_15127,N_14810,N_14850);
and U15128 (N_15128,N_14991,N_14915);
nor U15129 (N_15129,N_14800,N_14795);
and U15130 (N_15130,N_14912,N_14988);
and U15131 (N_15131,N_14775,N_14909);
nor U15132 (N_15132,N_14946,N_14797);
nand U15133 (N_15133,N_14803,N_14845);
and U15134 (N_15134,N_14945,N_14774);
xnor U15135 (N_15135,N_14923,N_14928);
and U15136 (N_15136,N_14856,N_14867);
and U15137 (N_15137,N_14839,N_14905);
nand U15138 (N_15138,N_14902,N_14755);
and U15139 (N_15139,N_14930,N_14976);
or U15140 (N_15140,N_14751,N_14947);
nor U15141 (N_15141,N_14798,N_14909);
or U15142 (N_15142,N_14797,N_14774);
xnor U15143 (N_15143,N_14759,N_14815);
and U15144 (N_15144,N_14830,N_14818);
nand U15145 (N_15145,N_14755,N_14868);
and U15146 (N_15146,N_14848,N_14975);
or U15147 (N_15147,N_14818,N_14882);
nand U15148 (N_15148,N_14952,N_14785);
and U15149 (N_15149,N_14818,N_14986);
nor U15150 (N_15150,N_14760,N_14927);
xor U15151 (N_15151,N_14781,N_14958);
and U15152 (N_15152,N_14986,N_14808);
nor U15153 (N_15153,N_14923,N_14756);
xnor U15154 (N_15154,N_14933,N_14864);
and U15155 (N_15155,N_14907,N_14751);
or U15156 (N_15156,N_14870,N_14963);
xor U15157 (N_15157,N_14753,N_14821);
or U15158 (N_15158,N_14775,N_14774);
or U15159 (N_15159,N_14797,N_14876);
nor U15160 (N_15160,N_14860,N_14800);
nand U15161 (N_15161,N_14759,N_14844);
or U15162 (N_15162,N_14916,N_14888);
and U15163 (N_15163,N_14950,N_14816);
or U15164 (N_15164,N_14771,N_14793);
nand U15165 (N_15165,N_14877,N_14868);
xnor U15166 (N_15166,N_14846,N_14848);
nand U15167 (N_15167,N_14991,N_14879);
xor U15168 (N_15168,N_14853,N_14757);
nand U15169 (N_15169,N_14796,N_14798);
or U15170 (N_15170,N_14914,N_14794);
nand U15171 (N_15171,N_14942,N_14892);
nor U15172 (N_15172,N_14845,N_14944);
nand U15173 (N_15173,N_14838,N_14836);
xor U15174 (N_15174,N_14868,N_14974);
and U15175 (N_15175,N_14813,N_14889);
and U15176 (N_15176,N_14869,N_14808);
or U15177 (N_15177,N_14926,N_14990);
nor U15178 (N_15178,N_14798,N_14980);
nand U15179 (N_15179,N_14750,N_14752);
and U15180 (N_15180,N_14991,N_14969);
nand U15181 (N_15181,N_14995,N_14778);
nor U15182 (N_15182,N_14874,N_14813);
nand U15183 (N_15183,N_14789,N_14923);
nor U15184 (N_15184,N_14990,N_14829);
nor U15185 (N_15185,N_14919,N_14971);
xnor U15186 (N_15186,N_14773,N_14924);
nor U15187 (N_15187,N_14864,N_14830);
and U15188 (N_15188,N_14914,N_14989);
and U15189 (N_15189,N_14981,N_14786);
and U15190 (N_15190,N_14773,N_14988);
nor U15191 (N_15191,N_14857,N_14896);
nor U15192 (N_15192,N_14774,N_14872);
nand U15193 (N_15193,N_14757,N_14913);
and U15194 (N_15194,N_14856,N_14936);
or U15195 (N_15195,N_14986,N_14990);
or U15196 (N_15196,N_14776,N_14760);
nand U15197 (N_15197,N_14959,N_14864);
nor U15198 (N_15198,N_14786,N_14853);
nor U15199 (N_15199,N_14938,N_14922);
nand U15200 (N_15200,N_14980,N_14930);
nand U15201 (N_15201,N_14765,N_14859);
or U15202 (N_15202,N_14786,N_14965);
and U15203 (N_15203,N_14763,N_14928);
and U15204 (N_15204,N_14984,N_14848);
xnor U15205 (N_15205,N_14972,N_14959);
and U15206 (N_15206,N_14828,N_14820);
and U15207 (N_15207,N_14966,N_14972);
and U15208 (N_15208,N_14772,N_14971);
xnor U15209 (N_15209,N_14946,N_14867);
or U15210 (N_15210,N_14763,N_14967);
nand U15211 (N_15211,N_14811,N_14841);
nor U15212 (N_15212,N_14897,N_14980);
and U15213 (N_15213,N_14770,N_14800);
and U15214 (N_15214,N_14970,N_14924);
xor U15215 (N_15215,N_14937,N_14925);
xor U15216 (N_15216,N_14969,N_14960);
and U15217 (N_15217,N_14915,N_14834);
and U15218 (N_15218,N_14857,N_14879);
nand U15219 (N_15219,N_14928,N_14852);
and U15220 (N_15220,N_14760,N_14921);
or U15221 (N_15221,N_14947,N_14785);
nor U15222 (N_15222,N_14945,N_14761);
nor U15223 (N_15223,N_14983,N_14755);
xnor U15224 (N_15224,N_14785,N_14932);
nand U15225 (N_15225,N_14984,N_14939);
or U15226 (N_15226,N_14983,N_14952);
nand U15227 (N_15227,N_14976,N_14888);
and U15228 (N_15228,N_14774,N_14754);
nand U15229 (N_15229,N_14934,N_14981);
xor U15230 (N_15230,N_14942,N_14824);
nand U15231 (N_15231,N_14820,N_14854);
nor U15232 (N_15232,N_14917,N_14867);
and U15233 (N_15233,N_14966,N_14871);
or U15234 (N_15234,N_14773,N_14855);
and U15235 (N_15235,N_14973,N_14778);
nand U15236 (N_15236,N_14780,N_14891);
and U15237 (N_15237,N_14784,N_14998);
nor U15238 (N_15238,N_14905,N_14775);
xnor U15239 (N_15239,N_14818,N_14909);
and U15240 (N_15240,N_14762,N_14907);
and U15241 (N_15241,N_14952,N_14809);
nand U15242 (N_15242,N_14986,N_14772);
or U15243 (N_15243,N_14874,N_14853);
xor U15244 (N_15244,N_14772,N_14764);
and U15245 (N_15245,N_14800,N_14956);
xnor U15246 (N_15246,N_14936,N_14829);
xnor U15247 (N_15247,N_14821,N_14954);
xnor U15248 (N_15248,N_14970,N_14922);
nand U15249 (N_15249,N_14841,N_14766);
nor U15250 (N_15250,N_15044,N_15038);
nand U15251 (N_15251,N_15099,N_15139);
and U15252 (N_15252,N_15002,N_15178);
nor U15253 (N_15253,N_15046,N_15027);
and U15254 (N_15254,N_15228,N_15180);
and U15255 (N_15255,N_15152,N_15213);
or U15256 (N_15256,N_15215,N_15132);
xor U15257 (N_15257,N_15047,N_15086);
and U15258 (N_15258,N_15185,N_15042);
xor U15259 (N_15259,N_15013,N_15202);
xor U15260 (N_15260,N_15140,N_15123);
xor U15261 (N_15261,N_15175,N_15081);
or U15262 (N_15262,N_15217,N_15201);
and U15263 (N_15263,N_15238,N_15231);
xnor U15264 (N_15264,N_15097,N_15067);
xnor U15265 (N_15265,N_15075,N_15190);
or U15266 (N_15266,N_15035,N_15028);
nand U15267 (N_15267,N_15151,N_15120);
and U15268 (N_15268,N_15025,N_15051);
or U15269 (N_15269,N_15003,N_15017);
nand U15270 (N_15270,N_15012,N_15198);
nand U15271 (N_15271,N_15143,N_15080);
or U15272 (N_15272,N_15076,N_15235);
nand U15273 (N_15273,N_15052,N_15216);
and U15274 (N_15274,N_15021,N_15144);
and U15275 (N_15275,N_15242,N_15107);
xnor U15276 (N_15276,N_15095,N_15244);
nand U15277 (N_15277,N_15210,N_15134);
and U15278 (N_15278,N_15094,N_15045);
nand U15279 (N_15279,N_15059,N_15219);
and U15280 (N_15280,N_15005,N_15089);
xnor U15281 (N_15281,N_15241,N_15162);
or U15282 (N_15282,N_15166,N_15204);
nand U15283 (N_15283,N_15225,N_15179);
xnor U15284 (N_15284,N_15088,N_15148);
or U15285 (N_15285,N_15010,N_15009);
nor U15286 (N_15286,N_15066,N_15114);
nand U15287 (N_15287,N_15174,N_15194);
and U15288 (N_15288,N_15065,N_15177);
and U15289 (N_15289,N_15187,N_15049);
nand U15290 (N_15290,N_15159,N_15040);
or U15291 (N_15291,N_15138,N_15237);
or U15292 (N_15292,N_15248,N_15023);
or U15293 (N_15293,N_15087,N_15041);
xnor U15294 (N_15294,N_15110,N_15034);
and U15295 (N_15295,N_15083,N_15048);
and U15296 (N_15296,N_15186,N_15208);
and U15297 (N_15297,N_15207,N_15188);
nand U15298 (N_15298,N_15043,N_15109);
nor U15299 (N_15299,N_15163,N_15016);
xnor U15300 (N_15300,N_15155,N_15195);
nand U15301 (N_15301,N_15221,N_15243);
nor U15302 (N_15302,N_15226,N_15211);
nor U15303 (N_15303,N_15061,N_15032);
nand U15304 (N_15304,N_15230,N_15150);
and U15305 (N_15305,N_15183,N_15102);
nor U15306 (N_15306,N_15117,N_15121);
and U15307 (N_15307,N_15036,N_15006);
and U15308 (N_15308,N_15118,N_15018);
xnor U15309 (N_15309,N_15160,N_15029);
nor U15310 (N_15310,N_15167,N_15020);
nor U15311 (N_15311,N_15232,N_15037);
xor U15312 (N_15312,N_15014,N_15004);
xor U15313 (N_15313,N_15074,N_15068);
or U15314 (N_15314,N_15113,N_15193);
nand U15315 (N_15315,N_15101,N_15070);
and U15316 (N_15316,N_15209,N_15000);
xor U15317 (N_15317,N_15220,N_15153);
xor U15318 (N_15318,N_15098,N_15077);
nand U15319 (N_15319,N_15031,N_15057);
xnor U15320 (N_15320,N_15096,N_15136);
and U15321 (N_15321,N_15227,N_15008);
or U15322 (N_15322,N_15001,N_15156);
or U15323 (N_15323,N_15203,N_15115);
xor U15324 (N_15324,N_15030,N_15093);
nor U15325 (N_15325,N_15126,N_15146);
nand U15326 (N_15326,N_15182,N_15022);
xnor U15327 (N_15327,N_15197,N_15119);
xor U15328 (N_15328,N_15073,N_15192);
xnor U15329 (N_15329,N_15060,N_15112);
or U15330 (N_15330,N_15124,N_15222);
xor U15331 (N_15331,N_15168,N_15145);
nor U15332 (N_15332,N_15085,N_15141);
nand U15333 (N_15333,N_15026,N_15082);
nor U15334 (N_15334,N_15196,N_15240);
nor U15335 (N_15335,N_15106,N_15050);
nand U15336 (N_15336,N_15246,N_15189);
nor U15337 (N_15337,N_15191,N_15053);
xor U15338 (N_15338,N_15129,N_15104);
nand U15339 (N_15339,N_15039,N_15071);
nor U15340 (N_15340,N_15170,N_15090);
nand U15341 (N_15341,N_15054,N_15111);
nand U15342 (N_15342,N_15116,N_15033);
nand U15343 (N_15343,N_15058,N_15069);
or U15344 (N_15344,N_15127,N_15214);
nor U15345 (N_15345,N_15135,N_15133);
xnor U15346 (N_15346,N_15245,N_15128);
xnor U15347 (N_15347,N_15165,N_15154);
nand U15348 (N_15348,N_15206,N_15100);
xnor U15349 (N_15349,N_15056,N_15091);
or U15350 (N_15350,N_15105,N_15015);
xor U15351 (N_15351,N_15236,N_15169);
and U15352 (N_15352,N_15072,N_15011);
and U15353 (N_15353,N_15024,N_15055);
nor U15354 (N_15354,N_15249,N_15218);
or U15355 (N_15355,N_15147,N_15161);
and U15356 (N_15356,N_15171,N_15131);
nor U15357 (N_15357,N_15158,N_15084);
or U15358 (N_15358,N_15064,N_15239);
and U15359 (N_15359,N_15062,N_15007);
nand U15360 (N_15360,N_15181,N_15164);
xnor U15361 (N_15361,N_15176,N_15103);
nand U15362 (N_15362,N_15229,N_15157);
nand U15363 (N_15363,N_15019,N_15078);
nor U15364 (N_15364,N_15172,N_15247);
nor U15365 (N_15365,N_15233,N_15125);
and U15366 (N_15366,N_15173,N_15122);
and U15367 (N_15367,N_15234,N_15212);
xnor U15368 (N_15368,N_15063,N_15142);
and U15369 (N_15369,N_15205,N_15092);
nand U15370 (N_15370,N_15223,N_15184);
or U15371 (N_15371,N_15108,N_15149);
and U15372 (N_15372,N_15224,N_15137);
xnor U15373 (N_15373,N_15199,N_15200);
nand U15374 (N_15374,N_15079,N_15130);
or U15375 (N_15375,N_15091,N_15166);
and U15376 (N_15376,N_15215,N_15185);
and U15377 (N_15377,N_15190,N_15247);
or U15378 (N_15378,N_15093,N_15151);
xnor U15379 (N_15379,N_15082,N_15033);
xnor U15380 (N_15380,N_15111,N_15167);
nor U15381 (N_15381,N_15249,N_15195);
and U15382 (N_15382,N_15093,N_15048);
and U15383 (N_15383,N_15055,N_15130);
xor U15384 (N_15384,N_15094,N_15208);
nor U15385 (N_15385,N_15152,N_15030);
xor U15386 (N_15386,N_15027,N_15099);
nand U15387 (N_15387,N_15239,N_15185);
or U15388 (N_15388,N_15044,N_15145);
and U15389 (N_15389,N_15244,N_15164);
nor U15390 (N_15390,N_15146,N_15218);
nand U15391 (N_15391,N_15244,N_15188);
and U15392 (N_15392,N_15062,N_15079);
xnor U15393 (N_15393,N_15137,N_15239);
or U15394 (N_15394,N_15244,N_15128);
and U15395 (N_15395,N_15042,N_15242);
xnor U15396 (N_15396,N_15075,N_15120);
and U15397 (N_15397,N_15229,N_15167);
nor U15398 (N_15398,N_15082,N_15120);
nand U15399 (N_15399,N_15034,N_15006);
nand U15400 (N_15400,N_15099,N_15082);
nor U15401 (N_15401,N_15199,N_15005);
nor U15402 (N_15402,N_15013,N_15095);
or U15403 (N_15403,N_15001,N_15025);
and U15404 (N_15404,N_15123,N_15061);
and U15405 (N_15405,N_15150,N_15007);
or U15406 (N_15406,N_15061,N_15119);
and U15407 (N_15407,N_15160,N_15087);
or U15408 (N_15408,N_15058,N_15111);
nand U15409 (N_15409,N_15184,N_15228);
or U15410 (N_15410,N_15067,N_15070);
or U15411 (N_15411,N_15246,N_15154);
xor U15412 (N_15412,N_15038,N_15092);
and U15413 (N_15413,N_15095,N_15202);
nor U15414 (N_15414,N_15088,N_15170);
nand U15415 (N_15415,N_15164,N_15153);
nand U15416 (N_15416,N_15122,N_15240);
and U15417 (N_15417,N_15185,N_15038);
or U15418 (N_15418,N_15101,N_15035);
nand U15419 (N_15419,N_15223,N_15069);
and U15420 (N_15420,N_15019,N_15217);
nor U15421 (N_15421,N_15053,N_15093);
nor U15422 (N_15422,N_15113,N_15199);
nor U15423 (N_15423,N_15134,N_15103);
nor U15424 (N_15424,N_15112,N_15005);
nor U15425 (N_15425,N_15134,N_15139);
nor U15426 (N_15426,N_15041,N_15150);
xor U15427 (N_15427,N_15132,N_15035);
nor U15428 (N_15428,N_15162,N_15087);
xor U15429 (N_15429,N_15158,N_15218);
and U15430 (N_15430,N_15103,N_15023);
xnor U15431 (N_15431,N_15041,N_15247);
xnor U15432 (N_15432,N_15039,N_15101);
xor U15433 (N_15433,N_15245,N_15226);
nand U15434 (N_15434,N_15172,N_15120);
nor U15435 (N_15435,N_15068,N_15079);
or U15436 (N_15436,N_15096,N_15207);
nor U15437 (N_15437,N_15133,N_15172);
or U15438 (N_15438,N_15194,N_15101);
nand U15439 (N_15439,N_15191,N_15083);
and U15440 (N_15440,N_15171,N_15139);
or U15441 (N_15441,N_15132,N_15067);
xnor U15442 (N_15442,N_15229,N_15207);
and U15443 (N_15443,N_15190,N_15189);
xor U15444 (N_15444,N_15120,N_15072);
nor U15445 (N_15445,N_15051,N_15249);
nor U15446 (N_15446,N_15249,N_15179);
or U15447 (N_15447,N_15036,N_15169);
nand U15448 (N_15448,N_15200,N_15124);
and U15449 (N_15449,N_15166,N_15011);
nor U15450 (N_15450,N_15245,N_15204);
or U15451 (N_15451,N_15175,N_15066);
or U15452 (N_15452,N_15118,N_15107);
nand U15453 (N_15453,N_15167,N_15003);
nand U15454 (N_15454,N_15169,N_15104);
and U15455 (N_15455,N_15216,N_15224);
nor U15456 (N_15456,N_15057,N_15170);
xnor U15457 (N_15457,N_15018,N_15136);
nor U15458 (N_15458,N_15086,N_15118);
nand U15459 (N_15459,N_15224,N_15058);
xor U15460 (N_15460,N_15118,N_15016);
nor U15461 (N_15461,N_15198,N_15073);
and U15462 (N_15462,N_15111,N_15239);
and U15463 (N_15463,N_15221,N_15179);
and U15464 (N_15464,N_15054,N_15110);
or U15465 (N_15465,N_15131,N_15071);
nand U15466 (N_15466,N_15091,N_15046);
and U15467 (N_15467,N_15155,N_15203);
nor U15468 (N_15468,N_15199,N_15019);
nor U15469 (N_15469,N_15193,N_15196);
nor U15470 (N_15470,N_15247,N_15217);
or U15471 (N_15471,N_15240,N_15183);
and U15472 (N_15472,N_15151,N_15048);
and U15473 (N_15473,N_15105,N_15153);
or U15474 (N_15474,N_15010,N_15005);
or U15475 (N_15475,N_15165,N_15157);
xnor U15476 (N_15476,N_15224,N_15118);
or U15477 (N_15477,N_15169,N_15132);
or U15478 (N_15478,N_15139,N_15194);
nand U15479 (N_15479,N_15038,N_15006);
and U15480 (N_15480,N_15187,N_15233);
and U15481 (N_15481,N_15164,N_15129);
xnor U15482 (N_15482,N_15173,N_15097);
and U15483 (N_15483,N_15153,N_15239);
nor U15484 (N_15484,N_15119,N_15045);
and U15485 (N_15485,N_15110,N_15175);
and U15486 (N_15486,N_15131,N_15039);
xnor U15487 (N_15487,N_15177,N_15154);
nor U15488 (N_15488,N_15105,N_15106);
or U15489 (N_15489,N_15110,N_15164);
xnor U15490 (N_15490,N_15081,N_15163);
and U15491 (N_15491,N_15146,N_15011);
nand U15492 (N_15492,N_15214,N_15181);
nor U15493 (N_15493,N_15043,N_15229);
or U15494 (N_15494,N_15207,N_15135);
or U15495 (N_15495,N_15113,N_15041);
nand U15496 (N_15496,N_15187,N_15218);
or U15497 (N_15497,N_15120,N_15181);
xnor U15498 (N_15498,N_15224,N_15226);
nand U15499 (N_15499,N_15054,N_15135);
xor U15500 (N_15500,N_15350,N_15473);
nor U15501 (N_15501,N_15351,N_15359);
and U15502 (N_15502,N_15325,N_15377);
and U15503 (N_15503,N_15460,N_15261);
and U15504 (N_15504,N_15362,N_15371);
and U15505 (N_15505,N_15487,N_15295);
or U15506 (N_15506,N_15331,N_15282);
nand U15507 (N_15507,N_15434,N_15318);
nand U15508 (N_15508,N_15453,N_15496);
xnor U15509 (N_15509,N_15286,N_15442);
nand U15510 (N_15510,N_15468,N_15431);
and U15511 (N_15511,N_15346,N_15361);
nand U15512 (N_15512,N_15255,N_15381);
and U15513 (N_15513,N_15312,N_15327);
nand U15514 (N_15514,N_15328,N_15333);
or U15515 (N_15515,N_15320,N_15317);
nand U15516 (N_15516,N_15304,N_15281);
xnor U15517 (N_15517,N_15298,N_15447);
xnor U15518 (N_15518,N_15276,N_15311);
or U15519 (N_15519,N_15402,N_15438);
nor U15520 (N_15520,N_15352,N_15372);
or U15521 (N_15521,N_15428,N_15388);
xnor U15522 (N_15522,N_15403,N_15278);
and U15523 (N_15523,N_15467,N_15396);
or U15524 (N_15524,N_15347,N_15287);
nand U15525 (N_15525,N_15477,N_15260);
and U15526 (N_15526,N_15257,N_15454);
xor U15527 (N_15527,N_15364,N_15455);
and U15528 (N_15528,N_15265,N_15400);
and U15529 (N_15529,N_15275,N_15335);
xor U15530 (N_15530,N_15369,N_15425);
nand U15531 (N_15531,N_15262,N_15417);
and U15532 (N_15532,N_15322,N_15370);
or U15533 (N_15533,N_15376,N_15291);
xor U15534 (N_15534,N_15380,N_15493);
xor U15535 (N_15535,N_15296,N_15269);
nand U15536 (N_15536,N_15332,N_15419);
and U15537 (N_15537,N_15285,N_15283);
nand U15538 (N_15538,N_15469,N_15337);
xnor U15539 (N_15539,N_15472,N_15259);
or U15540 (N_15540,N_15410,N_15432);
xnor U15541 (N_15541,N_15422,N_15349);
nor U15542 (N_15542,N_15484,N_15435);
or U15543 (N_15543,N_15436,N_15382);
nand U15544 (N_15544,N_15301,N_15268);
and U15545 (N_15545,N_15365,N_15358);
or U15546 (N_15546,N_15483,N_15448);
and U15547 (N_15547,N_15456,N_15492);
or U15548 (N_15548,N_15343,N_15280);
nor U15549 (N_15549,N_15408,N_15267);
nor U15550 (N_15550,N_15258,N_15273);
nand U15551 (N_15551,N_15452,N_15463);
nor U15552 (N_15552,N_15310,N_15314);
or U15553 (N_15553,N_15319,N_15475);
xnor U15554 (N_15554,N_15266,N_15489);
nand U15555 (N_15555,N_15451,N_15450);
nand U15556 (N_15556,N_15449,N_15412);
or U15557 (N_15557,N_15413,N_15383);
nor U15558 (N_15558,N_15446,N_15289);
xor U15559 (N_15559,N_15406,N_15354);
xnor U15560 (N_15560,N_15367,N_15409);
nor U15561 (N_15561,N_15480,N_15395);
or U15562 (N_15562,N_15445,N_15386);
nor U15563 (N_15563,N_15385,N_15437);
nor U15564 (N_15564,N_15379,N_15485);
xnor U15565 (N_15565,N_15326,N_15429);
nand U15566 (N_15566,N_15481,N_15300);
nand U15567 (N_15567,N_15405,N_15482);
nand U15568 (N_15568,N_15391,N_15421);
or U15569 (N_15569,N_15324,N_15290);
nor U15570 (N_15570,N_15415,N_15294);
or U15571 (N_15571,N_15478,N_15252);
nand U15572 (N_15572,N_15302,N_15497);
nand U15573 (N_15573,N_15279,N_15416);
and U15574 (N_15574,N_15253,N_15368);
or U15575 (N_15575,N_15345,N_15374);
nand U15576 (N_15576,N_15315,N_15474);
nand U15577 (N_15577,N_15389,N_15459);
or U15578 (N_15578,N_15307,N_15427);
nor U15579 (N_15579,N_15341,N_15423);
and U15580 (N_15580,N_15313,N_15270);
and U15581 (N_15581,N_15303,N_15339);
nor U15582 (N_15582,N_15397,N_15355);
and U15583 (N_15583,N_15441,N_15336);
nand U15584 (N_15584,N_15271,N_15338);
or U15585 (N_15585,N_15256,N_15342);
or U15586 (N_15586,N_15430,N_15363);
or U15587 (N_15587,N_15297,N_15274);
nand U15588 (N_15588,N_15323,N_15387);
nand U15589 (N_15589,N_15277,N_15378);
and U15590 (N_15590,N_15498,N_15264);
nor U15591 (N_15591,N_15494,N_15292);
and U15592 (N_15592,N_15420,N_15470);
nand U15593 (N_15593,N_15356,N_15272);
nor U15594 (N_15594,N_15418,N_15254);
xor U15595 (N_15595,N_15404,N_15305);
nand U15596 (N_15596,N_15366,N_15321);
and U15597 (N_15597,N_15476,N_15433);
xor U15598 (N_15598,N_15334,N_15439);
xnor U15599 (N_15599,N_15251,N_15495);
and U15600 (N_15600,N_15401,N_15424);
or U15601 (N_15601,N_15440,N_15263);
nor U15602 (N_15602,N_15461,N_15462);
nor U15603 (N_15603,N_15411,N_15330);
or U15604 (N_15604,N_15457,N_15399);
nand U15605 (N_15605,N_15344,N_15309);
nor U15606 (N_15606,N_15340,N_15288);
or U15607 (N_15607,N_15373,N_15479);
or U15608 (N_15608,N_15316,N_15486);
xnor U15609 (N_15609,N_15464,N_15306);
or U15610 (N_15610,N_15393,N_15284);
or U15611 (N_15611,N_15357,N_15488);
nand U15612 (N_15612,N_15491,N_15443);
xnor U15613 (N_15613,N_15375,N_15299);
nor U15614 (N_15614,N_15465,N_15407);
or U15615 (N_15615,N_15444,N_15353);
nor U15616 (N_15616,N_15458,N_15329);
or U15617 (N_15617,N_15384,N_15466);
nor U15618 (N_15618,N_15471,N_15390);
xnor U15619 (N_15619,N_15392,N_15360);
or U15620 (N_15620,N_15250,N_15398);
or U15621 (N_15621,N_15308,N_15499);
nor U15622 (N_15622,N_15293,N_15414);
nor U15623 (N_15623,N_15490,N_15348);
nor U15624 (N_15624,N_15394,N_15426);
xor U15625 (N_15625,N_15498,N_15391);
and U15626 (N_15626,N_15444,N_15495);
xnor U15627 (N_15627,N_15354,N_15269);
xor U15628 (N_15628,N_15424,N_15342);
and U15629 (N_15629,N_15425,N_15390);
xnor U15630 (N_15630,N_15301,N_15376);
nand U15631 (N_15631,N_15285,N_15325);
nand U15632 (N_15632,N_15386,N_15331);
xor U15633 (N_15633,N_15475,N_15343);
and U15634 (N_15634,N_15430,N_15315);
nor U15635 (N_15635,N_15374,N_15409);
nor U15636 (N_15636,N_15388,N_15284);
nand U15637 (N_15637,N_15292,N_15414);
nor U15638 (N_15638,N_15378,N_15441);
xnor U15639 (N_15639,N_15441,N_15269);
xor U15640 (N_15640,N_15338,N_15409);
or U15641 (N_15641,N_15487,N_15361);
or U15642 (N_15642,N_15414,N_15276);
or U15643 (N_15643,N_15373,N_15374);
and U15644 (N_15644,N_15314,N_15277);
xor U15645 (N_15645,N_15425,N_15277);
or U15646 (N_15646,N_15478,N_15443);
xor U15647 (N_15647,N_15478,N_15324);
or U15648 (N_15648,N_15327,N_15394);
or U15649 (N_15649,N_15308,N_15403);
xnor U15650 (N_15650,N_15491,N_15294);
and U15651 (N_15651,N_15342,N_15453);
nand U15652 (N_15652,N_15286,N_15479);
nor U15653 (N_15653,N_15260,N_15428);
nor U15654 (N_15654,N_15483,N_15273);
nand U15655 (N_15655,N_15373,N_15309);
nor U15656 (N_15656,N_15314,N_15433);
and U15657 (N_15657,N_15472,N_15301);
nand U15658 (N_15658,N_15442,N_15344);
and U15659 (N_15659,N_15342,N_15288);
nor U15660 (N_15660,N_15255,N_15316);
nor U15661 (N_15661,N_15485,N_15462);
nand U15662 (N_15662,N_15270,N_15417);
and U15663 (N_15663,N_15310,N_15416);
nand U15664 (N_15664,N_15467,N_15340);
nand U15665 (N_15665,N_15497,N_15266);
xnor U15666 (N_15666,N_15284,N_15376);
and U15667 (N_15667,N_15449,N_15295);
nor U15668 (N_15668,N_15258,N_15434);
and U15669 (N_15669,N_15445,N_15305);
nand U15670 (N_15670,N_15278,N_15301);
nand U15671 (N_15671,N_15476,N_15497);
nand U15672 (N_15672,N_15435,N_15393);
and U15673 (N_15673,N_15342,N_15381);
xor U15674 (N_15674,N_15425,N_15303);
nand U15675 (N_15675,N_15447,N_15395);
or U15676 (N_15676,N_15459,N_15395);
and U15677 (N_15677,N_15270,N_15322);
and U15678 (N_15678,N_15375,N_15318);
or U15679 (N_15679,N_15391,N_15258);
or U15680 (N_15680,N_15442,N_15411);
and U15681 (N_15681,N_15280,N_15292);
xnor U15682 (N_15682,N_15325,N_15367);
nor U15683 (N_15683,N_15353,N_15296);
or U15684 (N_15684,N_15441,N_15467);
xnor U15685 (N_15685,N_15283,N_15332);
nor U15686 (N_15686,N_15352,N_15279);
or U15687 (N_15687,N_15302,N_15275);
nor U15688 (N_15688,N_15272,N_15387);
or U15689 (N_15689,N_15423,N_15372);
nor U15690 (N_15690,N_15256,N_15429);
nor U15691 (N_15691,N_15434,N_15312);
or U15692 (N_15692,N_15409,N_15478);
xor U15693 (N_15693,N_15309,N_15422);
nand U15694 (N_15694,N_15383,N_15390);
nor U15695 (N_15695,N_15486,N_15411);
or U15696 (N_15696,N_15332,N_15256);
or U15697 (N_15697,N_15359,N_15446);
xor U15698 (N_15698,N_15396,N_15399);
nor U15699 (N_15699,N_15457,N_15257);
or U15700 (N_15700,N_15416,N_15298);
and U15701 (N_15701,N_15344,N_15458);
nor U15702 (N_15702,N_15320,N_15346);
nor U15703 (N_15703,N_15279,N_15472);
nand U15704 (N_15704,N_15260,N_15495);
or U15705 (N_15705,N_15273,N_15313);
nand U15706 (N_15706,N_15313,N_15311);
and U15707 (N_15707,N_15318,N_15392);
nand U15708 (N_15708,N_15372,N_15304);
or U15709 (N_15709,N_15499,N_15373);
and U15710 (N_15710,N_15434,N_15497);
and U15711 (N_15711,N_15498,N_15396);
and U15712 (N_15712,N_15479,N_15487);
or U15713 (N_15713,N_15308,N_15254);
nand U15714 (N_15714,N_15485,N_15491);
and U15715 (N_15715,N_15381,N_15439);
nor U15716 (N_15716,N_15259,N_15258);
nor U15717 (N_15717,N_15390,N_15413);
nand U15718 (N_15718,N_15479,N_15452);
xnor U15719 (N_15719,N_15271,N_15369);
nand U15720 (N_15720,N_15370,N_15382);
xnor U15721 (N_15721,N_15311,N_15344);
nor U15722 (N_15722,N_15419,N_15310);
or U15723 (N_15723,N_15331,N_15456);
and U15724 (N_15724,N_15351,N_15427);
nor U15725 (N_15725,N_15404,N_15343);
nand U15726 (N_15726,N_15385,N_15454);
and U15727 (N_15727,N_15369,N_15266);
nor U15728 (N_15728,N_15308,N_15357);
or U15729 (N_15729,N_15356,N_15426);
or U15730 (N_15730,N_15371,N_15403);
nor U15731 (N_15731,N_15349,N_15322);
nor U15732 (N_15732,N_15438,N_15361);
nand U15733 (N_15733,N_15323,N_15269);
xnor U15734 (N_15734,N_15286,N_15289);
and U15735 (N_15735,N_15344,N_15252);
or U15736 (N_15736,N_15333,N_15473);
xnor U15737 (N_15737,N_15423,N_15415);
nand U15738 (N_15738,N_15408,N_15479);
and U15739 (N_15739,N_15453,N_15275);
nand U15740 (N_15740,N_15251,N_15383);
nor U15741 (N_15741,N_15454,N_15498);
nand U15742 (N_15742,N_15422,N_15334);
nor U15743 (N_15743,N_15420,N_15252);
and U15744 (N_15744,N_15437,N_15358);
and U15745 (N_15745,N_15466,N_15299);
and U15746 (N_15746,N_15278,N_15440);
nor U15747 (N_15747,N_15294,N_15346);
or U15748 (N_15748,N_15360,N_15397);
nor U15749 (N_15749,N_15444,N_15270);
xnor U15750 (N_15750,N_15587,N_15623);
or U15751 (N_15751,N_15724,N_15669);
or U15752 (N_15752,N_15719,N_15523);
or U15753 (N_15753,N_15556,N_15679);
xor U15754 (N_15754,N_15699,N_15631);
nor U15755 (N_15755,N_15698,N_15546);
nor U15756 (N_15756,N_15501,N_15642);
or U15757 (N_15757,N_15648,N_15539);
and U15758 (N_15758,N_15637,N_15685);
and U15759 (N_15759,N_15639,N_15700);
nand U15760 (N_15760,N_15684,N_15668);
xnor U15761 (N_15761,N_15671,N_15504);
xnor U15762 (N_15762,N_15721,N_15599);
xor U15763 (N_15763,N_15554,N_15675);
xor U15764 (N_15764,N_15562,N_15712);
xnor U15765 (N_15765,N_15658,N_15583);
nor U15766 (N_15766,N_15686,N_15748);
and U15767 (N_15767,N_15688,N_15739);
and U15768 (N_15768,N_15503,N_15695);
xnor U15769 (N_15769,N_15530,N_15718);
or U15770 (N_15770,N_15536,N_15577);
or U15771 (N_15771,N_15713,N_15570);
nand U15772 (N_15772,N_15502,N_15550);
and U15773 (N_15773,N_15733,N_15507);
xor U15774 (N_15774,N_15618,N_15505);
xor U15775 (N_15775,N_15617,N_15532);
xor U15776 (N_15776,N_15666,N_15736);
nor U15777 (N_15777,N_15512,N_15552);
or U15778 (N_15778,N_15714,N_15627);
xor U15779 (N_15779,N_15542,N_15547);
nand U15780 (N_15780,N_15572,N_15726);
nand U15781 (N_15781,N_15659,N_15579);
xor U15782 (N_15782,N_15533,N_15731);
or U15783 (N_15783,N_15680,N_15635);
or U15784 (N_15784,N_15535,N_15591);
xnor U15785 (N_15785,N_15705,N_15519);
nand U15786 (N_15786,N_15506,N_15727);
nor U15787 (N_15787,N_15742,N_15697);
xnor U15788 (N_15788,N_15664,N_15551);
and U15789 (N_15789,N_15513,N_15691);
nand U15790 (N_15790,N_15683,N_15701);
xor U15791 (N_15791,N_15598,N_15749);
nand U15792 (N_15792,N_15508,N_15693);
or U15793 (N_15793,N_15611,N_15633);
or U15794 (N_15794,N_15704,N_15608);
or U15795 (N_15795,N_15741,N_15616);
nand U15796 (N_15796,N_15703,N_15560);
and U15797 (N_15797,N_15515,N_15612);
xnor U15798 (N_15798,N_15740,N_15606);
or U15799 (N_15799,N_15628,N_15594);
or U15800 (N_15800,N_15578,N_15640);
nor U15801 (N_15801,N_15672,N_15600);
or U15802 (N_15802,N_15604,N_15722);
xnor U15803 (N_15803,N_15730,N_15745);
and U15804 (N_15804,N_15571,N_15596);
xnor U15805 (N_15805,N_15595,N_15626);
or U15806 (N_15806,N_15555,N_15711);
or U15807 (N_15807,N_15743,N_15651);
nand U15808 (N_15808,N_15514,N_15568);
and U15809 (N_15809,N_15538,N_15661);
and U15810 (N_15810,N_15609,N_15621);
nor U15811 (N_15811,N_15581,N_15707);
nor U15812 (N_15812,N_15663,N_15567);
xor U15813 (N_15813,N_15682,N_15559);
and U15814 (N_15814,N_15602,N_15681);
or U15815 (N_15815,N_15629,N_15641);
xor U15816 (N_15816,N_15580,N_15603);
nand U15817 (N_15817,N_15574,N_15541);
nand U15818 (N_15818,N_15649,N_15723);
and U15819 (N_15819,N_15689,N_15638);
xnor U15820 (N_15820,N_15717,N_15660);
nand U15821 (N_15821,N_15563,N_15735);
nand U15822 (N_15822,N_15738,N_15747);
nand U15823 (N_15823,N_15696,N_15509);
nand U15824 (N_15824,N_15725,N_15511);
nand U15825 (N_15825,N_15647,N_15518);
nand U15826 (N_15826,N_15737,N_15636);
and U15827 (N_15827,N_15543,N_15549);
and U15828 (N_15828,N_15565,N_15566);
and U15829 (N_15829,N_15584,N_15561);
xnor U15830 (N_15830,N_15593,N_15615);
xnor U15831 (N_15831,N_15597,N_15706);
xor U15832 (N_15832,N_15522,N_15592);
or U15833 (N_15833,N_15564,N_15630);
or U15834 (N_15834,N_15527,N_15620);
xor U15835 (N_15835,N_15732,N_15605);
xor U15836 (N_15836,N_15510,N_15548);
nand U15837 (N_15837,N_15670,N_15526);
xnor U15838 (N_15838,N_15607,N_15710);
nor U15839 (N_15839,N_15619,N_15674);
or U15840 (N_15840,N_15694,N_15540);
and U15841 (N_15841,N_15744,N_15545);
nor U15842 (N_15842,N_15653,N_15589);
nand U15843 (N_15843,N_15654,N_15575);
or U15844 (N_15844,N_15709,N_15521);
or U15845 (N_15845,N_15517,N_15678);
and U15846 (N_15846,N_15676,N_15632);
or U15847 (N_15847,N_15657,N_15646);
xor U15848 (N_15848,N_15655,N_15729);
and U15849 (N_15849,N_15528,N_15534);
nand U15850 (N_15850,N_15673,N_15558);
or U15851 (N_15851,N_15610,N_15531);
nand U15852 (N_15852,N_15500,N_15728);
nor U15853 (N_15853,N_15715,N_15569);
or U15854 (N_15854,N_15590,N_15588);
and U15855 (N_15855,N_15716,N_15624);
or U15856 (N_15856,N_15720,N_15520);
nand U15857 (N_15857,N_15734,N_15573);
nor U15858 (N_15858,N_15692,N_15586);
nor U15859 (N_15859,N_15687,N_15665);
nor U15860 (N_15860,N_15544,N_15643);
xnor U15861 (N_15861,N_15652,N_15582);
and U15862 (N_15862,N_15650,N_15667);
nand U15863 (N_15863,N_15702,N_15677);
xor U15864 (N_15864,N_15622,N_15529);
nand U15865 (N_15865,N_15708,N_15690);
nor U15866 (N_15866,N_15576,N_15557);
nor U15867 (N_15867,N_15625,N_15524);
or U15868 (N_15868,N_15613,N_15601);
nand U15869 (N_15869,N_15644,N_15585);
nor U15870 (N_15870,N_15614,N_15537);
nor U15871 (N_15871,N_15645,N_15516);
xnor U15872 (N_15872,N_15634,N_15525);
xor U15873 (N_15873,N_15553,N_15662);
or U15874 (N_15874,N_15746,N_15656);
and U15875 (N_15875,N_15634,N_15654);
and U15876 (N_15876,N_15504,N_15648);
xor U15877 (N_15877,N_15552,N_15585);
or U15878 (N_15878,N_15713,N_15557);
or U15879 (N_15879,N_15575,N_15722);
or U15880 (N_15880,N_15598,N_15744);
xnor U15881 (N_15881,N_15654,N_15672);
nand U15882 (N_15882,N_15633,N_15593);
nor U15883 (N_15883,N_15639,N_15652);
nand U15884 (N_15884,N_15567,N_15741);
nor U15885 (N_15885,N_15564,N_15606);
nand U15886 (N_15886,N_15700,N_15634);
nor U15887 (N_15887,N_15671,N_15724);
or U15888 (N_15888,N_15715,N_15583);
nand U15889 (N_15889,N_15602,N_15637);
nand U15890 (N_15890,N_15668,N_15683);
nor U15891 (N_15891,N_15568,N_15645);
or U15892 (N_15892,N_15583,N_15741);
or U15893 (N_15893,N_15613,N_15690);
xor U15894 (N_15894,N_15604,N_15507);
xnor U15895 (N_15895,N_15588,N_15677);
xor U15896 (N_15896,N_15517,N_15577);
or U15897 (N_15897,N_15511,N_15747);
or U15898 (N_15898,N_15557,N_15682);
nand U15899 (N_15899,N_15532,N_15567);
nor U15900 (N_15900,N_15657,N_15690);
nand U15901 (N_15901,N_15650,N_15714);
xor U15902 (N_15902,N_15504,N_15530);
or U15903 (N_15903,N_15661,N_15652);
nor U15904 (N_15904,N_15722,N_15527);
nand U15905 (N_15905,N_15554,N_15741);
nor U15906 (N_15906,N_15747,N_15628);
nand U15907 (N_15907,N_15749,N_15717);
and U15908 (N_15908,N_15676,N_15654);
nor U15909 (N_15909,N_15593,N_15608);
and U15910 (N_15910,N_15690,N_15619);
nor U15911 (N_15911,N_15537,N_15580);
or U15912 (N_15912,N_15694,N_15513);
and U15913 (N_15913,N_15515,N_15537);
xor U15914 (N_15914,N_15721,N_15563);
nand U15915 (N_15915,N_15661,N_15645);
nand U15916 (N_15916,N_15524,N_15645);
nand U15917 (N_15917,N_15713,N_15725);
nor U15918 (N_15918,N_15585,N_15645);
nor U15919 (N_15919,N_15589,N_15558);
nor U15920 (N_15920,N_15653,N_15683);
xnor U15921 (N_15921,N_15565,N_15592);
or U15922 (N_15922,N_15675,N_15552);
and U15923 (N_15923,N_15694,N_15596);
or U15924 (N_15924,N_15689,N_15563);
or U15925 (N_15925,N_15527,N_15551);
or U15926 (N_15926,N_15525,N_15509);
or U15927 (N_15927,N_15681,N_15568);
nor U15928 (N_15928,N_15716,N_15591);
nor U15929 (N_15929,N_15563,N_15518);
or U15930 (N_15930,N_15515,N_15742);
nand U15931 (N_15931,N_15655,N_15675);
xnor U15932 (N_15932,N_15713,N_15729);
nand U15933 (N_15933,N_15531,N_15526);
or U15934 (N_15934,N_15538,N_15718);
xnor U15935 (N_15935,N_15738,N_15629);
nand U15936 (N_15936,N_15669,N_15604);
xnor U15937 (N_15937,N_15743,N_15656);
nor U15938 (N_15938,N_15510,N_15585);
nand U15939 (N_15939,N_15715,N_15604);
xor U15940 (N_15940,N_15595,N_15649);
xor U15941 (N_15941,N_15507,N_15610);
nand U15942 (N_15942,N_15525,N_15618);
xnor U15943 (N_15943,N_15542,N_15732);
nand U15944 (N_15944,N_15699,N_15648);
xor U15945 (N_15945,N_15712,N_15717);
nor U15946 (N_15946,N_15597,N_15747);
xnor U15947 (N_15947,N_15568,N_15676);
or U15948 (N_15948,N_15669,N_15594);
nand U15949 (N_15949,N_15671,N_15579);
xnor U15950 (N_15950,N_15529,N_15533);
xnor U15951 (N_15951,N_15673,N_15511);
or U15952 (N_15952,N_15663,N_15712);
nand U15953 (N_15953,N_15708,N_15720);
nor U15954 (N_15954,N_15549,N_15618);
and U15955 (N_15955,N_15530,N_15546);
or U15956 (N_15956,N_15657,N_15659);
nand U15957 (N_15957,N_15632,N_15718);
and U15958 (N_15958,N_15556,N_15544);
nor U15959 (N_15959,N_15676,N_15688);
or U15960 (N_15960,N_15703,N_15608);
or U15961 (N_15961,N_15569,N_15621);
or U15962 (N_15962,N_15733,N_15598);
xor U15963 (N_15963,N_15581,N_15703);
nand U15964 (N_15964,N_15728,N_15681);
or U15965 (N_15965,N_15705,N_15507);
nor U15966 (N_15966,N_15715,N_15540);
xnor U15967 (N_15967,N_15523,N_15650);
xnor U15968 (N_15968,N_15645,N_15699);
and U15969 (N_15969,N_15666,N_15668);
nand U15970 (N_15970,N_15640,N_15665);
nor U15971 (N_15971,N_15506,N_15665);
or U15972 (N_15972,N_15700,N_15631);
or U15973 (N_15973,N_15724,N_15703);
nor U15974 (N_15974,N_15525,N_15739);
and U15975 (N_15975,N_15606,N_15613);
nor U15976 (N_15976,N_15525,N_15578);
and U15977 (N_15977,N_15600,N_15539);
xor U15978 (N_15978,N_15625,N_15679);
and U15979 (N_15979,N_15579,N_15632);
nor U15980 (N_15980,N_15507,N_15640);
nand U15981 (N_15981,N_15684,N_15611);
xnor U15982 (N_15982,N_15583,N_15539);
nand U15983 (N_15983,N_15579,N_15580);
nand U15984 (N_15984,N_15694,N_15725);
xor U15985 (N_15985,N_15748,N_15620);
xnor U15986 (N_15986,N_15658,N_15519);
xnor U15987 (N_15987,N_15577,N_15707);
and U15988 (N_15988,N_15513,N_15608);
xnor U15989 (N_15989,N_15531,N_15575);
or U15990 (N_15990,N_15520,N_15530);
nand U15991 (N_15991,N_15681,N_15525);
nor U15992 (N_15992,N_15538,N_15649);
xor U15993 (N_15993,N_15715,N_15707);
and U15994 (N_15994,N_15662,N_15680);
nor U15995 (N_15995,N_15507,N_15653);
and U15996 (N_15996,N_15626,N_15596);
xor U15997 (N_15997,N_15595,N_15687);
nor U15998 (N_15998,N_15715,N_15742);
and U15999 (N_15999,N_15737,N_15571);
or U16000 (N_16000,N_15752,N_15848);
or U16001 (N_16001,N_15940,N_15840);
or U16002 (N_16002,N_15830,N_15825);
or U16003 (N_16003,N_15851,N_15989);
xor U16004 (N_16004,N_15810,N_15904);
xor U16005 (N_16005,N_15920,N_15950);
and U16006 (N_16006,N_15828,N_15844);
or U16007 (N_16007,N_15758,N_15806);
and U16008 (N_16008,N_15903,N_15843);
nor U16009 (N_16009,N_15857,N_15962);
xnor U16010 (N_16010,N_15885,N_15833);
or U16011 (N_16011,N_15964,N_15995);
and U16012 (N_16012,N_15864,N_15919);
and U16013 (N_16013,N_15789,N_15882);
and U16014 (N_16014,N_15967,N_15985);
nand U16015 (N_16015,N_15750,N_15970);
nand U16016 (N_16016,N_15767,N_15772);
xor U16017 (N_16017,N_15971,N_15974);
or U16018 (N_16018,N_15841,N_15947);
nor U16019 (N_16019,N_15937,N_15814);
and U16020 (N_16020,N_15861,N_15800);
nor U16021 (N_16021,N_15777,N_15880);
and U16022 (N_16022,N_15834,N_15948);
nor U16023 (N_16023,N_15860,N_15933);
nor U16024 (N_16024,N_15872,N_15794);
or U16025 (N_16025,N_15899,N_15957);
or U16026 (N_16026,N_15892,N_15979);
xnor U16027 (N_16027,N_15846,N_15781);
nand U16028 (N_16028,N_15775,N_15949);
nor U16029 (N_16029,N_15969,N_15922);
and U16030 (N_16030,N_15982,N_15910);
nand U16031 (N_16031,N_15818,N_15803);
nor U16032 (N_16032,N_15958,N_15845);
xor U16033 (N_16033,N_15918,N_15905);
xor U16034 (N_16034,N_15879,N_15997);
nor U16035 (N_16035,N_15779,N_15799);
nand U16036 (N_16036,N_15852,N_15894);
or U16037 (N_16037,N_15832,N_15801);
nand U16038 (N_16038,N_15981,N_15856);
nand U16039 (N_16039,N_15812,N_15932);
or U16040 (N_16040,N_15956,N_15805);
nor U16041 (N_16041,N_15798,N_15963);
nor U16042 (N_16042,N_15754,N_15944);
or U16043 (N_16043,N_15824,N_15916);
nand U16044 (N_16044,N_15959,N_15975);
nand U16045 (N_16045,N_15836,N_15931);
nor U16046 (N_16046,N_15761,N_15802);
and U16047 (N_16047,N_15816,N_15926);
nor U16048 (N_16048,N_15990,N_15782);
or U16049 (N_16049,N_15900,N_15924);
nor U16050 (N_16050,N_15788,N_15823);
nor U16051 (N_16051,N_15927,N_15925);
or U16052 (N_16052,N_15796,N_15917);
and U16053 (N_16053,N_15795,N_15888);
nor U16054 (N_16054,N_15776,N_15953);
xnor U16055 (N_16055,N_15943,N_15778);
xnor U16056 (N_16056,N_15991,N_15973);
and U16057 (N_16057,N_15793,N_15759);
or U16058 (N_16058,N_15804,N_15988);
xor U16059 (N_16059,N_15842,N_15780);
nand U16060 (N_16060,N_15952,N_15993);
or U16061 (N_16061,N_15809,N_15865);
xnor U16062 (N_16062,N_15898,N_15791);
xnor U16063 (N_16063,N_15983,N_15908);
and U16064 (N_16064,N_15853,N_15813);
xor U16065 (N_16065,N_15883,N_15762);
or U16066 (N_16066,N_15873,N_15786);
nand U16067 (N_16067,N_15942,N_15829);
nor U16068 (N_16068,N_15822,N_15902);
nand U16069 (N_16069,N_15870,N_15890);
and U16070 (N_16070,N_15797,N_15835);
xnor U16071 (N_16071,N_15886,N_15869);
and U16072 (N_16072,N_15751,N_15994);
or U16073 (N_16073,N_15895,N_15760);
xor U16074 (N_16074,N_15930,N_15763);
xor U16075 (N_16075,N_15838,N_15811);
nor U16076 (N_16076,N_15987,N_15855);
nor U16077 (N_16077,N_15935,N_15757);
nor U16078 (N_16078,N_15913,N_15901);
xor U16079 (N_16079,N_15911,N_15766);
xor U16080 (N_16080,N_15774,N_15887);
nand U16081 (N_16081,N_15907,N_15992);
or U16082 (N_16082,N_15819,N_15821);
nand U16083 (N_16083,N_15753,N_15929);
nor U16084 (N_16084,N_15909,N_15893);
or U16085 (N_16085,N_15977,N_15874);
or U16086 (N_16086,N_15889,N_15984);
or U16087 (N_16087,N_15875,N_15928);
or U16088 (N_16088,N_15976,N_15831);
or U16089 (N_16089,N_15849,N_15996);
or U16090 (N_16090,N_15764,N_15912);
and U16091 (N_16091,N_15980,N_15847);
and U16092 (N_16092,N_15938,N_15850);
or U16093 (N_16093,N_15951,N_15941);
nand U16094 (N_16094,N_15891,N_15968);
nand U16095 (N_16095,N_15858,N_15945);
or U16096 (N_16096,N_15936,N_15966);
xnor U16097 (N_16097,N_15770,N_15784);
and U16098 (N_16098,N_15978,N_15965);
nand U16099 (N_16099,N_15866,N_15755);
and U16100 (N_16100,N_15871,N_15790);
nor U16101 (N_16101,N_15815,N_15773);
or U16102 (N_16102,N_15765,N_15817);
nand U16103 (N_16103,N_15923,N_15807);
or U16104 (N_16104,N_15839,N_15859);
nand U16105 (N_16105,N_15808,N_15837);
xor U16106 (N_16106,N_15921,N_15939);
nand U16107 (N_16107,N_15867,N_15826);
xnor U16108 (N_16108,N_15787,N_15876);
nor U16109 (N_16109,N_15785,N_15960);
and U16110 (N_16110,N_15881,N_15771);
or U16111 (N_16111,N_15946,N_15863);
nor U16112 (N_16112,N_15986,N_15792);
xor U16113 (N_16113,N_15972,N_15999);
nor U16114 (N_16114,N_15868,N_15955);
or U16115 (N_16115,N_15769,N_15783);
xnor U16116 (N_16116,N_15906,N_15961);
nand U16117 (N_16117,N_15768,N_15914);
nand U16118 (N_16118,N_15854,N_15862);
nand U16119 (N_16119,N_15827,N_15878);
or U16120 (N_16120,N_15820,N_15897);
nand U16121 (N_16121,N_15896,N_15756);
xnor U16122 (N_16122,N_15877,N_15934);
nor U16123 (N_16123,N_15884,N_15998);
and U16124 (N_16124,N_15915,N_15954);
xor U16125 (N_16125,N_15897,N_15819);
nand U16126 (N_16126,N_15942,N_15809);
nand U16127 (N_16127,N_15900,N_15997);
xor U16128 (N_16128,N_15902,N_15906);
nand U16129 (N_16129,N_15865,N_15798);
and U16130 (N_16130,N_15754,N_15891);
and U16131 (N_16131,N_15850,N_15814);
and U16132 (N_16132,N_15782,N_15839);
or U16133 (N_16133,N_15781,N_15758);
nor U16134 (N_16134,N_15922,N_15911);
or U16135 (N_16135,N_15815,N_15972);
and U16136 (N_16136,N_15957,N_15759);
and U16137 (N_16137,N_15941,N_15799);
and U16138 (N_16138,N_15883,N_15888);
and U16139 (N_16139,N_15820,N_15944);
nor U16140 (N_16140,N_15793,N_15968);
nand U16141 (N_16141,N_15970,N_15949);
xnor U16142 (N_16142,N_15756,N_15829);
or U16143 (N_16143,N_15967,N_15872);
nand U16144 (N_16144,N_15756,N_15961);
nand U16145 (N_16145,N_15927,N_15886);
nor U16146 (N_16146,N_15953,N_15808);
and U16147 (N_16147,N_15970,N_15956);
nor U16148 (N_16148,N_15812,N_15865);
xnor U16149 (N_16149,N_15861,N_15754);
and U16150 (N_16150,N_15793,N_15904);
and U16151 (N_16151,N_15985,N_15873);
xor U16152 (N_16152,N_15952,N_15874);
or U16153 (N_16153,N_15952,N_15939);
and U16154 (N_16154,N_15992,N_15838);
nor U16155 (N_16155,N_15925,N_15841);
and U16156 (N_16156,N_15989,N_15804);
nor U16157 (N_16157,N_15853,N_15829);
nand U16158 (N_16158,N_15813,N_15774);
and U16159 (N_16159,N_15965,N_15782);
and U16160 (N_16160,N_15874,N_15822);
and U16161 (N_16161,N_15908,N_15968);
or U16162 (N_16162,N_15975,N_15987);
nor U16163 (N_16163,N_15867,N_15918);
xor U16164 (N_16164,N_15761,N_15999);
xnor U16165 (N_16165,N_15924,N_15796);
xnor U16166 (N_16166,N_15892,N_15805);
nand U16167 (N_16167,N_15881,N_15863);
nand U16168 (N_16168,N_15957,N_15891);
or U16169 (N_16169,N_15766,N_15834);
and U16170 (N_16170,N_15837,N_15994);
xor U16171 (N_16171,N_15901,N_15914);
xor U16172 (N_16172,N_15822,N_15786);
nor U16173 (N_16173,N_15884,N_15841);
nor U16174 (N_16174,N_15818,N_15783);
xor U16175 (N_16175,N_15804,N_15925);
and U16176 (N_16176,N_15892,N_15809);
and U16177 (N_16177,N_15971,N_15754);
nand U16178 (N_16178,N_15910,N_15832);
nor U16179 (N_16179,N_15802,N_15911);
nand U16180 (N_16180,N_15913,N_15968);
nand U16181 (N_16181,N_15780,N_15810);
or U16182 (N_16182,N_15874,N_15993);
and U16183 (N_16183,N_15816,N_15946);
and U16184 (N_16184,N_15873,N_15900);
nor U16185 (N_16185,N_15917,N_15997);
or U16186 (N_16186,N_15792,N_15804);
or U16187 (N_16187,N_15978,N_15940);
nand U16188 (N_16188,N_15894,N_15790);
nor U16189 (N_16189,N_15801,N_15951);
nor U16190 (N_16190,N_15938,N_15871);
nand U16191 (N_16191,N_15808,N_15752);
nor U16192 (N_16192,N_15930,N_15946);
nor U16193 (N_16193,N_15788,N_15883);
and U16194 (N_16194,N_15901,N_15829);
and U16195 (N_16195,N_15824,N_15818);
xor U16196 (N_16196,N_15978,N_15896);
or U16197 (N_16197,N_15952,N_15941);
nand U16198 (N_16198,N_15844,N_15769);
xor U16199 (N_16199,N_15808,N_15894);
and U16200 (N_16200,N_15843,N_15927);
xor U16201 (N_16201,N_15863,N_15918);
nor U16202 (N_16202,N_15924,N_15941);
xnor U16203 (N_16203,N_15949,N_15904);
nor U16204 (N_16204,N_15956,N_15757);
nand U16205 (N_16205,N_15968,N_15948);
or U16206 (N_16206,N_15963,N_15872);
or U16207 (N_16207,N_15868,N_15880);
or U16208 (N_16208,N_15932,N_15897);
xnor U16209 (N_16209,N_15870,N_15930);
nor U16210 (N_16210,N_15788,N_15770);
nor U16211 (N_16211,N_15990,N_15931);
nand U16212 (N_16212,N_15801,N_15921);
nor U16213 (N_16213,N_15910,N_15920);
or U16214 (N_16214,N_15787,N_15760);
or U16215 (N_16215,N_15940,N_15828);
nand U16216 (N_16216,N_15838,N_15879);
or U16217 (N_16217,N_15831,N_15830);
xnor U16218 (N_16218,N_15921,N_15875);
or U16219 (N_16219,N_15991,N_15755);
or U16220 (N_16220,N_15881,N_15862);
or U16221 (N_16221,N_15807,N_15996);
and U16222 (N_16222,N_15870,N_15956);
nor U16223 (N_16223,N_15791,N_15950);
nor U16224 (N_16224,N_15987,N_15925);
or U16225 (N_16225,N_15847,N_15984);
nand U16226 (N_16226,N_15824,N_15944);
xor U16227 (N_16227,N_15874,N_15918);
xor U16228 (N_16228,N_15800,N_15869);
nor U16229 (N_16229,N_15844,N_15893);
and U16230 (N_16230,N_15979,N_15814);
or U16231 (N_16231,N_15940,N_15903);
xnor U16232 (N_16232,N_15915,N_15848);
and U16233 (N_16233,N_15806,N_15909);
or U16234 (N_16234,N_15866,N_15809);
or U16235 (N_16235,N_15872,N_15847);
nor U16236 (N_16236,N_15825,N_15770);
or U16237 (N_16237,N_15856,N_15758);
and U16238 (N_16238,N_15876,N_15896);
xor U16239 (N_16239,N_15774,N_15825);
xor U16240 (N_16240,N_15895,N_15797);
xnor U16241 (N_16241,N_15888,N_15874);
nor U16242 (N_16242,N_15955,N_15863);
or U16243 (N_16243,N_15824,N_15908);
nor U16244 (N_16244,N_15862,N_15807);
or U16245 (N_16245,N_15997,N_15827);
and U16246 (N_16246,N_15895,N_15865);
nor U16247 (N_16247,N_15974,N_15938);
and U16248 (N_16248,N_15821,N_15868);
or U16249 (N_16249,N_15798,N_15966);
xnor U16250 (N_16250,N_16198,N_16079);
xor U16251 (N_16251,N_16049,N_16184);
xnor U16252 (N_16252,N_16164,N_16106);
xnor U16253 (N_16253,N_16135,N_16018);
xor U16254 (N_16254,N_16229,N_16157);
and U16255 (N_16255,N_16228,N_16212);
and U16256 (N_16256,N_16072,N_16071);
and U16257 (N_16257,N_16160,N_16122);
and U16258 (N_16258,N_16119,N_16065);
and U16259 (N_16259,N_16206,N_16100);
or U16260 (N_16260,N_16069,N_16218);
xor U16261 (N_16261,N_16078,N_16068);
nor U16262 (N_16262,N_16020,N_16153);
nor U16263 (N_16263,N_16156,N_16003);
nor U16264 (N_16264,N_16008,N_16052);
xor U16265 (N_16265,N_16015,N_16090);
nand U16266 (N_16266,N_16140,N_16217);
or U16267 (N_16267,N_16213,N_16014);
xor U16268 (N_16268,N_16026,N_16149);
nand U16269 (N_16269,N_16127,N_16031);
and U16270 (N_16270,N_16200,N_16097);
xnor U16271 (N_16271,N_16089,N_16115);
nor U16272 (N_16272,N_16032,N_16121);
or U16273 (N_16273,N_16028,N_16233);
xnor U16274 (N_16274,N_16033,N_16131);
nand U16275 (N_16275,N_16216,N_16120);
nand U16276 (N_16276,N_16047,N_16166);
and U16277 (N_16277,N_16150,N_16038);
nor U16278 (N_16278,N_16221,N_16141);
or U16279 (N_16279,N_16201,N_16134);
nor U16280 (N_16280,N_16171,N_16182);
xnor U16281 (N_16281,N_16136,N_16024);
nand U16282 (N_16282,N_16103,N_16054);
xnor U16283 (N_16283,N_16017,N_16023);
and U16284 (N_16284,N_16151,N_16016);
or U16285 (N_16285,N_16105,N_16142);
nand U16286 (N_16286,N_16067,N_16043);
and U16287 (N_16287,N_16183,N_16042);
xor U16288 (N_16288,N_16125,N_16178);
nor U16289 (N_16289,N_16027,N_16163);
nand U16290 (N_16290,N_16210,N_16118);
xnor U16291 (N_16291,N_16104,N_16245);
xnor U16292 (N_16292,N_16167,N_16138);
xor U16293 (N_16293,N_16040,N_16227);
and U16294 (N_16294,N_16108,N_16082);
xnor U16295 (N_16295,N_16235,N_16096);
nor U16296 (N_16296,N_16080,N_16062);
and U16297 (N_16297,N_16231,N_16092);
nand U16298 (N_16298,N_16061,N_16113);
nor U16299 (N_16299,N_16168,N_16075);
or U16300 (N_16300,N_16205,N_16145);
nor U16301 (N_16301,N_16222,N_16155);
nand U16302 (N_16302,N_16034,N_16013);
nor U16303 (N_16303,N_16177,N_16091);
nand U16304 (N_16304,N_16186,N_16109);
or U16305 (N_16305,N_16132,N_16191);
nand U16306 (N_16306,N_16226,N_16060);
or U16307 (N_16307,N_16051,N_16162);
nor U16308 (N_16308,N_16022,N_16006);
and U16309 (N_16309,N_16010,N_16035);
or U16310 (N_16310,N_16139,N_16190);
and U16311 (N_16311,N_16057,N_16137);
or U16312 (N_16312,N_16204,N_16159);
xnor U16313 (N_16313,N_16111,N_16173);
xnor U16314 (N_16314,N_16146,N_16143);
nor U16315 (N_16315,N_16238,N_16041);
or U16316 (N_16316,N_16181,N_16037);
or U16317 (N_16317,N_16246,N_16126);
nand U16318 (N_16318,N_16036,N_16225);
nor U16319 (N_16319,N_16058,N_16208);
or U16320 (N_16320,N_16209,N_16128);
xor U16321 (N_16321,N_16189,N_16081);
nor U16322 (N_16322,N_16211,N_16176);
or U16323 (N_16323,N_16207,N_16000);
and U16324 (N_16324,N_16188,N_16203);
or U16325 (N_16325,N_16077,N_16242);
and U16326 (N_16326,N_16165,N_16117);
nand U16327 (N_16327,N_16011,N_16107);
or U16328 (N_16328,N_16224,N_16232);
nor U16329 (N_16329,N_16002,N_16172);
and U16330 (N_16330,N_16086,N_16001);
xnor U16331 (N_16331,N_16088,N_16192);
nor U16332 (N_16332,N_16073,N_16196);
or U16333 (N_16333,N_16021,N_16187);
xor U16334 (N_16334,N_16070,N_16193);
nand U16335 (N_16335,N_16084,N_16243);
and U16336 (N_16336,N_16099,N_16130);
and U16337 (N_16337,N_16087,N_16179);
nor U16338 (N_16338,N_16056,N_16064);
nand U16339 (N_16339,N_16247,N_16029);
xor U16340 (N_16340,N_16019,N_16170);
and U16341 (N_16341,N_16116,N_16133);
or U16342 (N_16342,N_16180,N_16239);
xor U16343 (N_16343,N_16025,N_16129);
nor U16344 (N_16344,N_16110,N_16114);
nor U16345 (N_16345,N_16161,N_16102);
nor U16346 (N_16346,N_16152,N_16175);
nand U16347 (N_16347,N_16199,N_16147);
and U16348 (N_16348,N_16174,N_16240);
nor U16349 (N_16349,N_16220,N_16249);
nand U16350 (N_16350,N_16195,N_16059);
xor U16351 (N_16351,N_16053,N_16050);
xor U16352 (N_16352,N_16148,N_16074);
or U16353 (N_16353,N_16214,N_16158);
or U16354 (N_16354,N_16234,N_16197);
or U16355 (N_16355,N_16124,N_16083);
nor U16356 (N_16356,N_16045,N_16112);
or U16357 (N_16357,N_16215,N_16123);
nand U16358 (N_16358,N_16046,N_16007);
nor U16359 (N_16359,N_16185,N_16202);
nand U16360 (N_16360,N_16098,N_16244);
xnor U16361 (N_16361,N_16004,N_16237);
and U16362 (N_16362,N_16066,N_16241);
nor U16363 (N_16363,N_16223,N_16085);
nand U16364 (N_16364,N_16009,N_16154);
nand U16365 (N_16365,N_16230,N_16101);
nor U16366 (N_16366,N_16063,N_16055);
nand U16367 (N_16367,N_16236,N_16048);
nor U16368 (N_16368,N_16219,N_16093);
or U16369 (N_16369,N_16144,N_16030);
or U16370 (N_16370,N_16094,N_16005);
or U16371 (N_16371,N_16012,N_16044);
xor U16372 (N_16372,N_16076,N_16039);
or U16373 (N_16373,N_16248,N_16169);
nand U16374 (N_16374,N_16194,N_16095);
or U16375 (N_16375,N_16031,N_16207);
and U16376 (N_16376,N_16079,N_16141);
nor U16377 (N_16377,N_16094,N_16074);
or U16378 (N_16378,N_16235,N_16005);
or U16379 (N_16379,N_16051,N_16155);
or U16380 (N_16380,N_16199,N_16236);
and U16381 (N_16381,N_16143,N_16072);
nand U16382 (N_16382,N_16108,N_16016);
nand U16383 (N_16383,N_16197,N_16091);
and U16384 (N_16384,N_16028,N_16045);
xnor U16385 (N_16385,N_16150,N_16197);
and U16386 (N_16386,N_16007,N_16123);
nand U16387 (N_16387,N_16113,N_16121);
xnor U16388 (N_16388,N_16121,N_16145);
and U16389 (N_16389,N_16218,N_16180);
and U16390 (N_16390,N_16061,N_16129);
or U16391 (N_16391,N_16227,N_16096);
and U16392 (N_16392,N_16248,N_16098);
xor U16393 (N_16393,N_16179,N_16219);
nor U16394 (N_16394,N_16210,N_16101);
nand U16395 (N_16395,N_16237,N_16030);
xnor U16396 (N_16396,N_16068,N_16097);
or U16397 (N_16397,N_16161,N_16023);
nand U16398 (N_16398,N_16050,N_16037);
nor U16399 (N_16399,N_16237,N_16152);
nand U16400 (N_16400,N_16097,N_16247);
and U16401 (N_16401,N_16125,N_16030);
or U16402 (N_16402,N_16026,N_16218);
and U16403 (N_16403,N_16030,N_16018);
or U16404 (N_16404,N_16246,N_16205);
nor U16405 (N_16405,N_16040,N_16023);
nand U16406 (N_16406,N_16134,N_16074);
xor U16407 (N_16407,N_16200,N_16067);
and U16408 (N_16408,N_16203,N_16212);
and U16409 (N_16409,N_16161,N_16047);
nand U16410 (N_16410,N_16235,N_16112);
or U16411 (N_16411,N_16024,N_16230);
nand U16412 (N_16412,N_16139,N_16129);
and U16413 (N_16413,N_16181,N_16164);
or U16414 (N_16414,N_16121,N_16070);
or U16415 (N_16415,N_16120,N_16241);
or U16416 (N_16416,N_16006,N_16129);
nor U16417 (N_16417,N_16047,N_16035);
xnor U16418 (N_16418,N_16104,N_16004);
or U16419 (N_16419,N_16192,N_16175);
or U16420 (N_16420,N_16049,N_16066);
nor U16421 (N_16421,N_16092,N_16202);
and U16422 (N_16422,N_16141,N_16199);
or U16423 (N_16423,N_16058,N_16068);
or U16424 (N_16424,N_16057,N_16004);
and U16425 (N_16425,N_16237,N_16230);
xor U16426 (N_16426,N_16056,N_16099);
and U16427 (N_16427,N_16190,N_16238);
or U16428 (N_16428,N_16054,N_16219);
nand U16429 (N_16429,N_16198,N_16166);
nor U16430 (N_16430,N_16041,N_16017);
xor U16431 (N_16431,N_16217,N_16076);
or U16432 (N_16432,N_16016,N_16005);
xnor U16433 (N_16433,N_16074,N_16099);
and U16434 (N_16434,N_16080,N_16247);
or U16435 (N_16435,N_16217,N_16145);
xnor U16436 (N_16436,N_16122,N_16030);
or U16437 (N_16437,N_16139,N_16085);
nor U16438 (N_16438,N_16180,N_16048);
or U16439 (N_16439,N_16008,N_16027);
nor U16440 (N_16440,N_16164,N_16187);
or U16441 (N_16441,N_16094,N_16156);
or U16442 (N_16442,N_16019,N_16107);
and U16443 (N_16443,N_16111,N_16203);
nor U16444 (N_16444,N_16245,N_16185);
and U16445 (N_16445,N_16157,N_16187);
and U16446 (N_16446,N_16172,N_16234);
xor U16447 (N_16447,N_16222,N_16021);
xnor U16448 (N_16448,N_16238,N_16032);
and U16449 (N_16449,N_16078,N_16092);
xor U16450 (N_16450,N_16187,N_16194);
nor U16451 (N_16451,N_16028,N_16135);
xor U16452 (N_16452,N_16183,N_16137);
and U16453 (N_16453,N_16103,N_16081);
xor U16454 (N_16454,N_16155,N_16024);
nand U16455 (N_16455,N_16157,N_16110);
nor U16456 (N_16456,N_16037,N_16030);
and U16457 (N_16457,N_16022,N_16192);
or U16458 (N_16458,N_16167,N_16065);
nor U16459 (N_16459,N_16181,N_16245);
xor U16460 (N_16460,N_16124,N_16134);
and U16461 (N_16461,N_16234,N_16103);
nand U16462 (N_16462,N_16238,N_16146);
xnor U16463 (N_16463,N_16170,N_16165);
or U16464 (N_16464,N_16190,N_16145);
xor U16465 (N_16465,N_16001,N_16248);
nor U16466 (N_16466,N_16176,N_16101);
or U16467 (N_16467,N_16201,N_16017);
xnor U16468 (N_16468,N_16005,N_16035);
nor U16469 (N_16469,N_16248,N_16074);
nand U16470 (N_16470,N_16084,N_16187);
nand U16471 (N_16471,N_16098,N_16023);
nand U16472 (N_16472,N_16236,N_16220);
and U16473 (N_16473,N_16132,N_16124);
xnor U16474 (N_16474,N_16016,N_16064);
or U16475 (N_16475,N_16211,N_16021);
nor U16476 (N_16476,N_16079,N_16108);
nor U16477 (N_16477,N_16173,N_16148);
nor U16478 (N_16478,N_16114,N_16078);
nor U16479 (N_16479,N_16179,N_16188);
nand U16480 (N_16480,N_16016,N_16053);
and U16481 (N_16481,N_16100,N_16187);
and U16482 (N_16482,N_16192,N_16154);
or U16483 (N_16483,N_16030,N_16119);
or U16484 (N_16484,N_16004,N_16002);
and U16485 (N_16485,N_16096,N_16005);
nand U16486 (N_16486,N_16022,N_16063);
or U16487 (N_16487,N_16236,N_16181);
and U16488 (N_16488,N_16102,N_16024);
nor U16489 (N_16489,N_16249,N_16164);
xnor U16490 (N_16490,N_16017,N_16249);
xnor U16491 (N_16491,N_16197,N_16214);
and U16492 (N_16492,N_16001,N_16099);
nor U16493 (N_16493,N_16177,N_16090);
nor U16494 (N_16494,N_16159,N_16157);
and U16495 (N_16495,N_16148,N_16054);
or U16496 (N_16496,N_16139,N_16200);
and U16497 (N_16497,N_16099,N_16196);
nand U16498 (N_16498,N_16099,N_16146);
nor U16499 (N_16499,N_16014,N_16237);
nor U16500 (N_16500,N_16266,N_16393);
or U16501 (N_16501,N_16488,N_16495);
nand U16502 (N_16502,N_16477,N_16387);
nor U16503 (N_16503,N_16327,N_16290);
xnor U16504 (N_16504,N_16317,N_16499);
nand U16505 (N_16505,N_16255,N_16334);
nand U16506 (N_16506,N_16490,N_16275);
xor U16507 (N_16507,N_16367,N_16457);
nand U16508 (N_16508,N_16383,N_16453);
and U16509 (N_16509,N_16464,N_16368);
xnor U16510 (N_16510,N_16376,N_16395);
nor U16511 (N_16511,N_16330,N_16372);
nand U16512 (N_16512,N_16413,N_16469);
and U16513 (N_16513,N_16314,N_16468);
nand U16514 (N_16514,N_16251,N_16265);
and U16515 (N_16515,N_16373,N_16284);
nor U16516 (N_16516,N_16369,N_16320);
or U16517 (N_16517,N_16305,N_16342);
nor U16518 (N_16518,N_16482,N_16260);
or U16519 (N_16519,N_16288,N_16353);
and U16520 (N_16520,N_16461,N_16313);
xnor U16521 (N_16521,N_16474,N_16388);
xor U16522 (N_16522,N_16385,N_16308);
nand U16523 (N_16523,N_16358,N_16448);
nor U16524 (N_16524,N_16264,N_16311);
and U16525 (N_16525,N_16422,N_16412);
nand U16526 (N_16526,N_16401,N_16352);
nand U16527 (N_16527,N_16269,N_16476);
nand U16528 (N_16528,N_16390,N_16472);
and U16529 (N_16529,N_16494,N_16470);
or U16530 (N_16530,N_16431,N_16278);
nor U16531 (N_16531,N_16392,N_16487);
nand U16532 (N_16532,N_16349,N_16359);
and U16533 (N_16533,N_16415,N_16440);
and U16534 (N_16534,N_16366,N_16295);
and U16535 (N_16535,N_16259,N_16449);
nor U16536 (N_16536,N_16341,N_16414);
xor U16537 (N_16537,N_16492,N_16460);
xor U16538 (N_16538,N_16377,N_16426);
nand U16539 (N_16539,N_16454,N_16261);
xor U16540 (N_16540,N_16362,N_16384);
xnor U16541 (N_16541,N_16346,N_16434);
or U16542 (N_16542,N_16455,N_16458);
xor U16543 (N_16543,N_16445,N_16354);
xor U16544 (N_16544,N_16298,N_16277);
nor U16545 (N_16545,N_16273,N_16348);
nor U16546 (N_16546,N_16361,N_16439);
and U16547 (N_16547,N_16322,N_16340);
or U16548 (N_16548,N_16452,N_16436);
or U16549 (N_16549,N_16344,N_16382);
nor U16550 (N_16550,N_16258,N_16296);
xor U16551 (N_16551,N_16307,N_16420);
and U16552 (N_16552,N_16299,N_16312);
and U16553 (N_16553,N_16475,N_16425);
nand U16554 (N_16554,N_16355,N_16394);
nor U16555 (N_16555,N_16432,N_16318);
or U16556 (N_16556,N_16337,N_16428);
nand U16557 (N_16557,N_16484,N_16329);
or U16558 (N_16558,N_16302,N_16315);
nor U16559 (N_16559,N_16467,N_16304);
nand U16560 (N_16560,N_16316,N_16252);
nand U16561 (N_16561,N_16417,N_16423);
nand U16562 (N_16562,N_16250,N_16292);
or U16563 (N_16563,N_16380,N_16424);
xnor U16564 (N_16564,N_16447,N_16410);
or U16565 (N_16565,N_16291,N_16399);
xor U16566 (N_16566,N_16371,N_16491);
and U16567 (N_16567,N_16286,N_16324);
and U16568 (N_16568,N_16350,N_16381);
or U16569 (N_16569,N_16407,N_16360);
nand U16570 (N_16570,N_16421,N_16272);
nor U16571 (N_16571,N_16374,N_16450);
nor U16572 (N_16572,N_16441,N_16282);
or U16573 (N_16573,N_16435,N_16416);
or U16574 (N_16574,N_16486,N_16325);
and U16575 (N_16575,N_16283,N_16375);
and U16576 (N_16576,N_16333,N_16411);
nor U16577 (N_16577,N_16306,N_16444);
or U16578 (N_16578,N_16293,N_16479);
or U16579 (N_16579,N_16338,N_16336);
nor U16580 (N_16580,N_16357,N_16498);
nand U16581 (N_16581,N_16281,N_16285);
xor U16582 (N_16582,N_16271,N_16493);
and U16583 (N_16583,N_16427,N_16267);
xnor U16584 (N_16584,N_16268,N_16321);
nor U16585 (N_16585,N_16347,N_16465);
nor U16586 (N_16586,N_16398,N_16339);
nand U16587 (N_16587,N_16433,N_16300);
xnor U16588 (N_16588,N_16456,N_16473);
or U16589 (N_16589,N_16309,N_16471);
or U16590 (N_16590,N_16262,N_16451);
nand U16591 (N_16591,N_16328,N_16345);
or U16592 (N_16592,N_16481,N_16497);
nor U16593 (N_16593,N_16326,N_16364);
nor U16594 (N_16594,N_16496,N_16378);
nand U16595 (N_16595,N_16438,N_16332);
xnor U16596 (N_16596,N_16405,N_16463);
xnor U16597 (N_16597,N_16418,N_16370);
nand U16598 (N_16598,N_16301,N_16396);
or U16599 (N_16599,N_16442,N_16429);
nor U16600 (N_16600,N_16403,N_16483);
and U16601 (N_16601,N_16256,N_16404);
and U16602 (N_16602,N_16386,N_16419);
nand U16603 (N_16603,N_16446,N_16489);
nor U16604 (N_16604,N_16279,N_16485);
nand U16605 (N_16605,N_16294,N_16356);
xnor U16606 (N_16606,N_16257,N_16287);
or U16607 (N_16607,N_16319,N_16303);
xor U16608 (N_16608,N_16466,N_16408);
and U16609 (N_16609,N_16443,N_16430);
nor U16610 (N_16610,N_16363,N_16343);
nor U16611 (N_16611,N_16274,N_16402);
xnor U16612 (N_16612,N_16437,N_16406);
xnor U16613 (N_16613,N_16254,N_16389);
and U16614 (N_16614,N_16310,N_16379);
xnor U16615 (N_16615,N_16478,N_16459);
or U16616 (N_16616,N_16297,N_16397);
and U16617 (N_16617,N_16331,N_16253);
xor U16618 (N_16618,N_16365,N_16280);
xor U16619 (N_16619,N_16289,N_16462);
and U16620 (N_16620,N_16351,N_16276);
nand U16621 (N_16621,N_16391,N_16323);
xnor U16622 (N_16622,N_16409,N_16270);
nand U16623 (N_16623,N_16480,N_16335);
xnor U16624 (N_16624,N_16400,N_16263);
or U16625 (N_16625,N_16268,N_16257);
or U16626 (N_16626,N_16311,N_16396);
xor U16627 (N_16627,N_16312,N_16297);
nor U16628 (N_16628,N_16407,N_16379);
xor U16629 (N_16629,N_16398,N_16271);
xor U16630 (N_16630,N_16274,N_16319);
nand U16631 (N_16631,N_16485,N_16381);
nand U16632 (N_16632,N_16486,N_16438);
xor U16633 (N_16633,N_16434,N_16464);
nor U16634 (N_16634,N_16325,N_16438);
or U16635 (N_16635,N_16463,N_16387);
xnor U16636 (N_16636,N_16294,N_16329);
xnor U16637 (N_16637,N_16286,N_16414);
nor U16638 (N_16638,N_16289,N_16493);
nand U16639 (N_16639,N_16250,N_16366);
and U16640 (N_16640,N_16314,N_16382);
or U16641 (N_16641,N_16435,N_16384);
or U16642 (N_16642,N_16426,N_16340);
nand U16643 (N_16643,N_16259,N_16453);
nand U16644 (N_16644,N_16383,N_16488);
nor U16645 (N_16645,N_16477,N_16461);
or U16646 (N_16646,N_16283,N_16367);
nand U16647 (N_16647,N_16333,N_16425);
or U16648 (N_16648,N_16420,N_16261);
and U16649 (N_16649,N_16342,N_16445);
nand U16650 (N_16650,N_16333,N_16364);
and U16651 (N_16651,N_16424,N_16463);
nand U16652 (N_16652,N_16439,N_16314);
and U16653 (N_16653,N_16349,N_16469);
or U16654 (N_16654,N_16373,N_16418);
nor U16655 (N_16655,N_16468,N_16389);
xnor U16656 (N_16656,N_16275,N_16277);
xor U16657 (N_16657,N_16474,N_16410);
nor U16658 (N_16658,N_16291,N_16390);
or U16659 (N_16659,N_16256,N_16350);
nor U16660 (N_16660,N_16329,N_16358);
nor U16661 (N_16661,N_16364,N_16431);
nor U16662 (N_16662,N_16458,N_16414);
or U16663 (N_16663,N_16264,N_16282);
and U16664 (N_16664,N_16251,N_16330);
nand U16665 (N_16665,N_16250,N_16489);
or U16666 (N_16666,N_16331,N_16345);
or U16667 (N_16667,N_16456,N_16463);
nor U16668 (N_16668,N_16284,N_16422);
nor U16669 (N_16669,N_16252,N_16319);
nor U16670 (N_16670,N_16388,N_16393);
and U16671 (N_16671,N_16326,N_16436);
xnor U16672 (N_16672,N_16385,N_16432);
and U16673 (N_16673,N_16466,N_16393);
nor U16674 (N_16674,N_16302,N_16272);
and U16675 (N_16675,N_16451,N_16271);
xnor U16676 (N_16676,N_16344,N_16427);
and U16677 (N_16677,N_16465,N_16381);
xnor U16678 (N_16678,N_16397,N_16283);
nand U16679 (N_16679,N_16451,N_16351);
nand U16680 (N_16680,N_16407,N_16384);
nor U16681 (N_16681,N_16388,N_16305);
xor U16682 (N_16682,N_16309,N_16469);
or U16683 (N_16683,N_16388,N_16259);
xnor U16684 (N_16684,N_16351,N_16491);
nor U16685 (N_16685,N_16450,N_16329);
nor U16686 (N_16686,N_16361,N_16408);
or U16687 (N_16687,N_16499,N_16253);
or U16688 (N_16688,N_16314,N_16263);
or U16689 (N_16689,N_16324,N_16451);
and U16690 (N_16690,N_16296,N_16489);
and U16691 (N_16691,N_16370,N_16459);
or U16692 (N_16692,N_16413,N_16292);
or U16693 (N_16693,N_16321,N_16299);
and U16694 (N_16694,N_16458,N_16262);
and U16695 (N_16695,N_16395,N_16265);
or U16696 (N_16696,N_16265,N_16432);
or U16697 (N_16697,N_16323,N_16404);
or U16698 (N_16698,N_16327,N_16392);
and U16699 (N_16699,N_16346,N_16292);
nand U16700 (N_16700,N_16283,N_16494);
nor U16701 (N_16701,N_16447,N_16281);
and U16702 (N_16702,N_16276,N_16284);
nand U16703 (N_16703,N_16315,N_16499);
or U16704 (N_16704,N_16447,N_16437);
and U16705 (N_16705,N_16437,N_16486);
xor U16706 (N_16706,N_16465,N_16487);
nor U16707 (N_16707,N_16416,N_16362);
xor U16708 (N_16708,N_16430,N_16384);
or U16709 (N_16709,N_16367,N_16424);
or U16710 (N_16710,N_16293,N_16290);
nand U16711 (N_16711,N_16404,N_16271);
nor U16712 (N_16712,N_16327,N_16467);
nand U16713 (N_16713,N_16492,N_16253);
xor U16714 (N_16714,N_16285,N_16339);
xor U16715 (N_16715,N_16404,N_16259);
nor U16716 (N_16716,N_16456,N_16387);
nand U16717 (N_16717,N_16429,N_16415);
nand U16718 (N_16718,N_16445,N_16317);
nand U16719 (N_16719,N_16272,N_16429);
and U16720 (N_16720,N_16470,N_16359);
nand U16721 (N_16721,N_16425,N_16458);
nand U16722 (N_16722,N_16423,N_16449);
nand U16723 (N_16723,N_16387,N_16346);
nand U16724 (N_16724,N_16284,N_16281);
and U16725 (N_16725,N_16307,N_16436);
nand U16726 (N_16726,N_16403,N_16433);
nand U16727 (N_16727,N_16310,N_16262);
xnor U16728 (N_16728,N_16472,N_16316);
nand U16729 (N_16729,N_16327,N_16494);
nor U16730 (N_16730,N_16411,N_16379);
nand U16731 (N_16731,N_16335,N_16281);
xor U16732 (N_16732,N_16336,N_16293);
nand U16733 (N_16733,N_16260,N_16308);
xor U16734 (N_16734,N_16485,N_16368);
and U16735 (N_16735,N_16302,N_16402);
nand U16736 (N_16736,N_16377,N_16491);
nand U16737 (N_16737,N_16482,N_16371);
and U16738 (N_16738,N_16488,N_16448);
nor U16739 (N_16739,N_16273,N_16349);
and U16740 (N_16740,N_16488,N_16355);
xor U16741 (N_16741,N_16255,N_16268);
and U16742 (N_16742,N_16456,N_16496);
or U16743 (N_16743,N_16497,N_16392);
or U16744 (N_16744,N_16349,N_16252);
nor U16745 (N_16745,N_16488,N_16362);
xnor U16746 (N_16746,N_16280,N_16389);
and U16747 (N_16747,N_16327,N_16490);
xor U16748 (N_16748,N_16254,N_16293);
and U16749 (N_16749,N_16368,N_16477);
or U16750 (N_16750,N_16643,N_16538);
and U16751 (N_16751,N_16715,N_16630);
nand U16752 (N_16752,N_16682,N_16558);
and U16753 (N_16753,N_16541,N_16520);
or U16754 (N_16754,N_16650,N_16598);
or U16755 (N_16755,N_16585,N_16512);
xnor U16756 (N_16756,N_16664,N_16610);
nor U16757 (N_16757,N_16724,N_16572);
and U16758 (N_16758,N_16640,N_16513);
nor U16759 (N_16759,N_16644,N_16668);
or U16760 (N_16760,N_16613,N_16564);
nand U16761 (N_16761,N_16674,N_16569);
nor U16762 (N_16762,N_16661,N_16626);
nor U16763 (N_16763,N_16500,N_16739);
nand U16764 (N_16764,N_16575,N_16502);
nor U16765 (N_16765,N_16718,N_16593);
nor U16766 (N_16766,N_16720,N_16628);
nor U16767 (N_16767,N_16709,N_16698);
nand U16768 (N_16768,N_16607,N_16605);
and U16769 (N_16769,N_16586,N_16740);
nor U16770 (N_16770,N_16537,N_16536);
nand U16771 (N_16771,N_16527,N_16596);
xnor U16772 (N_16772,N_16648,N_16702);
nor U16773 (N_16773,N_16595,N_16686);
nand U16774 (N_16774,N_16691,N_16620);
nor U16775 (N_16775,N_16559,N_16714);
or U16776 (N_16776,N_16694,N_16529);
nand U16777 (N_16777,N_16647,N_16567);
nand U16778 (N_16778,N_16562,N_16649);
xnor U16779 (N_16779,N_16543,N_16684);
and U16780 (N_16780,N_16568,N_16514);
nand U16781 (N_16781,N_16723,N_16540);
nor U16782 (N_16782,N_16518,N_16544);
nor U16783 (N_16783,N_16515,N_16574);
or U16784 (N_16784,N_16652,N_16546);
nor U16785 (N_16785,N_16528,N_16534);
nor U16786 (N_16786,N_16573,N_16614);
nand U16787 (N_16787,N_16659,N_16639);
or U16788 (N_16788,N_16676,N_16744);
xor U16789 (N_16789,N_16632,N_16616);
nor U16790 (N_16790,N_16594,N_16547);
nor U16791 (N_16791,N_16505,N_16622);
nand U16792 (N_16792,N_16583,N_16557);
and U16793 (N_16793,N_16703,N_16654);
and U16794 (N_16794,N_16587,N_16716);
or U16795 (N_16795,N_16539,N_16623);
and U16796 (N_16796,N_16734,N_16641);
or U16797 (N_16797,N_16592,N_16705);
nand U16798 (N_16798,N_16679,N_16732);
and U16799 (N_16799,N_16629,N_16693);
nor U16800 (N_16800,N_16591,N_16516);
or U16801 (N_16801,N_16609,N_16554);
nand U16802 (N_16802,N_16600,N_16657);
or U16803 (N_16803,N_16711,N_16524);
and U16804 (N_16804,N_16503,N_16566);
nand U16805 (N_16805,N_16669,N_16673);
nor U16806 (N_16806,N_16701,N_16531);
and U16807 (N_16807,N_16656,N_16655);
nor U16808 (N_16808,N_16606,N_16700);
nor U16809 (N_16809,N_16506,N_16633);
and U16810 (N_16810,N_16725,N_16533);
xnor U16811 (N_16811,N_16508,N_16627);
nor U16812 (N_16812,N_16581,N_16578);
and U16813 (N_16813,N_16662,N_16667);
or U16814 (N_16814,N_16548,N_16708);
nor U16815 (N_16815,N_16742,N_16617);
nand U16816 (N_16816,N_16707,N_16683);
xnor U16817 (N_16817,N_16729,N_16571);
and U16818 (N_16818,N_16728,N_16699);
and U16819 (N_16819,N_16730,N_16560);
nand U16820 (N_16820,N_16618,N_16638);
xor U16821 (N_16821,N_16511,N_16692);
nand U16822 (N_16822,N_16553,N_16748);
nand U16823 (N_16823,N_16577,N_16555);
or U16824 (N_16824,N_16672,N_16646);
and U16825 (N_16825,N_16717,N_16675);
or U16826 (N_16826,N_16678,N_16565);
or U16827 (N_16827,N_16526,N_16521);
xor U16828 (N_16828,N_16738,N_16625);
and U16829 (N_16829,N_16525,N_16731);
nor U16830 (N_16830,N_16608,N_16737);
and U16831 (N_16831,N_16645,N_16580);
nor U16832 (N_16832,N_16597,N_16712);
xnor U16833 (N_16833,N_16749,N_16636);
or U16834 (N_16834,N_16519,N_16615);
or U16835 (N_16835,N_16579,N_16576);
xor U16836 (N_16836,N_16582,N_16552);
nor U16837 (N_16837,N_16726,N_16687);
nor U16838 (N_16838,N_16589,N_16670);
and U16839 (N_16839,N_16680,N_16507);
and U16840 (N_16840,N_16671,N_16721);
and U16841 (N_16841,N_16556,N_16660);
or U16842 (N_16842,N_16745,N_16601);
and U16843 (N_16843,N_16743,N_16746);
and U16844 (N_16844,N_16689,N_16619);
or U16845 (N_16845,N_16612,N_16602);
nand U16846 (N_16846,N_16570,N_16501);
nor U16847 (N_16847,N_16747,N_16510);
and U16848 (N_16848,N_16697,N_16706);
xnor U16849 (N_16849,N_16663,N_16517);
nand U16850 (N_16850,N_16713,N_16530);
nand U16851 (N_16851,N_16635,N_16685);
xnor U16852 (N_16852,N_16621,N_16523);
or U16853 (N_16853,N_16653,N_16551);
nor U16854 (N_16854,N_16532,N_16561);
nor U16855 (N_16855,N_16603,N_16563);
xnor U16856 (N_16856,N_16722,N_16509);
xnor U16857 (N_16857,N_16666,N_16611);
or U16858 (N_16858,N_16665,N_16677);
nor U16859 (N_16859,N_16658,N_16704);
nor U16860 (N_16860,N_16549,N_16634);
xor U16861 (N_16861,N_16642,N_16542);
nand U16862 (N_16862,N_16736,N_16624);
nand U16863 (N_16863,N_16599,N_16545);
and U16864 (N_16864,N_16604,N_16584);
or U16865 (N_16865,N_16631,N_16695);
nand U16866 (N_16866,N_16535,N_16504);
xnor U16867 (N_16867,N_16588,N_16550);
or U16868 (N_16868,N_16719,N_16733);
nor U16869 (N_16869,N_16522,N_16590);
nand U16870 (N_16870,N_16710,N_16727);
nand U16871 (N_16871,N_16681,N_16690);
nand U16872 (N_16872,N_16735,N_16651);
nand U16873 (N_16873,N_16637,N_16688);
or U16874 (N_16874,N_16741,N_16696);
nand U16875 (N_16875,N_16516,N_16712);
xor U16876 (N_16876,N_16659,N_16629);
nand U16877 (N_16877,N_16663,N_16666);
or U16878 (N_16878,N_16509,N_16556);
nor U16879 (N_16879,N_16728,N_16616);
or U16880 (N_16880,N_16728,N_16736);
nand U16881 (N_16881,N_16600,N_16585);
nand U16882 (N_16882,N_16562,N_16605);
xor U16883 (N_16883,N_16702,N_16518);
nand U16884 (N_16884,N_16668,N_16608);
nor U16885 (N_16885,N_16652,N_16506);
nand U16886 (N_16886,N_16617,N_16509);
and U16887 (N_16887,N_16510,N_16592);
or U16888 (N_16888,N_16682,N_16582);
or U16889 (N_16889,N_16661,N_16629);
xnor U16890 (N_16890,N_16539,N_16525);
and U16891 (N_16891,N_16528,N_16501);
xnor U16892 (N_16892,N_16719,N_16579);
nand U16893 (N_16893,N_16513,N_16611);
nor U16894 (N_16894,N_16700,N_16506);
nand U16895 (N_16895,N_16687,N_16539);
nor U16896 (N_16896,N_16642,N_16572);
nor U16897 (N_16897,N_16589,N_16689);
or U16898 (N_16898,N_16709,N_16599);
or U16899 (N_16899,N_16631,N_16579);
nand U16900 (N_16900,N_16735,N_16629);
and U16901 (N_16901,N_16544,N_16607);
nor U16902 (N_16902,N_16744,N_16535);
nor U16903 (N_16903,N_16607,N_16529);
and U16904 (N_16904,N_16739,N_16591);
or U16905 (N_16905,N_16614,N_16744);
xnor U16906 (N_16906,N_16696,N_16543);
xnor U16907 (N_16907,N_16707,N_16501);
and U16908 (N_16908,N_16582,N_16658);
and U16909 (N_16909,N_16540,N_16642);
nand U16910 (N_16910,N_16667,N_16535);
nor U16911 (N_16911,N_16540,N_16665);
and U16912 (N_16912,N_16611,N_16644);
nand U16913 (N_16913,N_16589,N_16681);
nand U16914 (N_16914,N_16609,N_16584);
nor U16915 (N_16915,N_16550,N_16743);
or U16916 (N_16916,N_16549,N_16511);
or U16917 (N_16917,N_16536,N_16735);
xor U16918 (N_16918,N_16710,N_16736);
nand U16919 (N_16919,N_16530,N_16546);
or U16920 (N_16920,N_16662,N_16527);
nand U16921 (N_16921,N_16577,N_16511);
nor U16922 (N_16922,N_16615,N_16678);
or U16923 (N_16923,N_16575,N_16726);
nor U16924 (N_16924,N_16588,N_16505);
xnor U16925 (N_16925,N_16708,N_16616);
nor U16926 (N_16926,N_16635,N_16519);
and U16927 (N_16927,N_16530,N_16584);
or U16928 (N_16928,N_16624,N_16552);
and U16929 (N_16929,N_16639,N_16669);
or U16930 (N_16930,N_16715,N_16742);
and U16931 (N_16931,N_16726,N_16724);
xnor U16932 (N_16932,N_16570,N_16705);
xor U16933 (N_16933,N_16666,N_16505);
nand U16934 (N_16934,N_16594,N_16722);
and U16935 (N_16935,N_16662,N_16608);
or U16936 (N_16936,N_16730,N_16599);
or U16937 (N_16937,N_16530,N_16601);
nor U16938 (N_16938,N_16666,N_16732);
nor U16939 (N_16939,N_16513,N_16658);
nand U16940 (N_16940,N_16719,N_16611);
nor U16941 (N_16941,N_16629,N_16707);
or U16942 (N_16942,N_16569,N_16714);
nand U16943 (N_16943,N_16666,N_16653);
xor U16944 (N_16944,N_16629,N_16634);
nor U16945 (N_16945,N_16588,N_16548);
xor U16946 (N_16946,N_16708,N_16505);
or U16947 (N_16947,N_16525,N_16642);
nand U16948 (N_16948,N_16626,N_16588);
and U16949 (N_16949,N_16519,N_16569);
and U16950 (N_16950,N_16501,N_16622);
nor U16951 (N_16951,N_16683,N_16657);
or U16952 (N_16952,N_16649,N_16695);
nand U16953 (N_16953,N_16635,N_16554);
nand U16954 (N_16954,N_16547,N_16608);
and U16955 (N_16955,N_16515,N_16712);
or U16956 (N_16956,N_16665,N_16512);
nand U16957 (N_16957,N_16525,N_16655);
or U16958 (N_16958,N_16671,N_16716);
or U16959 (N_16959,N_16640,N_16712);
xor U16960 (N_16960,N_16644,N_16607);
nand U16961 (N_16961,N_16683,N_16623);
nand U16962 (N_16962,N_16597,N_16675);
nand U16963 (N_16963,N_16617,N_16584);
nor U16964 (N_16964,N_16505,N_16690);
xnor U16965 (N_16965,N_16584,N_16662);
and U16966 (N_16966,N_16578,N_16686);
nor U16967 (N_16967,N_16541,N_16596);
nor U16968 (N_16968,N_16727,N_16611);
nor U16969 (N_16969,N_16510,N_16624);
and U16970 (N_16970,N_16661,N_16638);
or U16971 (N_16971,N_16565,N_16525);
xor U16972 (N_16972,N_16545,N_16558);
and U16973 (N_16973,N_16515,N_16682);
nand U16974 (N_16974,N_16578,N_16501);
xnor U16975 (N_16975,N_16617,N_16657);
or U16976 (N_16976,N_16697,N_16669);
nor U16977 (N_16977,N_16693,N_16624);
nor U16978 (N_16978,N_16673,N_16594);
or U16979 (N_16979,N_16663,N_16725);
and U16980 (N_16980,N_16605,N_16689);
xor U16981 (N_16981,N_16704,N_16620);
or U16982 (N_16982,N_16579,N_16745);
nor U16983 (N_16983,N_16568,N_16596);
nand U16984 (N_16984,N_16545,N_16560);
nor U16985 (N_16985,N_16737,N_16643);
or U16986 (N_16986,N_16630,N_16614);
and U16987 (N_16987,N_16684,N_16719);
and U16988 (N_16988,N_16660,N_16732);
or U16989 (N_16989,N_16685,N_16576);
xor U16990 (N_16990,N_16645,N_16615);
nand U16991 (N_16991,N_16694,N_16625);
xor U16992 (N_16992,N_16747,N_16558);
xor U16993 (N_16993,N_16695,N_16591);
or U16994 (N_16994,N_16598,N_16622);
and U16995 (N_16995,N_16715,N_16594);
or U16996 (N_16996,N_16748,N_16596);
nor U16997 (N_16997,N_16717,N_16524);
nor U16998 (N_16998,N_16554,N_16630);
nand U16999 (N_16999,N_16662,N_16594);
nand U17000 (N_17000,N_16802,N_16902);
nand U17001 (N_17001,N_16848,N_16897);
or U17002 (N_17002,N_16823,N_16800);
xor U17003 (N_17003,N_16986,N_16791);
or U17004 (N_17004,N_16813,N_16868);
and U17005 (N_17005,N_16947,N_16876);
xor U17006 (N_17006,N_16935,N_16937);
xnor U17007 (N_17007,N_16967,N_16846);
xor U17008 (N_17008,N_16932,N_16908);
or U17009 (N_17009,N_16867,N_16941);
or U17010 (N_17010,N_16923,N_16826);
nor U17011 (N_17011,N_16784,N_16753);
and U17012 (N_17012,N_16883,N_16994);
nand U17013 (N_17013,N_16936,N_16871);
and U17014 (N_17014,N_16801,N_16840);
and U17015 (N_17015,N_16879,N_16922);
nand U17016 (N_17016,N_16804,N_16837);
xnor U17017 (N_17017,N_16755,N_16828);
or U17018 (N_17018,N_16835,N_16825);
nor U17019 (N_17019,N_16955,N_16851);
and U17020 (N_17020,N_16914,N_16767);
nor U17021 (N_17021,N_16796,N_16950);
and U17022 (N_17022,N_16906,N_16963);
and U17023 (N_17023,N_16841,N_16987);
nand U17024 (N_17024,N_16903,N_16972);
nor U17025 (N_17025,N_16974,N_16977);
nor U17026 (N_17026,N_16930,N_16996);
nand U17027 (N_17027,N_16939,N_16872);
nand U17028 (N_17028,N_16949,N_16905);
and U17029 (N_17029,N_16777,N_16888);
and U17030 (N_17030,N_16951,N_16958);
nand U17031 (N_17031,N_16991,N_16865);
nor U17032 (N_17032,N_16863,N_16975);
nor U17033 (N_17033,N_16807,N_16772);
xnor U17034 (N_17034,N_16971,N_16790);
nand U17035 (N_17035,N_16761,N_16766);
nand U17036 (N_17036,N_16757,N_16944);
nand U17037 (N_17037,N_16797,N_16995);
and U17038 (N_17038,N_16833,N_16962);
and U17039 (N_17039,N_16758,N_16836);
or U17040 (N_17040,N_16857,N_16943);
xnor U17041 (N_17041,N_16893,N_16961);
nor U17042 (N_17042,N_16889,N_16969);
xor U17043 (N_17043,N_16859,N_16899);
nand U17044 (N_17044,N_16882,N_16829);
nor U17045 (N_17045,N_16763,N_16966);
or U17046 (N_17046,N_16811,N_16901);
or U17047 (N_17047,N_16979,N_16960);
nand U17048 (N_17048,N_16844,N_16860);
nand U17049 (N_17049,N_16822,N_16850);
nand U17050 (N_17050,N_16988,N_16843);
xor U17051 (N_17051,N_16812,N_16938);
nor U17052 (N_17052,N_16916,N_16895);
nand U17053 (N_17053,N_16849,N_16997);
and U17054 (N_17054,N_16983,N_16847);
and U17055 (N_17055,N_16978,N_16959);
and U17056 (N_17056,N_16984,N_16990);
and U17057 (N_17057,N_16752,N_16970);
or U17058 (N_17058,N_16781,N_16933);
xor U17059 (N_17059,N_16919,N_16892);
xor U17060 (N_17060,N_16830,N_16957);
xnor U17061 (N_17061,N_16915,N_16884);
nand U17062 (N_17062,N_16803,N_16946);
nor U17063 (N_17063,N_16779,N_16799);
or U17064 (N_17064,N_16775,N_16981);
or U17065 (N_17065,N_16982,N_16940);
nand U17066 (N_17066,N_16788,N_16819);
nor U17067 (N_17067,N_16810,N_16861);
nand U17068 (N_17068,N_16808,N_16998);
nor U17069 (N_17069,N_16900,N_16780);
xor U17070 (N_17070,N_16989,N_16824);
nor U17071 (N_17071,N_16934,N_16862);
xnor U17072 (N_17072,N_16965,N_16776);
or U17073 (N_17073,N_16818,N_16993);
nor U17074 (N_17074,N_16976,N_16948);
nand U17075 (N_17075,N_16855,N_16778);
or U17076 (N_17076,N_16842,N_16869);
or U17077 (N_17077,N_16853,N_16870);
nand U17078 (N_17078,N_16917,N_16792);
xnor U17079 (N_17079,N_16913,N_16839);
nor U17080 (N_17080,N_16890,N_16771);
nor U17081 (N_17081,N_16877,N_16827);
nor U17082 (N_17082,N_16911,N_16864);
nor U17083 (N_17083,N_16794,N_16815);
and U17084 (N_17084,N_16832,N_16785);
nor U17085 (N_17085,N_16821,N_16782);
nand U17086 (N_17086,N_16793,N_16956);
or U17087 (N_17087,N_16898,N_16927);
xor U17088 (N_17088,N_16954,N_16920);
or U17089 (N_17089,N_16945,N_16789);
nor U17090 (N_17090,N_16891,N_16968);
and U17091 (N_17091,N_16964,N_16931);
xnor U17092 (N_17092,N_16907,N_16875);
xor U17093 (N_17093,N_16786,N_16952);
or U17094 (N_17094,N_16760,N_16756);
nand U17095 (N_17095,N_16816,N_16754);
nand U17096 (N_17096,N_16904,N_16762);
and U17097 (N_17097,N_16838,N_16878);
nor U17098 (N_17098,N_16834,N_16942);
nand U17099 (N_17099,N_16874,N_16770);
nor U17100 (N_17100,N_16866,N_16924);
xnor U17101 (N_17101,N_16831,N_16751);
and U17102 (N_17102,N_16820,N_16980);
nor U17103 (N_17103,N_16929,N_16845);
xor U17104 (N_17104,N_16759,N_16928);
xor U17105 (N_17105,N_16881,N_16773);
nor U17106 (N_17106,N_16887,N_16910);
xor U17107 (N_17107,N_16750,N_16852);
nor U17108 (N_17108,N_16783,N_16894);
or U17109 (N_17109,N_16798,N_16774);
or U17110 (N_17110,N_16768,N_16953);
nor U17111 (N_17111,N_16896,N_16921);
xor U17112 (N_17112,N_16918,N_16814);
nand U17113 (N_17113,N_16912,N_16764);
and U17114 (N_17114,N_16854,N_16787);
nor U17115 (N_17115,N_16886,N_16858);
xnor U17116 (N_17116,N_16992,N_16909);
xor U17117 (N_17117,N_16925,N_16880);
nor U17118 (N_17118,N_16817,N_16806);
and U17119 (N_17119,N_16809,N_16973);
nor U17120 (N_17120,N_16885,N_16795);
or U17121 (N_17121,N_16765,N_16805);
xor U17122 (N_17122,N_16873,N_16999);
nand U17123 (N_17123,N_16926,N_16856);
xor U17124 (N_17124,N_16985,N_16769);
and U17125 (N_17125,N_16967,N_16924);
nand U17126 (N_17126,N_16987,N_16976);
and U17127 (N_17127,N_16811,N_16871);
nor U17128 (N_17128,N_16784,N_16904);
xor U17129 (N_17129,N_16819,N_16760);
and U17130 (N_17130,N_16945,N_16851);
or U17131 (N_17131,N_16835,N_16974);
and U17132 (N_17132,N_16988,N_16893);
xor U17133 (N_17133,N_16842,N_16838);
nand U17134 (N_17134,N_16934,N_16987);
xor U17135 (N_17135,N_16753,N_16866);
or U17136 (N_17136,N_16855,N_16875);
nand U17137 (N_17137,N_16984,N_16823);
xnor U17138 (N_17138,N_16915,N_16837);
xor U17139 (N_17139,N_16933,N_16777);
xnor U17140 (N_17140,N_16752,N_16814);
xnor U17141 (N_17141,N_16934,N_16851);
and U17142 (N_17142,N_16894,N_16983);
or U17143 (N_17143,N_16927,N_16903);
xnor U17144 (N_17144,N_16924,N_16938);
and U17145 (N_17145,N_16938,N_16877);
and U17146 (N_17146,N_16873,N_16842);
nor U17147 (N_17147,N_16974,N_16905);
nand U17148 (N_17148,N_16879,N_16877);
and U17149 (N_17149,N_16943,N_16833);
nor U17150 (N_17150,N_16996,N_16862);
nor U17151 (N_17151,N_16955,N_16951);
and U17152 (N_17152,N_16938,N_16927);
nand U17153 (N_17153,N_16939,N_16929);
xor U17154 (N_17154,N_16751,N_16885);
nand U17155 (N_17155,N_16843,N_16753);
xor U17156 (N_17156,N_16760,N_16863);
xnor U17157 (N_17157,N_16985,N_16823);
nor U17158 (N_17158,N_16997,N_16787);
or U17159 (N_17159,N_16785,N_16762);
xnor U17160 (N_17160,N_16963,N_16986);
xor U17161 (N_17161,N_16836,N_16904);
xnor U17162 (N_17162,N_16903,N_16957);
nor U17163 (N_17163,N_16818,N_16847);
nor U17164 (N_17164,N_16893,N_16867);
nand U17165 (N_17165,N_16919,N_16873);
nor U17166 (N_17166,N_16959,N_16818);
or U17167 (N_17167,N_16945,N_16817);
or U17168 (N_17168,N_16819,N_16853);
nand U17169 (N_17169,N_16869,N_16822);
xnor U17170 (N_17170,N_16834,N_16754);
xor U17171 (N_17171,N_16983,N_16941);
xor U17172 (N_17172,N_16766,N_16782);
nor U17173 (N_17173,N_16775,N_16786);
nor U17174 (N_17174,N_16816,N_16812);
nand U17175 (N_17175,N_16879,N_16785);
and U17176 (N_17176,N_16906,N_16846);
xnor U17177 (N_17177,N_16900,N_16987);
nand U17178 (N_17178,N_16833,N_16891);
or U17179 (N_17179,N_16833,N_16960);
or U17180 (N_17180,N_16871,N_16843);
or U17181 (N_17181,N_16790,N_16874);
xor U17182 (N_17182,N_16904,N_16997);
nand U17183 (N_17183,N_16924,N_16878);
xor U17184 (N_17184,N_16924,N_16850);
xnor U17185 (N_17185,N_16860,N_16758);
nor U17186 (N_17186,N_16820,N_16764);
and U17187 (N_17187,N_16910,N_16999);
and U17188 (N_17188,N_16915,N_16865);
nor U17189 (N_17189,N_16967,N_16921);
nand U17190 (N_17190,N_16884,N_16788);
and U17191 (N_17191,N_16935,N_16932);
and U17192 (N_17192,N_16882,N_16769);
xnor U17193 (N_17193,N_16901,N_16825);
nor U17194 (N_17194,N_16939,N_16976);
and U17195 (N_17195,N_16884,N_16772);
nand U17196 (N_17196,N_16934,N_16947);
xor U17197 (N_17197,N_16986,N_16750);
xnor U17198 (N_17198,N_16988,N_16875);
and U17199 (N_17199,N_16992,N_16785);
and U17200 (N_17200,N_16857,N_16848);
and U17201 (N_17201,N_16758,N_16791);
xor U17202 (N_17202,N_16989,N_16832);
nand U17203 (N_17203,N_16806,N_16871);
nand U17204 (N_17204,N_16941,N_16963);
or U17205 (N_17205,N_16842,N_16798);
or U17206 (N_17206,N_16915,N_16876);
nand U17207 (N_17207,N_16762,N_16796);
nor U17208 (N_17208,N_16850,N_16864);
nand U17209 (N_17209,N_16926,N_16769);
and U17210 (N_17210,N_16754,N_16896);
nand U17211 (N_17211,N_16870,N_16767);
or U17212 (N_17212,N_16914,N_16897);
nand U17213 (N_17213,N_16860,N_16871);
nand U17214 (N_17214,N_16836,N_16973);
nor U17215 (N_17215,N_16966,N_16832);
and U17216 (N_17216,N_16927,N_16886);
xnor U17217 (N_17217,N_16966,N_16783);
xor U17218 (N_17218,N_16773,N_16996);
xor U17219 (N_17219,N_16761,N_16770);
nand U17220 (N_17220,N_16760,N_16826);
or U17221 (N_17221,N_16816,N_16792);
or U17222 (N_17222,N_16751,N_16897);
xnor U17223 (N_17223,N_16909,N_16935);
xor U17224 (N_17224,N_16943,N_16826);
or U17225 (N_17225,N_16868,N_16801);
and U17226 (N_17226,N_16945,N_16850);
nor U17227 (N_17227,N_16794,N_16885);
xnor U17228 (N_17228,N_16918,N_16886);
or U17229 (N_17229,N_16911,N_16990);
or U17230 (N_17230,N_16937,N_16865);
and U17231 (N_17231,N_16850,N_16853);
and U17232 (N_17232,N_16755,N_16883);
or U17233 (N_17233,N_16945,N_16773);
or U17234 (N_17234,N_16772,N_16938);
nor U17235 (N_17235,N_16883,N_16995);
xnor U17236 (N_17236,N_16859,N_16952);
nand U17237 (N_17237,N_16817,N_16784);
and U17238 (N_17238,N_16928,N_16914);
or U17239 (N_17239,N_16938,N_16907);
xor U17240 (N_17240,N_16975,N_16756);
nand U17241 (N_17241,N_16867,N_16778);
xnor U17242 (N_17242,N_16791,N_16909);
xnor U17243 (N_17243,N_16976,N_16990);
xor U17244 (N_17244,N_16756,N_16944);
or U17245 (N_17245,N_16840,N_16954);
nor U17246 (N_17246,N_16916,N_16898);
nand U17247 (N_17247,N_16847,N_16778);
and U17248 (N_17248,N_16914,N_16789);
nand U17249 (N_17249,N_16914,N_16972);
and U17250 (N_17250,N_17053,N_17083);
xor U17251 (N_17251,N_17071,N_17206);
and U17252 (N_17252,N_17043,N_17248);
nor U17253 (N_17253,N_17190,N_17135);
xnor U17254 (N_17254,N_17088,N_17130);
nor U17255 (N_17255,N_17243,N_17075);
nand U17256 (N_17256,N_17225,N_17042);
nand U17257 (N_17257,N_17133,N_17119);
or U17258 (N_17258,N_17184,N_17163);
nand U17259 (N_17259,N_17087,N_17217);
nor U17260 (N_17260,N_17113,N_17047);
and U17261 (N_17261,N_17147,N_17199);
and U17262 (N_17262,N_17028,N_17126);
xor U17263 (N_17263,N_17162,N_17137);
nand U17264 (N_17264,N_17122,N_17139);
and U17265 (N_17265,N_17143,N_17121);
xnor U17266 (N_17266,N_17192,N_17068);
xnor U17267 (N_17267,N_17002,N_17213);
and U17268 (N_17268,N_17127,N_17156);
nor U17269 (N_17269,N_17164,N_17009);
nand U17270 (N_17270,N_17233,N_17165);
xor U17271 (N_17271,N_17107,N_17200);
xor U17272 (N_17272,N_17101,N_17161);
nor U17273 (N_17273,N_17040,N_17228);
nand U17274 (N_17274,N_17004,N_17136);
nor U17275 (N_17275,N_17021,N_17219);
and U17276 (N_17276,N_17099,N_17030);
nor U17277 (N_17277,N_17066,N_17237);
nor U17278 (N_17278,N_17058,N_17116);
xnor U17279 (N_17279,N_17191,N_17212);
nor U17280 (N_17280,N_17074,N_17044);
and U17281 (N_17281,N_17031,N_17017);
nand U17282 (N_17282,N_17229,N_17109);
and U17283 (N_17283,N_17026,N_17175);
nand U17284 (N_17284,N_17240,N_17239);
nand U17285 (N_17285,N_17020,N_17152);
or U17286 (N_17286,N_17061,N_17069);
or U17287 (N_17287,N_17179,N_17117);
nand U17288 (N_17288,N_17128,N_17157);
nor U17289 (N_17289,N_17180,N_17039);
nand U17290 (N_17290,N_17029,N_17102);
or U17291 (N_17291,N_17211,N_17096);
nor U17292 (N_17292,N_17059,N_17168);
and U17293 (N_17293,N_17106,N_17045);
nor U17294 (N_17294,N_17203,N_17024);
nand U17295 (N_17295,N_17145,N_17129);
nand U17296 (N_17296,N_17006,N_17226);
nand U17297 (N_17297,N_17158,N_17073);
nand U17298 (N_17298,N_17245,N_17110);
and U17299 (N_17299,N_17159,N_17111);
and U17300 (N_17300,N_17005,N_17100);
xnor U17301 (N_17301,N_17052,N_17064);
or U17302 (N_17302,N_17197,N_17124);
xnor U17303 (N_17303,N_17003,N_17172);
nand U17304 (N_17304,N_17085,N_17012);
xor U17305 (N_17305,N_17169,N_17167);
and U17306 (N_17306,N_17097,N_17132);
or U17307 (N_17307,N_17041,N_17019);
and U17308 (N_17308,N_17193,N_17105);
xor U17309 (N_17309,N_17176,N_17092);
nor U17310 (N_17310,N_17185,N_17247);
nor U17311 (N_17311,N_17234,N_17181);
nand U17312 (N_17312,N_17142,N_17242);
xor U17313 (N_17313,N_17236,N_17218);
xor U17314 (N_17314,N_17010,N_17013);
and U17315 (N_17315,N_17027,N_17151);
nand U17316 (N_17316,N_17249,N_17155);
nand U17317 (N_17317,N_17120,N_17238);
nor U17318 (N_17318,N_17186,N_17048);
xnor U17319 (N_17319,N_17008,N_17204);
or U17320 (N_17320,N_17150,N_17063);
xnor U17321 (N_17321,N_17050,N_17149);
or U17322 (N_17322,N_17207,N_17093);
nand U17323 (N_17323,N_17223,N_17138);
or U17324 (N_17324,N_17195,N_17216);
nand U17325 (N_17325,N_17174,N_17095);
or U17326 (N_17326,N_17070,N_17221);
nor U17327 (N_17327,N_17182,N_17170);
xnor U17328 (N_17328,N_17046,N_17015);
nand U17329 (N_17329,N_17177,N_17072);
xnor U17330 (N_17330,N_17079,N_17062);
and U17331 (N_17331,N_17224,N_17115);
nor U17332 (N_17332,N_17194,N_17057);
nor U17333 (N_17333,N_17104,N_17210);
nor U17334 (N_17334,N_17077,N_17188);
nand U17335 (N_17335,N_17198,N_17108);
nor U17336 (N_17336,N_17160,N_17178);
nand U17337 (N_17337,N_17067,N_17140);
and U17338 (N_17338,N_17022,N_17166);
and U17339 (N_17339,N_17246,N_17000);
nand U17340 (N_17340,N_17094,N_17034);
nand U17341 (N_17341,N_17011,N_17227);
xor U17342 (N_17342,N_17001,N_17146);
nor U17343 (N_17343,N_17016,N_17038);
or U17344 (N_17344,N_17018,N_17214);
nor U17345 (N_17345,N_17084,N_17209);
xnor U17346 (N_17346,N_17208,N_17118);
and U17347 (N_17347,N_17196,N_17187);
nor U17348 (N_17348,N_17103,N_17076);
or U17349 (N_17349,N_17037,N_17086);
nor U17350 (N_17350,N_17056,N_17241);
or U17351 (N_17351,N_17141,N_17078);
nor U17352 (N_17352,N_17089,N_17035);
xnor U17353 (N_17353,N_17205,N_17049);
xor U17354 (N_17354,N_17183,N_17114);
nor U17355 (N_17355,N_17014,N_17222);
or U17356 (N_17356,N_17082,N_17051);
nor U17357 (N_17357,N_17230,N_17144);
or U17358 (N_17358,N_17033,N_17007);
or U17359 (N_17359,N_17060,N_17131);
nand U17360 (N_17360,N_17215,N_17134);
or U17361 (N_17361,N_17153,N_17081);
nand U17362 (N_17362,N_17080,N_17202);
or U17363 (N_17363,N_17171,N_17148);
and U17364 (N_17364,N_17025,N_17231);
and U17365 (N_17365,N_17189,N_17090);
xnor U17366 (N_17366,N_17123,N_17244);
and U17367 (N_17367,N_17112,N_17055);
nand U17368 (N_17368,N_17154,N_17235);
nand U17369 (N_17369,N_17232,N_17201);
nand U17370 (N_17370,N_17091,N_17036);
and U17371 (N_17371,N_17023,N_17173);
nand U17372 (N_17372,N_17098,N_17220);
and U17373 (N_17373,N_17065,N_17054);
nand U17374 (N_17374,N_17125,N_17032);
and U17375 (N_17375,N_17139,N_17131);
or U17376 (N_17376,N_17011,N_17190);
nand U17377 (N_17377,N_17064,N_17106);
nand U17378 (N_17378,N_17107,N_17242);
nand U17379 (N_17379,N_17081,N_17072);
and U17380 (N_17380,N_17102,N_17062);
or U17381 (N_17381,N_17084,N_17241);
or U17382 (N_17382,N_17223,N_17242);
or U17383 (N_17383,N_17197,N_17105);
nand U17384 (N_17384,N_17078,N_17006);
nand U17385 (N_17385,N_17086,N_17057);
and U17386 (N_17386,N_17010,N_17046);
nand U17387 (N_17387,N_17030,N_17206);
xnor U17388 (N_17388,N_17239,N_17111);
nand U17389 (N_17389,N_17140,N_17061);
and U17390 (N_17390,N_17021,N_17172);
nor U17391 (N_17391,N_17133,N_17232);
or U17392 (N_17392,N_17052,N_17133);
nor U17393 (N_17393,N_17194,N_17188);
nand U17394 (N_17394,N_17153,N_17050);
nand U17395 (N_17395,N_17078,N_17191);
nand U17396 (N_17396,N_17041,N_17029);
and U17397 (N_17397,N_17010,N_17223);
and U17398 (N_17398,N_17036,N_17216);
nor U17399 (N_17399,N_17098,N_17160);
nand U17400 (N_17400,N_17070,N_17184);
or U17401 (N_17401,N_17037,N_17090);
and U17402 (N_17402,N_17142,N_17182);
nor U17403 (N_17403,N_17036,N_17094);
nand U17404 (N_17404,N_17234,N_17129);
and U17405 (N_17405,N_17013,N_17206);
xor U17406 (N_17406,N_17124,N_17193);
xor U17407 (N_17407,N_17008,N_17174);
or U17408 (N_17408,N_17164,N_17016);
nor U17409 (N_17409,N_17226,N_17048);
and U17410 (N_17410,N_17192,N_17179);
and U17411 (N_17411,N_17075,N_17047);
nor U17412 (N_17412,N_17034,N_17224);
xnor U17413 (N_17413,N_17142,N_17016);
nand U17414 (N_17414,N_17107,N_17168);
xor U17415 (N_17415,N_17163,N_17002);
or U17416 (N_17416,N_17114,N_17065);
xnor U17417 (N_17417,N_17171,N_17036);
or U17418 (N_17418,N_17244,N_17234);
nor U17419 (N_17419,N_17246,N_17051);
and U17420 (N_17420,N_17013,N_17181);
xor U17421 (N_17421,N_17219,N_17049);
and U17422 (N_17422,N_17113,N_17007);
xnor U17423 (N_17423,N_17222,N_17013);
or U17424 (N_17424,N_17166,N_17181);
nor U17425 (N_17425,N_17132,N_17174);
xor U17426 (N_17426,N_17079,N_17149);
nor U17427 (N_17427,N_17230,N_17097);
nand U17428 (N_17428,N_17197,N_17031);
nand U17429 (N_17429,N_17114,N_17244);
and U17430 (N_17430,N_17176,N_17118);
and U17431 (N_17431,N_17243,N_17109);
nor U17432 (N_17432,N_17138,N_17170);
nand U17433 (N_17433,N_17088,N_17193);
nand U17434 (N_17434,N_17019,N_17207);
or U17435 (N_17435,N_17171,N_17238);
xnor U17436 (N_17436,N_17039,N_17190);
nor U17437 (N_17437,N_17112,N_17080);
or U17438 (N_17438,N_17165,N_17060);
xnor U17439 (N_17439,N_17080,N_17233);
nor U17440 (N_17440,N_17145,N_17209);
or U17441 (N_17441,N_17213,N_17107);
nor U17442 (N_17442,N_17198,N_17022);
nand U17443 (N_17443,N_17002,N_17231);
nor U17444 (N_17444,N_17013,N_17131);
or U17445 (N_17445,N_17174,N_17138);
or U17446 (N_17446,N_17104,N_17083);
and U17447 (N_17447,N_17231,N_17135);
nor U17448 (N_17448,N_17194,N_17149);
or U17449 (N_17449,N_17079,N_17241);
nor U17450 (N_17450,N_17209,N_17184);
and U17451 (N_17451,N_17198,N_17214);
nor U17452 (N_17452,N_17051,N_17218);
nand U17453 (N_17453,N_17086,N_17087);
and U17454 (N_17454,N_17026,N_17130);
nand U17455 (N_17455,N_17188,N_17212);
or U17456 (N_17456,N_17113,N_17180);
nor U17457 (N_17457,N_17006,N_17245);
nand U17458 (N_17458,N_17120,N_17093);
nand U17459 (N_17459,N_17066,N_17159);
and U17460 (N_17460,N_17147,N_17022);
nor U17461 (N_17461,N_17065,N_17213);
and U17462 (N_17462,N_17052,N_17099);
nand U17463 (N_17463,N_17045,N_17007);
nor U17464 (N_17464,N_17030,N_17231);
or U17465 (N_17465,N_17067,N_17079);
xnor U17466 (N_17466,N_17231,N_17039);
nor U17467 (N_17467,N_17238,N_17138);
nor U17468 (N_17468,N_17154,N_17132);
or U17469 (N_17469,N_17035,N_17224);
and U17470 (N_17470,N_17143,N_17133);
and U17471 (N_17471,N_17056,N_17116);
nor U17472 (N_17472,N_17240,N_17060);
or U17473 (N_17473,N_17102,N_17232);
nand U17474 (N_17474,N_17115,N_17114);
nand U17475 (N_17475,N_17063,N_17161);
and U17476 (N_17476,N_17024,N_17076);
nand U17477 (N_17477,N_17144,N_17033);
or U17478 (N_17478,N_17138,N_17080);
xor U17479 (N_17479,N_17212,N_17178);
or U17480 (N_17480,N_17057,N_17246);
and U17481 (N_17481,N_17206,N_17149);
xnor U17482 (N_17482,N_17025,N_17018);
nand U17483 (N_17483,N_17246,N_17134);
and U17484 (N_17484,N_17024,N_17064);
or U17485 (N_17485,N_17153,N_17105);
or U17486 (N_17486,N_17167,N_17205);
or U17487 (N_17487,N_17044,N_17198);
or U17488 (N_17488,N_17098,N_17218);
or U17489 (N_17489,N_17047,N_17142);
nand U17490 (N_17490,N_17120,N_17060);
nor U17491 (N_17491,N_17050,N_17229);
and U17492 (N_17492,N_17034,N_17051);
nor U17493 (N_17493,N_17002,N_17126);
nand U17494 (N_17494,N_17223,N_17169);
or U17495 (N_17495,N_17204,N_17091);
or U17496 (N_17496,N_17237,N_17111);
and U17497 (N_17497,N_17069,N_17177);
or U17498 (N_17498,N_17057,N_17092);
xnor U17499 (N_17499,N_17029,N_17131);
nor U17500 (N_17500,N_17299,N_17348);
and U17501 (N_17501,N_17254,N_17333);
nand U17502 (N_17502,N_17335,N_17327);
nand U17503 (N_17503,N_17337,N_17362);
xnor U17504 (N_17504,N_17295,N_17436);
or U17505 (N_17505,N_17417,N_17435);
nand U17506 (N_17506,N_17264,N_17270);
and U17507 (N_17507,N_17431,N_17399);
xor U17508 (N_17508,N_17446,N_17411);
nand U17509 (N_17509,N_17463,N_17458);
nand U17510 (N_17510,N_17284,N_17483);
nor U17511 (N_17511,N_17386,N_17484);
nor U17512 (N_17512,N_17412,N_17360);
nor U17513 (N_17513,N_17317,N_17278);
xnor U17514 (N_17514,N_17404,N_17267);
or U17515 (N_17515,N_17387,N_17488);
nor U17516 (N_17516,N_17394,N_17340);
nand U17517 (N_17517,N_17376,N_17416);
or U17518 (N_17518,N_17457,N_17426);
nor U17519 (N_17519,N_17467,N_17425);
xor U17520 (N_17520,N_17379,N_17437);
nand U17521 (N_17521,N_17305,N_17345);
nor U17522 (N_17522,N_17468,N_17304);
or U17523 (N_17523,N_17498,N_17350);
nor U17524 (N_17524,N_17427,N_17357);
and U17525 (N_17525,N_17447,N_17341);
and U17526 (N_17526,N_17401,N_17328);
and U17527 (N_17527,N_17453,N_17429);
nor U17528 (N_17528,N_17253,N_17480);
nor U17529 (N_17529,N_17410,N_17441);
xnor U17530 (N_17530,N_17332,N_17450);
and U17531 (N_17531,N_17297,N_17359);
nand U17532 (N_17532,N_17396,N_17257);
nor U17533 (N_17533,N_17403,N_17300);
xnor U17534 (N_17534,N_17369,N_17384);
or U17535 (N_17535,N_17449,N_17489);
nor U17536 (N_17536,N_17288,N_17413);
and U17537 (N_17537,N_17378,N_17279);
and U17538 (N_17538,N_17409,N_17260);
nor U17539 (N_17539,N_17298,N_17481);
or U17540 (N_17540,N_17444,N_17255);
nor U17541 (N_17541,N_17302,N_17448);
nand U17542 (N_17542,N_17265,N_17497);
or U17543 (N_17543,N_17324,N_17277);
xor U17544 (N_17544,N_17296,N_17469);
and U17545 (N_17545,N_17308,N_17293);
or U17546 (N_17546,N_17287,N_17363);
and U17547 (N_17547,N_17455,N_17486);
and U17548 (N_17548,N_17310,N_17274);
and U17549 (N_17549,N_17276,N_17474);
xnor U17550 (N_17550,N_17268,N_17487);
xor U17551 (N_17551,N_17263,N_17492);
and U17552 (N_17552,N_17471,N_17459);
nor U17553 (N_17553,N_17347,N_17452);
xnor U17554 (N_17554,N_17424,N_17356);
xor U17555 (N_17555,N_17322,N_17490);
or U17556 (N_17556,N_17400,N_17285);
and U17557 (N_17557,N_17313,N_17323);
or U17558 (N_17558,N_17301,N_17389);
and U17559 (N_17559,N_17361,N_17418);
nor U17560 (N_17560,N_17314,N_17461);
nand U17561 (N_17561,N_17303,N_17368);
xor U17562 (N_17562,N_17491,N_17414);
nor U17563 (N_17563,N_17273,N_17405);
or U17564 (N_17564,N_17321,N_17259);
and U17565 (N_17565,N_17434,N_17421);
and U17566 (N_17566,N_17250,N_17432);
nand U17567 (N_17567,N_17419,N_17352);
or U17568 (N_17568,N_17364,N_17262);
nor U17569 (N_17569,N_17343,N_17466);
or U17570 (N_17570,N_17383,N_17460);
nor U17571 (N_17571,N_17261,N_17377);
or U17572 (N_17572,N_17355,N_17309);
nor U17573 (N_17573,N_17472,N_17294);
xor U17574 (N_17574,N_17477,N_17499);
nand U17575 (N_17575,N_17326,N_17318);
xor U17576 (N_17576,N_17439,N_17388);
nor U17577 (N_17577,N_17428,N_17430);
or U17578 (N_17578,N_17408,N_17464);
nor U17579 (N_17579,N_17272,N_17269);
or U17580 (N_17580,N_17251,N_17380);
nand U17581 (N_17581,N_17445,N_17456);
and U17582 (N_17582,N_17433,N_17398);
and U17583 (N_17583,N_17373,N_17256);
and U17584 (N_17584,N_17479,N_17342);
xor U17585 (N_17585,N_17306,N_17375);
nand U17586 (N_17586,N_17381,N_17358);
or U17587 (N_17587,N_17307,N_17454);
or U17588 (N_17588,N_17330,N_17353);
and U17589 (N_17589,N_17271,N_17370);
and U17590 (N_17590,N_17275,N_17266);
xor U17591 (N_17591,N_17280,N_17283);
nand U17592 (N_17592,N_17349,N_17494);
nor U17593 (N_17593,N_17382,N_17311);
nand U17594 (N_17594,N_17485,N_17312);
and U17595 (N_17595,N_17496,N_17366);
or U17596 (N_17596,N_17367,N_17319);
xnor U17597 (N_17597,N_17422,N_17393);
nor U17598 (N_17598,N_17397,N_17391);
and U17599 (N_17599,N_17291,N_17351);
nand U17600 (N_17600,N_17344,N_17407);
nand U17601 (N_17601,N_17372,N_17442);
nor U17602 (N_17602,N_17493,N_17371);
xor U17603 (N_17603,N_17315,N_17406);
xor U17604 (N_17604,N_17475,N_17420);
nand U17605 (N_17605,N_17392,N_17415);
nand U17606 (N_17606,N_17292,N_17316);
nand U17607 (N_17607,N_17465,N_17443);
or U17608 (N_17608,N_17289,N_17495);
or U17609 (N_17609,N_17462,N_17374);
and U17610 (N_17610,N_17252,N_17482);
nor U17611 (N_17611,N_17320,N_17258);
nand U17612 (N_17612,N_17385,N_17346);
or U17613 (N_17613,N_17290,N_17440);
xor U17614 (N_17614,N_17281,N_17423);
or U17615 (N_17615,N_17438,N_17470);
and U17616 (N_17616,N_17476,N_17329);
nor U17617 (N_17617,N_17334,N_17325);
or U17618 (N_17618,N_17336,N_17365);
nand U17619 (N_17619,N_17354,N_17478);
nand U17620 (N_17620,N_17331,N_17286);
nand U17621 (N_17621,N_17338,N_17451);
nor U17622 (N_17622,N_17339,N_17395);
xor U17623 (N_17623,N_17473,N_17402);
xnor U17624 (N_17624,N_17390,N_17282);
nand U17625 (N_17625,N_17457,N_17314);
and U17626 (N_17626,N_17491,N_17256);
nand U17627 (N_17627,N_17284,N_17383);
nand U17628 (N_17628,N_17298,N_17445);
and U17629 (N_17629,N_17449,N_17395);
and U17630 (N_17630,N_17341,N_17477);
and U17631 (N_17631,N_17490,N_17457);
or U17632 (N_17632,N_17414,N_17493);
xnor U17633 (N_17633,N_17443,N_17416);
nand U17634 (N_17634,N_17293,N_17300);
or U17635 (N_17635,N_17349,N_17398);
xor U17636 (N_17636,N_17294,N_17459);
and U17637 (N_17637,N_17334,N_17491);
xnor U17638 (N_17638,N_17439,N_17343);
nand U17639 (N_17639,N_17384,N_17312);
xor U17640 (N_17640,N_17489,N_17497);
xor U17641 (N_17641,N_17402,N_17454);
or U17642 (N_17642,N_17269,N_17399);
xor U17643 (N_17643,N_17303,N_17389);
xnor U17644 (N_17644,N_17455,N_17493);
or U17645 (N_17645,N_17335,N_17272);
or U17646 (N_17646,N_17386,N_17403);
or U17647 (N_17647,N_17466,N_17416);
nand U17648 (N_17648,N_17417,N_17428);
xor U17649 (N_17649,N_17492,N_17448);
nor U17650 (N_17650,N_17379,N_17363);
xnor U17651 (N_17651,N_17405,N_17449);
nor U17652 (N_17652,N_17297,N_17279);
nor U17653 (N_17653,N_17311,N_17265);
or U17654 (N_17654,N_17300,N_17398);
nor U17655 (N_17655,N_17332,N_17422);
and U17656 (N_17656,N_17406,N_17320);
or U17657 (N_17657,N_17382,N_17296);
and U17658 (N_17658,N_17434,N_17262);
and U17659 (N_17659,N_17325,N_17351);
xor U17660 (N_17660,N_17336,N_17482);
nand U17661 (N_17661,N_17265,N_17282);
or U17662 (N_17662,N_17320,N_17479);
xnor U17663 (N_17663,N_17470,N_17426);
nor U17664 (N_17664,N_17289,N_17283);
and U17665 (N_17665,N_17309,N_17364);
and U17666 (N_17666,N_17258,N_17382);
xor U17667 (N_17667,N_17367,N_17300);
or U17668 (N_17668,N_17410,N_17292);
nor U17669 (N_17669,N_17479,N_17275);
xnor U17670 (N_17670,N_17377,N_17251);
xor U17671 (N_17671,N_17356,N_17315);
or U17672 (N_17672,N_17499,N_17376);
nand U17673 (N_17673,N_17377,N_17420);
and U17674 (N_17674,N_17392,N_17290);
xor U17675 (N_17675,N_17259,N_17436);
and U17676 (N_17676,N_17336,N_17312);
and U17677 (N_17677,N_17259,N_17460);
nand U17678 (N_17678,N_17388,N_17456);
nor U17679 (N_17679,N_17420,N_17329);
and U17680 (N_17680,N_17476,N_17347);
nand U17681 (N_17681,N_17317,N_17267);
and U17682 (N_17682,N_17291,N_17492);
nand U17683 (N_17683,N_17370,N_17482);
nor U17684 (N_17684,N_17284,N_17387);
or U17685 (N_17685,N_17300,N_17256);
or U17686 (N_17686,N_17425,N_17420);
or U17687 (N_17687,N_17454,N_17361);
xnor U17688 (N_17688,N_17395,N_17260);
or U17689 (N_17689,N_17309,N_17261);
nor U17690 (N_17690,N_17312,N_17253);
or U17691 (N_17691,N_17266,N_17441);
or U17692 (N_17692,N_17486,N_17367);
nand U17693 (N_17693,N_17264,N_17258);
and U17694 (N_17694,N_17482,N_17325);
or U17695 (N_17695,N_17315,N_17275);
or U17696 (N_17696,N_17275,N_17324);
or U17697 (N_17697,N_17303,N_17484);
nand U17698 (N_17698,N_17434,N_17309);
nor U17699 (N_17699,N_17412,N_17490);
and U17700 (N_17700,N_17325,N_17275);
nand U17701 (N_17701,N_17324,N_17336);
and U17702 (N_17702,N_17381,N_17332);
nand U17703 (N_17703,N_17462,N_17412);
or U17704 (N_17704,N_17477,N_17439);
nor U17705 (N_17705,N_17292,N_17327);
nand U17706 (N_17706,N_17281,N_17311);
and U17707 (N_17707,N_17260,N_17258);
or U17708 (N_17708,N_17455,N_17412);
nor U17709 (N_17709,N_17416,N_17407);
nand U17710 (N_17710,N_17396,N_17416);
nor U17711 (N_17711,N_17401,N_17464);
nor U17712 (N_17712,N_17309,N_17483);
xnor U17713 (N_17713,N_17334,N_17370);
or U17714 (N_17714,N_17304,N_17496);
and U17715 (N_17715,N_17301,N_17418);
nand U17716 (N_17716,N_17393,N_17439);
nand U17717 (N_17717,N_17318,N_17417);
nand U17718 (N_17718,N_17459,N_17463);
or U17719 (N_17719,N_17360,N_17276);
or U17720 (N_17720,N_17341,N_17260);
xor U17721 (N_17721,N_17253,N_17448);
xor U17722 (N_17722,N_17401,N_17430);
and U17723 (N_17723,N_17375,N_17252);
or U17724 (N_17724,N_17339,N_17342);
xnor U17725 (N_17725,N_17387,N_17360);
or U17726 (N_17726,N_17447,N_17404);
or U17727 (N_17727,N_17455,N_17492);
nor U17728 (N_17728,N_17477,N_17433);
nand U17729 (N_17729,N_17422,N_17439);
and U17730 (N_17730,N_17287,N_17368);
or U17731 (N_17731,N_17310,N_17495);
nor U17732 (N_17732,N_17429,N_17282);
nor U17733 (N_17733,N_17328,N_17414);
and U17734 (N_17734,N_17256,N_17357);
and U17735 (N_17735,N_17460,N_17490);
or U17736 (N_17736,N_17474,N_17292);
or U17737 (N_17737,N_17421,N_17261);
or U17738 (N_17738,N_17402,N_17275);
and U17739 (N_17739,N_17393,N_17309);
and U17740 (N_17740,N_17410,N_17409);
or U17741 (N_17741,N_17352,N_17305);
or U17742 (N_17742,N_17366,N_17294);
xor U17743 (N_17743,N_17459,N_17485);
nand U17744 (N_17744,N_17440,N_17364);
nor U17745 (N_17745,N_17426,N_17482);
or U17746 (N_17746,N_17442,N_17417);
nor U17747 (N_17747,N_17274,N_17431);
nor U17748 (N_17748,N_17420,N_17261);
and U17749 (N_17749,N_17285,N_17261);
nor U17750 (N_17750,N_17561,N_17500);
and U17751 (N_17751,N_17726,N_17590);
nor U17752 (N_17752,N_17646,N_17715);
and U17753 (N_17753,N_17506,N_17734);
nor U17754 (N_17754,N_17632,N_17635);
nor U17755 (N_17755,N_17505,N_17507);
and U17756 (N_17756,N_17552,N_17584);
nand U17757 (N_17757,N_17524,N_17730);
xor U17758 (N_17758,N_17703,N_17652);
and U17759 (N_17759,N_17565,N_17607);
and U17760 (N_17760,N_17623,N_17711);
and U17761 (N_17761,N_17585,N_17609);
nor U17762 (N_17762,N_17658,N_17731);
and U17763 (N_17763,N_17605,N_17667);
and U17764 (N_17764,N_17621,N_17697);
or U17765 (N_17765,N_17574,N_17695);
nor U17766 (N_17766,N_17696,N_17688);
xor U17767 (N_17767,N_17745,N_17555);
or U17768 (N_17768,N_17698,N_17663);
xnor U17769 (N_17769,N_17662,N_17580);
nand U17770 (N_17770,N_17577,N_17626);
nand U17771 (N_17771,N_17625,N_17606);
xor U17772 (N_17772,N_17553,N_17729);
nand U17773 (N_17773,N_17710,N_17690);
nand U17774 (N_17774,N_17655,N_17593);
and U17775 (N_17775,N_17651,N_17549);
nor U17776 (N_17776,N_17747,N_17633);
or U17777 (N_17777,N_17707,N_17741);
and U17778 (N_17778,N_17589,N_17738);
xor U17779 (N_17779,N_17743,N_17749);
nand U17780 (N_17780,N_17597,N_17583);
or U17781 (N_17781,N_17504,N_17684);
nor U17782 (N_17782,N_17724,N_17706);
nand U17783 (N_17783,N_17642,N_17515);
or U17784 (N_17784,N_17599,N_17518);
and U17785 (N_17785,N_17675,N_17714);
nand U17786 (N_17786,N_17670,N_17512);
nor U17787 (N_17787,N_17579,N_17689);
xor U17788 (N_17788,N_17575,N_17554);
nor U17789 (N_17789,N_17532,N_17622);
nand U17790 (N_17790,N_17564,N_17535);
nor U17791 (N_17791,N_17647,N_17576);
nor U17792 (N_17792,N_17680,N_17668);
and U17793 (N_17793,N_17664,N_17719);
or U17794 (N_17794,N_17570,N_17666);
nor U17795 (N_17795,N_17727,N_17661);
xnor U17796 (N_17796,N_17627,N_17644);
and U17797 (N_17797,N_17608,N_17669);
or U17798 (N_17798,N_17694,N_17657);
and U17799 (N_17799,N_17619,N_17519);
nand U17800 (N_17800,N_17540,N_17679);
nor U17801 (N_17801,N_17620,N_17572);
xnor U17802 (N_17802,N_17536,N_17596);
nand U17803 (N_17803,N_17722,N_17602);
nor U17804 (N_17804,N_17582,N_17613);
and U17805 (N_17805,N_17617,N_17681);
nand U17806 (N_17806,N_17521,N_17693);
or U17807 (N_17807,N_17648,N_17742);
or U17808 (N_17808,N_17636,N_17514);
xor U17809 (N_17809,N_17713,N_17691);
nand U17810 (N_17810,N_17740,N_17685);
and U17811 (N_17811,N_17629,N_17721);
and U17812 (N_17812,N_17525,N_17520);
or U17813 (N_17813,N_17723,N_17601);
nor U17814 (N_17814,N_17557,N_17656);
xnor U17815 (N_17815,N_17587,N_17522);
or U17816 (N_17816,N_17598,N_17566);
or U17817 (N_17817,N_17737,N_17573);
and U17818 (N_17818,N_17538,N_17526);
xor U17819 (N_17819,N_17614,N_17702);
or U17820 (N_17820,N_17508,N_17611);
or U17821 (N_17821,N_17643,N_17531);
xnor U17822 (N_17822,N_17650,N_17682);
xor U17823 (N_17823,N_17541,N_17717);
xnor U17824 (N_17824,N_17733,N_17547);
nand U17825 (N_17825,N_17624,N_17728);
nor U17826 (N_17826,N_17513,N_17604);
and U17827 (N_17827,N_17529,N_17692);
nand U17828 (N_17828,N_17618,N_17704);
nor U17829 (N_17829,N_17708,N_17527);
xor U17830 (N_17830,N_17603,N_17739);
and U17831 (N_17831,N_17595,N_17503);
nand U17832 (N_17832,N_17533,N_17592);
xnor U17833 (N_17833,N_17659,N_17628);
nor U17834 (N_17834,N_17586,N_17581);
xnor U17835 (N_17835,N_17560,N_17530);
or U17836 (N_17836,N_17558,N_17687);
xor U17837 (N_17837,N_17534,N_17509);
xor U17838 (N_17838,N_17563,N_17545);
and U17839 (N_17839,N_17568,N_17649);
xor U17840 (N_17840,N_17701,N_17502);
nand U17841 (N_17841,N_17523,N_17612);
nand U17842 (N_17842,N_17716,N_17516);
and U17843 (N_17843,N_17700,N_17591);
and U17844 (N_17844,N_17528,N_17676);
nand U17845 (N_17845,N_17539,N_17748);
or U17846 (N_17846,N_17537,N_17654);
and U17847 (N_17847,N_17683,N_17674);
or U17848 (N_17848,N_17567,N_17544);
nor U17849 (N_17849,N_17594,N_17725);
or U17850 (N_17850,N_17665,N_17638);
nand U17851 (N_17851,N_17641,N_17640);
and U17852 (N_17852,N_17543,N_17610);
or U17853 (N_17853,N_17639,N_17578);
nor U17854 (N_17854,N_17660,N_17732);
nand U17855 (N_17855,N_17546,N_17615);
and U17856 (N_17856,N_17600,N_17616);
nor U17857 (N_17857,N_17637,N_17671);
nor U17858 (N_17858,N_17712,N_17709);
xor U17859 (N_17859,N_17634,N_17630);
nand U17860 (N_17860,N_17699,N_17735);
xnor U17861 (N_17861,N_17556,N_17736);
xor U17862 (N_17862,N_17645,N_17673);
nor U17863 (N_17863,N_17571,N_17510);
or U17864 (N_17864,N_17744,N_17588);
xor U17865 (N_17865,N_17501,N_17517);
and U17866 (N_17866,N_17677,N_17551);
xnor U17867 (N_17867,N_17720,N_17562);
and U17868 (N_17868,N_17631,N_17569);
or U17869 (N_17869,N_17653,N_17746);
and U17870 (N_17870,N_17686,N_17511);
nor U17871 (N_17871,N_17718,N_17542);
or U17872 (N_17872,N_17548,N_17705);
or U17873 (N_17873,N_17550,N_17672);
and U17874 (N_17874,N_17559,N_17678);
and U17875 (N_17875,N_17535,N_17628);
and U17876 (N_17876,N_17518,N_17701);
and U17877 (N_17877,N_17656,N_17716);
nor U17878 (N_17878,N_17745,N_17668);
and U17879 (N_17879,N_17611,N_17739);
and U17880 (N_17880,N_17743,N_17675);
nor U17881 (N_17881,N_17510,N_17645);
or U17882 (N_17882,N_17741,N_17650);
nand U17883 (N_17883,N_17740,N_17708);
nor U17884 (N_17884,N_17563,N_17502);
or U17885 (N_17885,N_17557,N_17595);
nor U17886 (N_17886,N_17615,N_17663);
nor U17887 (N_17887,N_17588,N_17638);
nor U17888 (N_17888,N_17644,N_17715);
and U17889 (N_17889,N_17660,N_17577);
nor U17890 (N_17890,N_17684,N_17742);
xnor U17891 (N_17891,N_17565,N_17725);
and U17892 (N_17892,N_17728,N_17654);
nor U17893 (N_17893,N_17518,N_17503);
nand U17894 (N_17894,N_17666,N_17658);
nor U17895 (N_17895,N_17720,N_17603);
nand U17896 (N_17896,N_17673,N_17518);
nand U17897 (N_17897,N_17572,N_17623);
or U17898 (N_17898,N_17607,N_17592);
nor U17899 (N_17899,N_17536,N_17666);
and U17900 (N_17900,N_17614,N_17744);
xor U17901 (N_17901,N_17604,N_17622);
nor U17902 (N_17902,N_17626,N_17507);
or U17903 (N_17903,N_17528,N_17719);
xor U17904 (N_17904,N_17574,N_17650);
or U17905 (N_17905,N_17568,N_17689);
and U17906 (N_17906,N_17557,N_17655);
or U17907 (N_17907,N_17621,N_17713);
nand U17908 (N_17908,N_17626,N_17529);
and U17909 (N_17909,N_17747,N_17713);
xnor U17910 (N_17910,N_17739,N_17561);
or U17911 (N_17911,N_17655,N_17734);
xnor U17912 (N_17912,N_17681,N_17587);
or U17913 (N_17913,N_17715,N_17642);
or U17914 (N_17914,N_17510,N_17597);
nor U17915 (N_17915,N_17736,N_17539);
and U17916 (N_17916,N_17511,N_17676);
or U17917 (N_17917,N_17749,N_17511);
nor U17918 (N_17918,N_17516,N_17719);
nor U17919 (N_17919,N_17614,N_17637);
or U17920 (N_17920,N_17747,N_17688);
and U17921 (N_17921,N_17709,N_17634);
nor U17922 (N_17922,N_17678,N_17680);
nor U17923 (N_17923,N_17717,N_17609);
or U17924 (N_17924,N_17630,N_17670);
xnor U17925 (N_17925,N_17662,N_17550);
and U17926 (N_17926,N_17678,N_17642);
nor U17927 (N_17927,N_17549,N_17707);
xor U17928 (N_17928,N_17607,N_17729);
xor U17929 (N_17929,N_17631,N_17545);
nand U17930 (N_17930,N_17728,N_17549);
and U17931 (N_17931,N_17544,N_17619);
and U17932 (N_17932,N_17585,N_17680);
and U17933 (N_17933,N_17530,N_17709);
nor U17934 (N_17934,N_17579,N_17635);
and U17935 (N_17935,N_17714,N_17676);
and U17936 (N_17936,N_17537,N_17738);
and U17937 (N_17937,N_17520,N_17725);
nand U17938 (N_17938,N_17714,N_17589);
and U17939 (N_17939,N_17691,N_17704);
nand U17940 (N_17940,N_17574,N_17599);
xnor U17941 (N_17941,N_17718,N_17677);
nand U17942 (N_17942,N_17736,N_17504);
and U17943 (N_17943,N_17668,N_17707);
nor U17944 (N_17944,N_17643,N_17674);
or U17945 (N_17945,N_17591,N_17586);
and U17946 (N_17946,N_17669,N_17524);
nor U17947 (N_17947,N_17648,N_17618);
or U17948 (N_17948,N_17674,N_17679);
nand U17949 (N_17949,N_17560,N_17599);
and U17950 (N_17950,N_17633,N_17552);
nor U17951 (N_17951,N_17619,N_17621);
nor U17952 (N_17952,N_17741,N_17744);
xor U17953 (N_17953,N_17734,N_17677);
and U17954 (N_17954,N_17526,N_17531);
and U17955 (N_17955,N_17621,N_17723);
or U17956 (N_17956,N_17523,N_17660);
and U17957 (N_17957,N_17662,N_17581);
nor U17958 (N_17958,N_17696,N_17563);
and U17959 (N_17959,N_17692,N_17596);
or U17960 (N_17960,N_17557,N_17521);
xnor U17961 (N_17961,N_17657,N_17594);
and U17962 (N_17962,N_17539,N_17749);
nor U17963 (N_17963,N_17713,N_17563);
or U17964 (N_17964,N_17594,N_17636);
and U17965 (N_17965,N_17669,N_17654);
or U17966 (N_17966,N_17531,N_17713);
or U17967 (N_17967,N_17523,N_17639);
and U17968 (N_17968,N_17503,N_17691);
or U17969 (N_17969,N_17584,N_17583);
xor U17970 (N_17970,N_17554,N_17735);
xor U17971 (N_17971,N_17641,N_17732);
or U17972 (N_17972,N_17595,N_17609);
nand U17973 (N_17973,N_17564,N_17650);
nor U17974 (N_17974,N_17649,N_17655);
nand U17975 (N_17975,N_17597,N_17587);
nor U17976 (N_17976,N_17570,N_17605);
and U17977 (N_17977,N_17625,N_17619);
nor U17978 (N_17978,N_17523,N_17688);
nor U17979 (N_17979,N_17644,N_17580);
and U17980 (N_17980,N_17633,N_17640);
nor U17981 (N_17981,N_17603,N_17656);
nand U17982 (N_17982,N_17741,N_17708);
nand U17983 (N_17983,N_17580,N_17747);
or U17984 (N_17984,N_17614,N_17733);
nor U17985 (N_17985,N_17673,N_17628);
xnor U17986 (N_17986,N_17731,N_17596);
nand U17987 (N_17987,N_17685,N_17610);
nand U17988 (N_17988,N_17611,N_17678);
and U17989 (N_17989,N_17668,N_17729);
and U17990 (N_17990,N_17734,N_17612);
nor U17991 (N_17991,N_17706,N_17610);
xor U17992 (N_17992,N_17674,N_17566);
nor U17993 (N_17993,N_17712,N_17675);
or U17994 (N_17994,N_17742,N_17645);
xnor U17995 (N_17995,N_17677,N_17524);
or U17996 (N_17996,N_17658,N_17594);
and U17997 (N_17997,N_17632,N_17651);
xnor U17998 (N_17998,N_17544,N_17680);
nor U17999 (N_17999,N_17548,N_17646);
and U18000 (N_18000,N_17908,N_17934);
nand U18001 (N_18001,N_17875,N_17805);
xor U18002 (N_18002,N_17791,N_17995);
xor U18003 (N_18003,N_17971,N_17784);
nand U18004 (N_18004,N_17782,N_17996);
nor U18005 (N_18005,N_17994,N_17983);
xnor U18006 (N_18006,N_17786,N_17915);
xnor U18007 (N_18007,N_17894,N_17970);
xor U18008 (N_18008,N_17937,N_17959);
xnor U18009 (N_18009,N_17867,N_17756);
nor U18010 (N_18010,N_17837,N_17865);
nand U18011 (N_18011,N_17785,N_17905);
and U18012 (N_18012,N_17774,N_17869);
xnor U18013 (N_18013,N_17797,N_17892);
nand U18014 (N_18014,N_17977,N_17826);
and U18015 (N_18015,N_17918,N_17808);
xor U18016 (N_18016,N_17888,N_17821);
nor U18017 (N_18017,N_17763,N_17890);
xor U18018 (N_18018,N_17861,N_17945);
or U18019 (N_18019,N_17991,N_17832);
and U18020 (N_18020,N_17943,N_17876);
xor U18021 (N_18021,N_17897,N_17795);
nor U18022 (N_18022,N_17925,N_17758);
nand U18023 (N_18023,N_17884,N_17771);
nand U18024 (N_18024,N_17950,N_17985);
and U18025 (N_18025,N_17778,N_17789);
or U18026 (N_18026,N_17843,N_17962);
nor U18027 (N_18027,N_17834,N_17998);
nor U18028 (N_18028,N_17916,N_17831);
or U18029 (N_18029,N_17801,N_17761);
or U18030 (N_18030,N_17858,N_17928);
xnor U18031 (N_18031,N_17799,N_17811);
nor U18032 (N_18032,N_17856,N_17804);
or U18033 (N_18033,N_17929,N_17933);
xor U18034 (N_18034,N_17987,N_17988);
nor U18035 (N_18035,N_17790,N_17978);
xor U18036 (N_18036,N_17770,N_17841);
nor U18037 (N_18037,N_17823,N_17932);
nor U18038 (N_18038,N_17752,N_17939);
xnor U18039 (N_18039,N_17825,N_17850);
xor U18040 (N_18040,N_17907,N_17765);
nand U18041 (N_18041,N_17922,N_17931);
and U18042 (N_18042,N_17842,N_17768);
xor U18043 (N_18043,N_17776,N_17762);
xor U18044 (N_18044,N_17901,N_17935);
xor U18045 (N_18045,N_17948,N_17775);
nand U18046 (N_18046,N_17859,N_17904);
nor U18047 (N_18047,N_17838,N_17800);
or U18048 (N_18048,N_17819,N_17817);
or U18049 (N_18049,N_17913,N_17899);
and U18050 (N_18050,N_17847,N_17878);
nor U18051 (N_18051,N_17802,N_17990);
nand U18052 (N_18052,N_17952,N_17967);
and U18053 (N_18053,N_17984,N_17751);
xor U18054 (N_18054,N_17941,N_17912);
and U18055 (N_18055,N_17940,N_17997);
nand U18056 (N_18056,N_17871,N_17764);
xor U18057 (N_18057,N_17853,N_17862);
nand U18058 (N_18058,N_17860,N_17844);
xnor U18059 (N_18059,N_17927,N_17914);
or U18060 (N_18060,N_17975,N_17972);
nor U18061 (N_18061,N_17852,N_17814);
or U18062 (N_18062,N_17957,N_17783);
or U18063 (N_18063,N_17921,N_17911);
nor U18064 (N_18064,N_17849,N_17777);
or U18065 (N_18065,N_17796,N_17886);
nand U18066 (N_18066,N_17779,N_17963);
nor U18067 (N_18067,N_17855,N_17794);
nand U18068 (N_18068,N_17999,N_17836);
nor U18069 (N_18069,N_17760,N_17816);
nand U18070 (N_18070,N_17924,N_17829);
nor U18071 (N_18071,N_17767,N_17750);
and U18072 (N_18072,N_17891,N_17974);
xor U18073 (N_18073,N_17902,N_17961);
xor U18074 (N_18074,N_17828,N_17906);
xnor U18075 (N_18075,N_17936,N_17887);
xor U18076 (N_18076,N_17981,N_17840);
or U18077 (N_18077,N_17960,N_17864);
nand U18078 (N_18078,N_17900,N_17813);
xor U18079 (N_18079,N_17755,N_17986);
or U18080 (N_18080,N_17873,N_17772);
nor U18081 (N_18081,N_17893,N_17976);
nand U18082 (N_18082,N_17980,N_17926);
nand U18083 (N_18083,N_17930,N_17910);
nor U18084 (N_18084,N_17954,N_17880);
nand U18085 (N_18085,N_17958,N_17964);
nor U18086 (N_18086,N_17883,N_17848);
and U18087 (N_18087,N_17879,N_17803);
or U18088 (N_18088,N_17857,N_17810);
and U18089 (N_18089,N_17917,N_17798);
and U18090 (N_18090,N_17973,N_17992);
nand U18091 (N_18091,N_17872,N_17788);
and U18092 (N_18092,N_17903,N_17868);
xnor U18093 (N_18093,N_17773,N_17898);
and U18094 (N_18094,N_17835,N_17827);
nor U18095 (N_18095,N_17949,N_17877);
and U18096 (N_18096,N_17965,N_17909);
nand U18097 (N_18097,N_17809,N_17919);
and U18098 (N_18098,N_17846,N_17989);
nor U18099 (N_18099,N_17870,N_17956);
nand U18100 (N_18100,N_17874,N_17969);
nor U18101 (N_18101,N_17993,N_17889);
nor U18102 (N_18102,N_17830,N_17955);
nor U18103 (N_18103,N_17979,N_17754);
and U18104 (N_18104,N_17966,N_17938);
and U18105 (N_18105,N_17982,N_17851);
or U18106 (N_18106,N_17895,N_17845);
and U18107 (N_18107,N_17753,N_17863);
and U18108 (N_18108,N_17812,N_17953);
and U18109 (N_18109,N_17781,N_17818);
or U18110 (N_18110,N_17944,N_17806);
xor U18111 (N_18111,N_17759,N_17793);
nor U18112 (N_18112,N_17780,N_17881);
or U18113 (N_18113,N_17920,N_17882);
nor U18114 (N_18114,N_17820,N_17947);
xnor U18115 (N_18115,N_17757,N_17792);
or U18116 (N_18116,N_17942,N_17968);
and U18117 (N_18117,N_17766,N_17896);
nor U18118 (N_18118,N_17833,N_17854);
or U18119 (N_18119,N_17951,N_17807);
and U18120 (N_18120,N_17787,N_17839);
nor U18121 (N_18121,N_17824,N_17769);
xnor U18122 (N_18122,N_17923,N_17885);
xor U18123 (N_18123,N_17815,N_17822);
nor U18124 (N_18124,N_17866,N_17946);
nor U18125 (N_18125,N_17757,N_17974);
or U18126 (N_18126,N_17804,N_17830);
nor U18127 (N_18127,N_17909,N_17913);
nor U18128 (N_18128,N_17925,N_17914);
nor U18129 (N_18129,N_17995,N_17830);
nand U18130 (N_18130,N_17751,N_17790);
or U18131 (N_18131,N_17919,N_17843);
nor U18132 (N_18132,N_17851,N_17805);
nor U18133 (N_18133,N_17904,N_17908);
or U18134 (N_18134,N_17884,N_17760);
and U18135 (N_18135,N_17902,N_17891);
xnor U18136 (N_18136,N_17751,N_17889);
or U18137 (N_18137,N_17783,N_17997);
nand U18138 (N_18138,N_17840,N_17973);
xnor U18139 (N_18139,N_17877,N_17878);
and U18140 (N_18140,N_17845,N_17835);
nor U18141 (N_18141,N_17995,N_17901);
nor U18142 (N_18142,N_17865,N_17969);
or U18143 (N_18143,N_17848,N_17806);
and U18144 (N_18144,N_17882,N_17886);
nand U18145 (N_18145,N_17869,N_17879);
xnor U18146 (N_18146,N_17905,N_17936);
xor U18147 (N_18147,N_17876,N_17794);
xnor U18148 (N_18148,N_17780,N_17800);
nor U18149 (N_18149,N_17999,N_17801);
nand U18150 (N_18150,N_17752,N_17859);
nor U18151 (N_18151,N_17882,N_17774);
and U18152 (N_18152,N_17818,N_17907);
xnor U18153 (N_18153,N_17927,N_17917);
or U18154 (N_18154,N_17926,N_17814);
and U18155 (N_18155,N_17994,N_17926);
nand U18156 (N_18156,N_17790,N_17997);
nor U18157 (N_18157,N_17760,N_17951);
nor U18158 (N_18158,N_17910,N_17788);
and U18159 (N_18159,N_17972,N_17814);
and U18160 (N_18160,N_17871,N_17870);
or U18161 (N_18161,N_17927,N_17961);
xnor U18162 (N_18162,N_17828,N_17787);
nor U18163 (N_18163,N_17991,N_17888);
and U18164 (N_18164,N_17825,N_17903);
or U18165 (N_18165,N_17755,N_17781);
nand U18166 (N_18166,N_17758,N_17949);
xor U18167 (N_18167,N_17805,N_17970);
and U18168 (N_18168,N_17881,N_17787);
or U18169 (N_18169,N_17795,N_17972);
or U18170 (N_18170,N_17800,N_17896);
xor U18171 (N_18171,N_17901,N_17907);
nand U18172 (N_18172,N_17911,N_17889);
nor U18173 (N_18173,N_17903,N_17824);
or U18174 (N_18174,N_17940,N_17865);
or U18175 (N_18175,N_17839,N_17871);
xnor U18176 (N_18176,N_17883,N_17826);
nand U18177 (N_18177,N_17907,N_17882);
and U18178 (N_18178,N_17882,N_17859);
or U18179 (N_18179,N_17887,N_17995);
or U18180 (N_18180,N_17961,N_17781);
nand U18181 (N_18181,N_17751,N_17993);
nor U18182 (N_18182,N_17854,N_17978);
xor U18183 (N_18183,N_17807,N_17832);
or U18184 (N_18184,N_17785,N_17884);
nand U18185 (N_18185,N_17925,N_17814);
xnor U18186 (N_18186,N_17903,N_17861);
nand U18187 (N_18187,N_17853,N_17926);
and U18188 (N_18188,N_17793,N_17830);
xor U18189 (N_18189,N_17886,N_17767);
and U18190 (N_18190,N_17972,N_17802);
nand U18191 (N_18191,N_17934,N_17997);
nand U18192 (N_18192,N_17779,N_17872);
or U18193 (N_18193,N_17956,N_17919);
and U18194 (N_18194,N_17806,N_17879);
or U18195 (N_18195,N_17802,N_17945);
nand U18196 (N_18196,N_17853,N_17944);
and U18197 (N_18197,N_17870,N_17820);
nand U18198 (N_18198,N_17875,N_17892);
and U18199 (N_18199,N_17757,N_17964);
xor U18200 (N_18200,N_17828,N_17997);
and U18201 (N_18201,N_17779,N_17819);
nor U18202 (N_18202,N_17793,N_17912);
or U18203 (N_18203,N_17999,N_17998);
xnor U18204 (N_18204,N_17832,N_17896);
and U18205 (N_18205,N_17914,N_17845);
xnor U18206 (N_18206,N_17992,N_17835);
and U18207 (N_18207,N_17905,N_17832);
nand U18208 (N_18208,N_17863,N_17947);
xor U18209 (N_18209,N_17883,N_17812);
or U18210 (N_18210,N_17908,N_17811);
and U18211 (N_18211,N_17911,N_17862);
nand U18212 (N_18212,N_17928,N_17974);
and U18213 (N_18213,N_17908,N_17845);
nor U18214 (N_18214,N_17928,N_17822);
xor U18215 (N_18215,N_17863,N_17956);
xnor U18216 (N_18216,N_17818,N_17939);
xor U18217 (N_18217,N_17898,N_17839);
or U18218 (N_18218,N_17902,N_17753);
nand U18219 (N_18219,N_17941,N_17852);
nor U18220 (N_18220,N_17832,N_17958);
or U18221 (N_18221,N_17837,N_17845);
nor U18222 (N_18222,N_17766,N_17857);
nand U18223 (N_18223,N_17934,N_17995);
xnor U18224 (N_18224,N_17839,N_17825);
nand U18225 (N_18225,N_17904,N_17911);
nand U18226 (N_18226,N_17759,N_17782);
xor U18227 (N_18227,N_17904,N_17990);
and U18228 (N_18228,N_17765,N_17924);
xnor U18229 (N_18229,N_17796,N_17840);
nor U18230 (N_18230,N_17906,N_17972);
xor U18231 (N_18231,N_17892,N_17959);
nand U18232 (N_18232,N_17979,N_17936);
or U18233 (N_18233,N_17790,N_17758);
and U18234 (N_18234,N_17792,N_17797);
or U18235 (N_18235,N_17959,N_17863);
or U18236 (N_18236,N_17776,N_17949);
or U18237 (N_18237,N_17959,N_17971);
and U18238 (N_18238,N_17878,N_17873);
xor U18239 (N_18239,N_17807,N_17928);
or U18240 (N_18240,N_17854,N_17989);
or U18241 (N_18241,N_17934,N_17914);
nor U18242 (N_18242,N_17829,N_17950);
nor U18243 (N_18243,N_17934,N_17816);
or U18244 (N_18244,N_17991,N_17850);
nand U18245 (N_18245,N_17922,N_17841);
nor U18246 (N_18246,N_17988,N_17790);
or U18247 (N_18247,N_17990,N_17954);
nand U18248 (N_18248,N_17818,N_17956);
and U18249 (N_18249,N_17846,N_17789);
or U18250 (N_18250,N_18230,N_18194);
nand U18251 (N_18251,N_18066,N_18239);
xnor U18252 (N_18252,N_18127,N_18229);
and U18253 (N_18253,N_18045,N_18064);
and U18254 (N_18254,N_18035,N_18008);
nor U18255 (N_18255,N_18163,N_18214);
or U18256 (N_18256,N_18181,N_18168);
and U18257 (N_18257,N_18177,N_18201);
and U18258 (N_18258,N_18139,N_18134);
and U18259 (N_18259,N_18243,N_18028);
nor U18260 (N_18260,N_18207,N_18026);
or U18261 (N_18261,N_18149,N_18096);
xor U18262 (N_18262,N_18224,N_18056);
nor U18263 (N_18263,N_18082,N_18037);
nor U18264 (N_18264,N_18129,N_18154);
and U18265 (N_18265,N_18241,N_18137);
nand U18266 (N_18266,N_18180,N_18121);
nor U18267 (N_18267,N_18038,N_18093);
nor U18268 (N_18268,N_18101,N_18222);
nand U18269 (N_18269,N_18019,N_18090);
or U18270 (N_18270,N_18059,N_18080);
xnor U18271 (N_18271,N_18218,N_18020);
nand U18272 (N_18272,N_18015,N_18021);
and U18273 (N_18273,N_18004,N_18244);
nor U18274 (N_18274,N_18073,N_18076);
nor U18275 (N_18275,N_18012,N_18133);
or U18276 (N_18276,N_18072,N_18063);
xor U18277 (N_18277,N_18226,N_18125);
nand U18278 (N_18278,N_18046,N_18071);
nor U18279 (N_18279,N_18116,N_18246);
nand U18280 (N_18280,N_18210,N_18171);
xor U18281 (N_18281,N_18086,N_18043);
xnor U18282 (N_18282,N_18123,N_18013);
and U18283 (N_18283,N_18184,N_18196);
nand U18284 (N_18284,N_18113,N_18213);
and U18285 (N_18285,N_18176,N_18029);
and U18286 (N_18286,N_18088,N_18234);
xor U18287 (N_18287,N_18248,N_18105);
xnor U18288 (N_18288,N_18006,N_18153);
nand U18289 (N_18289,N_18040,N_18077);
or U18290 (N_18290,N_18068,N_18204);
and U18291 (N_18291,N_18011,N_18039);
or U18292 (N_18292,N_18122,N_18051);
xor U18293 (N_18293,N_18156,N_18164);
nor U18294 (N_18294,N_18014,N_18136);
or U18295 (N_18295,N_18069,N_18190);
xor U18296 (N_18296,N_18148,N_18049);
nand U18297 (N_18297,N_18114,N_18245);
nand U18298 (N_18298,N_18099,N_18107);
and U18299 (N_18299,N_18198,N_18216);
nor U18300 (N_18300,N_18085,N_18124);
and U18301 (N_18301,N_18159,N_18078);
nand U18302 (N_18302,N_18007,N_18233);
xnor U18303 (N_18303,N_18146,N_18165);
and U18304 (N_18304,N_18131,N_18092);
nor U18305 (N_18305,N_18065,N_18200);
xnor U18306 (N_18306,N_18000,N_18211);
xor U18307 (N_18307,N_18160,N_18016);
nor U18308 (N_18308,N_18178,N_18001);
nor U18309 (N_18309,N_18120,N_18174);
xnor U18310 (N_18310,N_18054,N_18023);
or U18311 (N_18311,N_18158,N_18030);
nor U18312 (N_18312,N_18034,N_18217);
xor U18313 (N_18313,N_18130,N_18002);
nand U18314 (N_18314,N_18195,N_18132);
xor U18315 (N_18315,N_18236,N_18084);
nor U18316 (N_18316,N_18151,N_18227);
and U18317 (N_18317,N_18033,N_18141);
xor U18318 (N_18318,N_18138,N_18018);
or U18319 (N_18319,N_18097,N_18193);
and U18320 (N_18320,N_18017,N_18205);
nand U18321 (N_18321,N_18240,N_18183);
nor U18322 (N_18322,N_18118,N_18050);
xor U18323 (N_18323,N_18208,N_18155);
nor U18324 (N_18324,N_18188,N_18094);
nand U18325 (N_18325,N_18247,N_18157);
nor U18326 (N_18326,N_18061,N_18238);
nand U18327 (N_18327,N_18025,N_18206);
xnor U18328 (N_18328,N_18009,N_18228);
or U18329 (N_18329,N_18182,N_18098);
or U18330 (N_18330,N_18242,N_18058);
nor U18331 (N_18331,N_18167,N_18110);
or U18332 (N_18332,N_18108,N_18215);
or U18333 (N_18333,N_18111,N_18103);
nor U18334 (N_18334,N_18219,N_18135);
xor U18335 (N_18335,N_18191,N_18152);
and U18336 (N_18336,N_18022,N_18143);
and U18337 (N_18337,N_18209,N_18170);
or U18338 (N_18338,N_18232,N_18150);
nor U18339 (N_18339,N_18032,N_18142);
nand U18340 (N_18340,N_18199,N_18117);
or U18341 (N_18341,N_18042,N_18081);
nor U18342 (N_18342,N_18075,N_18145);
and U18343 (N_18343,N_18024,N_18074);
xor U18344 (N_18344,N_18048,N_18052);
and U18345 (N_18345,N_18189,N_18237);
or U18346 (N_18346,N_18166,N_18100);
nor U18347 (N_18347,N_18060,N_18161);
and U18348 (N_18348,N_18053,N_18144);
nand U18349 (N_18349,N_18179,N_18087);
and U18350 (N_18350,N_18126,N_18115);
xor U18351 (N_18351,N_18031,N_18102);
nand U18352 (N_18352,N_18225,N_18041);
nand U18353 (N_18353,N_18221,N_18055);
or U18354 (N_18354,N_18010,N_18112);
nand U18355 (N_18355,N_18220,N_18047);
nor U18356 (N_18356,N_18091,N_18119);
xor U18357 (N_18357,N_18162,N_18128);
nor U18358 (N_18358,N_18186,N_18223);
or U18359 (N_18359,N_18083,N_18003);
nor U18360 (N_18360,N_18089,N_18140);
and U18361 (N_18361,N_18036,N_18104);
xor U18362 (N_18362,N_18109,N_18027);
or U18363 (N_18363,N_18095,N_18067);
nand U18364 (N_18364,N_18044,N_18235);
and U18365 (N_18365,N_18005,N_18172);
nor U18366 (N_18366,N_18212,N_18249);
xnor U18367 (N_18367,N_18192,N_18147);
and U18368 (N_18368,N_18197,N_18175);
xnor U18369 (N_18369,N_18203,N_18106);
xnor U18370 (N_18370,N_18202,N_18173);
nor U18371 (N_18371,N_18169,N_18187);
nor U18372 (N_18372,N_18231,N_18062);
and U18373 (N_18373,N_18079,N_18057);
nand U18374 (N_18374,N_18185,N_18070);
nor U18375 (N_18375,N_18218,N_18181);
nor U18376 (N_18376,N_18124,N_18045);
xor U18377 (N_18377,N_18225,N_18204);
and U18378 (N_18378,N_18138,N_18175);
nand U18379 (N_18379,N_18176,N_18213);
xor U18380 (N_18380,N_18184,N_18012);
xnor U18381 (N_18381,N_18010,N_18193);
and U18382 (N_18382,N_18235,N_18007);
xnor U18383 (N_18383,N_18167,N_18080);
nor U18384 (N_18384,N_18020,N_18004);
nand U18385 (N_18385,N_18206,N_18208);
nand U18386 (N_18386,N_18145,N_18142);
nand U18387 (N_18387,N_18059,N_18062);
nor U18388 (N_18388,N_18137,N_18232);
nor U18389 (N_18389,N_18067,N_18021);
xor U18390 (N_18390,N_18207,N_18171);
nor U18391 (N_18391,N_18115,N_18162);
xor U18392 (N_18392,N_18200,N_18171);
and U18393 (N_18393,N_18173,N_18214);
xor U18394 (N_18394,N_18027,N_18091);
nor U18395 (N_18395,N_18039,N_18171);
or U18396 (N_18396,N_18246,N_18063);
xnor U18397 (N_18397,N_18084,N_18143);
nand U18398 (N_18398,N_18021,N_18181);
and U18399 (N_18399,N_18244,N_18146);
nor U18400 (N_18400,N_18128,N_18117);
xor U18401 (N_18401,N_18105,N_18141);
nor U18402 (N_18402,N_18118,N_18110);
or U18403 (N_18403,N_18184,N_18078);
and U18404 (N_18404,N_18040,N_18246);
nor U18405 (N_18405,N_18235,N_18202);
or U18406 (N_18406,N_18093,N_18166);
and U18407 (N_18407,N_18077,N_18186);
nand U18408 (N_18408,N_18180,N_18077);
xor U18409 (N_18409,N_18119,N_18209);
xor U18410 (N_18410,N_18247,N_18046);
and U18411 (N_18411,N_18003,N_18089);
and U18412 (N_18412,N_18167,N_18213);
or U18413 (N_18413,N_18241,N_18052);
nand U18414 (N_18414,N_18037,N_18239);
and U18415 (N_18415,N_18227,N_18184);
and U18416 (N_18416,N_18178,N_18156);
or U18417 (N_18417,N_18191,N_18049);
nor U18418 (N_18418,N_18229,N_18177);
nor U18419 (N_18419,N_18126,N_18001);
nand U18420 (N_18420,N_18060,N_18072);
and U18421 (N_18421,N_18198,N_18079);
xor U18422 (N_18422,N_18161,N_18211);
xor U18423 (N_18423,N_18102,N_18234);
and U18424 (N_18424,N_18149,N_18204);
and U18425 (N_18425,N_18066,N_18181);
nand U18426 (N_18426,N_18011,N_18181);
xnor U18427 (N_18427,N_18091,N_18097);
nand U18428 (N_18428,N_18035,N_18243);
and U18429 (N_18429,N_18248,N_18097);
and U18430 (N_18430,N_18232,N_18069);
xnor U18431 (N_18431,N_18060,N_18141);
xnor U18432 (N_18432,N_18070,N_18229);
or U18433 (N_18433,N_18018,N_18184);
nor U18434 (N_18434,N_18240,N_18031);
or U18435 (N_18435,N_18128,N_18100);
or U18436 (N_18436,N_18071,N_18242);
and U18437 (N_18437,N_18005,N_18215);
nor U18438 (N_18438,N_18146,N_18045);
and U18439 (N_18439,N_18111,N_18135);
nand U18440 (N_18440,N_18047,N_18028);
nor U18441 (N_18441,N_18129,N_18082);
and U18442 (N_18442,N_18006,N_18032);
nand U18443 (N_18443,N_18090,N_18147);
nand U18444 (N_18444,N_18132,N_18071);
nand U18445 (N_18445,N_18106,N_18080);
nor U18446 (N_18446,N_18195,N_18178);
or U18447 (N_18447,N_18244,N_18166);
nand U18448 (N_18448,N_18240,N_18214);
nand U18449 (N_18449,N_18221,N_18009);
and U18450 (N_18450,N_18094,N_18200);
and U18451 (N_18451,N_18180,N_18022);
and U18452 (N_18452,N_18176,N_18055);
nand U18453 (N_18453,N_18152,N_18026);
nor U18454 (N_18454,N_18094,N_18129);
and U18455 (N_18455,N_18105,N_18210);
xor U18456 (N_18456,N_18181,N_18222);
nor U18457 (N_18457,N_18163,N_18096);
xnor U18458 (N_18458,N_18216,N_18233);
and U18459 (N_18459,N_18041,N_18080);
nor U18460 (N_18460,N_18157,N_18095);
or U18461 (N_18461,N_18126,N_18168);
or U18462 (N_18462,N_18207,N_18035);
nand U18463 (N_18463,N_18233,N_18184);
nor U18464 (N_18464,N_18178,N_18021);
nand U18465 (N_18465,N_18006,N_18089);
nor U18466 (N_18466,N_18176,N_18024);
and U18467 (N_18467,N_18026,N_18008);
xnor U18468 (N_18468,N_18223,N_18099);
nand U18469 (N_18469,N_18085,N_18076);
nor U18470 (N_18470,N_18180,N_18108);
nand U18471 (N_18471,N_18052,N_18029);
or U18472 (N_18472,N_18078,N_18026);
nand U18473 (N_18473,N_18075,N_18219);
nor U18474 (N_18474,N_18007,N_18037);
and U18475 (N_18475,N_18161,N_18080);
nor U18476 (N_18476,N_18209,N_18151);
xnor U18477 (N_18477,N_18011,N_18050);
and U18478 (N_18478,N_18123,N_18107);
or U18479 (N_18479,N_18213,N_18029);
nor U18480 (N_18480,N_18185,N_18157);
nor U18481 (N_18481,N_18081,N_18207);
xnor U18482 (N_18482,N_18029,N_18196);
and U18483 (N_18483,N_18219,N_18023);
nor U18484 (N_18484,N_18143,N_18133);
xor U18485 (N_18485,N_18104,N_18093);
nand U18486 (N_18486,N_18005,N_18109);
and U18487 (N_18487,N_18031,N_18215);
or U18488 (N_18488,N_18132,N_18140);
nand U18489 (N_18489,N_18090,N_18186);
nor U18490 (N_18490,N_18162,N_18062);
and U18491 (N_18491,N_18088,N_18029);
xor U18492 (N_18492,N_18118,N_18160);
and U18493 (N_18493,N_18231,N_18242);
or U18494 (N_18494,N_18157,N_18173);
nor U18495 (N_18495,N_18040,N_18117);
or U18496 (N_18496,N_18195,N_18139);
xnor U18497 (N_18497,N_18124,N_18216);
nor U18498 (N_18498,N_18073,N_18025);
xor U18499 (N_18499,N_18062,N_18125);
nor U18500 (N_18500,N_18402,N_18338);
or U18501 (N_18501,N_18364,N_18434);
xnor U18502 (N_18502,N_18444,N_18340);
xor U18503 (N_18503,N_18292,N_18428);
or U18504 (N_18504,N_18264,N_18381);
or U18505 (N_18505,N_18328,N_18351);
xnor U18506 (N_18506,N_18360,N_18394);
nor U18507 (N_18507,N_18337,N_18412);
nor U18508 (N_18508,N_18332,N_18398);
nor U18509 (N_18509,N_18466,N_18485);
and U18510 (N_18510,N_18469,N_18354);
nor U18511 (N_18511,N_18317,N_18288);
and U18512 (N_18512,N_18278,N_18293);
and U18513 (N_18513,N_18311,N_18445);
nand U18514 (N_18514,N_18322,N_18251);
nor U18515 (N_18515,N_18393,N_18496);
nand U18516 (N_18516,N_18489,N_18345);
xnor U18517 (N_18517,N_18438,N_18309);
nor U18518 (N_18518,N_18255,N_18250);
nand U18519 (N_18519,N_18291,N_18478);
or U18520 (N_18520,N_18352,N_18376);
nor U18521 (N_18521,N_18396,N_18480);
and U18522 (N_18522,N_18481,N_18477);
and U18523 (N_18523,N_18454,N_18363);
nor U18524 (N_18524,N_18353,N_18372);
nor U18525 (N_18525,N_18474,N_18410);
xor U18526 (N_18526,N_18308,N_18463);
xnor U18527 (N_18527,N_18304,N_18423);
xor U18528 (N_18528,N_18327,N_18273);
or U18529 (N_18529,N_18325,N_18303);
or U18530 (N_18530,N_18349,N_18447);
and U18531 (N_18531,N_18287,N_18290);
nand U18532 (N_18532,N_18275,N_18407);
xor U18533 (N_18533,N_18295,N_18421);
and U18534 (N_18534,N_18446,N_18417);
nand U18535 (N_18535,N_18461,N_18470);
and U18536 (N_18536,N_18358,N_18483);
and U18537 (N_18537,N_18413,N_18348);
or U18538 (N_18538,N_18310,N_18263);
or U18539 (N_18539,N_18261,N_18324);
xor U18540 (N_18540,N_18335,N_18448);
and U18541 (N_18541,N_18462,N_18355);
nand U18542 (N_18542,N_18280,N_18371);
xor U18543 (N_18543,N_18331,N_18406);
and U18544 (N_18544,N_18440,N_18418);
nand U18545 (N_18545,N_18476,N_18374);
or U18546 (N_18546,N_18258,N_18386);
and U18547 (N_18547,N_18299,N_18464);
nand U18548 (N_18548,N_18395,N_18443);
nand U18549 (N_18549,N_18276,N_18254);
or U18550 (N_18550,N_18387,N_18404);
nor U18551 (N_18551,N_18384,N_18424);
and U18552 (N_18552,N_18366,N_18377);
nor U18553 (N_18553,N_18260,N_18419);
and U18554 (N_18554,N_18495,N_18433);
nand U18555 (N_18555,N_18294,N_18493);
or U18556 (N_18556,N_18257,N_18449);
nor U18557 (N_18557,N_18334,N_18341);
and U18558 (N_18558,N_18465,N_18343);
xnor U18559 (N_18559,N_18467,N_18427);
or U18560 (N_18560,N_18456,N_18475);
nor U18561 (N_18561,N_18442,N_18432);
nor U18562 (N_18562,N_18297,N_18326);
nand U18563 (N_18563,N_18488,N_18459);
nand U18564 (N_18564,N_18356,N_18460);
and U18565 (N_18565,N_18498,N_18411);
and U18566 (N_18566,N_18468,N_18473);
xor U18567 (N_18567,N_18379,N_18430);
nand U18568 (N_18568,N_18408,N_18270);
nand U18569 (N_18569,N_18262,N_18415);
nand U18570 (N_18570,N_18450,N_18333);
nand U18571 (N_18571,N_18370,N_18472);
xnor U18572 (N_18572,N_18329,N_18347);
nand U18573 (N_18573,N_18405,N_18367);
nand U18574 (N_18574,N_18330,N_18401);
and U18575 (N_18575,N_18274,N_18296);
nor U18576 (N_18576,N_18316,N_18437);
nand U18577 (N_18577,N_18256,N_18390);
nand U18578 (N_18578,N_18494,N_18455);
or U18579 (N_18579,N_18383,N_18409);
or U18580 (N_18580,N_18365,N_18298);
nand U18581 (N_18581,N_18361,N_18499);
and U18582 (N_18582,N_18458,N_18319);
nand U18583 (N_18583,N_18300,N_18312);
nand U18584 (N_18584,N_18403,N_18441);
nor U18585 (N_18585,N_18416,N_18429);
or U18586 (N_18586,N_18487,N_18368);
and U18587 (N_18587,N_18373,N_18267);
nand U18588 (N_18588,N_18350,N_18399);
nand U18589 (N_18589,N_18285,N_18482);
nor U18590 (N_18590,N_18359,N_18382);
and U18591 (N_18591,N_18321,N_18388);
nor U18592 (N_18592,N_18265,N_18271);
and U18593 (N_18593,N_18431,N_18397);
and U18594 (N_18594,N_18344,N_18385);
xor U18595 (N_18595,N_18305,N_18479);
and U18596 (N_18596,N_18490,N_18252);
xnor U18597 (N_18597,N_18272,N_18277);
and U18598 (N_18598,N_18497,N_18471);
xnor U18599 (N_18599,N_18253,N_18318);
xor U18600 (N_18600,N_18268,N_18457);
xor U18601 (N_18601,N_18284,N_18313);
nand U18602 (N_18602,N_18422,N_18378);
xnor U18603 (N_18603,N_18289,N_18269);
nand U18604 (N_18604,N_18420,N_18314);
nand U18605 (N_18605,N_18266,N_18369);
nor U18606 (N_18606,N_18439,N_18484);
xor U18607 (N_18607,N_18339,N_18491);
and U18608 (N_18608,N_18342,N_18323);
or U18609 (N_18609,N_18389,N_18453);
and U18610 (N_18610,N_18306,N_18286);
xnor U18611 (N_18611,N_18302,N_18283);
xnor U18612 (N_18612,N_18357,N_18336);
nand U18613 (N_18613,N_18380,N_18452);
nor U18614 (N_18614,N_18392,N_18301);
nor U18615 (N_18615,N_18436,N_18451);
and U18616 (N_18616,N_18426,N_18375);
or U18617 (N_18617,N_18362,N_18282);
nand U18618 (N_18618,N_18414,N_18279);
nor U18619 (N_18619,N_18259,N_18492);
or U18620 (N_18620,N_18281,N_18400);
or U18621 (N_18621,N_18435,N_18486);
and U18622 (N_18622,N_18425,N_18315);
xnor U18623 (N_18623,N_18307,N_18320);
and U18624 (N_18624,N_18346,N_18391);
nor U18625 (N_18625,N_18408,N_18254);
nor U18626 (N_18626,N_18254,N_18438);
or U18627 (N_18627,N_18285,N_18493);
xnor U18628 (N_18628,N_18418,N_18307);
xnor U18629 (N_18629,N_18379,N_18475);
nor U18630 (N_18630,N_18378,N_18434);
xor U18631 (N_18631,N_18387,N_18424);
nor U18632 (N_18632,N_18474,N_18335);
and U18633 (N_18633,N_18395,N_18432);
nor U18634 (N_18634,N_18382,N_18299);
or U18635 (N_18635,N_18379,N_18259);
xnor U18636 (N_18636,N_18466,N_18440);
or U18637 (N_18637,N_18352,N_18320);
xor U18638 (N_18638,N_18408,N_18483);
xor U18639 (N_18639,N_18260,N_18380);
xnor U18640 (N_18640,N_18251,N_18389);
and U18641 (N_18641,N_18276,N_18376);
xor U18642 (N_18642,N_18484,N_18449);
and U18643 (N_18643,N_18326,N_18497);
xor U18644 (N_18644,N_18265,N_18422);
and U18645 (N_18645,N_18282,N_18453);
nand U18646 (N_18646,N_18442,N_18429);
or U18647 (N_18647,N_18286,N_18362);
nand U18648 (N_18648,N_18278,N_18433);
nor U18649 (N_18649,N_18455,N_18261);
or U18650 (N_18650,N_18254,N_18454);
nand U18651 (N_18651,N_18367,N_18340);
nand U18652 (N_18652,N_18343,N_18319);
and U18653 (N_18653,N_18303,N_18422);
nor U18654 (N_18654,N_18335,N_18338);
nor U18655 (N_18655,N_18352,N_18375);
nor U18656 (N_18656,N_18264,N_18327);
and U18657 (N_18657,N_18311,N_18484);
nand U18658 (N_18658,N_18473,N_18414);
or U18659 (N_18659,N_18388,N_18259);
nand U18660 (N_18660,N_18305,N_18499);
nand U18661 (N_18661,N_18343,N_18442);
xnor U18662 (N_18662,N_18350,N_18377);
nor U18663 (N_18663,N_18268,N_18412);
and U18664 (N_18664,N_18253,N_18379);
nor U18665 (N_18665,N_18370,N_18366);
nor U18666 (N_18666,N_18251,N_18279);
xnor U18667 (N_18667,N_18366,N_18312);
xnor U18668 (N_18668,N_18441,N_18339);
nor U18669 (N_18669,N_18384,N_18391);
nand U18670 (N_18670,N_18384,N_18315);
and U18671 (N_18671,N_18312,N_18422);
or U18672 (N_18672,N_18491,N_18278);
or U18673 (N_18673,N_18298,N_18483);
nand U18674 (N_18674,N_18407,N_18256);
nor U18675 (N_18675,N_18383,N_18333);
xor U18676 (N_18676,N_18374,N_18391);
and U18677 (N_18677,N_18380,N_18358);
nand U18678 (N_18678,N_18402,N_18495);
and U18679 (N_18679,N_18397,N_18354);
xor U18680 (N_18680,N_18364,N_18312);
nand U18681 (N_18681,N_18490,N_18416);
nor U18682 (N_18682,N_18464,N_18476);
or U18683 (N_18683,N_18455,N_18349);
nand U18684 (N_18684,N_18376,N_18416);
nand U18685 (N_18685,N_18381,N_18346);
nand U18686 (N_18686,N_18302,N_18427);
and U18687 (N_18687,N_18251,N_18329);
nand U18688 (N_18688,N_18460,N_18254);
and U18689 (N_18689,N_18347,N_18290);
and U18690 (N_18690,N_18427,N_18376);
nand U18691 (N_18691,N_18285,N_18454);
nand U18692 (N_18692,N_18423,N_18275);
or U18693 (N_18693,N_18432,N_18436);
and U18694 (N_18694,N_18439,N_18442);
xor U18695 (N_18695,N_18383,N_18323);
xnor U18696 (N_18696,N_18345,N_18284);
xnor U18697 (N_18697,N_18384,N_18357);
nor U18698 (N_18698,N_18303,N_18265);
nand U18699 (N_18699,N_18261,N_18433);
nand U18700 (N_18700,N_18404,N_18451);
nor U18701 (N_18701,N_18283,N_18351);
nand U18702 (N_18702,N_18425,N_18342);
or U18703 (N_18703,N_18369,N_18409);
nand U18704 (N_18704,N_18329,N_18446);
or U18705 (N_18705,N_18279,N_18327);
or U18706 (N_18706,N_18294,N_18295);
nand U18707 (N_18707,N_18391,N_18269);
xor U18708 (N_18708,N_18278,N_18485);
or U18709 (N_18709,N_18297,N_18391);
xnor U18710 (N_18710,N_18293,N_18440);
or U18711 (N_18711,N_18300,N_18438);
nor U18712 (N_18712,N_18476,N_18275);
and U18713 (N_18713,N_18254,N_18252);
nor U18714 (N_18714,N_18360,N_18407);
or U18715 (N_18715,N_18398,N_18472);
or U18716 (N_18716,N_18380,N_18459);
nand U18717 (N_18717,N_18305,N_18460);
nor U18718 (N_18718,N_18401,N_18443);
and U18719 (N_18719,N_18381,N_18387);
nor U18720 (N_18720,N_18341,N_18484);
and U18721 (N_18721,N_18265,N_18285);
and U18722 (N_18722,N_18417,N_18381);
nor U18723 (N_18723,N_18478,N_18321);
nor U18724 (N_18724,N_18390,N_18458);
xnor U18725 (N_18725,N_18464,N_18258);
nor U18726 (N_18726,N_18414,N_18462);
or U18727 (N_18727,N_18407,N_18295);
or U18728 (N_18728,N_18465,N_18397);
and U18729 (N_18729,N_18470,N_18253);
or U18730 (N_18730,N_18452,N_18297);
and U18731 (N_18731,N_18468,N_18397);
or U18732 (N_18732,N_18258,N_18331);
and U18733 (N_18733,N_18303,N_18299);
and U18734 (N_18734,N_18373,N_18347);
or U18735 (N_18735,N_18465,N_18327);
xor U18736 (N_18736,N_18321,N_18411);
or U18737 (N_18737,N_18423,N_18357);
or U18738 (N_18738,N_18294,N_18335);
and U18739 (N_18739,N_18350,N_18295);
nor U18740 (N_18740,N_18433,N_18460);
xnor U18741 (N_18741,N_18273,N_18462);
or U18742 (N_18742,N_18357,N_18315);
nor U18743 (N_18743,N_18407,N_18291);
nor U18744 (N_18744,N_18463,N_18323);
nor U18745 (N_18745,N_18370,N_18377);
xor U18746 (N_18746,N_18326,N_18383);
xor U18747 (N_18747,N_18408,N_18496);
or U18748 (N_18748,N_18384,N_18271);
nand U18749 (N_18749,N_18410,N_18308);
xnor U18750 (N_18750,N_18593,N_18709);
nor U18751 (N_18751,N_18700,N_18620);
and U18752 (N_18752,N_18743,N_18587);
or U18753 (N_18753,N_18534,N_18515);
and U18754 (N_18754,N_18637,N_18598);
and U18755 (N_18755,N_18522,N_18726);
nor U18756 (N_18756,N_18652,N_18705);
nor U18757 (N_18757,N_18591,N_18514);
nand U18758 (N_18758,N_18539,N_18551);
xor U18759 (N_18759,N_18579,N_18502);
xnor U18760 (N_18760,N_18675,N_18578);
nor U18761 (N_18761,N_18524,N_18537);
and U18762 (N_18762,N_18626,N_18692);
xnor U18763 (N_18763,N_18658,N_18544);
and U18764 (N_18764,N_18733,N_18684);
nand U18765 (N_18765,N_18546,N_18582);
and U18766 (N_18766,N_18623,N_18628);
nand U18767 (N_18767,N_18670,N_18633);
nor U18768 (N_18768,N_18535,N_18569);
or U18769 (N_18769,N_18563,N_18744);
nor U18770 (N_18770,N_18717,N_18636);
or U18771 (N_18771,N_18559,N_18560);
xnor U18772 (N_18772,N_18592,N_18666);
xnor U18773 (N_18773,N_18523,N_18631);
or U18774 (N_18774,N_18727,N_18568);
and U18775 (N_18775,N_18525,N_18610);
or U18776 (N_18776,N_18635,N_18695);
nand U18777 (N_18777,N_18708,N_18714);
or U18778 (N_18778,N_18629,N_18528);
nand U18779 (N_18779,N_18734,N_18698);
or U18780 (N_18780,N_18682,N_18580);
xor U18781 (N_18781,N_18719,N_18701);
nor U18782 (N_18782,N_18645,N_18651);
and U18783 (N_18783,N_18543,N_18596);
nand U18784 (N_18784,N_18737,N_18627);
and U18785 (N_18785,N_18672,N_18589);
xnor U18786 (N_18786,N_18606,N_18527);
nand U18787 (N_18787,N_18621,N_18601);
or U18788 (N_18788,N_18731,N_18664);
xor U18789 (N_18789,N_18736,N_18584);
nor U18790 (N_18790,N_18630,N_18595);
nand U18791 (N_18791,N_18632,N_18558);
and U18792 (N_18792,N_18583,N_18590);
xnor U18793 (N_18793,N_18740,N_18653);
or U18794 (N_18794,N_18696,N_18639);
xnor U18795 (N_18795,N_18612,N_18564);
nand U18796 (N_18796,N_18641,N_18570);
or U18797 (N_18797,N_18644,N_18713);
nand U18798 (N_18798,N_18691,N_18741);
nor U18799 (N_18799,N_18616,N_18575);
nand U18800 (N_18800,N_18510,N_18536);
or U18801 (N_18801,N_18723,N_18566);
and U18802 (N_18802,N_18573,N_18724);
nand U18803 (N_18803,N_18619,N_18703);
nor U18804 (N_18804,N_18683,N_18605);
nand U18805 (N_18805,N_18561,N_18694);
xor U18806 (N_18806,N_18676,N_18607);
nor U18807 (N_18807,N_18702,N_18681);
nand U18808 (N_18808,N_18690,N_18716);
nor U18809 (N_18809,N_18545,N_18625);
nand U18810 (N_18810,N_18665,N_18687);
nand U18811 (N_18811,N_18688,N_18655);
nor U18812 (N_18812,N_18745,N_18618);
nand U18813 (N_18813,N_18585,N_18686);
nand U18814 (N_18814,N_18728,N_18549);
nor U18815 (N_18815,N_18624,N_18602);
xor U18816 (N_18816,N_18507,N_18689);
xor U18817 (N_18817,N_18553,N_18519);
or U18818 (N_18818,N_18503,N_18597);
or U18819 (N_18819,N_18529,N_18646);
xnor U18820 (N_18820,N_18574,N_18746);
xor U18821 (N_18821,N_18600,N_18648);
or U18822 (N_18822,N_18656,N_18530);
nand U18823 (N_18823,N_18729,N_18643);
nor U18824 (N_18824,N_18667,N_18715);
nor U18825 (N_18825,N_18697,N_18538);
nor U18826 (N_18826,N_18571,N_18506);
or U18827 (N_18827,N_18581,N_18668);
or U18828 (N_18828,N_18532,N_18622);
nor U18829 (N_18829,N_18547,N_18517);
xnor U18830 (N_18830,N_18699,N_18604);
nand U18831 (N_18831,N_18548,N_18680);
xor U18832 (N_18832,N_18674,N_18611);
xnor U18833 (N_18833,N_18640,N_18603);
or U18834 (N_18834,N_18642,N_18531);
nand U18835 (N_18835,N_18725,N_18511);
nor U18836 (N_18836,N_18660,N_18533);
or U18837 (N_18837,N_18565,N_18710);
nand U18838 (N_18838,N_18718,N_18613);
xnor U18839 (N_18839,N_18671,N_18673);
nor U18840 (N_18840,N_18550,N_18540);
nor U18841 (N_18841,N_18742,N_18541);
nand U18842 (N_18842,N_18730,N_18614);
or U18843 (N_18843,N_18738,N_18512);
and U18844 (N_18844,N_18526,N_18685);
or U18845 (N_18845,N_18654,N_18693);
xnor U18846 (N_18846,N_18501,N_18707);
and U18847 (N_18847,N_18554,N_18748);
nand U18848 (N_18848,N_18555,N_18678);
or U18849 (N_18849,N_18749,N_18594);
and U18850 (N_18850,N_18567,N_18706);
nor U18851 (N_18851,N_18513,N_18663);
xnor U18852 (N_18852,N_18552,N_18588);
nor U18853 (N_18853,N_18609,N_18577);
xnor U18854 (N_18854,N_18679,N_18721);
or U18855 (N_18855,N_18557,N_18661);
and U18856 (N_18856,N_18556,N_18650);
nor U18857 (N_18857,N_18516,N_18608);
and U18858 (N_18858,N_18562,N_18634);
xor U18859 (N_18859,N_18732,N_18662);
nor U18860 (N_18860,N_18711,N_18504);
and U18861 (N_18861,N_18500,N_18647);
xor U18862 (N_18862,N_18720,N_18586);
nor U18863 (N_18863,N_18712,N_18704);
and U18864 (N_18864,N_18722,N_18669);
or U18865 (N_18865,N_18572,N_18508);
nor U18866 (N_18866,N_18657,N_18520);
nand U18867 (N_18867,N_18542,N_18599);
or U18868 (N_18868,N_18617,N_18649);
and U18869 (N_18869,N_18518,N_18659);
or U18870 (N_18870,N_18638,N_18615);
and U18871 (N_18871,N_18735,N_18576);
nor U18872 (N_18872,N_18677,N_18521);
xor U18873 (N_18873,N_18509,N_18739);
nor U18874 (N_18874,N_18505,N_18747);
or U18875 (N_18875,N_18593,N_18526);
nand U18876 (N_18876,N_18578,N_18595);
or U18877 (N_18877,N_18637,N_18742);
and U18878 (N_18878,N_18704,N_18692);
or U18879 (N_18879,N_18608,N_18661);
xnor U18880 (N_18880,N_18594,N_18688);
or U18881 (N_18881,N_18709,N_18665);
and U18882 (N_18882,N_18649,N_18521);
or U18883 (N_18883,N_18560,N_18639);
nand U18884 (N_18884,N_18723,N_18647);
xor U18885 (N_18885,N_18718,N_18736);
or U18886 (N_18886,N_18519,N_18712);
nor U18887 (N_18887,N_18538,N_18708);
xnor U18888 (N_18888,N_18510,N_18513);
or U18889 (N_18889,N_18620,N_18558);
and U18890 (N_18890,N_18710,N_18661);
and U18891 (N_18891,N_18739,N_18719);
nand U18892 (N_18892,N_18528,N_18668);
xnor U18893 (N_18893,N_18676,N_18643);
nand U18894 (N_18894,N_18684,N_18602);
and U18895 (N_18895,N_18744,N_18537);
and U18896 (N_18896,N_18688,N_18724);
xnor U18897 (N_18897,N_18715,N_18568);
nand U18898 (N_18898,N_18630,N_18662);
or U18899 (N_18899,N_18673,N_18586);
nor U18900 (N_18900,N_18585,N_18506);
and U18901 (N_18901,N_18694,N_18714);
xnor U18902 (N_18902,N_18669,N_18681);
and U18903 (N_18903,N_18639,N_18541);
nand U18904 (N_18904,N_18500,N_18540);
and U18905 (N_18905,N_18527,N_18630);
nand U18906 (N_18906,N_18625,N_18662);
nor U18907 (N_18907,N_18580,N_18541);
nor U18908 (N_18908,N_18562,N_18686);
or U18909 (N_18909,N_18501,N_18646);
nor U18910 (N_18910,N_18522,N_18619);
xnor U18911 (N_18911,N_18628,N_18532);
xor U18912 (N_18912,N_18532,N_18650);
nor U18913 (N_18913,N_18575,N_18675);
nor U18914 (N_18914,N_18535,N_18542);
and U18915 (N_18915,N_18540,N_18717);
nor U18916 (N_18916,N_18715,N_18612);
nand U18917 (N_18917,N_18625,N_18675);
nor U18918 (N_18918,N_18551,N_18700);
and U18919 (N_18919,N_18742,N_18728);
and U18920 (N_18920,N_18535,N_18520);
xnor U18921 (N_18921,N_18563,N_18737);
and U18922 (N_18922,N_18599,N_18645);
nor U18923 (N_18923,N_18586,N_18744);
or U18924 (N_18924,N_18569,N_18584);
or U18925 (N_18925,N_18625,N_18524);
nor U18926 (N_18926,N_18564,N_18580);
and U18927 (N_18927,N_18647,N_18524);
or U18928 (N_18928,N_18574,N_18505);
or U18929 (N_18929,N_18530,N_18592);
nand U18930 (N_18930,N_18644,N_18679);
xnor U18931 (N_18931,N_18547,N_18522);
xor U18932 (N_18932,N_18511,N_18661);
nor U18933 (N_18933,N_18502,N_18566);
nor U18934 (N_18934,N_18612,N_18676);
nand U18935 (N_18935,N_18651,N_18646);
xnor U18936 (N_18936,N_18540,N_18591);
or U18937 (N_18937,N_18546,N_18649);
or U18938 (N_18938,N_18659,N_18712);
nand U18939 (N_18939,N_18528,N_18611);
and U18940 (N_18940,N_18738,N_18560);
nor U18941 (N_18941,N_18602,N_18697);
xnor U18942 (N_18942,N_18561,N_18566);
or U18943 (N_18943,N_18604,N_18520);
xnor U18944 (N_18944,N_18572,N_18709);
nand U18945 (N_18945,N_18514,N_18641);
nand U18946 (N_18946,N_18666,N_18564);
and U18947 (N_18947,N_18670,N_18731);
nand U18948 (N_18948,N_18669,N_18619);
nor U18949 (N_18949,N_18742,N_18679);
nand U18950 (N_18950,N_18555,N_18693);
and U18951 (N_18951,N_18619,N_18583);
or U18952 (N_18952,N_18521,N_18672);
or U18953 (N_18953,N_18740,N_18643);
and U18954 (N_18954,N_18608,N_18522);
nor U18955 (N_18955,N_18707,N_18503);
xor U18956 (N_18956,N_18642,N_18737);
nand U18957 (N_18957,N_18554,N_18651);
and U18958 (N_18958,N_18723,N_18636);
or U18959 (N_18959,N_18528,N_18686);
or U18960 (N_18960,N_18694,N_18553);
and U18961 (N_18961,N_18541,N_18661);
xor U18962 (N_18962,N_18720,N_18684);
and U18963 (N_18963,N_18598,N_18711);
and U18964 (N_18964,N_18748,N_18501);
nor U18965 (N_18965,N_18650,N_18573);
nand U18966 (N_18966,N_18651,N_18696);
or U18967 (N_18967,N_18598,N_18594);
nor U18968 (N_18968,N_18573,N_18709);
and U18969 (N_18969,N_18679,N_18526);
and U18970 (N_18970,N_18653,N_18635);
xor U18971 (N_18971,N_18677,N_18704);
and U18972 (N_18972,N_18727,N_18636);
nand U18973 (N_18973,N_18740,N_18512);
nand U18974 (N_18974,N_18552,N_18562);
nor U18975 (N_18975,N_18603,N_18505);
nand U18976 (N_18976,N_18707,N_18591);
nor U18977 (N_18977,N_18565,N_18604);
and U18978 (N_18978,N_18557,N_18643);
nand U18979 (N_18979,N_18704,N_18676);
nor U18980 (N_18980,N_18655,N_18630);
or U18981 (N_18981,N_18647,N_18711);
or U18982 (N_18982,N_18672,N_18607);
nor U18983 (N_18983,N_18588,N_18665);
nand U18984 (N_18984,N_18685,N_18670);
or U18985 (N_18985,N_18592,N_18509);
xor U18986 (N_18986,N_18608,N_18518);
or U18987 (N_18987,N_18557,N_18686);
and U18988 (N_18988,N_18691,N_18556);
xor U18989 (N_18989,N_18654,N_18713);
nor U18990 (N_18990,N_18500,N_18723);
and U18991 (N_18991,N_18697,N_18521);
and U18992 (N_18992,N_18622,N_18698);
or U18993 (N_18993,N_18657,N_18578);
nand U18994 (N_18994,N_18620,N_18516);
and U18995 (N_18995,N_18565,N_18636);
or U18996 (N_18996,N_18612,N_18607);
and U18997 (N_18997,N_18569,N_18739);
or U18998 (N_18998,N_18711,N_18674);
and U18999 (N_18999,N_18613,N_18554);
and U19000 (N_19000,N_18902,N_18907);
nor U19001 (N_19001,N_18955,N_18937);
or U19002 (N_19002,N_18842,N_18914);
and U19003 (N_19003,N_18910,N_18808);
nand U19004 (N_19004,N_18767,N_18807);
and U19005 (N_19005,N_18828,N_18831);
nor U19006 (N_19006,N_18980,N_18860);
or U19007 (N_19007,N_18809,N_18838);
or U19008 (N_19008,N_18965,N_18868);
or U19009 (N_19009,N_18909,N_18953);
xor U19010 (N_19010,N_18879,N_18781);
xnor U19011 (N_19011,N_18834,N_18755);
nor U19012 (N_19012,N_18815,N_18797);
nor U19013 (N_19013,N_18811,N_18950);
xor U19014 (N_19014,N_18986,N_18863);
or U19015 (N_19015,N_18941,N_18867);
or U19016 (N_19016,N_18787,N_18819);
nand U19017 (N_19017,N_18888,N_18946);
xor U19018 (N_19018,N_18821,N_18843);
and U19019 (N_19019,N_18794,N_18785);
nand U19020 (N_19020,N_18874,N_18939);
and U19021 (N_19021,N_18938,N_18885);
nor U19022 (N_19022,N_18791,N_18964);
xnor U19023 (N_19023,N_18873,N_18792);
and U19024 (N_19024,N_18833,N_18816);
nor U19025 (N_19025,N_18884,N_18793);
nand U19026 (N_19026,N_18853,N_18890);
nor U19027 (N_19027,N_18927,N_18799);
and U19028 (N_19028,N_18786,N_18775);
xnor U19029 (N_19029,N_18958,N_18857);
nand U19030 (N_19030,N_18948,N_18957);
and U19031 (N_19031,N_18920,N_18998);
and U19032 (N_19032,N_18855,N_18766);
and U19033 (N_19033,N_18974,N_18899);
nand U19034 (N_19034,N_18844,N_18881);
and U19035 (N_19035,N_18795,N_18764);
and U19036 (N_19036,N_18829,N_18915);
nand U19037 (N_19037,N_18901,N_18886);
or U19038 (N_19038,N_18825,N_18897);
xnor U19039 (N_19039,N_18753,N_18973);
nand U19040 (N_19040,N_18782,N_18960);
xnor U19041 (N_19041,N_18846,N_18845);
nand U19042 (N_19042,N_18759,N_18994);
or U19043 (N_19043,N_18752,N_18878);
xnor U19044 (N_19044,N_18985,N_18898);
or U19045 (N_19045,N_18977,N_18911);
or U19046 (N_19046,N_18757,N_18996);
or U19047 (N_19047,N_18817,N_18944);
nor U19048 (N_19048,N_18943,N_18850);
or U19049 (N_19049,N_18959,N_18777);
nor U19050 (N_19050,N_18771,N_18923);
or U19051 (N_19051,N_18913,N_18989);
nand U19052 (N_19052,N_18768,N_18999);
and U19053 (N_19053,N_18983,N_18796);
or U19054 (N_19054,N_18991,N_18990);
or U19055 (N_19055,N_18848,N_18849);
and U19056 (N_19056,N_18905,N_18904);
and U19057 (N_19057,N_18967,N_18952);
nor U19058 (N_19058,N_18949,N_18981);
nor U19059 (N_19059,N_18798,N_18827);
nand U19060 (N_19060,N_18945,N_18880);
xnor U19061 (N_19061,N_18803,N_18876);
nor U19062 (N_19062,N_18887,N_18783);
nor U19063 (N_19063,N_18954,N_18971);
nand U19064 (N_19064,N_18784,N_18839);
and U19065 (N_19065,N_18751,N_18818);
and U19066 (N_19066,N_18925,N_18963);
nor U19067 (N_19067,N_18832,N_18896);
nand U19068 (N_19068,N_18922,N_18800);
and U19069 (N_19069,N_18758,N_18988);
nor U19070 (N_19070,N_18822,N_18810);
xnor U19071 (N_19071,N_18979,N_18956);
and U19072 (N_19072,N_18864,N_18856);
nor U19073 (N_19073,N_18987,N_18840);
xnor U19074 (N_19074,N_18761,N_18961);
and U19075 (N_19075,N_18760,N_18895);
nor U19076 (N_19076,N_18984,N_18823);
and U19077 (N_19077,N_18916,N_18847);
xnor U19078 (N_19078,N_18893,N_18936);
or U19079 (N_19079,N_18778,N_18789);
nand U19080 (N_19080,N_18870,N_18892);
nand U19081 (N_19081,N_18804,N_18756);
or U19082 (N_19082,N_18773,N_18862);
and U19083 (N_19083,N_18851,N_18805);
nor U19084 (N_19084,N_18866,N_18951);
or U19085 (N_19085,N_18982,N_18933);
or U19086 (N_19086,N_18934,N_18801);
nand U19087 (N_19087,N_18770,N_18932);
xnor U19088 (N_19088,N_18772,N_18894);
or U19089 (N_19089,N_18820,N_18869);
or U19090 (N_19090,N_18776,N_18877);
nor U19091 (N_19091,N_18774,N_18969);
or U19092 (N_19092,N_18763,N_18872);
or U19093 (N_19093,N_18802,N_18917);
nand U19094 (N_19094,N_18900,N_18995);
nand U19095 (N_19095,N_18769,N_18812);
nand U19096 (N_19096,N_18930,N_18972);
nand U19097 (N_19097,N_18826,N_18942);
xnor U19098 (N_19098,N_18806,N_18931);
or U19099 (N_19099,N_18889,N_18968);
xnor U19100 (N_19100,N_18765,N_18908);
nand U19101 (N_19101,N_18762,N_18919);
or U19102 (N_19102,N_18871,N_18830);
nor U19103 (N_19103,N_18858,N_18940);
and U19104 (N_19104,N_18935,N_18859);
or U19105 (N_19105,N_18924,N_18854);
nor U19106 (N_19106,N_18836,N_18962);
nor U19107 (N_19107,N_18978,N_18918);
nor U19108 (N_19108,N_18837,N_18790);
or U19109 (N_19109,N_18966,N_18906);
or U19110 (N_19110,N_18813,N_18992);
xor U19111 (N_19111,N_18865,N_18947);
or U19112 (N_19112,N_18835,N_18921);
nor U19113 (N_19113,N_18882,N_18852);
and U19114 (N_19114,N_18754,N_18780);
xnor U19115 (N_19115,N_18875,N_18975);
nor U19116 (N_19116,N_18997,N_18861);
nor U19117 (N_19117,N_18976,N_18824);
nor U19118 (N_19118,N_18993,N_18928);
nor U19119 (N_19119,N_18779,N_18814);
or U19120 (N_19120,N_18841,N_18929);
nand U19121 (N_19121,N_18903,N_18891);
nor U19122 (N_19122,N_18970,N_18788);
nor U19123 (N_19123,N_18912,N_18750);
xnor U19124 (N_19124,N_18926,N_18883);
nand U19125 (N_19125,N_18967,N_18905);
and U19126 (N_19126,N_18974,N_18996);
xnor U19127 (N_19127,N_18981,N_18857);
or U19128 (N_19128,N_18798,N_18797);
and U19129 (N_19129,N_18924,N_18869);
nor U19130 (N_19130,N_18753,N_18880);
nand U19131 (N_19131,N_18884,N_18860);
xor U19132 (N_19132,N_18889,N_18883);
nor U19133 (N_19133,N_18946,N_18986);
xnor U19134 (N_19134,N_18845,N_18955);
nand U19135 (N_19135,N_18805,N_18912);
nor U19136 (N_19136,N_18849,N_18863);
or U19137 (N_19137,N_18948,N_18905);
nor U19138 (N_19138,N_18751,N_18972);
nor U19139 (N_19139,N_18963,N_18779);
and U19140 (N_19140,N_18924,N_18754);
and U19141 (N_19141,N_18938,N_18972);
and U19142 (N_19142,N_18981,N_18816);
or U19143 (N_19143,N_18894,N_18933);
and U19144 (N_19144,N_18776,N_18887);
nand U19145 (N_19145,N_18839,N_18769);
or U19146 (N_19146,N_18821,N_18924);
nor U19147 (N_19147,N_18752,N_18818);
xnor U19148 (N_19148,N_18945,N_18926);
nand U19149 (N_19149,N_18877,N_18910);
nand U19150 (N_19150,N_18778,N_18850);
nor U19151 (N_19151,N_18947,N_18768);
or U19152 (N_19152,N_18787,N_18785);
nand U19153 (N_19153,N_18906,N_18891);
nor U19154 (N_19154,N_18836,N_18878);
xor U19155 (N_19155,N_18960,N_18827);
xnor U19156 (N_19156,N_18822,N_18959);
or U19157 (N_19157,N_18914,N_18958);
xor U19158 (N_19158,N_18948,N_18865);
or U19159 (N_19159,N_18751,N_18900);
nand U19160 (N_19160,N_18852,N_18867);
and U19161 (N_19161,N_18802,N_18913);
and U19162 (N_19162,N_18836,N_18928);
xor U19163 (N_19163,N_18766,N_18794);
or U19164 (N_19164,N_18995,N_18758);
xnor U19165 (N_19165,N_18863,N_18950);
xor U19166 (N_19166,N_18830,N_18934);
and U19167 (N_19167,N_18894,N_18958);
xnor U19168 (N_19168,N_18838,N_18881);
nand U19169 (N_19169,N_18916,N_18767);
or U19170 (N_19170,N_18844,N_18823);
and U19171 (N_19171,N_18922,N_18830);
and U19172 (N_19172,N_18779,N_18941);
xor U19173 (N_19173,N_18821,N_18770);
nand U19174 (N_19174,N_18829,N_18751);
xnor U19175 (N_19175,N_18799,N_18868);
or U19176 (N_19176,N_18804,N_18848);
or U19177 (N_19177,N_18827,N_18935);
nor U19178 (N_19178,N_18916,N_18869);
nand U19179 (N_19179,N_18807,N_18768);
and U19180 (N_19180,N_18883,N_18971);
or U19181 (N_19181,N_18901,N_18750);
or U19182 (N_19182,N_18945,N_18752);
nor U19183 (N_19183,N_18827,N_18816);
or U19184 (N_19184,N_18997,N_18983);
nand U19185 (N_19185,N_18889,N_18879);
and U19186 (N_19186,N_18930,N_18948);
xnor U19187 (N_19187,N_18849,N_18795);
nand U19188 (N_19188,N_18812,N_18815);
or U19189 (N_19189,N_18826,N_18754);
nor U19190 (N_19190,N_18887,N_18922);
nand U19191 (N_19191,N_18926,N_18859);
or U19192 (N_19192,N_18803,N_18787);
and U19193 (N_19193,N_18923,N_18897);
nor U19194 (N_19194,N_18914,N_18946);
nor U19195 (N_19195,N_18791,N_18877);
and U19196 (N_19196,N_18869,N_18939);
nand U19197 (N_19197,N_18812,N_18954);
nor U19198 (N_19198,N_18755,N_18851);
and U19199 (N_19199,N_18872,N_18842);
nor U19200 (N_19200,N_18804,N_18968);
xnor U19201 (N_19201,N_18835,N_18931);
nor U19202 (N_19202,N_18885,N_18784);
or U19203 (N_19203,N_18974,N_18808);
nor U19204 (N_19204,N_18965,N_18892);
or U19205 (N_19205,N_18963,N_18958);
or U19206 (N_19206,N_18811,N_18933);
nor U19207 (N_19207,N_18823,N_18882);
xnor U19208 (N_19208,N_18786,N_18827);
or U19209 (N_19209,N_18784,N_18755);
nor U19210 (N_19210,N_18756,N_18900);
and U19211 (N_19211,N_18909,N_18880);
and U19212 (N_19212,N_18840,N_18829);
or U19213 (N_19213,N_18891,N_18867);
nand U19214 (N_19214,N_18955,N_18886);
xor U19215 (N_19215,N_18771,N_18909);
nand U19216 (N_19216,N_18793,N_18824);
and U19217 (N_19217,N_18846,N_18914);
nor U19218 (N_19218,N_18846,N_18858);
xnor U19219 (N_19219,N_18837,N_18912);
and U19220 (N_19220,N_18850,N_18950);
xor U19221 (N_19221,N_18970,N_18847);
and U19222 (N_19222,N_18816,N_18962);
nand U19223 (N_19223,N_18856,N_18800);
xor U19224 (N_19224,N_18760,N_18818);
nor U19225 (N_19225,N_18765,N_18800);
and U19226 (N_19226,N_18775,N_18974);
and U19227 (N_19227,N_18850,N_18802);
and U19228 (N_19228,N_18957,N_18893);
xor U19229 (N_19229,N_18839,N_18876);
nand U19230 (N_19230,N_18849,N_18905);
nand U19231 (N_19231,N_18874,N_18955);
nor U19232 (N_19232,N_18774,N_18962);
or U19233 (N_19233,N_18823,N_18750);
or U19234 (N_19234,N_18943,N_18817);
xor U19235 (N_19235,N_18796,N_18856);
or U19236 (N_19236,N_18845,N_18921);
xnor U19237 (N_19237,N_18981,N_18946);
xnor U19238 (N_19238,N_18870,N_18824);
nand U19239 (N_19239,N_18989,N_18948);
nand U19240 (N_19240,N_18920,N_18760);
nand U19241 (N_19241,N_18788,N_18960);
and U19242 (N_19242,N_18793,N_18870);
xor U19243 (N_19243,N_18800,N_18987);
nand U19244 (N_19244,N_18765,N_18780);
xnor U19245 (N_19245,N_18909,N_18924);
or U19246 (N_19246,N_18950,N_18916);
nor U19247 (N_19247,N_18911,N_18947);
nand U19248 (N_19248,N_18860,N_18890);
nand U19249 (N_19249,N_18960,N_18932);
xor U19250 (N_19250,N_19204,N_19085);
xnor U19251 (N_19251,N_19239,N_19091);
nor U19252 (N_19252,N_19128,N_19212);
xnor U19253 (N_19253,N_19063,N_19077);
or U19254 (N_19254,N_19156,N_19025);
and U19255 (N_19255,N_19233,N_19097);
and U19256 (N_19256,N_19140,N_19051);
or U19257 (N_19257,N_19163,N_19093);
or U19258 (N_19258,N_19169,N_19226);
nor U19259 (N_19259,N_19065,N_19027);
or U19260 (N_19260,N_19146,N_19058);
and U19261 (N_19261,N_19249,N_19104);
and U19262 (N_19262,N_19033,N_19121);
nor U19263 (N_19263,N_19147,N_19072);
xor U19264 (N_19264,N_19073,N_19122);
or U19265 (N_19265,N_19192,N_19167);
and U19266 (N_19266,N_19139,N_19062);
xnor U19267 (N_19267,N_19029,N_19083);
nor U19268 (N_19268,N_19030,N_19057);
nand U19269 (N_19269,N_19217,N_19056);
xor U19270 (N_19270,N_19246,N_19081);
nand U19271 (N_19271,N_19235,N_19069);
nor U19272 (N_19272,N_19215,N_19173);
and U19273 (N_19273,N_19092,N_19106);
and U19274 (N_19274,N_19149,N_19130);
xor U19275 (N_19275,N_19059,N_19195);
or U19276 (N_19276,N_19236,N_19196);
nand U19277 (N_19277,N_19043,N_19135);
nand U19278 (N_19278,N_19018,N_19222);
and U19279 (N_19279,N_19165,N_19209);
nand U19280 (N_19280,N_19011,N_19129);
nand U19281 (N_19281,N_19203,N_19151);
or U19282 (N_19282,N_19199,N_19098);
and U19283 (N_19283,N_19157,N_19002);
or U19284 (N_19284,N_19118,N_19080);
nor U19285 (N_19285,N_19008,N_19017);
nand U19286 (N_19286,N_19112,N_19108);
nor U19287 (N_19287,N_19116,N_19144);
or U19288 (N_19288,N_19187,N_19075);
nand U19289 (N_19289,N_19188,N_19225);
nand U19290 (N_19290,N_19004,N_19031);
and U19291 (N_19291,N_19096,N_19229);
nand U19292 (N_19292,N_19055,N_19170);
nor U19293 (N_19293,N_19078,N_19003);
or U19294 (N_19294,N_19000,N_19207);
or U19295 (N_19295,N_19099,N_19105);
xnor U19296 (N_19296,N_19037,N_19124);
or U19297 (N_19297,N_19119,N_19224);
or U19298 (N_19298,N_19131,N_19016);
or U19299 (N_19299,N_19114,N_19023);
or U19300 (N_19300,N_19164,N_19090);
nand U19301 (N_19301,N_19176,N_19041);
nor U19302 (N_19302,N_19185,N_19039);
nor U19303 (N_19303,N_19134,N_19158);
and U19304 (N_19304,N_19107,N_19198);
xor U19305 (N_19305,N_19221,N_19145);
nand U19306 (N_19306,N_19136,N_19237);
nor U19307 (N_19307,N_19210,N_19049);
and U19308 (N_19308,N_19159,N_19168);
and U19309 (N_19309,N_19101,N_19184);
nor U19310 (N_19310,N_19022,N_19028);
xor U19311 (N_19311,N_19171,N_19174);
xor U19312 (N_19312,N_19143,N_19162);
nor U19313 (N_19313,N_19230,N_19197);
nand U19314 (N_19314,N_19042,N_19227);
or U19315 (N_19315,N_19154,N_19153);
nand U19316 (N_19316,N_19047,N_19040);
and U19317 (N_19317,N_19111,N_19232);
or U19318 (N_19318,N_19206,N_19223);
and U19319 (N_19319,N_19218,N_19208);
nand U19320 (N_19320,N_19006,N_19228);
xnor U19321 (N_19321,N_19240,N_19005);
nor U19322 (N_19322,N_19061,N_19200);
nand U19323 (N_19323,N_19234,N_19150);
nand U19324 (N_19324,N_19180,N_19007);
and U19325 (N_19325,N_19087,N_19179);
nor U19326 (N_19326,N_19046,N_19088);
or U19327 (N_19327,N_19248,N_19067);
and U19328 (N_19328,N_19216,N_19127);
and U19329 (N_19329,N_19183,N_19095);
or U19330 (N_19330,N_19021,N_19054);
or U19331 (N_19331,N_19019,N_19070);
or U19332 (N_19332,N_19202,N_19175);
nor U19333 (N_19333,N_19053,N_19120);
nand U19334 (N_19334,N_19133,N_19194);
nor U19335 (N_19335,N_19242,N_19084);
nand U19336 (N_19336,N_19213,N_19068);
or U19337 (N_19337,N_19238,N_19193);
and U19338 (N_19338,N_19032,N_19102);
nand U19339 (N_19339,N_19132,N_19001);
nor U19340 (N_19340,N_19048,N_19066);
nor U19341 (N_19341,N_19244,N_19214);
or U19342 (N_19342,N_19211,N_19082);
xor U19343 (N_19343,N_19141,N_19178);
and U19344 (N_19344,N_19100,N_19034);
nand U19345 (N_19345,N_19117,N_19020);
or U19346 (N_19346,N_19182,N_19012);
nor U19347 (N_19347,N_19115,N_19137);
and U19348 (N_19348,N_19024,N_19189);
xnor U19349 (N_19349,N_19126,N_19191);
or U19350 (N_19350,N_19086,N_19241);
or U19351 (N_19351,N_19036,N_19245);
or U19352 (N_19352,N_19015,N_19045);
nand U19353 (N_19353,N_19060,N_19071);
or U19354 (N_19354,N_19110,N_19014);
nand U19355 (N_19355,N_19125,N_19220);
nand U19356 (N_19356,N_19201,N_19089);
and U19357 (N_19357,N_19219,N_19205);
and U19358 (N_19358,N_19148,N_19247);
xor U19359 (N_19359,N_19123,N_19177);
xnor U19360 (N_19360,N_19186,N_19160);
and U19361 (N_19361,N_19190,N_19109);
nand U19362 (N_19362,N_19231,N_19152);
and U19363 (N_19363,N_19161,N_19035);
or U19364 (N_19364,N_19103,N_19113);
or U19365 (N_19365,N_19138,N_19010);
or U19366 (N_19366,N_19026,N_19142);
and U19367 (N_19367,N_19044,N_19052);
nor U19368 (N_19368,N_19076,N_19094);
xnor U19369 (N_19369,N_19172,N_19181);
and U19370 (N_19370,N_19155,N_19243);
nand U19371 (N_19371,N_19064,N_19050);
nor U19372 (N_19372,N_19074,N_19166);
and U19373 (N_19373,N_19013,N_19038);
and U19374 (N_19374,N_19009,N_19079);
or U19375 (N_19375,N_19161,N_19112);
nand U19376 (N_19376,N_19158,N_19180);
or U19377 (N_19377,N_19237,N_19028);
nand U19378 (N_19378,N_19110,N_19205);
xor U19379 (N_19379,N_19188,N_19129);
nand U19380 (N_19380,N_19203,N_19163);
nor U19381 (N_19381,N_19185,N_19155);
and U19382 (N_19382,N_19078,N_19025);
xnor U19383 (N_19383,N_19183,N_19066);
nor U19384 (N_19384,N_19183,N_19180);
xor U19385 (N_19385,N_19124,N_19201);
nor U19386 (N_19386,N_19177,N_19140);
nand U19387 (N_19387,N_19172,N_19051);
nor U19388 (N_19388,N_19132,N_19095);
nand U19389 (N_19389,N_19096,N_19017);
or U19390 (N_19390,N_19181,N_19199);
xnor U19391 (N_19391,N_19088,N_19125);
or U19392 (N_19392,N_19171,N_19141);
and U19393 (N_19393,N_19120,N_19248);
nor U19394 (N_19394,N_19085,N_19037);
xnor U19395 (N_19395,N_19120,N_19243);
and U19396 (N_19396,N_19034,N_19098);
or U19397 (N_19397,N_19230,N_19102);
nand U19398 (N_19398,N_19115,N_19034);
and U19399 (N_19399,N_19154,N_19232);
nand U19400 (N_19400,N_19038,N_19164);
nor U19401 (N_19401,N_19205,N_19007);
and U19402 (N_19402,N_19003,N_19144);
xnor U19403 (N_19403,N_19164,N_19074);
nor U19404 (N_19404,N_19111,N_19064);
and U19405 (N_19405,N_19044,N_19158);
xor U19406 (N_19406,N_19133,N_19171);
and U19407 (N_19407,N_19076,N_19203);
nor U19408 (N_19408,N_19222,N_19229);
nor U19409 (N_19409,N_19246,N_19002);
nor U19410 (N_19410,N_19200,N_19002);
and U19411 (N_19411,N_19202,N_19079);
or U19412 (N_19412,N_19048,N_19133);
xnor U19413 (N_19413,N_19214,N_19199);
nor U19414 (N_19414,N_19004,N_19239);
nand U19415 (N_19415,N_19237,N_19211);
and U19416 (N_19416,N_19191,N_19100);
and U19417 (N_19417,N_19052,N_19168);
nand U19418 (N_19418,N_19219,N_19118);
or U19419 (N_19419,N_19024,N_19152);
and U19420 (N_19420,N_19065,N_19101);
and U19421 (N_19421,N_19198,N_19190);
xnor U19422 (N_19422,N_19177,N_19212);
nand U19423 (N_19423,N_19068,N_19095);
nand U19424 (N_19424,N_19210,N_19015);
xor U19425 (N_19425,N_19014,N_19063);
nor U19426 (N_19426,N_19033,N_19145);
nand U19427 (N_19427,N_19202,N_19094);
xnor U19428 (N_19428,N_19191,N_19028);
nand U19429 (N_19429,N_19145,N_19200);
or U19430 (N_19430,N_19191,N_19163);
xor U19431 (N_19431,N_19248,N_19180);
xnor U19432 (N_19432,N_19136,N_19087);
or U19433 (N_19433,N_19026,N_19060);
nor U19434 (N_19434,N_19185,N_19051);
nor U19435 (N_19435,N_19114,N_19059);
or U19436 (N_19436,N_19053,N_19001);
nor U19437 (N_19437,N_19163,N_19066);
nor U19438 (N_19438,N_19045,N_19226);
nand U19439 (N_19439,N_19037,N_19129);
nor U19440 (N_19440,N_19070,N_19104);
nand U19441 (N_19441,N_19010,N_19058);
and U19442 (N_19442,N_19172,N_19048);
or U19443 (N_19443,N_19052,N_19162);
nand U19444 (N_19444,N_19082,N_19200);
xor U19445 (N_19445,N_19162,N_19171);
nor U19446 (N_19446,N_19230,N_19219);
or U19447 (N_19447,N_19190,N_19071);
nand U19448 (N_19448,N_19099,N_19221);
nor U19449 (N_19449,N_19073,N_19217);
and U19450 (N_19450,N_19239,N_19120);
xnor U19451 (N_19451,N_19067,N_19206);
nor U19452 (N_19452,N_19076,N_19011);
or U19453 (N_19453,N_19188,N_19247);
or U19454 (N_19454,N_19201,N_19037);
xor U19455 (N_19455,N_19043,N_19142);
nand U19456 (N_19456,N_19088,N_19200);
or U19457 (N_19457,N_19154,N_19165);
xnor U19458 (N_19458,N_19187,N_19192);
or U19459 (N_19459,N_19187,N_19070);
or U19460 (N_19460,N_19203,N_19124);
xor U19461 (N_19461,N_19103,N_19077);
xnor U19462 (N_19462,N_19213,N_19176);
nor U19463 (N_19463,N_19101,N_19089);
nor U19464 (N_19464,N_19068,N_19097);
or U19465 (N_19465,N_19070,N_19139);
or U19466 (N_19466,N_19176,N_19145);
nand U19467 (N_19467,N_19005,N_19198);
or U19468 (N_19468,N_19113,N_19221);
nand U19469 (N_19469,N_19168,N_19031);
or U19470 (N_19470,N_19003,N_19147);
nand U19471 (N_19471,N_19014,N_19249);
nand U19472 (N_19472,N_19159,N_19237);
nand U19473 (N_19473,N_19149,N_19027);
xnor U19474 (N_19474,N_19167,N_19041);
and U19475 (N_19475,N_19030,N_19018);
and U19476 (N_19476,N_19087,N_19172);
or U19477 (N_19477,N_19164,N_19234);
nand U19478 (N_19478,N_19179,N_19003);
or U19479 (N_19479,N_19108,N_19234);
nor U19480 (N_19480,N_19065,N_19009);
or U19481 (N_19481,N_19238,N_19057);
or U19482 (N_19482,N_19023,N_19080);
nand U19483 (N_19483,N_19070,N_19082);
xor U19484 (N_19484,N_19108,N_19161);
and U19485 (N_19485,N_19110,N_19041);
nor U19486 (N_19486,N_19128,N_19061);
nor U19487 (N_19487,N_19150,N_19018);
or U19488 (N_19488,N_19181,N_19146);
or U19489 (N_19489,N_19125,N_19079);
and U19490 (N_19490,N_19139,N_19016);
or U19491 (N_19491,N_19187,N_19180);
xor U19492 (N_19492,N_19089,N_19097);
and U19493 (N_19493,N_19188,N_19230);
or U19494 (N_19494,N_19110,N_19156);
xor U19495 (N_19495,N_19058,N_19181);
xor U19496 (N_19496,N_19197,N_19068);
nand U19497 (N_19497,N_19248,N_19187);
xor U19498 (N_19498,N_19114,N_19020);
nand U19499 (N_19499,N_19134,N_19039);
nand U19500 (N_19500,N_19447,N_19393);
nand U19501 (N_19501,N_19301,N_19368);
xnor U19502 (N_19502,N_19288,N_19443);
or U19503 (N_19503,N_19431,N_19488);
or U19504 (N_19504,N_19277,N_19337);
nand U19505 (N_19505,N_19265,N_19294);
xor U19506 (N_19506,N_19302,N_19261);
xor U19507 (N_19507,N_19293,N_19339);
nand U19508 (N_19508,N_19309,N_19434);
xor U19509 (N_19509,N_19410,N_19405);
xnor U19510 (N_19510,N_19433,N_19442);
or U19511 (N_19511,N_19499,N_19336);
and U19512 (N_19512,N_19348,N_19358);
or U19513 (N_19513,N_19425,N_19338);
xnor U19514 (N_19514,N_19260,N_19334);
nor U19515 (N_19515,N_19355,N_19283);
nor U19516 (N_19516,N_19392,N_19446);
nand U19517 (N_19517,N_19484,N_19373);
xor U19518 (N_19518,N_19417,N_19490);
or U19519 (N_19519,N_19333,N_19310);
or U19520 (N_19520,N_19426,N_19388);
nand U19521 (N_19521,N_19395,N_19450);
xnor U19522 (N_19522,N_19292,N_19376);
xnor U19523 (N_19523,N_19432,N_19295);
nor U19524 (N_19524,N_19491,N_19315);
nand U19525 (N_19525,N_19360,N_19251);
nand U19526 (N_19526,N_19359,N_19275);
or U19527 (N_19527,N_19390,N_19342);
xor U19528 (N_19528,N_19252,N_19391);
and U19529 (N_19529,N_19280,N_19285);
nor U19530 (N_19530,N_19341,N_19329);
nand U19531 (N_19531,N_19335,N_19418);
nand U19532 (N_19532,N_19435,N_19367);
nor U19533 (N_19533,N_19469,N_19462);
or U19534 (N_19534,N_19445,N_19250);
and U19535 (N_19535,N_19455,N_19382);
nor U19536 (N_19536,N_19386,N_19403);
xnor U19537 (N_19537,N_19350,N_19254);
nand U19538 (N_19538,N_19489,N_19317);
or U19539 (N_19539,N_19492,N_19378);
nor U19540 (N_19540,N_19374,N_19476);
xor U19541 (N_19541,N_19344,N_19316);
or U19542 (N_19542,N_19354,N_19456);
or U19543 (N_19543,N_19286,N_19424);
or U19544 (N_19544,N_19276,N_19467);
nor U19545 (N_19545,N_19311,N_19497);
and U19546 (N_19546,N_19493,N_19379);
xnor U19547 (N_19547,N_19279,N_19304);
nand U19548 (N_19548,N_19300,N_19389);
nand U19549 (N_19549,N_19299,N_19253);
or U19550 (N_19550,N_19298,N_19290);
and U19551 (N_19551,N_19262,N_19330);
nand U19552 (N_19552,N_19287,N_19412);
nor U19553 (N_19553,N_19414,N_19481);
nor U19554 (N_19554,N_19474,N_19364);
nand U19555 (N_19555,N_19256,N_19461);
or U19556 (N_19556,N_19327,N_19346);
and U19557 (N_19557,N_19413,N_19479);
xor U19558 (N_19558,N_19271,N_19406);
nand U19559 (N_19559,N_19255,N_19291);
or U19560 (N_19560,N_19483,N_19257);
and U19561 (N_19561,N_19480,N_19454);
xnor U19562 (N_19562,N_19420,N_19259);
and U19563 (N_19563,N_19486,N_19281);
nor U19564 (N_19564,N_19487,N_19421);
or U19565 (N_19565,N_19284,N_19377);
or U19566 (N_19566,N_19282,N_19363);
or U19567 (N_19567,N_19305,N_19345);
or U19568 (N_19568,N_19466,N_19495);
or U19569 (N_19569,N_19473,N_19464);
nand U19570 (N_19570,N_19258,N_19401);
or U19571 (N_19571,N_19369,N_19452);
nand U19572 (N_19572,N_19325,N_19314);
or U19573 (N_19573,N_19268,N_19384);
or U19574 (N_19574,N_19353,N_19303);
or U19575 (N_19575,N_19270,N_19470);
nor U19576 (N_19576,N_19404,N_19349);
or U19577 (N_19577,N_19396,N_19444);
or U19578 (N_19578,N_19331,N_19460);
nand U19579 (N_19579,N_19320,N_19313);
or U19580 (N_19580,N_19267,N_19263);
nor U19581 (N_19581,N_19326,N_19416);
or U19582 (N_19582,N_19423,N_19428);
or U19583 (N_19583,N_19352,N_19296);
nand U19584 (N_19584,N_19411,N_19289);
nand U19585 (N_19585,N_19278,N_19394);
nand U19586 (N_19586,N_19272,N_19387);
and U19587 (N_19587,N_19318,N_19471);
nand U19588 (N_19588,N_19371,N_19436);
nor U19589 (N_19589,N_19370,N_19306);
nand U19590 (N_19590,N_19472,N_19328);
or U19591 (N_19591,N_19324,N_19266);
nand U19592 (N_19592,N_19312,N_19458);
nor U19593 (N_19593,N_19437,N_19449);
nor U19594 (N_19594,N_19477,N_19332);
xnor U19595 (N_19595,N_19356,N_19430);
and U19596 (N_19596,N_19468,N_19415);
and U19597 (N_19597,N_19494,N_19399);
nand U19598 (N_19598,N_19496,N_19408);
xnor U19599 (N_19599,N_19482,N_19448);
xor U19600 (N_19600,N_19319,N_19429);
xor U19601 (N_19601,N_19343,N_19419);
or U19602 (N_19602,N_19340,N_19365);
and U19603 (N_19603,N_19402,N_19380);
and U19604 (N_19604,N_19465,N_19357);
xnor U19605 (N_19605,N_19273,N_19400);
nand U19606 (N_19606,N_19459,N_19308);
nand U19607 (N_19607,N_19427,N_19385);
nand U19608 (N_19608,N_19397,N_19361);
and U19609 (N_19609,N_19439,N_19269);
nand U19610 (N_19610,N_19475,N_19441);
xor U19611 (N_19611,N_19485,N_19372);
nand U19612 (N_19612,N_19297,N_19322);
and U19613 (N_19613,N_19422,N_19407);
and U19614 (N_19614,N_19478,N_19274);
nor U19615 (N_19615,N_19453,N_19438);
and U19616 (N_19616,N_19457,N_19351);
or U19617 (N_19617,N_19323,N_19307);
xor U19618 (N_19618,N_19398,N_19381);
nor U19619 (N_19619,N_19409,N_19347);
xnor U19620 (N_19620,N_19498,N_19362);
xnor U19621 (N_19621,N_19440,N_19366);
xor U19622 (N_19622,N_19264,N_19321);
nor U19623 (N_19623,N_19375,N_19383);
or U19624 (N_19624,N_19451,N_19463);
or U19625 (N_19625,N_19324,N_19310);
xnor U19626 (N_19626,N_19320,N_19343);
and U19627 (N_19627,N_19364,N_19336);
nor U19628 (N_19628,N_19385,N_19299);
or U19629 (N_19629,N_19482,N_19308);
xor U19630 (N_19630,N_19462,N_19384);
nand U19631 (N_19631,N_19393,N_19252);
or U19632 (N_19632,N_19311,N_19417);
or U19633 (N_19633,N_19358,N_19494);
and U19634 (N_19634,N_19322,N_19397);
or U19635 (N_19635,N_19474,N_19457);
nand U19636 (N_19636,N_19390,N_19460);
and U19637 (N_19637,N_19279,N_19471);
nand U19638 (N_19638,N_19347,N_19449);
nor U19639 (N_19639,N_19343,N_19412);
xor U19640 (N_19640,N_19331,N_19440);
nor U19641 (N_19641,N_19426,N_19292);
nor U19642 (N_19642,N_19445,N_19453);
and U19643 (N_19643,N_19289,N_19313);
or U19644 (N_19644,N_19377,N_19283);
nand U19645 (N_19645,N_19481,N_19463);
nand U19646 (N_19646,N_19268,N_19266);
nand U19647 (N_19647,N_19265,N_19282);
xnor U19648 (N_19648,N_19374,N_19277);
xor U19649 (N_19649,N_19252,N_19301);
nand U19650 (N_19650,N_19427,N_19424);
or U19651 (N_19651,N_19322,N_19398);
xnor U19652 (N_19652,N_19488,N_19341);
and U19653 (N_19653,N_19424,N_19275);
nor U19654 (N_19654,N_19489,N_19331);
and U19655 (N_19655,N_19461,N_19426);
nor U19656 (N_19656,N_19274,N_19324);
and U19657 (N_19657,N_19498,N_19270);
or U19658 (N_19658,N_19444,N_19342);
or U19659 (N_19659,N_19457,N_19399);
nor U19660 (N_19660,N_19300,N_19387);
xnor U19661 (N_19661,N_19452,N_19289);
nand U19662 (N_19662,N_19499,N_19328);
nand U19663 (N_19663,N_19379,N_19350);
nor U19664 (N_19664,N_19304,N_19328);
and U19665 (N_19665,N_19442,N_19331);
nand U19666 (N_19666,N_19443,N_19400);
xnor U19667 (N_19667,N_19285,N_19493);
nand U19668 (N_19668,N_19499,N_19263);
nor U19669 (N_19669,N_19430,N_19470);
and U19670 (N_19670,N_19423,N_19421);
and U19671 (N_19671,N_19363,N_19418);
nor U19672 (N_19672,N_19364,N_19316);
nand U19673 (N_19673,N_19316,N_19410);
and U19674 (N_19674,N_19460,N_19378);
xor U19675 (N_19675,N_19398,N_19383);
xnor U19676 (N_19676,N_19356,N_19378);
nor U19677 (N_19677,N_19270,N_19399);
nand U19678 (N_19678,N_19469,N_19389);
nand U19679 (N_19679,N_19361,N_19472);
or U19680 (N_19680,N_19328,N_19341);
or U19681 (N_19681,N_19303,N_19446);
nor U19682 (N_19682,N_19302,N_19431);
or U19683 (N_19683,N_19372,N_19461);
and U19684 (N_19684,N_19348,N_19451);
or U19685 (N_19685,N_19325,N_19470);
or U19686 (N_19686,N_19398,N_19459);
xor U19687 (N_19687,N_19466,N_19298);
nand U19688 (N_19688,N_19332,N_19315);
nand U19689 (N_19689,N_19345,N_19277);
xor U19690 (N_19690,N_19284,N_19416);
nor U19691 (N_19691,N_19376,N_19405);
and U19692 (N_19692,N_19485,N_19352);
xnor U19693 (N_19693,N_19357,N_19307);
xor U19694 (N_19694,N_19435,N_19490);
xor U19695 (N_19695,N_19404,N_19451);
or U19696 (N_19696,N_19318,N_19262);
or U19697 (N_19697,N_19380,N_19444);
xnor U19698 (N_19698,N_19261,N_19251);
nand U19699 (N_19699,N_19495,N_19398);
nor U19700 (N_19700,N_19375,N_19392);
or U19701 (N_19701,N_19344,N_19427);
nor U19702 (N_19702,N_19339,N_19409);
or U19703 (N_19703,N_19480,N_19431);
nand U19704 (N_19704,N_19352,N_19373);
nor U19705 (N_19705,N_19366,N_19373);
xor U19706 (N_19706,N_19454,N_19443);
xor U19707 (N_19707,N_19379,N_19374);
nand U19708 (N_19708,N_19250,N_19287);
nand U19709 (N_19709,N_19250,N_19403);
or U19710 (N_19710,N_19389,N_19424);
xnor U19711 (N_19711,N_19445,N_19270);
nand U19712 (N_19712,N_19280,N_19270);
or U19713 (N_19713,N_19483,N_19446);
and U19714 (N_19714,N_19492,N_19348);
or U19715 (N_19715,N_19267,N_19383);
nor U19716 (N_19716,N_19250,N_19475);
or U19717 (N_19717,N_19336,N_19432);
xor U19718 (N_19718,N_19270,N_19429);
and U19719 (N_19719,N_19283,N_19416);
or U19720 (N_19720,N_19390,N_19444);
nor U19721 (N_19721,N_19291,N_19288);
or U19722 (N_19722,N_19310,N_19463);
nor U19723 (N_19723,N_19492,N_19439);
nand U19724 (N_19724,N_19387,N_19298);
nand U19725 (N_19725,N_19438,N_19364);
xnor U19726 (N_19726,N_19481,N_19333);
and U19727 (N_19727,N_19266,N_19253);
nand U19728 (N_19728,N_19253,N_19443);
and U19729 (N_19729,N_19375,N_19430);
and U19730 (N_19730,N_19250,N_19441);
and U19731 (N_19731,N_19332,N_19355);
or U19732 (N_19732,N_19355,N_19413);
and U19733 (N_19733,N_19425,N_19297);
or U19734 (N_19734,N_19284,N_19453);
or U19735 (N_19735,N_19276,N_19487);
nor U19736 (N_19736,N_19477,N_19434);
xor U19737 (N_19737,N_19298,N_19305);
and U19738 (N_19738,N_19309,N_19319);
or U19739 (N_19739,N_19367,N_19318);
xnor U19740 (N_19740,N_19364,N_19403);
nand U19741 (N_19741,N_19472,N_19451);
xnor U19742 (N_19742,N_19479,N_19437);
or U19743 (N_19743,N_19306,N_19331);
nor U19744 (N_19744,N_19453,N_19398);
xnor U19745 (N_19745,N_19283,N_19292);
and U19746 (N_19746,N_19492,N_19446);
nand U19747 (N_19747,N_19499,N_19479);
nand U19748 (N_19748,N_19371,N_19393);
xnor U19749 (N_19749,N_19392,N_19434);
xor U19750 (N_19750,N_19591,N_19742);
and U19751 (N_19751,N_19656,N_19532);
nand U19752 (N_19752,N_19579,N_19657);
nor U19753 (N_19753,N_19562,N_19640);
xor U19754 (N_19754,N_19634,N_19523);
or U19755 (N_19755,N_19552,N_19658);
or U19756 (N_19756,N_19527,N_19625);
xor U19757 (N_19757,N_19568,N_19633);
or U19758 (N_19758,N_19596,N_19593);
and U19759 (N_19759,N_19585,N_19538);
xor U19760 (N_19760,N_19639,N_19668);
xor U19761 (N_19761,N_19711,N_19533);
xnor U19762 (N_19762,N_19748,N_19644);
nand U19763 (N_19763,N_19715,N_19655);
nand U19764 (N_19764,N_19580,N_19602);
nand U19765 (N_19765,N_19537,N_19745);
and U19766 (N_19766,N_19652,N_19605);
or U19767 (N_19767,N_19623,N_19674);
nor U19768 (N_19768,N_19528,N_19685);
and U19769 (N_19769,N_19660,N_19524);
and U19770 (N_19770,N_19555,N_19522);
nor U19771 (N_19771,N_19693,N_19735);
nor U19772 (N_19772,N_19720,N_19502);
nor U19773 (N_19773,N_19675,N_19719);
and U19774 (N_19774,N_19646,N_19567);
and U19775 (N_19775,N_19628,N_19520);
or U19776 (N_19776,N_19511,N_19558);
nor U19777 (N_19777,N_19615,N_19738);
nand U19778 (N_19778,N_19647,N_19728);
nor U19779 (N_19779,N_19603,N_19565);
xor U19780 (N_19780,N_19598,N_19687);
or U19781 (N_19781,N_19515,N_19561);
nor U19782 (N_19782,N_19667,N_19546);
xnor U19783 (N_19783,N_19671,N_19648);
and U19784 (N_19784,N_19590,N_19686);
nand U19785 (N_19785,N_19730,N_19588);
and U19786 (N_19786,N_19582,N_19570);
nor U19787 (N_19787,N_19717,N_19526);
xnor U19788 (N_19788,N_19747,N_19684);
nor U19789 (N_19789,N_19698,N_19697);
xnor U19790 (N_19790,N_19610,N_19581);
nor U19791 (N_19791,N_19514,N_19606);
nand U19792 (N_19792,N_19741,N_19551);
or U19793 (N_19793,N_19519,N_19732);
or U19794 (N_19794,N_19553,N_19702);
and U19795 (N_19795,N_19535,N_19680);
xnor U19796 (N_19796,N_19575,N_19716);
xnor U19797 (N_19797,N_19682,N_19681);
or U19798 (N_19798,N_19649,N_19584);
xnor U19799 (N_19799,N_19540,N_19700);
nor U19800 (N_19800,N_19589,N_19729);
and U19801 (N_19801,N_19577,N_19677);
or U19802 (N_19802,N_19616,N_19501);
and U19803 (N_19803,N_19594,N_19612);
nor U19804 (N_19804,N_19572,N_19614);
nor U19805 (N_19805,N_19542,N_19642);
xnor U19806 (N_19806,N_19661,N_19638);
xor U19807 (N_19807,N_19713,N_19544);
and U19808 (N_19808,N_19506,N_19683);
nand U19809 (N_19809,N_19613,N_19564);
and U19810 (N_19810,N_19726,N_19550);
nor U19811 (N_19811,N_19529,N_19679);
xnor U19812 (N_19812,N_19556,N_19691);
or U19813 (N_19813,N_19643,N_19508);
or U19814 (N_19814,N_19721,N_19695);
xor U19815 (N_19815,N_19694,N_19641);
or U19816 (N_19816,N_19517,N_19688);
nand U19817 (N_19817,N_19731,N_19611);
or U19818 (N_19818,N_19626,N_19712);
xnor U19819 (N_19819,N_19513,N_19505);
and U19820 (N_19820,N_19601,N_19531);
nand U19821 (N_19821,N_19653,N_19663);
xor U19822 (N_19822,N_19736,N_19709);
xor U19823 (N_19823,N_19664,N_19743);
nand U19824 (N_19824,N_19586,N_19666);
and U19825 (N_19825,N_19510,N_19737);
or U19826 (N_19826,N_19587,N_19650);
nor U19827 (N_19827,N_19718,N_19722);
nor U19828 (N_19828,N_19662,N_19500);
or U19829 (N_19829,N_19704,N_19618);
and U19830 (N_19830,N_19701,N_19706);
nand U19831 (N_19831,N_19690,N_19576);
or U19832 (N_19832,N_19543,N_19609);
and U19833 (N_19833,N_19516,N_19504);
nand U19834 (N_19834,N_19563,N_19723);
or U19835 (N_19835,N_19699,N_19600);
and U19836 (N_19836,N_19678,N_19632);
nor U19837 (N_19837,N_19503,N_19707);
and U19838 (N_19838,N_19733,N_19740);
nor U19839 (N_19839,N_19659,N_19607);
nor U19840 (N_19840,N_19714,N_19620);
xnor U19841 (N_19841,N_19554,N_19608);
or U19842 (N_19842,N_19566,N_19569);
xnor U19843 (N_19843,N_19597,N_19617);
xor U19844 (N_19844,N_19622,N_19676);
and U19845 (N_19845,N_19705,N_19692);
or U19846 (N_19846,N_19549,N_19595);
nand U19847 (N_19847,N_19548,N_19530);
xnor U19848 (N_19848,N_19725,N_19673);
nor U19849 (N_19849,N_19512,N_19749);
xor U19850 (N_19850,N_19509,N_19574);
nand U19851 (N_19851,N_19604,N_19637);
nor U19852 (N_19852,N_19631,N_19536);
and U19853 (N_19853,N_19696,N_19592);
and U19854 (N_19854,N_19539,N_19645);
and U19855 (N_19855,N_19734,N_19619);
nor U19856 (N_19856,N_19651,N_19571);
and U19857 (N_19857,N_19557,N_19703);
and U19858 (N_19858,N_19525,N_19583);
or U19859 (N_19859,N_19727,N_19665);
and U19860 (N_19860,N_19599,N_19627);
nor U19861 (N_19861,N_19672,N_19669);
xnor U19862 (N_19862,N_19739,N_19573);
xor U19863 (N_19863,N_19724,N_19559);
nor U19864 (N_19864,N_19630,N_19710);
xnor U19865 (N_19865,N_19621,N_19746);
or U19866 (N_19866,N_19578,N_19744);
and U19867 (N_19867,N_19708,N_19545);
xnor U19868 (N_19868,N_19507,N_19547);
xnor U19869 (N_19869,N_19689,N_19635);
and U19870 (N_19870,N_19629,N_19636);
nand U19871 (N_19871,N_19521,N_19560);
xor U19872 (N_19872,N_19624,N_19518);
and U19873 (N_19873,N_19534,N_19654);
or U19874 (N_19874,N_19670,N_19541);
nor U19875 (N_19875,N_19502,N_19715);
nor U19876 (N_19876,N_19614,N_19637);
or U19877 (N_19877,N_19664,N_19688);
nand U19878 (N_19878,N_19555,N_19737);
nand U19879 (N_19879,N_19665,N_19645);
and U19880 (N_19880,N_19648,N_19692);
and U19881 (N_19881,N_19714,N_19664);
nand U19882 (N_19882,N_19696,N_19715);
nand U19883 (N_19883,N_19506,N_19619);
and U19884 (N_19884,N_19632,N_19640);
or U19885 (N_19885,N_19665,N_19556);
or U19886 (N_19886,N_19591,N_19650);
or U19887 (N_19887,N_19562,N_19536);
or U19888 (N_19888,N_19620,N_19670);
or U19889 (N_19889,N_19558,N_19591);
and U19890 (N_19890,N_19585,N_19524);
nand U19891 (N_19891,N_19705,N_19686);
or U19892 (N_19892,N_19503,N_19705);
nor U19893 (N_19893,N_19690,N_19679);
xor U19894 (N_19894,N_19623,N_19718);
or U19895 (N_19895,N_19579,N_19724);
xor U19896 (N_19896,N_19657,N_19549);
xnor U19897 (N_19897,N_19662,N_19627);
nor U19898 (N_19898,N_19653,N_19636);
nand U19899 (N_19899,N_19692,N_19592);
nor U19900 (N_19900,N_19746,N_19505);
and U19901 (N_19901,N_19707,N_19530);
nand U19902 (N_19902,N_19534,N_19726);
nand U19903 (N_19903,N_19593,N_19620);
nor U19904 (N_19904,N_19570,N_19548);
nand U19905 (N_19905,N_19734,N_19531);
nand U19906 (N_19906,N_19694,N_19564);
nor U19907 (N_19907,N_19629,N_19716);
and U19908 (N_19908,N_19559,N_19699);
nor U19909 (N_19909,N_19542,N_19728);
or U19910 (N_19910,N_19642,N_19603);
and U19911 (N_19911,N_19588,N_19748);
nor U19912 (N_19912,N_19731,N_19730);
or U19913 (N_19913,N_19592,N_19504);
or U19914 (N_19914,N_19523,N_19516);
nor U19915 (N_19915,N_19594,N_19511);
and U19916 (N_19916,N_19702,N_19700);
and U19917 (N_19917,N_19643,N_19533);
nor U19918 (N_19918,N_19561,N_19744);
or U19919 (N_19919,N_19640,N_19512);
nor U19920 (N_19920,N_19712,N_19703);
nand U19921 (N_19921,N_19619,N_19626);
nor U19922 (N_19922,N_19740,N_19657);
nand U19923 (N_19923,N_19564,N_19532);
and U19924 (N_19924,N_19552,N_19649);
nand U19925 (N_19925,N_19699,N_19605);
and U19926 (N_19926,N_19579,N_19509);
nor U19927 (N_19927,N_19619,N_19589);
and U19928 (N_19928,N_19567,N_19591);
or U19929 (N_19929,N_19730,N_19542);
nor U19930 (N_19930,N_19607,N_19510);
and U19931 (N_19931,N_19689,N_19734);
or U19932 (N_19932,N_19506,N_19640);
and U19933 (N_19933,N_19671,N_19739);
and U19934 (N_19934,N_19541,N_19608);
nor U19935 (N_19935,N_19540,N_19708);
and U19936 (N_19936,N_19585,N_19505);
xnor U19937 (N_19937,N_19746,N_19587);
or U19938 (N_19938,N_19588,N_19708);
and U19939 (N_19939,N_19656,N_19705);
xor U19940 (N_19940,N_19738,N_19630);
or U19941 (N_19941,N_19520,N_19745);
nor U19942 (N_19942,N_19691,N_19569);
nand U19943 (N_19943,N_19575,N_19605);
nand U19944 (N_19944,N_19526,N_19537);
nor U19945 (N_19945,N_19547,N_19515);
nor U19946 (N_19946,N_19665,N_19634);
or U19947 (N_19947,N_19622,N_19698);
nand U19948 (N_19948,N_19692,N_19633);
nand U19949 (N_19949,N_19520,N_19728);
and U19950 (N_19950,N_19657,N_19518);
or U19951 (N_19951,N_19742,N_19710);
and U19952 (N_19952,N_19531,N_19663);
or U19953 (N_19953,N_19678,N_19744);
and U19954 (N_19954,N_19658,N_19581);
xnor U19955 (N_19955,N_19745,N_19589);
nor U19956 (N_19956,N_19519,N_19653);
nand U19957 (N_19957,N_19708,N_19641);
and U19958 (N_19958,N_19645,N_19669);
or U19959 (N_19959,N_19637,N_19732);
or U19960 (N_19960,N_19625,N_19656);
nor U19961 (N_19961,N_19568,N_19508);
and U19962 (N_19962,N_19571,N_19556);
nand U19963 (N_19963,N_19648,N_19520);
and U19964 (N_19964,N_19518,N_19741);
nand U19965 (N_19965,N_19640,N_19518);
nor U19966 (N_19966,N_19641,N_19583);
and U19967 (N_19967,N_19587,N_19531);
or U19968 (N_19968,N_19655,N_19559);
xnor U19969 (N_19969,N_19730,N_19650);
or U19970 (N_19970,N_19652,N_19651);
and U19971 (N_19971,N_19656,N_19677);
and U19972 (N_19972,N_19664,N_19518);
and U19973 (N_19973,N_19643,N_19579);
nor U19974 (N_19974,N_19708,N_19519);
and U19975 (N_19975,N_19519,N_19557);
nor U19976 (N_19976,N_19573,N_19696);
nor U19977 (N_19977,N_19747,N_19717);
or U19978 (N_19978,N_19619,N_19637);
or U19979 (N_19979,N_19543,N_19534);
nand U19980 (N_19980,N_19512,N_19634);
nor U19981 (N_19981,N_19701,N_19605);
nand U19982 (N_19982,N_19607,N_19705);
and U19983 (N_19983,N_19742,N_19575);
xor U19984 (N_19984,N_19591,N_19634);
and U19985 (N_19985,N_19704,N_19747);
and U19986 (N_19986,N_19733,N_19703);
nor U19987 (N_19987,N_19699,N_19731);
and U19988 (N_19988,N_19746,N_19663);
or U19989 (N_19989,N_19647,N_19651);
nor U19990 (N_19990,N_19665,N_19738);
nand U19991 (N_19991,N_19541,N_19556);
nor U19992 (N_19992,N_19733,N_19618);
nand U19993 (N_19993,N_19547,N_19693);
nand U19994 (N_19994,N_19671,N_19614);
or U19995 (N_19995,N_19715,N_19620);
nor U19996 (N_19996,N_19692,N_19738);
nand U19997 (N_19997,N_19502,N_19558);
or U19998 (N_19998,N_19719,N_19637);
xor U19999 (N_19999,N_19725,N_19592);
nand UO_0 (O_0,N_19922,N_19973);
nor UO_1 (O_1,N_19985,N_19909);
xor UO_2 (O_2,N_19960,N_19787);
or UO_3 (O_3,N_19886,N_19987);
nor UO_4 (O_4,N_19945,N_19926);
nand UO_5 (O_5,N_19750,N_19829);
or UO_6 (O_6,N_19967,N_19870);
nor UO_7 (O_7,N_19887,N_19836);
and UO_8 (O_8,N_19760,N_19785);
and UO_9 (O_9,N_19939,N_19768);
nand UO_10 (O_10,N_19869,N_19981);
and UO_11 (O_11,N_19952,N_19881);
nand UO_12 (O_12,N_19825,N_19810);
xor UO_13 (O_13,N_19853,N_19899);
xnor UO_14 (O_14,N_19898,N_19989);
xnor UO_15 (O_15,N_19924,N_19790);
or UO_16 (O_16,N_19902,N_19934);
nor UO_17 (O_17,N_19997,N_19873);
nor UO_18 (O_18,N_19995,N_19859);
xnor UO_19 (O_19,N_19980,N_19978);
xor UO_20 (O_20,N_19867,N_19818);
and UO_21 (O_21,N_19916,N_19851);
nand UO_22 (O_22,N_19868,N_19937);
and UO_23 (O_23,N_19765,N_19771);
xor UO_24 (O_24,N_19796,N_19969);
nor UO_25 (O_25,N_19932,N_19863);
nor UO_26 (O_26,N_19862,N_19848);
or UO_27 (O_27,N_19882,N_19976);
nor UO_28 (O_28,N_19963,N_19806);
or UO_29 (O_29,N_19782,N_19849);
and UO_30 (O_30,N_19817,N_19752);
xnor UO_31 (O_31,N_19766,N_19884);
nand UO_32 (O_32,N_19778,N_19865);
nand UO_33 (O_33,N_19991,N_19993);
or UO_34 (O_34,N_19927,N_19895);
nor UO_35 (O_35,N_19828,N_19809);
and UO_36 (O_36,N_19928,N_19835);
or UO_37 (O_37,N_19858,N_19918);
and UO_38 (O_38,N_19875,N_19802);
nand UO_39 (O_39,N_19794,N_19821);
nand UO_40 (O_40,N_19994,N_19948);
xnor UO_41 (O_41,N_19938,N_19880);
nor UO_42 (O_42,N_19779,N_19826);
nand UO_43 (O_43,N_19972,N_19775);
and UO_44 (O_44,N_19944,N_19955);
nand UO_45 (O_45,N_19906,N_19761);
and UO_46 (O_46,N_19846,N_19824);
xor UO_47 (O_47,N_19834,N_19767);
and UO_48 (O_48,N_19893,N_19908);
or UO_49 (O_49,N_19954,N_19946);
nand UO_50 (O_50,N_19907,N_19891);
nor UO_51 (O_51,N_19781,N_19959);
and UO_52 (O_52,N_19819,N_19943);
nand UO_53 (O_53,N_19979,N_19757);
nand UO_54 (O_54,N_19996,N_19795);
and UO_55 (O_55,N_19990,N_19776);
and UO_56 (O_56,N_19904,N_19970);
xnor UO_57 (O_57,N_19805,N_19983);
nand UO_58 (O_58,N_19772,N_19803);
nor UO_59 (O_59,N_19892,N_19897);
nand UO_60 (O_60,N_19827,N_19951);
xor UO_61 (O_61,N_19888,N_19911);
nand UO_62 (O_62,N_19903,N_19956);
nor UO_63 (O_63,N_19832,N_19874);
and UO_64 (O_64,N_19855,N_19759);
nand UO_65 (O_65,N_19808,N_19929);
xor UO_66 (O_66,N_19798,N_19807);
xnor UO_67 (O_67,N_19962,N_19811);
nand UO_68 (O_68,N_19949,N_19812);
nor UO_69 (O_69,N_19947,N_19964);
nor UO_70 (O_70,N_19936,N_19879);
and UO_71 (O_71,N_19861,N_19921);
or UO_72 (O_72,N_19910,N_19751);
nand UO_73 (O_73,N_19942,N_19982);
or UO_74 (O_74,N_19999,N_19844);
and UO_75 (O_75,N_19974,N_19913);
xnor UO_76 (O_76,N_19815,N_19877);
or UO_77 (O_77,N_19901,N_19860);
and UO_78 (O_78,N_19753,N_19847);
nor UO_79 (O_79,N_19833,N_19770);
nand UO_80 (O_80,N_19842,N_19883);
and UO_81 (O_81,N_19793,N_19769);
nor UO_82 (O_82,N_19998,N_19852);
nor UO_83 (O_83,N_19965,N_19839);
nor UO_84 (O_84,N_19977,N_19801);
nand UO_85 (O_85,N_19923,N_19762);
and UO_86 (O_86,N_19838,N_19777);
and UO_87 (O_87,N_19864,N_19890);
or UO_88 (O_88,N_19961,N_19837);
nand UO_89 (O_89,N_19784,N_19786);
or UO_90 (O_90,N_19933,N_19984);
nand UO_91 (O_91,N_19764,N_19788);
nor UO_92 (O_92,N_19935,N_19845);
xnor UO_93 (O_93,N_19917,N_19968);
xnor UO_94 (O_94,N_19878,N_19774);
or UO_95 (O_95,N_19866,N_19988);
or UO_96 (O_96,N_19941,N_19905);
nand UO_97 (O_97,N_19780,N_19919);
nor UO_98 (O_98,N_19843,N_19814);
nand UO_99 (O_99,N_19914,N_19797);
or UO_100 (O_100,N_19958,N_19915);
or UO_101 (O_101,N_19763,N_19966);
nor UO_102 (O_102,N_19940,N_19800);
or UO_103 (O_103,N_19854,N_19975);
or UO_104 (O_104,N_19871,N_19841);
xnor UO_105 (O_105,N_19900,N_19889);
and UO_106 (O_106,N_19754,N_19756);
nor UO_107 (O_107,N_19804,N_19813);
and UO_108 (O_108,N_19816,N_19755);
xor UO_109 (O_109,N_19992,N_19791);
and UO_110 (O_110,N_19799,N_19820);
and UO_111 (O_111,N_19953,N_19792);
nand UO_112 (O_112,N_19840,N_19758);
nor UO_113 (O_113,N_19789,N_19822);
or UO_114 (O_114,N_19850,N_19823);
nor UO_115 (O_115,N_19872,N_19896);
or UO_116 (O_116,N_19931,N_19856);
and UO_117 (O_117,N_19957,N_19876);
and UO_118 (O_118,N_19950,N_19773);
nor UO_119 (O_119,N_19912,N_19857);
xor UO_120 (O_120,N_19783,N_19830);
or UO_121 (O_121,N_19986,N_19971);
xor UO_122 (O_122,N_19925,N_19894);
or UO_123 (O_123,N_19885,N_19930);
and UO_124 (O_124,N_19831,N_19920);
xor UO_125 (O_125,N_19986,N_19942);
nand UO_126 (O_126,N_19789,N_19829);
nand UO_127 (O_127,N_19936,N_19812);
or UO_128 (O_128,N_19967,N_19797);
or UO_129 (O_129,N_19836,N_19970);
nand UO_130 (O_130,N_19960,N_19773);
xor UO_131 (O_131,N_19842,N_19803);
xor UO_132 (O_132,N_19829,N_19889);
or UO_133 (O_133,N_19885,N_19843);
nor UO_134 (O_134,N_19784,N_19940);
xor UO_135 (O_135,N_19985,N_19764);
nor UO_136 (O_136,N_19958,N_19788);
or UO_137 (O_137,N_19789,N_19867);
or UO_138 (O_138,N_19925,N_19963);
and UO_139 (O_139,N_19883,N_19759);
nand UO_140 (O_140,N_19905,N_19862);
and UO_141 (O_141,N_19979,N_19798);
nor UO_142 (O_142,N_19929,N_19852);
and UO_143 (O_143,N_19951,N_19883);
nor UO_144 (O_144,N_19848,N_19884);
or UO_145 (O_145,N_19929,N_19807);
xor UO_146 (O_146,N_19790,N_19837);
nand UO_147 (O_147,N_19914,N_19989);
xnor UO_148 (O_148,N_19940,N_19760);
or UO_149 (O_149,N_19971,N_19804);
xor UO_150 (O_150,N_19995,N_19757);
or UO_151 (O_151,N_19799,N_19796);
nor UO_152 (O_152,N_19868,N_19872);
nor UO_153 (O_153,N_19820,N_19898);
nor UO_154 (O_154,N_19758,N_19787);
and UO_155 (O_155,N_19771,N_19913);
nand UO_156 (O_156,N_19933,N_19946);
nor UO_157 (O_157,N_19780,N_19930);
nand UO_158 (O_158,N_19931,N_19804);
or UO_159 (O_159,N_19848,N_19854);
and UO_160 (O_160,N_19823,N_19994);
and UO_161 (O_161,N_19932,N_19938);
nor UO_162 (O_162,N_19897,N_19769);
nor UO_163 (O_163,N_19787,N_19962);
or UO_164 (O_164,N_19967,N_19928);
xnor UO_165 (O_165,N_19944,N_19952);
nor UO_166 (O_166,N_19948,N_19935);
nor UO_167 (O_167,N_19826,N_19882);
or UO_168 (O_168,N_19788,N_19780);
nand UO_169 (O_169,N_19951,N_19874);
xor UO_170 (O_170,N_19906,N_19921);
and UO_171 (O_171,N_19860,N_19790);
nor UO_172 (O_172,N_19985,N_19961);
nor UO_173 (O_173,N_19907,N_19877);
nor UO_174 (O_174,N_19879,N_19763);
nand UO_175 (O_175,N_19758,N_19776);
nand UO_176 (O_176,N_19790,N_19980);
xnor UO_177 (O_177,N_19899,N_19863);
or UO_178 (O_178,N_19859,N_19993);
nand UO_179 (O_179,N_19752,N_19820);
nand UO_180 (O_180,N_19756,N_19970);
and UO_181 (O_181,N_19934,N_19933);
and UO_182 (O_182,N_19780,N_19820);
or UO_183 (O_183,N_19901,N_19759);
and UO_184 (O_184,N_19830,N_19839);
nor UO_185 (O_185,N_19962,N_19987);
nand UO_186 (O_186,N_19899,N_19848);
or UO_187 (O_187,N_19877,N_19892);
nor UO_188 (O_188,N_19904,N_19787);
xnor UO_189 (O_189,N_19865,N_19962);
xor UO_190 (O_190,N_19927,N_19841);
nor UO_191 (O_191,N_19825,N_19765);
or UO_192 (O_192,N_19898,N_19831);
or UO_193 (O_193,N_19884,N_19893);
nor UO_194 (O_194,N_19772,N_19827);
or UO_195 (O_195,N_19898,N_19841);
and UO_196 (O_196,N_19895,N_19779);
nand UO_197 (O_197,N_19966,N_19832);
nand UO_198 (O_198,N_19975,N_19836);
or UO_199 (O_199,N_19752,N_19809);
nand UO_200 (O_200,N_19918,N_19903);
and UO_201 (O_201,N_19883,N_19853);
nand UO_202 (O_202,N_19952,N_19911);
and UO_203 (O_203,N_19826,N_19816);
nand UO_204 (O_204,N_19769,N_19950);
and UO_205 (O_205,N_19981,N_19923);
and UO_206 (O_206,N_19931,N_19932);
and UO_207 (O_207,N_19837,N_19817);
and UO_208 (O_208,N_19879,N_19949);
and UO_209 (O_209,N_19809,N_19958);
nand UO_210 (O_210,N_19976,N_19779);
nand UO_211 (O_211,N_19799,N_19986);
nor UO_212 (O_212,N_19773,N_19945);
and UO_213 (O_213,N_19772,N_19974);
nor UO_214 (O_214,N_19805,N_19840);
nand UO_215 (O_215,N_19767,N_19755);
nor UO_216 (O_216,N_19915,N_19836);
nor UO_217 (O_217,N_19915,N_19752);
xor UO_218 (O_218,N_19876,N_19947);
xnor UO_219 (O_219,N_19835,N_19804);
xnor UO_220 (O_220,N_19848,N_19913);
nor UO_221 (O_221,N_19753,N_19757);
nand UO_222 (O_222,N_19987,N_19815);
or UO_223 (O_223,N_19877,N_19848);
xor UO_224 (O_224,N_19878,N_19826);
nor UO_225 (O_225,N_19935,N_19870);
and UO_226 (O_226,N_19752,N_19891);
or UO_227 (O_227,N_19998,N_19993);
or UO_228 (O_228,N_19902,N_19858);
nand UO_229 (O_229,N_19952,N_19810);
nor UO_230 (O_230,N_19903,N_19848);
nand UO_231 (O_231,N_19893,N_19824);
and UO_232 (O_232,N_19969,N_19890);
xnor UO_233 (O_233,N_19993,N_19866);
nor UO_234 (O_234,N_19780,N_19827);
nand UO_235 (O_235,N_19978,N_19984);
xor UO_236 (O_236,N_19972,N_19793);
nor UO_237 (O_237,N_19860,N_19826);
nand UO_238 (O_238,N_19994,N_19763);
or UO_239 (O_239,N_19914,N_19761);
and UO_240 (O_240,N_19894,N_19868);
nor UO_241 (O_241,N_19763,N_19987);
and UO_242 (O_242,N_19807,N_19992);
nor UO_243 (O_243,N_19933,N_19771);
nand UO_244 (O_244,N_19862,N_19873);
and UO_245 (O_245,N_19756,N_19888);
nor UO_246 (O_246,N_19815,N_19871);
nand UO_247 (O_247,N_19840,N_19752);
nor UO_248 (O_248,N_19788,N_19997);
or UO_249 (O_249,N_19981,N_19952);
nand UO_250 (O_250,N_19852,N_19985);
nand UO_251 (O_251,N_19957,N_19974);
or UO_252 (O_252,N_19756,N_19764);
nor UO_253 (O_253,N_19864,N_19880);
and UO_254 (O_254,N_19869,N_19847);
xor UO_255 (O_255,N_19780,N_19834);
nand UO_256 (O_256,N_19844,N_19839);
xor UO_257 (O_257,N_19876,N_19788);
nor UO_258 (O_258,N_19778,N_19976);
nand UO_259 (O_259,N_19777,N_19906);
and UO_260 (O_260,N_19818,N_19771);
xnor UO_261 (O_261,N_19827,N_19777);
nor UO_262 (O_262,N_19900,N_19838);
and UO_263 (O_263,N_19960,N_19929);
and UO_264 (O_264,N_19759,N_19811);
nor UO_265 (O_265,N_19807,N_19752);
xnor UO_266 (O_266,N_19894,N_19952);
xor UO_267 (O_267,N_19933,N_19770);
xor UO_268 (O_268,N_19964,N_19817);
nand UO_269 (O_269,N_19878,N_19819);
nand UO_270 (O_270,N_19945,N_19985);
xor UO_271 (O_271,N_19767,N_19842);
xor UO_272 (O_272,N_19778,N_19935);
nand UO_273 (O_273,N_19927,N_19962);
nor UO_274 (O_274,N_19772,N_19832);
or UO_275 (O_275,N_19963,N_19814);
nor UO_276 (O_276,N_19758,N_19838);
nor UO_277 (O_277,N_19835,N_19943);
and UO_278 (O_278,N_19876,N_19985);
and UO_279 (O_279,N_19822,N_19834);
nand UO_280 (O_280,N_19956,N_19868);
nor UO_281 (O_281,N_19916,N_19772);
and UO_282 (O_282,N_19794,N_19990);
and UO_283 (O_283,N_19894,N_19962);
and UO_284 (O_284,N_19794,N_19882);
xnor UO_285 (O_285,N_19887,N_19893);
nand UO_286 (O_286,N_19762,N_19906);
nand UO_287 (O_287,N_19845,N_19823);
or UO_288 (O_288,N_19951,N_19982);
or UO_289 (O_289,N_19931,N_19781);
or UO_290 (O_290,N_19968,N_19803);
or UO_291 (O_291,N_19841,N_19981);
and UO_292 (O_292,N_19905,N_19978);
or UO_293 (O_293,N_19978,N_19947);
xor UO_294 (O_294,N_19898,N_19855);
or UO_295 (O_295,N_19804,N_19975);
nor UO_296 (O_296,N_19841,N_19917);
or UO_297 (O_297,N_19889,N_19801);
nand UO_298 (O_298,N_19852,N_19815);
and UO_299 (O_299,N_19943,N_19895);
or UO_300 (O_300,N_19888,N_19837);
nand UO_301 (O_301,N_19904,N_19879);
and UO_302 (O_302,N_19897,N_19760);
nand UO_303 (O_303,N_19769,N_19923);
nor UO_304 (O_304,N_19998,N_19896);
nor UO_305 (O_305,N_19838,N_19875);
xor UO_306 (O_306,N_19795,N_19973);
and UO_307 (O_307,N_19767,N_19817);
xor UO_308 (O_308,N_19854,N_19947);
and UO_309 (O_309,N_19987,N_19806);
xnor UO_310 (O_310,N_19894,N_19775);
nor UO_311 (O_311,N_19967,N_19907);
nor UO_312 (O_312,N_19900,N_19924);
nand UO_313 (O_313,N_19993,N_19792);
xnor UO_314 (O_314,N_19823,N_19920);
xnor UO_315 (O_315,N_19851,N_19881);
or UO_316 (O_316,N_19966,N_19810);
nor UO_317 (O_317,N_19789,N_19941);
nand UO_318 (O_318,N_19799,N_19928);
nor UO_319 (O_319,N_19753,N_19832);
xor UO_320 (O_320,N_19777,N_19946);
nand UO_321 (O_321,N_19824,N_19946);
and UO_322 (O_322,N_19771,N_19904);
or UO_323 (O_323,N_19770,N_19854);
nand UO_324 (O_324,N_19930,N_19771);
and UO_325 (O_325,N_19861,N_19953);
and UO_326 (O_326,N_19954,N_19924);
nand UO_327 (O_327,N_19764,N_19894);
and UO_328 (O_328,N_19977,N_19892);
nand UO_329 (O_329,N_19809,N_19967);
nand UO_330 (O_330,N_19975,N_19893);
nand UO_331 (O_331,N_19828,N_19852);
nand UO_332 (O_332,N_19956,N_19776);
or UO_333 (O_333,N_19887,N_19968);
nor UO_334 (O_334,N_19904,N_19936);
xor UO_335 (O_335,N_19911,N_19949);
nand UO_336 (O_336,N_19821,N_19895);
or UO_337 (O_337,N_19821,N_19943);
nor UO_338 (O_338,N_19930,N_19770);
and UO_339 (O_339,N_19877,N_19768);
nand UO_340 (O_340,N_19868,N_19890);
xnor UO_341 (O_341,N_19859,N_19982);
xnor UO_342 (O_342,N_19856,N_19764);
nor UO_343 (O_343,N_19803,N_19850);
xnor UO_344 (O_344,N_19855,N_19893);
xnor UO_345 (O_345,N_19893,N_19821);
and UO_346 (O_346,N_19830,N_19782);
nand UO_347 (O_347,N_19885,N_19868);
or UO_348 (O_348,N_19817,N_19810);
xnor UO_349 (O_349,N_19922,N_19964);
and UO_350 (O_350,N_19928,N_19929);
or UO_351 (O_351,N_19973,N_19813);
nor UO_352 (O_352,N_19880,N_19921);
or UO_353 (O_353,N_19846,N_19803);
xnor UO_354 (O_354,N_19971,N_19949);
or UO_355 (O_355,N_19858,N_19876);
and UO_356 (O_356,N_19861,N_19922);
and UO_357 (O_357,N_19822,N_19949);
and UO_358 (O_358,N_19900,N_19987);
nor UO_359 (O_359,N_19766,N_19997);
or UO_360 (O_360,N_19887,N_19961);
and UO_361 (O_361,N_19848,N_19963);
nand UO_362 (O_362,N_19889,N_19860);
or UO_363 (O_363,N_19900,N_19858);
and UO_364 (O_364,N_19912,N_19811);
nor UO_365 (O_365,N_19983,N_19799);
and UO_366 (O_366,N_19915,N_19960);
xor UO_367 (O_367,N_19754,N_19995);
nor UO_368 (O_368,N_19929,N_19878);
or UO_369 (O_369,N_19823,N_19832);
and UO_370 (O_370,N_19775,N_19909);
and UO_371 (O_371,N_19970,N_19945);
or UO_372 (O_372,N_19804,N_19809);
xnor UO_373 (O_373,N_19825,N_19783);
nand UO_374 (O_374,N_19806,N_19772);
and UO_375 (O_375,N_19874,N_19883);
or UO_376 (O_376,N_19796,N_19840);
nor UO_377 (O_377,N_19917,N_19801);
xor UO_378 (O_378,N_19883,N_19880);
xnor UO_379 (O_379,N_19838,N_19776);
or UO_380 (O_380,N_19969,N_19812);
nor UO_381 (O_381,N_19977,N_19922);
nand UO_382 (O_382,N_19789,N_19948);
or UO_383 (O_383,N_19753,N_19771);
and UO_384 (O_384,N_19819,N_19753);
nor UO_385 (O_385,N_19805,N_19828);
or UO_386 (O_386,N_19801,N_19896);
xor UO_387 (O_387,N_19777,N_19867);
or UO_388 (O_388,N_19875,N_19987);
nor UO_389 (O_389,N_19886,N_19982);
nand UO_390 (O_390,N_19979,N_19801);
and UO_391 (O_391,N_19959,N_19946);
nand UO_392 (O_392,N_19848,N_19999);
or UO_393 (O_393,N_19768,N_19760);
nand UO_394 (O_394,N_19858,N_19767);
and UO_395 (O_395,N_19999,N_19775);
nand UO_396 (O_396,N_19754,N_19917);
and UO_397 (O_397,N_19786,N_19982);
or UO_398 (O_398,N_19980,N_19761);
xnor UO_399 (O_399,N_19987,N_19780);
and UO_400 (O_400,N_19849,N_19825);
or UO_401 (O_401,N_19965,N_19961);
nand UO_402 (O_402,N_19852,N_19814);
nor UO_403 (O_403,N_19955,N_19864);
or UO_404 (O_404,N_19948,N_19782);
xnor UO_405 (O_405,N_19817,N_19797);
and UO_406 (O_406,N_19923,N_19966);
or UO_407 (O_407,N_19905,N_19848);
xor UO_408 (O_408,N_19856,N_19791);
xnor UO_409 (O_409,N_19908,N_19822);
nor UO_410 (O_410,N_19809,N_19998);
or UO_411 (O_411,N_19808,N_19877);
or UO_412 (O_412,N_19992,N_19753);
nand UO_413 (O_413,N_19844,N_19804);
xnor UO_414 (O_414,N_19979,N_19888);
xnor UO_415 (O_415,N_19797,N_19808);
nand UO_416 (O_416,N_19869,N_19856);
nor UO_417 (O_417,N_19876,N_19937);
nor UO_418 (O_418,N_19829,N_19882);
or UO_419 (O_419,N_19761,N_19916);
and UO_420 (O_420,N_19809,N_19794);
or UO_421 (O_421,N_19788,N_19915);
and UO_422 (O_422,N_19935,N_19754);
or UO_423 (O_423,N_19913,N_19783);
xnor UO_424 (O_424,N_19902,N_19801);
xor UO_425 (O_425,N_19993,N_19924);
and UO_426 (O_426,N_19918,N_19910);
and UO_427 (O_427,N_19927,N_19810);
or UO_428 (O_428,N_19777,N_19908);
nor UO_429 (O_429,N_19824,N_19786);
nand UO_430 (O_430,N_19762,N_19819);
nor UO_431 (O_431,N_19966,N_19856);
nor UO_432 (O_432,N_19993,N_19811);
nor UO_433 (O_433,N_19826,N_19784);
nor UO_434 (O_434,N_19754,N_19933);
or UO_435 (O_435,N_19872,N_19845);
and UO_436 (O_436,N_19862,N_19783);
xnor UO_437 (O_437,N_19959,N_19953);
nand UO_438 (O_438,N_19821,N_19853);
nor UO_439 (O_439,N_19755,N_19969);
xor UO_440 (O_440,N_19911,N_19773);
and UO_441 (O_441,N_19915,N_19860);
and UO_442 (O_442,N_19800,N_19773);
nand UO_443 (O_443,N_19888,N_19912);
nor UO_444 (O_444,N_19926,N_19753);
nand UO_445 (O_445,N_19997,N_19880);
nand UO_446 (O_446,N_19786,N_19783);
nor UO_447 (O_447,N_19863,N_19807);
nor UO_448 (O_448,N_19990,N_19807);
nor UO_449 (O_449,N_19840,N_19834);
nor UO_450 (O_450,N_19930,N_19848);
and UO_451 (O_451,N_19772,N_19769);
or UO_452 (O_452,N_19778,N_19822);
xnor UO_453 (O_453,N_19951,N_19958);
or UO_454 (O_454,N_19963,N_19922);
or UO_455 (O_455,N_19900,N_19881);
nand UO_456 (O_456,N_19928,N_19801);
or UO_457 (O_457,N_19768,N_19779);
or UO_458 (O_458,N_19861,N_19909);
or UO_459 (O_459,N_19842,N_19775);
xnor UO_460 (O_460,N_19988,N_19901);
and UO_461 (O_461,N_19930,N_19988);
xnor UO_462 (O_462,N_19807,N_19813);
and UO_463 (O_463,N_19954,N_19932);
or UO_464 (O_464,N_19973,N_19869);
and UO_465 (O_465,N_19827,N_19858);
xor UO_466 (O_466,N_19837,N_19905);
nand UO_467 (O_467,N_19910,N_19993);
nand UO_468 (O_468,N_19806,N_19785);
xor UO_469 (O_469,N_19781,N_19761);
nor UO_470 (O_470,N_19974,N_19773);
xor UO_471 (O_471,N_19986,N_19907);
and UO_472 (O_472,N_19765,N_19836);
and UO_473 (O_473,N_19768,N_19808);
xor UO_474 (O_474,N_19878,N_19901);
or UO_475 (O_475,N_19841,N_19914);
or UO_476 (O_476,N_19819,N_19811);
and UO_477 (O_477,N_19913,N_19885);
and UO_478 (O_478,N_19960,N_19812);
nand UO_479 (O_479,N_19946,N_19828);
or UO_480 (O_480,N_19791,N_19803);
or UO_481 (O_481,N_19754,N_19908);
xor UO_482 (O_482,N_19766,N_19883);
nor UO_483 (O_483,N_19915,N_19810);
or UO_484 (O_484,N_19876,N_19949);
nor UO_485 (O_485,N_19832,N_19927);
and UO_486 (O_486,N_19898,N_19977);
xnor UO_487 (O_487,N_19826,N_19991);
nand UO_488 (O_488,N_19940,N_19877);
nand UO_489 (O_489,N_19850,N_19871);
xor UO_490 (O_490,N_19794,N_19984);
nand UO_491 (O_491,N_19815,N_19854);
or UO_492 (O_492,N_19829,N_19950);
and UO_493 (O_493,N_19872,N_19806);
or UO_494 (O_494,N_19810,N_19845);
or UO_495 (O_495,N_19944,N_19921);
and UO_496 (O_496,N_19879,N_19848);
and UO_497 (O_497,N_19920,N_19796);
and UO_498 (O_498,N_19994,N_19910);
nor UO_499 (O_499,N_19831,N_19862);
or UO_500 (O_500,N_19752,N_19907);
nand UO_501 (O_501,N_19988,N_19801);
nor UO_502 (O_502,N_19971,N_19995);
and UO_503 (O_503,N_19884,N_19987);
nor UO_504 (O_504,N_19931,N_19951);
or UO_505 (O_505,N_19956,N_19812);
and UO_506 (O_506,N_19925,N_19835);
nor UO_507 (O_507,N_19897,N_19926);
and UO_508 (O_508,N_19894,N_19990);
nand UO_509 (O_509,N_19845,N_19765);
nand UO_510 (O_510,N_19976,N_19832);
nand UO_511 (O_511,N_19801,N_19796);
and UO_512 (O_512,N_19935,N_19889);
or UO_513 (O_513,N_19766,N_19767);
nand UO_514 (O_514,N_19857,N_19854);
and UO_515 (O_515,N_19902,N_19875);
nor UO_516 (O_516,N_19840,N_19961);
or UO_517 (O_517,N_19770,N_19909);
xnor UO_518 (O_518,N_19985,N_19815);
xor UO_519 (O_519,N_19809,N_19899);
or UO_520 (O_520,N_19772,N_19787);
xor UO_521 (O_521,N_19816,N_19881);
xor UO_522 (O_522,N_19950,N_19894);
nand UO_523 (O_523,N_19936,N_19817);
xor UO_524 (O_524,N_19906,N_19779);
nand UO_525 (O_525,N_19982,N_19958);
xnor UO_526 (O_526,N_19943,N_19978);
nor UO_527 (O_527,N_19895,N_19991);
nor UO_528 (O_528,N_19818,N_19871);
xor UO_529 (O_529,N_19802,N_19954);
xor UO_530 (O_530,N_19986,N_19976);
nand UO_531 (O_531,N_19843,N_19964);
xor UO_532 (O_532,N_19755,N_19986);
or UO_533 (O_533,N_19919,N_19927);
or UO_534 (O_534,N_19787,N_19883);
or UO_535 (O_535,N_19792,N_19957);
and UO_536 (O_536,N_19887,N_19891);
nand UO_537 (O_537,N_19910,N_19809);
or UO_538 (O_538,N_19838,N_19865);
nand UO_539 (O_539,N_19753,N_19985);
or UO_540 (O_540,N_19807,N_19848);
or UO_541 (O_541,N_19893,N_19873);
nor UO_542 (O_542,N_19896,N_19797);
and UO_543 (O_543,N_19919,N_19974);
xor UO_544 (O_544,N_19826,N_19975);
and UO_545 (O_545,N_19917,N_19810);
nor UO_546 (O_546,N_19823,N_19842);
nor UO_547 (O_547,N_19908,N_19805);
or UO_548 (O_548,N_19940,N_19765);
xnor UO_549 (O_549,N_19751,N_19842);
or UO_550 (O_550,N_19753,N_19856);
xor UO_551 (O_551,N_19918,N_19971);
or UO_552 (O_552,N_19910,N_19967);
nand UO_553 (O_553,N_19900,N_19752);
nor UO_554 (O_554,N_19860,N_19975);
nor UO_555 (O_555,N_19992,N_19982);
nand UO_556 (O_556,N_19816,N_19754);
nor UO_557 (O_557,N_19905,N_19947);
and UO_558 (O_558,N_19786,N_19927);
nand UO_559 (O_559,N_19761,N_19897);
and UO_560 (O_560,N_19934,N_19910);
nand UO_561 (O_561,N_19804,N_19986);
or UO_562 (O_562,N_19951,N_19922);
xor UO_563 (O_563,N_19847,N_19854);
nand UO_564 (O_564,N_19840,N_19973);
nor UO_565 (O_565,N_19920,N_19930);
nor UO_566 (O_566,N_19930,N_19814);
nor UO_567 (O_567,N_19947,N_19778);
xor UO_568 (O_568,N_19920,N_19924);
xor UO_569 (O_569,N_19827,N_19954);
nor UO_570 (O_570,N_19957,N_19905);
nor UO_571 (O_571,N_19893,N_19776);
nand UO_572 (O_572,N_19979,N_19978);
nor UO_573 (O_573,N_19997,N_19952);
nor UO_574 (O_574,N_19921,N_19852);
nor UO_575 (O_575,N_19823,N_19865);
nand UO_576 (O_576,N_19784,N_19899);
xnor UO_577 (O_577,N_19941,N_19880);
or UO_578 (O_578,N_19890,N_19924);
nor UO_579 (O_579,N_19823,N_19809);
or UO_580 (O_580,N_19819,N_19774);
nor UO_581 (O_581,N_19833,N_19856);
nor UO_582 (O_582,N_19840,N_19855);
nor UO_583 (O_583,N_19961,N_19753);
or UO_584 (O_584,N_19976,N_19907);
and UO_585 (O_585,N_19809,N_19813);
and UO_586 (O_586,N_19860,N_19781);
or UO_587 (O_587,N_19892,N_19896);
nand UO_588 (O_588,N_19763,N_19883);
nand UO_589 (O_589,N_19925,N_19814);
or UO_590 (O_590,N_19987,N_19994);
or UO_591 (O_591,N_19930,N_19971);
nand UO_592 (O_592,N_19767,N_19814);
and UO_593 (O_593,N_19870,N_19766);
xnor UO_594 (O_594,N_19860,N_19821);
or UO_595 (O_595,N_19864,N_19812);
xnor UO_596 (O_596,N_19941,N_19824);
xnor UO_597 (O_597,N_19767,N_19913);
nand UO_598 (O_598,N_19814,N_19824);
nand UO_599 (O_599,N_19893,N_19864);
and UO_600 (O_600,N_19770,N_19931);
or UO_601 (O_601,N_19947,N_19990);
nand UO_602 (O_602,N_19942,N_19844);
xnor UO_603 (O_603,N_19813,N_19914);
nand UO_604 (O_604,N_19922,N_19944);
nand UO_605 (O_605,N_19941,N_19957);
and UO_606 (O_606,N_19770,N_19822);
nor UO_607 (O_607,N_19844,N_19808);
nand UO_608 (O_608,N_19845,N_19928);
nor UO_609 (O_609,N_19977,N_19995);
xnor UO_610 (O_610,N_19885,N_19892);
nor UO_611 (O_611,N_19891,N_19995);
or UO_612 (O_612,N_19838,N_19799);
or UO_613 (O_613,N_19949,N_19801);
xor UO_614 (O_614,N_19869,N_19791);
and UO_615 (O_615,N_19768,N_19837);
nor UO_616 (O_616,N_19923,N_19795);
nand UO_617 (O_617,N_19851,N_19866);
xor UO_618 (O_618,N_19793,N_19896);
nor UO_619 (O_619,N_19776,N_19826);
or UO_620 (O_620,N_19797,N_19867);
nand UO_621 (O_621,N_19885,N_19773);
and UO_622 (O_622,N_19810,N_19928);
and UO_623 (O_623,N_19848,N_19869);
nand UO_624 (O_624,N_19978,N_19925);
nand UO_625 (O_625,N_19761,N_19772);
and UO_626 (O_626,N_19977,N_19862);
xor UO_627 (O_627,N_19962,N_19776);
and UO_628 (O_628,N_19896,N_19826);
xnor UO_629 (O_629,N_19895,N_19808);
xor UO_630 (O_630,N_19891,N_19826);
and UO_631 (O_631,N_19823,N_19775);
or UO_632 (O_632,N_19948,N_19867);
nor UO_633 (O_633,N_19754,N_19888);
xor UO_634 (O_634,N_19904,N_19786);
and UO_635 (O_635,N_19810,N_19980);
nor UO_636 (O_636,N_19923,N_19977);
and UO_637 (O_637,N_19920,N_19808);
xor UO_638 (O_638,N_19779,N_19876);
xor UO_639 (O_639,N_19922,N_19871);
and UO_640 (O_640,N_19882,N_19751);
xnor UO_641 (O_641,N_19767,N_19792);
and UO_642 (O_642,N_19906,N_19865);
nor UO_643 (O_643,N_19861,N_19789);
and UO_644 (O_644,N_19912,N_19867);
or UO_645 (O_645,N_19821,N_19875);
nor UO_646 (O_646,N_19920,N_19864);
xor UO_647 (O_647,N_19752,N_19929);
nor UO_648 (O_648,N_19977,N_19822);
xnor UO_649 (O_649,N_19816,N_19771);
nor UO_650 (O_650,N_19813,N_19917);
or UO_651 (O_651,N_19846,N_19761);
nor UO_652 (O_652,N_19899,N_19937);
or UO_653 (O_653,N_19756,N_19837);
nor UO_654 (O_654,N_19981,N_19792);
nor UO_655 (O_655,N_19986,N_19974);
and UO_656 (O_656,N_19826,N_19785);
xor UO_657 (O_657,N_19921,N_19926);
and UO_658 (O_658,N_19850,N_19811);
nor UO_659 (O_659,N_19783,N_19973);
xnor UO_660 (O_660,N_19983,N_19766);
or UO_661 (O_661,N_19814,N_19774);
or UO_662 (O_662,N_19860,N_19817);
or UO_663 (O_663,N_19821,N_19954);
nor UO_664 (O_664,N_19849,N_19750);
or UO_665 (O_665,N_19852,N_19915);
or UO_666 (O_666,N_19975,N_19923);
nand UO_667 (O_667,N_19873,N_19776);
xnor UO_668 (O_668,N_19999,N_19916);
xor UO_669 (O_669,N_19903,N_19895);
xnor UO_670 (O_670,N_19758,N_19817);
and UO_671 (O_671,N_19888,N_19971);
or UO_672 (O_672,N_19904,N_19777);
or UO_673 (O_673,N_19996,N_19865);
nand UO_674 (O_674,N_19764,N_19817);
and UO_675 (O_675,N_19924,N_19917);
or UO_676 (O_676,N_19808,N_19913);
nand UO_677 (O_677,N_19793,N_19981);
nand UO_678 (O_678,N_19858,N_19927);
or UO_679 (O_679,N_19903,N_19768);
nand UO_680 (O_680,N_19875,N_19767);
nand UO_681 (O_681,N_19863,N_19991);
and UO_682 (O_682,N_19838,N_19797);
nand UO_683 (O_683,N_19788,N_19864);
and UO_684 (O_684,N_19831,N_19968);
and UO_685 (O_685,N_19966,N_19976);
or UO_686 (O_686,N_19908,N_19860);
nand UO_687 (O_687,N_19834,N_19982);
or UO_688 (O_688,N_19839,N_19988);
and UO_689 (O_689,N_19937,N_19961);
or UO_690 (O_690,N_19796,N_19874);
nand UO_691 (O_691,N_19940,N_19985);
nand UO_692 (O_692,N_19828,N_19810);
xor UO_693 (O_693,N_19773,N_19774);
nand UO_694 (O_694,N_19918,N_19833);
and UO_695 (O_695,N_19943,N_19949);
nor UO_696 (O_696,N_19962,N_19846);
xor UO_697 (O_697,N_19849,N_19882);
nor UO_698 (O_698,N_19935,N_19784);
nand UO_699 (O_699,N_19947,N_19805);
nand UO_700 (O_700,N_19762,N_19820);
and UO_701 (O_701,N_19992,N_19785);
nor UO_702 (O_702,N_19971,N_19760);
or UO_703 (O_703,N_19881,N_19999);
nor UO_704 (O_704,N_19862,N_19941);
or UO_705 (O_705,N_19930,N_19871);
xor UO_706 (O_706,N_19900,N_19963);
or UO_707 (O_707,N_19821,N_19871);
or UO_708 (O_708,N_19932,N_19831);
or UO_709 (O_709,N_19945,N_19761);
or UO_710 (O_710,N_19791,N_19906);
nand UO_711 (O_711,N_19783,N_19883);
or UO_712 (O_712,N_19876,N_19938);
and UO_713 (O_713,N_19959,N_19882);
or UO_714 (O_714,N_19834,N_19771);
nand UO_715 (O_715,N_19935,N_19836);
nand UO_716 (O_716,N_19904,N_19750);
or UO_717 (O_717,N_19906,N_19852);
nand UO_718 (O_718,N_19823,N_19867);
nand UO_719 (O_719,N_19861,N_19796);
nor UO_720 (O_720,N_19881,N_19930);
nand UO_721 (O_721,N_19795,N_19863);
or UO_722 (O_722,N_19832,N_19850);
nand UO_723 (O_723,N_19829,N_19874);
and UO_724 (O_724,N_19825,N_19790);
nand UO_725 (O_725,N_19810,N_19958);
and UO_726 (O_726,N_19932,N_19884);
or UO_727 (O_727,N_19825,N_19818);
xnor UO_728 (O_728,N_19770,N_19844);
nand UO_729 (O_729,N_19825,N_19778);
xor UO_730 (O_730,N_19900,N_19792);
nor UO_731 (O_731,N_19775,N_19813);
nand UO_732 (O_732,N_19937,N_19932);
xor UO_733 (O_733,N_19994,N_19938);
or UO_734 (O_734,N_19986,N_19857);
xnor UO_735 (O_735,N_19800,N_19918);
and UO_736 (O_736,N_19815,N_19975);
xnor UO_737 (O_737,N_19931,N_19810);
or UO_738 (O_738,N_19914,N_19826);
or UO_739 (O_739,N_19760,N_19956);
or UO_740 (O_740,N_19750,N_19757);
or UO_741 (O_741,N_19881,N_19772);
nor UO_742 (O_742,N_19947,N_19930);
xor UO_743 (O_743,N_19760,N_19966);
nand UO_744 (O_744,N_19985,N_19750);
nand UO_745 (O_745,N_19807,N_19906);
nand UO_746 (O_746,N_19832,N_19901);
and UO_747 (O_747,N_19961,N_19892);
xor UO_748 (O_748,N_19825,N_19837);
nor UO_749 (O_749,N_19810,N_19856);
nor UO_750 (O_750,N_19987,N_19799);
nor UO_751 (O_751,N_19829,N_19957);
or UO_752 (O_752,N_19805,N_19757);
and UO_753 (O_753,N_19805,N_19891);
nor UO_754 (O_754,N_19905,N_19784);
or UO_755 (O_755,N_19869,N_19785);
or UO_756 (O_756,N_19874,N_19970);
and UO_757 (O_757,N_19907,N_19761);
and UO_758 (O_758,N_19791,N_19990);
nand UO_759 (O_759,N_19819,N_19798);
xnor UO_760 (O_760,N_19753,N_19910);
xnor UO_761 (O_761,N_19775,N_19889);
xor UO_762 (O_762,N_19911,N_19787);
nor UO_763 (O_763,N_19889,N_19972);
or UO_764 (O_764,N_19820,N_19958);
or UO_765 (O_765,N_19798,N_19783);
nor UO_766 (O_766,N_19825,N_19961);
nor UO_767 (O_767,N_19994,N_19820);
xnor UO_768 (O_768,N_19766,N_19829);
or UO_769 (O_769,N_19900,N_19761);
and UO_770 (O_770,N_19756,N_19982);
nor UO_771 (O_771,N_19795,N_19955);
nor UO_772 (O_772,N_19944,N_19844);
nor UO_773 (O_773,N_19759,N_19879);
and UO_774 (O_774,N_19845,N_19757);
nor UO_775 (O_775,N_19909,N_19881);
or UO_776 (O_776,N_19860,N_19807);
and UO_777 (O_777,N_19845,N_19956);
xor UO_778 (O_778,N_19922,N_19900);
nor UO_779 (O_779,N_19754,N_19903);
nand UO_780 (O_780,N_19801,N_19831);
nand UO_781 (O_781,N_19929,N_19955);
xor UO_782 (O_782,N_19771,N_19810);
nand UO_783 (O_783,N_19763,N_19799);
nand UO_784 (O_784,N_19859,N_19780);
nor UO_785 (O_785,N_19915,N_19774);
or UO_786 (O_786,N_19845,N_19832);
nor UO_787 (O_787,N_19894,N_19842);
or UO_788 (O_788,N_19793,N_19903);
nor UO_789 (O_789,N_19785,N_19979);
xnor UO_790 (O_790,N_19891,N_19843);
xnor UO_791 (O_791,N_19827,N_19901);
nand UO_792 (O_792,N_19762,N_19902);
xor UO_793 (O_793,N_19792,N_19859);
and UO_794 (O_794,N_19800,N_19779);
nor UO_795 (O_795,N_19935,N_19829);
or UO_796 (O_796,N_19800,N_19950);
or UO_797 (O_797,N_19853,N_19906);
xnor UO_798 (O_798,N_19898,N_19854);
nor UO_799 (O_799,N_19777,N_19951);
xor UO_800 (O_800,N_19794,N_19918);
nand UO_801 (O_801,N_19871,N_19896);
and UO_802 (O_802,N_19928,N_19893);
and UO_803 (O_803,N_19993,N_19832);
or UO_804 (O_804,N_19882,N_19845);
or UO_805 (O_805,N_19914,N_19794);
or UO_806 (O_806,N_19894,N_19889);
nand UO_807 (O_807,N_19820,N_19867);
xor UO_808 (O_808,N_19820,N_19817);
or UO_809 (O_809,N_19961,N_19936);
nor UO_810 (O_810,N_19798,N_19835);
nand UO_811 (O_811,N_19751,N_19902);
or UO_812 (O_812,N_19995,N_19976);
nand UO_813 (O_813,N_19994,N_19898);
nor UO_814 (O_814,N_19927,N_19875);
or UO_815 (O_815,N_19817,N_19876);
xor UO_816 (O_816,N_19947,N_19767);
nand UO_817 (O_817,N_19862,N_19838);
or UO_818 (O_818,N_19924,N_19901);
or UO_819 (O_819,N_19873,N_19784);
xnor UO_820 (O_820,N_19961,N_19967);
or UO_821 (O_821,N_19881,N_19870);
nand UO_822 (O_822,N_19777,N_19826);
nor UO_823 (O_823,N_19872,N_19844);
nand UO_824 (O_824,N_19804,N_19818);
xnor UO_825 (O_825,N_19888,N_19897);
nor UO_826 (O_826,N_19919,N_19990);
nand UO_827 (O_827,N_19905,N_19952);
or UO_828 (O_828,N_19885,N_19757);
nor UO_829 (O_829,N_19793,N_19806);
xor UO_830 (O_830,N_19893,N_19866);
nand UO_831 (O_831,N_19784,N_19780);
or UO_832 (O_832,N_19900,N_19890);
nor UO_833 (O_833,N_19790,N_19804);
and UO_834 (O_834,N_19813,N_19810);
or UO_835 (O_835,N_19811,N_19851);
and UO_836 (O_836,N_19880,N_19792);
and UO_837 (O_837,N_19954,N_19934);
xnor UO_838 (O_838,N_19894,N_19966);
nand UO_839 (O_839,N_19845,N_19955);
and UO_840 (O_840,N_19989,N_19799);
and UO_841 (O_841,N_19803,N_19832);
or UO_842 (O_842,N_19802,N_19950);
or UO_843 (O_843,N_19956,N_19958);
nor UO_844 (O_844,N_19994,N_19801);
nand UO_845 (O_845,N_19918,N_19808);
or UO_846 (O_846,N_19817,N_19898);
and UO_847 (O_847,N_19784,N_19833);
or UO_848 (O_848,N_19872,N_19949);
nor UO_849 (O_849,N_19969,N_19795);
xnor UO_850 (O_850,N_19824,N_19935);
nor UO_851 (O_851,N_19939,N_19934);
or UO_852 (O_852,N_19875,N_19811);
and UO_853 (O_853,N_19994,N_19844);
or UO_854 (O_854,N_19917,N_19820);
and UO_855 (O_855,N_19933,N_19978);
xnor UO_856 (O_856,N_19996,N_19910);
and UO_857 (O_857,N_19982,N_19903);
and UO_858 (O_858,N_19995,N_19914);
xor UO_859 (O_859,N_19789,N_19888);
nand UO_860 (O_860,N_19844,N_19961);
nor UO_861 (O_861,N_19777,N_19760);
and UO_862 (O_862,N_19757,N_19906);
nor UO_863 (O_863,N_19803,N_19859);
xnor UO_864 (O_864,N_19864,N_19939);
and UO_865 (O_865,N_19807,N_19945);
or UO_866 (O_866,N_19764,N_19876);
and UO_867 (O_867,N_19964,N_19762);
or UO_868 (O_868,N_19805,N_19780);
nand UO_869 (O_869,N_19834,N_19927);
nor UO_870 (O_870,N_19817,N_19967);
xnor UO_871 (O_871,N_19792,N_19896);
nand UO_872 (O_872,N_19795,N_19966);
nor UO_873 (O_873,N_19990,N_19870);
and UO_874 (O_874,N_19786,N_19787);
or UO_875 (O_875,N_19816,N_19791);
xnor UO_876 (O_876,N_19780,N_19929);
or UO_877 (O_877,N_19765,N_19786);
and UO_878 (O_878,N_19757,N_19976);
nor UO_879 (O_879,N_19827,N_19884);
or UO_880 (O_880,N_19876,N_19991);
nand UO_881 (O_881,N_19846,N_19837);
or UO_882 (O_882,N_19793,N_19804);
and UO_883 (O_883,N_19873,N_19962);
or UO_884 (O_884,N_19874,N_19906);
and UO_885 (O_885,N_19819,N_19767);
nand UO_886 (O_886,N_19919,N_19827);
or UO_887 (O_887,N_19958,N_19961);
and UO_888 (O_888,N_19903,N_19821);
or UO_889 (O_889,N_19789,N_19981);
nand UO_890 (O_890,N_19899,N_19761);
or UO_891 (O_891,N_19912,N_19756);
nor UO_892 (O_892,N_19803,N_19978);
nand UO_893 (O_893,N_19841,N_19845);
xnor UO_894 (O_894,N_19967,N_19933);
and UO_895 (O_895,N_19867,N_19956);
nor UO_896 (O_896,N_19780,N_19843);
xor UO_897 (O_897,N_19769,N_19829);
or UO_898 (O_898,N_19949,N_19901);
or UO_899 (O_899,N_19990,N_19991);
nor UO_900 (O_900,N_19781,N_19979);
and UO_901 (O_901,N_19896,N_19802);
nand UO_902 (O_902,N_19866,N_19945);
and UO_903 (O_903,N_19753,N_19790);
or UO_904 (O_904,N_19997,N_19936);
nor UO_905 (O_905,N_19877,N_19813);
nand UO_906 (O_906,N_19896,N_19757);
xnor UO_907 (O_907,N_19890,N_19753);
or UO_908 (O_908,N_19939,N_19990);
nand UO_909 (O_909,N_19924,N_19973);
and UO_910 (O_910,N_19836,N_19876);
nor UO_911 (O_911,N_19758,N_19879);
xor UO_912 (O_912,N_19781,N_19768);
or UO_913 (O_913,N_19871,N_19829);
nor UO_914 (O_914,N_19767,N_19894);
or UO_915 (O_915,N_19841,N_19936);
and UO_916 (O_916,N_19855,N_19811);
xnor UO_917 (O_917,N_19856,N_19817);
or UO_918 (O_918,N_19947,N_19835);
and UO_919 (O_919,N_19970,N_19941);
or UO_920 (O_920,N_19797,N_19791);
or UO_921 (O_921,N_19785,N_19751);
and UO_922 (O_922,N_19828,N_19897);
nor UO_923 (O_923,N_19994,N_19808);
or UO_924 (O_924,N_19861,N_19993);
nor UO_925 (O_925,N_19932,N_19927);
nand UO_926 (O_926,N_19845,N_19751);
and UO_927 (O_927,N_19892,N_19909);
and UO_928 (O_928,N_19957,N_19842);
nand UO_929 (O_929,N_19997,N_19761);
nand UO_930 (O_930,N_19893,N_19833);
and UO_931 (O_931,N_19791,N_19783);
nor UO_932 (O_932,N_19846,N_19956);
nor UO_933 (O_933,N_19773,N_19931);
nand UO_934 (O_934,N_19780,N_19931);
and UO_935 (O_935,N_19780,N_19926);
nand UO_936 (O_936,N_19916,N_19797);
and UO_937 (O_937,N_19794,N_19884);
and UO_938 (O_938,N_19756,N_19789);
xor UO_939 (O_939,N_19887,N_19755);
nand UO_940 (O_940,N_19941,N_19759);
or UO_941 (O_941,N_19852,N_19807);
or UO_942 (O_942,N_19900,N_19839);
and UO_943 (O_943,N_19843,N_19954);
xor UO_944 (O_944,N_19862,N_19843);
and UO_945 (O_945,N_19962,N_19772);
nand UO_946 (O_946,N_19781,N_19940);
nand UO_947 (O_947,N_19812,N_19891);
and UO_948 (O_948,N_19995,N_19810);
nor UO_949 (O_949,N_19997,N_19852);
nand UO_950 (O_950,N_19885,N_19834);
or UO_951 (O_951,N_19795,N_19810);
nor UO_952 (O_952,N_19911,N_19965);
nor UO_953 (O_953,N_19799,N_19906);
nand UO_954 (O_954,N_19841,N_19786);
and UO_955 (O_955,N_19821,N_19923);
or UO_956 (O_956,N_19854,N_19927);
nor UO_957 (O_957,N_19797,N_19789);
nor UO_958 (O_958,N_19977,N_19770);
xor UO_959 (O_959,N_19873,N_19774);
and UO_960 (O_960,N_19807,N_19887);
nand UO_961 (O_961,N_19825,N_19922);
nor UO_962 (O_962,N_19784,N_19773);
nand UO_963 (O_963,N_19809,N_19773);
xor UO_964 (O_964,N_19873,N_19832);
or UO_965 (O_965,N_19998,N_19754);
xnor UO_966 (O_966,N_19767,N_19836);
xor UO_967 (O_967,N_19830,N_19785);
and UO_968 (O_968,N_19804,N_19765);
and UO_969 (O_969,N_19935,N_19897);
nor UO_970 (O_970,N_19961,N_19989);
xnor UO_971 (O_971,N_19793,N_19897);
and UO_972 (O_972,N_19920,N_19876);
nand UO_973 (O_973,N_19780,N_19941);
xor UO_974 (O_974,N_19989,N_19800);
nor UO_975 (O_975,N_19916,N_19856);
or UO_976 (O_976,N_19824,N_19959);
or UO_977 (O_977,N_19850,N_19970);
and UO_978 (O_978,N_19847,N_19918);
or UO_979 (O_979,N_19999,N_19885);
xor UO_980 (O_980,N_19991,N_19977);
nand UO_981 (O_981,N_19793,N_19866);
xor UO_982 (O_982,N_19828,N_19804);
nand UO_983 (O_983,N_19915,N_19907);
xnor UO_984 (O_984,N_19869,N_19790);
xor UO_985 (O_985,N_19957,N_19841);
or UO_986 (O_986,N_19805,N_19969);
xor UO_987 (O_987,N_19913,N_19858);
xor UO_988 (O_988,N_19963,N_19899);
and UO_989 (O_989,N_19906,N_19892);
nand UO_990 (O_990,N_19861,N_19979);
nand UO_991 (O_991,N_19882,N_19942);
xnor UO_992 (O_992,N_19938,N_19768);
or UO_993 (O_993,N_19833,N_19837);
or UO_994 (O_994,N_19928,N_19942);
nand UO_995 (O_995,N_19966,N_19922);
or UO_996 (O_996,N_19861,N_19932);
or UO_997 (O_997,N_19888,N_19927);
nor UO_998 (O_998,N_19958,N_19866);
nand UO_999 (O_999,N_19841,N_19810);
or UO_1000 (O_1000,N_19927,N_19905);
or UO_1001 (O_1001,N_19940,N_19887);
or UO_1002 (O_1002,N_19971,N_19968);
nor UO_1003 (O_1003,N_19962,N_19967);
xor UO_1004 (O_1004,N_19835,N_19783);
nor UO_1005 (O_1005,N_19963,N_19843);
or UO_1006 (O_1006,N_19822,N_19821);
nor UO_1007 (O_1007,N_19785,N_19927);
and UO_1008 (O_1008,N_19812,N_19769);
xor UO_1009 (O_1009,N_19751,N_19826);
xor UO_1010 (O_1010,N_19871,N_19839);
and UO_1011 (O_1011,N_19780,N_19786);
xnor UO_1012 (O_1012,N_19991,N_19855);
nand UO_1013 (O_1013,N_19827,N_19935);
xnor UO_1014 (O_1014,N_19753,N_19798);
or UO_1015 (O_1015,N_19835,N_19789);
and UO_1016 (O_1016,N_19776,N_19886);
nor UO_1017 (O_1017,N_19952,N_19860);
nor UO_1018 (O_1018,N_19811,N_19784);
nand UO_1019 (O_1019,N_19831,N_19830);
or UO_1020 (O_1020,N_19936,N_19895);
or UO_1021 (O_1021,N_19987,N_19866);
nor UO_1022 (O_1022,N_19782,N_19916);
nand UO_1023 (O_1023,N_19761,N_19948);
nor UO_1024 (O_1024,N_19915,N_19976);
or UO_1025 (O_1025,N_19755,N_19823);
xor UO_1026 (O_1026,N_19885,N_19852);
nand UO_1027 (O_1027,N_19781,N_19759);
nor UO_1028 (O_1028,N_19870,N_19936);
and UO_1029 (O_1029,N_19838,N_19886);
or UO_1030 (O_1030,N_19928,N_19790);
and UO_1031 (O_1031,N_19846,N_19771);
nand UO_1032 (O_1032,N_19778,N_19960);
or UO_1033 (O_1033,N_19904,N_19842);
and UO_1034 (O_1034,N_19997,N_19862);
or UO_1035 (O_1035,N_19776,N_19903);
and UO_1036 (O_1036,N_19832,N_19782);
nor UO_1037 (O_1037,N_19843,N_19961);
or UO_1038 (O_1038,N_19930,N_19811);
or UO_1039 (O_1039,N_19772,N_19936);
nor UO_1040 (O_1040,N_19964,N_19884);
nor UO_1041 (O_1041,N_19874,N_19921);
nor UO_1042 (O_1042,N_19837,N_19859);
nor UO_1043 (O_1043,N_19818,N_19831);
or UO_1044 (O_1044,N_19854,N_19914);
nand UO_1045 (O_1045,N_19974,N_19795);
xor UO_1046 (O_1046,N_19770,N_19876);
xor UO_1047 (O_1047,N_19850,N_19797);
nor UO_1048 (O_1048,N_19940,N_19949);
and UO_1049 (O_1049,N_19898,N_19987);
nor UO_1050 (O_1050,N_19859,N_19933);
xnor UO_1051 (O_1051,N_19851,N_19973);
xor UO_1052 (O_1052,N_19951,N_19997);
nand UO_1053 (O_1053,N_19897,N_19934);
xor UO_1054 (O_1054,N_19920,N_19874);
and UO_1055 (O_1055,N_19970,N_19788);
xnor UO_1056 (O_1056,N_19757,N_19821);
or UO_1057 (O_1057,N_19913,N_19976);
and UO_1058 (O_1058,N_19829,N_19893);
nand UO_1059 (O_1059,N_19905,N_19883);
nand UO_1060 (O_1060,N_19971,N_19853);
nand UO_1061 (O_1061,N_19919,N_19851);
nand UO_1062 (O_1062,N_19986,N_19966);
nand UO_1063 (O_1063,N_19801,N_19850);
and UO_1064 (O_1064,N_19943,N_19908);
and UO_1065 (O_1065,N_19943,N_19874);
nand UO_1066 (O_1066,N_19847,N_19917);
nor UO_1067 (O_1067,N_19972,N_19902);
or UO_1068 (O_1068,N_19950,N_19893);
and UO_1069 (O_1069,N_19822,N_19860);
or UO_1070 (O_1070,N_19846,N_19769);
or UO_1071 (O_1071,N_19755,N_19797);
nand UO_1072 (O_1072,N_19867,N_19825);
xor UO_1073 (O_1073,N_19891,N_19947);
and UO_1074 (O_1074,N_19859,N_19900);
nor UO_1075 (O_1075,N_19868,N_19772);
xnor UO_1076 (O_1076,N_19850,N_19849);
nor UO_1077 (O_1077,N_19960,N_19935);
nand UO_1078 (O_1078,N_19988,N_19993);
or UO_1079 (O_1079,N_19929,N_19951);
and UO_1080 (O_1080,N_19993,N_19879);
and UO_1081 (O_1081,N_19911,N_19861);
and UO_1082 (O_1082,N_19779,N_19758);
nand UO_1083 (O_1083,N_19978,N_19903);
and UO_1084 (O_1084,N_19910,N_19959);
and UO_1085 (O_1085,N_19816,N_19768);
nor UO_1086 (O_1086,N_19985,N_19856);
xor UO_1087 (O_1087,N_19902,N_19764);
and UO_1088 (O_1088,N_19902,N_19913);
xor UO_1089 (O_1089,N_19789,N_19970);
nand UO_1090 (O_1090,N_19785,N_19863);
nand UO_1091 (O_1091,N_19969,N_19950);
nand UO_1092 (O_1092,N_19973,N_19756);
or UO_1093 (O_1093,N_19758,N_19856);
xor UO_1094 (O_1094,N_19883,N_19999);
nand UO_1095 (O_1095,N_19807,N_19971);
or UO_1096 (O_1096,N_19883,N_19885);
or UO_1097 (O_1097,N_19800,N_19924);
or UO_1098 (O_1098,N_19881,N_19760);
xnor UO_1099 (O_1099,N_19925,N_19811);
or UO_1100 (O_1100,N_19980,N_19884);
and UO_1101 (O_1101,N_19765,N_19979);
or UO_1102 (O_1102,N_19876,N_19820);
xor UO_1103 (O_1103,N_19866,N_19767);
nor UO_1104 (O_1104,N_19912,N_19877);
xor UO_1105 (O_1105,N_19845,N_19768);
or UO_1106 (O_1106,N_19917,N_19933);
nand UO_1107 (O_1107,N_19980,N_19842);
or UO_1108 (O_1108,N_19963,N_19983);
or UO_1109 (O_1109,N_19787,N_19861);
or UO_1110 (O_1110,N_19762,N_19945);
nor UO_1111 (O_1111,N_19994,N_19906);
or UO_1112 (O_1112,N_19805,N_19791);
or UO_1113 (O_1113,N_19782,N_19949);
nor UO_1114 (O_1114,N_19828,N_19801);
and UO_1115 (O_1115,N_19877,N_19871);
xor UO_1116 (O_1116,N_19846,N_19991);
xnor UO_1117 (O_1117,N_19751,N_19951);
or UO_1118 (O_1118,N_19881,N_19781);
and UO_1119 (O_1119,N_19853,N_19882);
xnor UO_1120 (O_1120,N_19925,N_19788);
xnor UO_1121 (O_1121,N_19824,N_19781);
xnor UO_1122 (O_1122,N_19899,N_19772);
xnor UO_1123 (O_1123,N_19848,N_19988);
and UO_1124 (O_1124,N_19979,N_19758);
xor UO_1125 (O_1125,N_19874,N_19754);
nor UO_1126 (O_1126,N_19949,N_19847);
or UO_1127 (O_1127,N_19765,N_19944);
and UO_1128 (O_1128,N_19849,N_19968);
nand UO_1129 (O_1129,N_19812,N_19771);
xor UO_1130 (O_1130,N_19814,N_19937);
nor UO_1131 (O_1131,N_19852,N_19911);
nor UO_1132 (O_1132,N_19752,N_19936);
nand UO_1133 (O_1133,N_19881,N_19922);
nor UO_1134 (O_1134,N_19803,N_19995);
and UO_1135 (O_1135,N_19986,N_19788);
nor UO_1136 (O_1136,N_19816,N_19885);
nand UO_1137 (O_1137,N_19834,N_19908);
xor UO_1138 (O_1138,N_19902,N_19956);
and UO_1139 (O_1139,N_19786,N_19985);
nor UO_1140 (O_1140,N_19919,N_19900);
and UO_1141 (O_1141,N_19827,N_19852);
nand UO_1142 (O_1142,N_19987,N_19818);
or UO_1143 (O_1143,N_19953,N_19806);
nor UO_1144 (O_1144,N_19859,N_19819);
and UO_1145 (O_1145,N_19792,N_19788);
nor UO_1146 (O_1146,N_19786,N_19878);
nor UO_1147 (O_1147,N_19976,N_19940);
or UO_1148 (O_1148,N_19789,N_19812);
and UO_1149 (O_1149,N_19788,N_19818);
nor UO_1150 (O_1150,N_19878,N_19956);
xor UO_1151 (O_1151,N_19866,N_19780);
nand UO_1152 (O_1152,N_19986,N_19874);
and UO_1153 (O_1153,N_19979,N_19887);
xor UO_1154 (O_1154,N_19798,N_19776);
and UO_1155 (O_1155,N_19991,N_19881);
nor UO_1156 (O_1156,N_19785,N_19787);
or UO_1157 (O_1157,N_19900,N_19847);
nand UO_1158 (O_1158,N_19815,N_19866);
xor UO_1159 (O_1159,N_19950,N_19883);
nand UO_1160 (O_1160,N_19905,N_19909);
or UO_1161 (O_1161,N_19889,N_19808);
or UO_1162 (O_1162,N_19787,N_19916);
nor UO_1163 (O_1163,N_19936,N_19950);
and UO_1164 (O_1164,N_19938,N_19837);
or UO_1165 (O_1165,N_19827,N_19891);
xor UO_1166 (O_1166,N_19784,N_19885);
nor UO_1167 (O_1167,N_19833,N_19804);
xor UO_1168 (O_1168,N_19810,N_19843);
xor UO_1169 (O_1169,N_19976,N_19916);
nand UO_1170 (O_1170,N_19801,N_19832);
xor UO_1171 (O_1171,N_19788,N_19964);
or UO_1172 (O_1172,N_19969,N_19903);
nand UO_1173 (O_1173,N_19939,N_19858);
and UO_1174 (O_1174,N_19907,N_19921);
and UO_1175 (O_1175,N_19951,N_19840);
and UO_1176 (O_1176,N_19846,N_19840);
and UO_1177 (O_1177,N_19947,N_19821);
or UO_1178 (O_1178,N_19863,N_19959);
nor UO_1179 (O_1179,N_19909,N_19866);
xor UO_1180 (O_1180,N_19940,N_19833);
and UO_1181 (O_1181,N_19888,N_19991);
nor UO_1182 (O_1182,N_19942,N_19892);
xnor UO_1183 (O_1183,N_19985,N_19834);
or UO_1184 (O_1184,N_19878,N_19823);
nand UO_1185 (O_1185,N_19999,N_19921);
or UO_1186 (O_1186,N_19855,N_19790);
or UO_1187 (O_1187,N_19801,N_19752);
and UO_1188 (O_1188,N_19881,N_19961);
nor UO_1189 (O_1189,N_19928,N_19808);
xnor UO_1190 (O_1190,N_19772,N_19991);
nor UO_1191 (O_1191,N_19889,N_19772);
nor UO_1192 (O_1192,N_19861,N_19841);
and UO_1193 (O_1193,N_19912,N_19814);
nand UO_1194 (O_1194,N_19855,N_19792);
or UO_1195 (O_1195,N_19925,N_19849);
nand UO_1196 (O_1196,N_19824,N_19878);
and UO_1197 (O_1197,N_19990,N_19756);
nor UO_1198 (O_1198,N_19893,N_19840);
and UO_1199 (O_1199,N_19973,N_19921);
nand UO_1200 (O_1200,N_19961,N_19912);
nor UO_1201 (O_1201,N_19763,N_19904);
nand UO_1202 (O_1202,N_19876,N_19975);
nor UO_1203 (O_1203,N_19959,N_19891);
nand UO_1204 (O_1204,N_19913,N_19832);
xnor UO_1205 (O_1205,N_19790,N_19813);
xnor UO_1206 (O_1206,N_19818,N_19905);
nand UO_1207 (O_1207,N_19912,N_19764);
or UO_1208 (O_1208,N_19985,N_19974);
nand UO_1209 (O_1209,N_19815,N_19805);
nand UO_1210 (O_1210,N_19966,N_19984);
nand UO_1211 (O_1211,N_19989,N_19839);
nor UO_1212 (O_1212,N_19894,N_19817);
nand UO_1213 (O_1213,N_19860,N_19984);
and UO_1214 (O_1214,N_19776,N_19880);
xor UO_1215 (O_1215,N_19985,N_19841);
and UO_1216 (O_1216,N_19852,N_19884);
nand UO_1217 (O_1217,N_19946,N_19920);
and UO_1218 (O_1218,N_19834,N_19901);
or UO_1219 (O_1219,N_19836,N_19925);
xnor UO_1220 (O_1220,N_19826,N_19793);
or UO_1221 (O_1221,N_19764,N_19768);
nand UO_1222 (O_1222,N_19983,N_19783);
nor UO_1223 (O_1223,N_19989,N_19981);
nand UO_1224 (O_1224,N_19954,N_19956);
nand UO_1225 (O_1225,N_19897,N_19848);
and UO_1226 (O_1226,N_19797,N_19894);
xor UO_1227 (O_1227,N_19802,N_19884);
or UO_1228 (O_1228,N_19961,N_19773);
and UO_1229 (O_1229,N_19778,N_19879);
nor UO_1230 (O_1230,N_19831,N_19911);
xnor UO_1231 (O_1231,N_19973,N_19775);
and UO_1232 (O_1232,N_19875,N_19922);
or UO_1233 (O_1233,N_19859,N_19994);
or UO_1234 (O_1234,N_19974,N_19906);
nor UO_1235 (O_1235,N_19866,N_19825);
and UO_1236 (O_1236,N_19803,N_19921);
and UO_1237 (O_1237,N_19826,N_19935);
or UO_1238 (O_1238,N_19970,N_19943);
and UO_1239 (O_1239,N_19914,N_19962);
nand UO_1240 (O_1240,N_19929,N_19829);
xor UO_1241 (O_1241,N_19931,N_19882);
xnor UO_1242 (O_1242,N_19961,N_19857);
xor UO_1243 (O_1243,N_19850,N_19844);
or UO_1244 (O_1244,N_19921,N_19875);
and UO_1245 (O_1245,N_19757,N_19799);
xnor UO_1246 (O_1246,N_19797,N_19965);
nand UO_1247 (O_1247,N_19886,N_19873);
xnor UO_1248 (O_1248,N_19876,N_19974);
and UO_1249 (O_1249,N_19918,N_19781);
nor UO_1250 (O_1250,N_19983,N_19912);
xor UO_1251 (O_1251,N_19952,N_19967);
and UO_1252 (O_1252,N_19788,N_19793);
xnor UO_1253 (O_1253,N_19854,N_19965);
and UO_1254 (O_1254,N_19772,N_19934);
xnor UO_1255 (O_1255,N_19876,N_19793);
nor UO_1256 (O_1256,N_19963,N_19868);
nor UO_1257 (O_1257,N_19773,N_19953);
xor UO_1258 (O_1258,N_19962,N_19767);
or UO_1259 (O_1259,N_19852,N_19989);
and UO_1260 (O_1260,N_19995,N_19967);
nor UO_1261 (O_1261,N_19899,N_19767);
and UO_1262 (O_1262,N_19808,N_19805);
and UO_1263 (O_1263,N_19819,N_19766);
nand UO_1264 (O_1264,N_19941,N_19830);
xor UO_1265 (O_1265,N_19919,N_19969);
and UO_1266 (O_1266,N_19997,N_19779);
and UO_1267 (O_1267,N_19895,N_19925);
xnor UO_1268 (O_1268,N_19967,N_19949);
nor UO_1269 (O_1269,N_19785,N_19965);
nor UO_1270 (O_1270,N_19801,N_19837);
xnor UO_1271 (O_1271,N_19768,N_19922);
or UO_1272 (O_1272,N_19895,N_19971);
xor UO_1273 (O_1273,N_19795,N_19865);
nand UO_1274 (O_1274,N_19907,N_19770);
xor UO_1275 (O_1275,N_19927,N_19933);
or UO_1276 (O_1276,N_19993,N_19836);
nor UO_1277 (O_1277,N_19915,N_19770);
nor UO_1278 (O_1278,N_19757,N_19925);
nand UO_1279 (O_1279,N_19984,N_19918);
and UO_1280 (O_1280,N_19889,N_19903);
or UO_1281 (O_1281,N_19826,N_19911);
xnor UO_1282 (O_1282,N_19945,N_19869);
nor UO_1283 (O_1283,N_19969,N_19959);
nor UO_1284 (O_1284,N_19797,N_19959);
and UO_1285 (O_1285,N_19923,N_19995);
xnor UO_1286 (O_1286,N_19972,N_19768);
nor UO_1287 (O_1287,N_19959,N_19944);
and UO_1288 (O_1288,N_19877,N_19999);
or UO_1289 (O_1289,N_19895,N_19764);
or UO_1290 (O_1290,N_19755,N_19848);
or UO_1291 (O_1291,N_19799,N_19918);
xor UO_1292 (O_1292,N_19822,N_19858);
xnor UO_1293 (O_1293,N_19856,N_19968);
or UO_1294 (O_1294,N_19766,N_19835);
and UO_1295 (O_1295,N_19802,N_19837);
nor UO_1296 (O_1296,N_19953,N_19837);
nand UO_1297 (O_1297,N_19928,N_19862);
or UO_1298 (O_1298,N_19942,N_19797);
nand UO_1299 (O_1299,N_19961,N_19897);
and UO_1300 (O_1300,N_19784,N_19978);
nand UO_1301 (O_1301,N_19862,N_19958);
or UO_1302 (O_1302,N_19931,N_19834);
or UO_1303 (O_1303,N_19936,N_19757);
nand UO_1304 (O_1304,N_19930,N_19994);
xnor UO_1305 (O_1305,N_19769,N_19892);
and UO_1306 (O_1306,N_19994,N_19969);
or UO_1307 (O_1307,N_19769,N_19827);
nor UO_1308 (O_1308,N_19815,N_19884);
nand UO_1309 (O_1309,N_19852,N_19902);
xor UO_1310 (O_1310,N_19764,N_19917);
nand UO_1311 (O_1311,N_19891,N_19775);
nand UO_1312 (O_1312,N_19990,N_19801);
or UO_1313 (O_1313,N_19889,N_19768);
xnor UO_1314 (O_1314,N_19907,N_19902);
xor UO_1315 (O_1315,N_19983,N_19834);
xor UO_1316 (O_1316,N_19778,N_19990);
xnor UO_1317 (O_1317,N_19875,N_19961);
xnor UO_1318 (O_1318,N_19862,N_19888);
or UO_1319 (O_1319,N_19869,N_19934);
nand UO_1320 (O_1320,N_19809,N_19859);
and UO_1321 (O_1321,N_19922,N_19867);
and UO_1322 (O_1322,N_19857,N_19881);
nor UO_1323 (O_1323,N_19959,N_19876);
xor UO_1324 (O_1324,N_19772,N_19752);
nand UO_1325 (O_1325,N_19758,N_19951);
or UO_1326 (O_1326,N_19814,N_19795);
or UO_1327 (O_1327,N_19897,N_19996);
nand UO_1328 (O_1328,N_19773,N_19980);
nor UO_1329 (O_1329,N_19979,N_19807);
xor UO_1330 (O_1330,N_19825,N_19773);
and UO_1331 (O_1331,N_19762,N_19989);
or UO_1332 (O_1332,N_19870,N_19978);
and UO_1333 (O_1333,N_19828,N_19947);
nor UO_1334 (O_1334,N_19809,N_19853);
nand UO_1335 (O_1335,N_19764,N_19900);
nor UO_1336 (O_1336,N_19805,N_19798);
nor UO_1337 (O_1337,N_19897,N_19864);
nand UO_1338 (O_1338,N_19858,N_19988);
or UO_1339 (O_1339,N_19976,N_19795);
nand UO_1340 (O_1340,N_19879,N_19892);
xnor UO_1341 (O_1341,N_19781,N_19997);
or UO_1342 (O_1342,N_19881,N_19945);
nor UO_1343 (O_1343,N_19907,N_19768);
nand UO_1344 (O_1344,N_19848,N_19829);
nand UO_1345 (O_1345,N_19895,N_19871);
xnor UO_1346 (O_1346,N_19985,N_19941);
nand UO_1347 (O_1347,N_19978,N_19995);
and UO_1348 (O_1348,N_19956,N_19916);
and UO_1349 (O_1349,N_19895,N_19981);
nor UO_1350 (O_1350,N_19987,N_19810);
or UO_1351 (O_1351,N_19753,N_19899);
nand UO_1352 (O_1352,N_19996,N_19853);
nand UO_1353 (O_1353,N_19756,N_19858);
xnor UO_1354 (O_1354,N_19858,N_19982);
nor UO_1355 (O_1355,N_19926,N_19890);
and UO_1356 (O_1356,N_19982,N_19851);
nand UO_1357 (O_1357,N_19785,N_19964);
xnor UO_1358 (O_1358,N_19752,N_19790);
or UO_1359 (O_1359,N_19931,N_19798);
or UO_1360 (O_1360,N_19794,N_19973);
or UO_1361 (O_1361,N_19890,N_19874);
nor UO_1362 (O_1362,N_19976,N_19782);
xnor UO_1363 (O_1363,N_19837,N_19914);
nor UO_1364 (O_1364,N_19776,N_19872);
or UO_1365 (O_1365,N_19945,N_19813);
or UO_1366 (O_1366,N_19812,N_19901);
xor UO_1367 (O_1367,N_19908,N_19892);
or UO_1368 (O_1368,N_19872,N_19890);
nand UO_1369 (O_1369,N_19873,N_19942);
and UO_1370 (O_1370,N_19977,N_19921);
xnor UO_1371 (O_1371,N_19854,N_19993);
nand UO_1372 (O_1372,N_19860,N_19974);
xor UO_1373 (O_1373,N_19929,N_19776);
nor UO_1374 (O_1374,N_19811,N_19762);
xnor UO_1375 (O_1375,N_19937,N_19758);
xor UO_1376 (O_1376,N_19914,N_19952);
or UO_1377 (O_1377,N_19882,N_19909);
nand UO_1378 (O_1378,N_19856,N_19848);
xor UO_1379 (O_1379,N_19845,N_19986);
nor UO_1380 (O_1380,N_19921,N_19930);
nor UO_1381 (O_1381,N_19973,N_19980);
or UO_1382 (O_1382,N_19931,N_19809);
xnor UO_1383 (O_1383,N_19891,N_19784);
nor UO_1384 (O_1384,N_19961,N_19974);
nand UO_1385 (O_1385,N_19882,N_19968);
and UO_1386 (O_1386,N_19855,N_19942);
or UO_1387 (O_1387,N_19833,N_19895);
and UO_1388 (O_1388,N_19823,N_19808);
xor UO_1389 (O_1389,N_19915,N_19948);
or UO_1390 (O_1390,N_19933,N_19804);
xnor UO_1391 (O_1391,N_19810,N_19750);
and UO_1392 (O_1392,N_19752,N_19925);
nor UO_1393 (O_1393,N_19837,N_19947);
xor UO_1394 (O_1394,N_19971,N_19793);
xor UO_1395 (O_1395,N_19837,N_19838);
and UO_1396 (O_1396,N_19865,N_19890);
nand UO_1397 (O_1397,N_19949,N_19851);
nor UO_1398 (O_1398,N_19863,N_19913);
and UO_1399 (O_1399,N_19792,N_19832);
nor UO_1400 (O_1400,N_19816,N_19807);
nor UO_1401 (O_1401,N_19983,N_19821);
nand UO_1402 (O_1402,N_19803,N_19960);
xor UO_1403 (O_1403,N_19975,N_19996);
nand UO_1404 (O_1404,N_19996,N_19833);
nor UO_1405 (O_1405,N_19887,N_19783);
nor UO_1406 (O_1406,N_19827,N_19920);
xnor UO_1407 (O_1407,N_19926,N_19867);
nor UO_1408 (O_1408,N_19912,N_19806);
nand UO_1409 (O_1409,N_19813,N_19820);
and UO_1410 (O_1410,N_19926,N_19758);
nand UO_1411 (O_1411,N_19913,N_19895);
nor UO_1412 (O_1412,N_19760,N_19765);
nor UO_1413 (O_1413,N_19974,N_19847);
xor UO_1414 (O_1414,N_19843,N_19955);
or UO_1415 (O_1415,N_19946,N_19823);
nand UO_1416 (O_1416,N_19892,N_19994);
nor UO_1417 (O_1417,N_19840,N_19955);
xor UO_1418 (O_1418,N_19809,N_19802);
nor UO_1419 (O_1419,N_19918,N_19954);
xor UO_1420 (O_1420,N_19952,N_19805);
and UO_1421 (O_1421,N_19901,N_19983);
or UO_1422 (O_1422,N_19838,N_19906);
nor UO_1423 (O_1423,N_19811,N_19782);
or UO_1424 (O_1424,N_19884,N_19972);
or UO_1425 (O_1425,N_19940,N_19854);
or UO_1426 (O_1426,N_19905,N_19871);
nand UO_1427 (O_1427,N_19988,N_19790);
nand UO_1428 (O_1428,N_19860,N_19836);
and UO_1429 (O_1429,N_19863,N_19806);
and UO_1430 (O_1430,N_19757,N_19828);
xor UO_1431 (O_1431,N_19815,N_19921);
nor UO_1432 (O_1432,N_19773,N_19968);
xnor UO_1433 (O_1433,N_19816,N_19960);
nor UO_1434 (O_1434,N_19876,N_19995);
or UO_1435 (O_1435,N_19973,N_19984);
nor UO_1436 (O_1436,N_19966,N_19971);
nor UO_1437 (O_1437,N_19916,N_19966);
nand UO_1438 (O_1438,N_19814,N_19781);
or UO_1439 (O_1439,N_19788,N_19892);
xor UO_1440 (O_1440,N_19874,N_19792);
nor UO_1441 (O_1441,N_19982,N_19868);
and UO_1442 (O_1442,N_19845,N_19766);
xnor UO_1443 (O_1443,N_19791,N_19833);
xnor UO_1444 (O_1444,N_19986,N_19964);
nor UO_1445 (O_1445,N_19854,N_19794);
or UO_1446 (O_1446,N_19819,N_19973);
nand UO_1447 (O_1447,N_19777,N_19991);
and UO_1448 (O_1448,N_19948,N_19836);
or UO_1449 (O_1449,N_19785,N_19852);
nand UO_1450 (O_1450,N_19908,N_19961);
and UO_1451 (O_1451,N_19812,N_19781);
or UO_1452 (O_1452,N_19973,N_19888);
and UO_1453 (O_1453,N_19955,N_19758);
xnor UO_1454 (O_1454,N_19904,N_19906);
or UO_1455 (O_1455,N_19950,N_19816);
and UO_1456 (O_1456,N_19756,N_19821);
or UO_1457 (O_1457,N_19891,N_19888);
and UO_1458 (O_1458,N_19907,N_19811);
nor UO_1459 (O_1459,N_19835,N_19949);
or UO_1460 (O_1460,N_19780,N_19969);
or UO_1461 (O_1461,N_19874,N_19905);
xnor UO_1462 (O_1462,N_19905,N_19827);
or UO_1463 (O_1463,N_19812,N_19821);
xor UO_1464 (O_1464,N_19961,N_19971);
and UO_1465 (O_1465,N_19914,N_19792);
and UO_1466 (O_1466,N_19794,N_19799);
nor UO_1467 (O_1467,N_19897,N_19756);
or UO_1468 (O_1468,N_19820,N_19954);
or UO_1469 (O_1469,N_19812,N_19992);
xnor UO_1470 (O_1470,N_19786,N_19871);
xor UO_1471 (O_1471,N_19983,N_19937);
nor UO_1472 (O_1472,N_19858,N_19936);
or UO_1473 (O_1473,N_19835,N_19964);
or UO_1474 (O_1474,N_19919,N_19918);
nor UO_1475 (O_1475,N_19904,N_19800);
nand UO_1476 (O_1476,N_19894,N_19897);
xor UO_1477 (O_1477,N_19897,N_19790);
and UO_1478 (O_1478,N_19910,N_19800);
nand UO_1479 (O_1479,N_19796,N_19816);
nand UO_1480 (O_1480,N_19803,N_19790);
or UO_1481 (O_1481,N_19942,N_19840);
xnor UO_1482 (O_1482,N_19991,N_19844);
and UO_1483 (O_1483,N_19773,N_19998);
nand UO_1484 (O_1484,N_19751,N_19901);
xnor UO_1485 (O_1485,N_19838,N_19911);
xor UO_1486 (O_1486,N_19859,N_19999);
and UO_1487 (O_1487,N_19787,N_19792);
nor UO_1488 (O_1488,N_19965,N_19829);
xnor UO_1489 (O_1489,N_19942,N_19810);
nor UO_1490 (O_1490,N_19831,N_19977);
or UO_1491 (O_1491,N_19949,N_19951);
and UO_1492 (O_1492,N_19916,N_19806);
nor UO_1493 (O_1493,N_19904,N_19859);
nand UO_1494 (O_1494,N_19779,N_19945);
or UO_1495 (O_1495,N_19848,N_19764);
nand UO_1496 (O_1496,N_19974,N_19838);
nor UO_1497 (O_1497,N_19930,N_19797);
or UO_1498 (O_1498,N_19999,N_19979);
and UO_1499 (O_1499,N_19799,N_19888);
nand UO_1500 (O_1500,N_19830,N_19760);
nand UO_1501 (O_1501,N_19858,N_19991);
and UO_1502 (O_1502,N_19794,N_19885);
nand UO_1503 (O_1503,N_19809,N_19996);
xnor UO_1504 (O_1504,N_19780,N_19801);
nor UO_1505 (O_1505,N_19860,N_19789);
nand UO_1506 (O_1506,N_19877,N_19781);
or UO_1507 (O_1507,N_19763,N_19781);
or UO_1508 (O_1508,N_19874,N_19849);
and UO_1509 (O_1509,N_19927,N_19994);
and UO_1510 (O_1510,N_19762,N_19909);
nor UO_1511 (O_1511,N_19783,N_19992);
or UO_1512 (O_1512,N_19956,N_19880);
and UO_1513 (O_1513,N_19960,N_19764);
nor UO_1514 (O_1514,N_19862,N_19942);
nand UO_1515 (O_1515,N_19761,N_19901);
nor UO_1516 (O_1516,N_19850,N_19758);
or UO_1517 (O_1517,N_19976,N_19776);
or UO_1518 (O_1518,N_19875,N_19986);
nand UO_1519 (O_1519,N_19764,N_19808);
or UO_1520 (O_1520,N_19956,N_19822);
xor UO_1521 (O_1521,N_19769,N_19881);
nor UO_1522 (O_1522,N_19764,N_19959);
or UO_1523 (O_1523,N_19943,N_19882);
nor UO_1524 (O_1524,N_19855,N_19959);
or UO_1525 (O_1525,N_19919,N_19807);
xnor UO_1526 (O_1526,N_19816,N_19925);
nand UO_1527 (O_1527,N_19968,N_19878);
or UO_1528 (O_1528,N_19838,N_19766);
nor UO_1529 (O_1529,N_19756,N_19813);
or UO_1530 (O_1530,N_19917,N_19763);
or UO_1531 (O_1531,N_19752,N_19917);
or UO_1532 (O_1532,N_19768,N_19881);
or UO_1533 (O_1533,N_19824,N_19768);
nor UO_1534 (O_1534,N_19859,N_19885);
and UO_1535 (O_1535,N_19869,N_19924);
and UO_1536 (O_1536,N_19885,N_19950);
and UO_1537 (O_1537,N_19958,N_19923);
or UO_1538 (O_1538,N_19963,N_19891);
nor UO_1539 (O_1539,N_19899,N_19905);
or UO_1540 (O_1540,N_19947,N_19971);
or UO_1541 (O_1541,N_19804,N_19839);
xnor UO_1542 (O_1542,N_19961,N_19938);
nand UO_1543 (O_1543,N_19774,N_19957);
nand UO_1544 (O_1544,N_19784,N_19912);
or UO_1545 (O_1545,N_19819,N_19850);
or UO_1546 (O_1546,N_19951,N_19923);
and UO_1547 (O_1547,N_19883,N_19997);
xor UO_1548 (O_1548,N_19850,N_19809);
xnor UO_1549 (O_1549,N_19936,N_19809);
and UO_1550 (O_1550,N_19938,N_19964);
nor UO_1551 (O_1551,N_19962,N_19835);
nand UO_1552 (O_1552,N_19764,N_19784);
xnor UO_1553 (O_1553,N_19875,N_19911);
or UO_1554 (O_1554,N_19811,N_19838);
or UO_1555 (O_1555,N_19786,N_19933);
xor UO_1556 (O_1556,N_19958,N_19884);
xor UO_1557 (O_1557,N_19907,N_19913);
nor UO_1558 (O_1558,N_19752,N_19854);
xor UO_1559 (O_1559,N_19880,N_19902);
and UO_1560 (O_1560,N_19862,N_19902);
xnor UO_1561 (O_1561,N_19919,N_19902);
and UO_1562 (O_1562,N_19761,N_19771);
xor UO_1563 (O_1563,N_19981,N_19947);
or UO_1564 (O_1564,N_19824,N_19865);
or UO_1565 (O_1565,N_19932,N_19955);
or UO_1566 (O_1566,N_19829,N_19994);
nand UO_1567 (O_1567,N_19868,N_19926);
and UO_1568 (O_1568,N_19851,N_19852);
or UO_1569 (O_1569,N_19995,N_19937);
or UO_1570 (O_1570,N_19984,N_19829);
nor UO_1571 (O_1571,N_19854,N_19948);
or UO_1572 (O_1572,N_19957,N_19837);
and UO_1573 (O_1573,N_19981,N_19856);
nor UO_1574 (O_1574,N_19783,N_19811);
xnor UO_1575 (O_1575,N_19913,N_19780);
or UO_1576 (O_1576,N_19871,N_19770);
xor UO_1577 (O_1577,N_19763,N_19968);
nand UO_1578 (O_1578,N_19981,N_19906);
and UO_1579 (O_1579,N_19786,N_19819);
xnor UO_1580 (O_1580,N_19873,N_19845);
xor UO_1581 (O_1581,N_19756,N_19975);
or UO_1582 (O_1582,N_19897,N_19918);
nand UO_1583 (O_1583,N_19829,N_19863);
and UO_1584 (O_1584,N_19990,N_19954);
xor UO_1585 (O_1585,N_19980,N_19851);
or UO_1586 (O_1586,N_19814,N_19904);
xnor UO_1587 (O_1587,N_19977,N_19996);
and UO_1588 (O_1588,N_19993,N_19778);
or UO_1589 (O_1589,N_19839,N_19939);
and UO_1590 (O_1590,N_19850,N_19934);
nand UO_1591 (O_1591,N_19808,N_19822);
or UO_1592 (O_1592,N_19911,N_19759);
xor UO_1593 (O_1593,N_19946,N_19884);
xnor UO_1594 (O_1594,N_19989,N_19814);
or UO_1595 (O_1595,N_19917,N_19830);
nor UO_1596 (O_1596,N_19762,N_19973);
xnor UO_1597 (O_1597,N_19792,N_19813);
nor UO_1598 (O_1598,N_19940,N_19848);
nand UO_1599 (O_1599,N_19947,N_19893);
or UO_1600 (O_1600,N_19768,N_19821);
xnor UO_1601 (O_1601,N_19945,N_19814);
or UO_1602 (O_1602,N_19789,N_19764);
nor UO_1603 (O_1603,N_19943,N_19828);
nand UO_1604 (O_1604,N_19823,N_19863);
and UO_1605 (O_1605,N_19776,N_19945);
and UO_1606 (O_1606,N_19808,N_19856);
nor UO_1607 (O_1607,N_19959,N_19929);
and UO_1608 (O_1608,N_19826,N_19982);
xor UO_1609 (O_1609,N_19845,N_19807);
nand UO_1610 (O_1610,N_19886,N_19884);
or UO_1611 (O_1611,N_19796,N_19824);
nand UO_1612 (O_1612,N_19998,N_19763);
nor UO_1613 (O_1613,N_19965,N_19909);
xor UO_1614 (O_1614,N_19928,N_19792);
nand UO_1615 (O_1615,N_19892,N_19761);
nand UO_1616 (O_1616,N_19998,N_19830);
xor UO_1617 (O_1617,N_19810,N_19756);
and UO_1618 (O_1618,N_19868,N_19936);
xnor UO_1619 (O_1619,N_19944,N_19782);
nor UO_1620 (O_1620,N_19779,N_19931);
nand UO_1621 (O_1621,N_19892,N_19784);
nand UO_1622 (O_1622,N_19809,N_19976);
nand UO_1623 (O_1623,N_19940,N_19819);
and UO_1624 (O_1624,N_19934,N_19912);
and UO_1625 (O_1625,N_19990,N_19969);
xor UO_1626 (O_1626,N_19751,N_19839);
or UO_1627 (O_1627,N_19915,N_19914);
nand UO_1628 (O_1628,N_19779,N_19755);
nand UO_1629 (O_1629,N_19913,N_19915);
and UO_1630 (O_1630,N_19809,N_19879);
and UO_1631 (O_1631,N_19923,N_19953);
nor UO_1632 (O_1632,N_19781,N_19776);
and UO_1633 (O_1633,N_19997,N_19990);
nor UO_1634 (O_1634,N_19786,N_19886);
nor UO_1635 (O_1635,N_19895,N_19954);
or UO_1636 (O_1636,N_19811,N_19936);
nor UO_1637 (O_1637,N_19829,N_19826);
nand UO_1638 (O_1638,N_19913,N_19756);
nand UO_1639 (O_1639,N_19941,N_19932);
nor UO_1640 (O_1640,N_19945,N_19952);
and UO_1641 (O_1641,N_19849,N_19959);
or UO_1642 (O_1642,N_19809,N_19797);
and UO_1643 (O_1643,N_19847,N_19967);
nand UO_1644 (O_1644,N_19916,N_19991);
or UO_1645 (O_1645,N_19965,N_19844);
nand UO_1646 (O_1646,N_19792,N_19779);
nand UO_1647 (O_1647,N_19998,N_19909);
or UO_1648 (O_1648,N_19789,N_19900);
nor UO_1649 (O_1649,N_19769,N_19838);
and UO_1650 (O_1650,N_19793,N_19751);
nand UO_1651 (O_1651,N_19754,N_19792);
and UO_1652 (O_1652,N_19765,N_19951);
nor UO_1653 (O_1653,N_19767,N_19785);
or UO_1654 (O_1654,N_19759,N_19858);
or UO_1655 (O_1655,N_19855,N_19858);
or UO_1656 (O_1656,N_19837,N_19872);
xnor UO_1657 (O_1657,N_19750,N_19791);
nor UO_1658 (O_1658,N_19812,N_19788);
and UO_1659 (O_1659,N_19802,N_19830);
xor UO_1660 (O_1660,N_19953,N_19878);
xor UO_1661 (O_1661,N_19961,N_19933);
and UO_1662 (O_1662,N_19968,N_19780);
nand UO_1663 (O_1663,N_19859,N_19954);
nand UO_1664 (O_1664,N_19945,N_19855);
nor UO_1665 (O_1665,N_19814,N_19947);
or UO_1666 (O_1666,N_19842,N_19940);
xor UO_1667 (O_1667,N_19789,N_19909);
nand UO_1668 (O_1668,N_19778,N_19934);
and UO_1669 (O_1669,N_19949,N_19813);
xor UO_1670 (O_1670,N_19864,N_19964);
nor UO_1671 (O_1671,N_19849,N_19945);
xnor UO_1672 (O_1672,N_19952,N_19896);
nand UO_1673 (O_1673,N_19926,N_19995);
and UO_1674 (O_1674,N_19916,N_19974);
or UO_1675 (O_1675,N_19813,N_19857);
nor UO_1676 (O_1676,N_19870,N_19922);
nor UO_1677 (O_1677,N_19969,N_19962);
nand UO_1678 (O_1678,N_19821,N_19828);
nor UO_1679 (O_1679,N_19865,N_19914);
and UO_1680 (O_1680,N_19970,N_19828);
nor UO_1681 (O_1681,N_19836,N_19812);
and UO_1682 (O_1682,N_19827,N_19968);
and UO_1683 (O_1683,N_19938,N_19853);
nor UO_1684 (O_1684,N_19879,N_19903);
nor UO_1685 (O_1685,N_19779,N_19828);
xor UO_1686 (O_1686,N_19818,N_19817);
nand UO_1687 (O_1687,N_19909,N_19887);
xnor UO_1688 (O_1688,N_19923,N_19999);
xor UO_1689 (O_1689,N_19758,N_19966);
nand UO_1690 (O_1690,N_19956,N_19913);
xor UO_1691 (O_1691,N_19827,N_19861);
and UO_1692 (O_1692,N_19999,N_19990);
or UO_1693 (O_1693,N_19821,N_19960);
and UO_1694 (O_1694,N_19944,N_19819);
or UO_1695 (O_1695,N_19919,N_19845);
nor UO_1696 (O_1696,N_19774,N_19923);
or UO_1697 (O_1697,N_19910,N_19790);
nor UO_1698 (O_1698,N_19781,N_19906);
xnor UO_1699 (O_1699,N_19892,N_19786);
or UO_1700 (O_1700,N_19770,N_19834);
nand UO_1701 (O_1701,N_19838,N_19916);
xnor UO_1702 (O_1702,N_19874,N_19937);
and UO_1703 (O_1703,N_19868,N_19791);
nand UO_1704 (O_1704,N_19889,N_19840);
nand UO_1705 (O_1705,N_19817,N_19951);
nor UO_1706 (O_1706,N_19775,N_19940);
and UO_1707 (O_1707,N_19784,N_19785);
nor UO_1708 (O_1708,N_19753,N_19831);
nor UO_1709 (O_1709,N_19983,N_19811);
nor UO_1710 (O_1710,N_19916,N_19943);
and UO_1711 (O_1711,N_19972,N_19908);
nor UO_1712 (O_1712,N_19957,N_19791);
and UO_1713 (O_1713,N_19786,N_19990);
or UO_1714 (O_1714,N_19757,N_19915);
nor UO_1715 (O_1715,N_19895,N_19785);
nor UO_1716 (O_1716,N_19918,N_19958);
nand UO_1717 (O_1717,N_19777,N_19990);
or UO_1718 (O_1718,N_19986,N_19793);
or UO_1719 (O_1719,N_19864,N_19996);
and UO_1720 (O_1720,N_19787,N_19793);
and UO_1721 (O_1721,N_19900,N_19911);
nand UO_1722 (O_1722,N_19752,N_19913);
nor UO_1723 (O_1723,N_19887,N_19811);
or UO_1724 (O_1724,N_19868,N_19790);
xnor UO_1725 (O_1725,N_19801,N_19811);
nor UO_1726 (O_1726,N_19797,N_19951);
and UO_1727 (O_1727,N_19793,N_19780);
or UO_1728 (O_1728,N_19952,N_19824);
nor UO_1729 (O_1729,N_19967,N_19988);
nor UO_1730 (O_1730,N_19901,N_19911);
nor UO_1731 (O_1731,N_19990,N_19785);
nor UO_1732 (O_1732,N_19921,N_19981);
nor UO_1733 (O_1733,N_19915,N_19975);
nand UO_1734 (O_1734,N_19756,N_19892);
or UO_1735 (O_1735,N_19921,N_19958);
and UO_1736 (O_1736,N_19898,N_19805);
xnor UO_1737 (O_1737,N_19883,N_19952);
or UO_1738 (O_1738,N_19895,N_19984);
or UO_1739 (O_1739,N_19797,N_19854);
and UO_1740 (O_1740,N_19835,N_19853);
and UO_1741 (O_1741,N_19818,N_19993);
nor UO_1742 (O_1742,N_19802,N_19888);
xor UO_1743 (O_1743,N_19762,N_19942);
xnor UO_1744 (O_1744,N_19880,N_19987);
and UO_1745 (O_1745,N_19958,N_19949);
and UO_1746 (O_1746,N_19787,N_19819);
and UO_1747 (O_1747,N_19891,N_19806);
nand UO_1748 (O_1748,N_19832,N_19973);
and UO_1749 (O_1749,N_19990,N_19896);
nor UO_1750 (O_1750,N_19760,N_19974);
and UO_1751 (O_1751,N_19935,N_19971);
and UO_1752 (O_1752,N_19869,N_19888);
xor UO_1753 (O_1753,N_19798,N_19920);
nor UO_1754 (O_1754,N_19752,N_19901);
or UO_1755 (O_1755,N_19912,N_19989);
or UO_1756 (O_1756,N_19823,N_19830);
xor UO_1757 (O_1757,N_19849,N_19881);
or UO_1758 (O_1758,N_19843,N_19750);
nor UO_1759 (O_1759,N_19876,N_19762);
nor UO_1760 (O_1760,N_19873,N_19961);
and UO_1761 (O_1761,N_19905,N_19891);
and UO_1762 (O_1762,N_19775,N_19811);
nand UO_1763 (O_1763,N_19836,N_19892);
nor UO_1764 (O_1764,N_19966,N_19860);
and UO_1765 (O_1765,N_19752,N_19899);
or UO_1766 (O_1766,N_19898,N_19942);
or UO_1767 (O_1767,N_19924,N_19885);
or UO_1768 (O_1768,N_19784,N_19882);
or UO_1769 (O_1769,N_19918,N_19767);
or UO_1770 (O_1770,N_19878,N_19857);
or UO_1771 (O_1771,N_19943,N_19820);
nand UO_1772 (O_1772,N_19794,N_19898);
xnor UO_1773 (O_1773,N_19866,N_19818);
or UO_1774 (O_1774,N_19883,N_19919);
nor UO_1775 (O_1775,N_19819,N_19958);
or UO_1776 (O_1776,N_19904,N_19809);
or UO_1777 (O_1777,N_19938,N_19931);
or UO_1778 (O_1778,N_19975,N_19904);
and UO_1779 (O_1779,N_19982,N_19840);
nand UO_1780 (O_1780,N_19872,N_19898);
and UO_1781 (O_1781,N_19917,N_19890);
or UO_1782 (O_1782,N_19755,N_19980);
and UO_1783 (O_1783,N_19753,N_19876);
nor UO_1784 (O_1784,N_19980,N_19944);
xnor UO_1785 (O_1785,N_19811,N_19872);
nor UO_1786 (O_1786,N_19761,N_19919);
or UO_1787 (O_1787,N_19994,N_19853);
nand UO_1788 (O_1788,N_19905,N_19847);
nor UO_1789 (O_1789,N_19940,N_19924);
and UO_1790 (O_1790,N_19792,N_19943);
and UO_1791 (O_1791,N_19990,N_19863);
xnor UO_1792 (O_1792,N_19771,N_19831);
xnor UO_1793 (O_1793,N_19777,N_19786);
nor UO_1794 (O_1794,N_19827,N_19990);
or UO_1795 (O_1795,N_19916,N_19789);
xnor UO_1796 (O_1796,N_19922,N_19930);
nand UO_1797 (O_1797,N_19797,N_19866);
nand UO_1798 (O_1798,N_19791,N_19921);
xor UO_1799 (O_1799,N_19761,N_19874);
or UO_1800 (O_1800,N_19856,N_19929);
or UO_1801 (O_1801,N_19948,N_19848);
nand UO_1802 (O_1802,N_19954,N_19848);
nor UO_1803 (O_1803,N_19808,N_19763);
and UO_1804 (O_1804,N_19813,N_19853);
and UO_1805 (O_1805,N_19966,N_19912);
xnor UO_1806 (O_1806,N_19968,N_19902);
or UO_1807 (O_1807,N_19841,N_19813);
xor UO_1808 (O_1808,N_19927,N_19846);
and UO_1809 (O_1809,N_19902,N_19836);
nor UO_1810 (O_1810,N_19925,N_19959);
nor UO_1811 (O_1811,N_19851,N_19765);
or UO_1812 (O_1812,N_19804,N_19796);
and UO_1813 (O_1813,N_19852,N_19896);
nor UO_1814 (O_1814,N_19839,N_19890);
and UO_1815 (O_1815,N_19858,N_19804);
nand UO_1816 (O_1816,N_19913,N_19985);
nor UO_1817 (O_1817,N_19952,N_19985);
and UO_1818 (O_1818,N_19924,N_19792);
nand UO_1819 (O_1819,N_19754,N_19915);
or UO_1820 (O_1820,N_19836,N_19981);
or UO_1821 (O_1821,N_19770,N_19932);
nand UO_1822 (O_1822,N_19852,N_19925);
nand UO_1823 (O_1823,N_19820,N_19837);
and UO_1824 (O_1824,N_19770,N_19950);
nand UO_1825 (O_1825,N_19875,N_19853);
nand UO_1826 (O_1826,N_19781,N_19894);
xor UO_1827 (O_1827,N_19960,N_19899);
or UO_1828 (O_1828,N_19892,N_19953);
xnor UO_1829 (O_1829,N_19826,N_19781);
and UO_1830 (O_1830,N_19921,N_19904);
nand UO_1831 (O_1831,N_19848,N_19819);
or UO_1832 (O_1832,N_19896,N_19917);
or UO_1833 (O_1833,N_19756,N_19916);
xnor UO_1834 (O_1834,N_19827,N_19822);
nand UO_1835 (O_1835,N_19948,N_19776);
and UO_1836 (O_1836,N_19808,N_19975);
and UO_1837 (O_1837,N_19842,N_19869);
nor UO_1838 (O_1838,N_19913,N_19975);
or UO_1839 (O_1839,N_19942,N_19860);
and UO_1840 (O_1840,N_19851,N_19782);
or UO_1841 (O_1841,N_19886,N_19953);
nand UO_1842 (O_1842,N_19974,N_19914);
nand UO_1843 (O_1843,N_19818,N_19756);
nand UO_1844 (O_1844,N_19750,N_19898);
and UO_1845 (O_1845,N_19950,N_19820);
xnor UO_1846 (O_1846,N_19874,N_19924);
nor UO_1847 (O_1847,N_19919,N_19804);
nor UO_1848 (O_1848,N_19904,N_19792);
xnor UO_1849 (O_1849,N_19933,N_19812);
nand UO_1850 (O_1850,N_19966,N_19759);
and UO_1851 (O_1851,N_19807,N_19950);
nand UO_1852 (O_1852,N_19783,N_19963);
or UO_1853 (O_1853,N_19750,N_19835);
xnor UO_1854 (O_1854,N_19892,N_19866);
nor UO_1855 (O_1855,N_19924,N_19768);
nor UO_1856 (O_1856,N_19784,N_19964);
nor UO_1857 (O_1857,N_19766,N_19860);
nand UO_1858 (O_1858,N_19826,N_19780);
and UO_1859 (O_1859,N_19755,N_19845);
or UO_1860 (O_1860,N_19887,N_19856);
nand UO_1861 (O_1861,N_19994,N_19830);
nor UO_1862 (O_1862,N_19828,N_19984);
and UO_1863 (O_1863,N_19849,N_19816);
nor UO_1864 (O_1864,N_19965,N_19992);
nor UO_1865 (O_1865,N_19839,N_19856);
and UO_1866 (O_1866,N_19861,N_19985);
or UO_1867 (O_1867,N_19769,N_19988);
xor UO_1868 (O_1868,N_19801,N_19844);
xnor UO_1869 (O_1869,N_19754,N_19938);
nor UO_1870 (O_1870,N_19976,N_19792);
and UO_1871 (O_1871,N_19796,N_19991);
nand UO_1872 (O_1872,N_19912,N_19843);
nand UO_1873 (O_1873,N_19838,N_19834);
nor UO_1874 (O_1874,N_19954,N_19750);
or UO_1875 (O_1875,N_19793,N_19855);
xor UO_1876 (O_1876,N_19778,N_19981);
or UO_1877 (O_1877,N_19865,N_19896);
nand UO_1878 (O_1878,N_19840,N_19879);
nand UO_1879 (O_1879,N_19830,N_19961);
or UO_1880 (O_1880,N_19919,N_19808);
or UO_1881 (O_1881,N_19816,N_19970);
nand UO_1882 (O_1882,N_19807,N_19850);
or UO_1883 (O_1883,N_19796,N_19999);
xnor UO_1884 (O_1884,N_19762,N_19994);
xor UO_1885 (O_1885,N_19854,N_19806);
or UO_1886 (O_1886,N_19787,N_19969);
and UO_1887 (O_1887,N_19923,N_19940);
nand UO_1888 (O_1888,N_19942,N_19930);
or UO_1889 (O_1889,N_19795,N_19892);
and UO_1890 (O_1890,N_19783,N_19869);
xnor UO_1891 (O_1891,N_19776,N_19841);
nor UO_1892 (O_1892,N_19887,N_19768);
xor UO_1893 (O_1893,N_19788,N_19842);
and UO_1894 (O_1894,N_19970,N_19797);
or UO_1895 (O_1895,N_19877,N_19865);
xor UO_1896 (O_1896,N_19845,N_19969);
xor UO_1897 (O_1897,N_19931,N_19962);
xor UO_1898 (O_1898,N_19813,N_19953);
nor UO_1899 (O_1899,N_19901,N_19795);
nor UO_1900 (O_1900,N_19821,N_19834);
nand UO_1901 (O_1901,N_19904,N_19981);
and UO_1902 (O_1902,N_19918,N_19786);
nor UO_1903 (O_1903,N_19782,N_19894);
and UO_1904 (O_1904,N_19784,N_19985);
nor UO_1905 (O_1905,N_19965,N_19884);
nor UO_1906 (O_1906,N_19794,N_19893);
nor UO_1907 (O_1907,N_19968,N_19786);
and UO_1908 (O_1908,N_19761,N_19964);
and UO_1909 (O_1909,N_19804,N_19789);
xnor UO_1910 (O_1910,N_19844,N_19955);
and UO_1911 (O_1911,N_19802,N_19959);
xor UO_1912 (O_1912,N_19904,N_19882);
xor UO_1913 (O_1913,N_19994,N_19936);
or UO_1914 (O_1914,N_19923,N_19760);
and UO_1915 (O_1915,N_19941,N_19811);
nand UO_1916 (O_1916,N_19923,N_19871);
nor UO_1917 (O_1917,N_19916,N_19954);
nor UO_1918 (O_1918,N_19881,N_19779);
nor UO_1919 (O_1919,N_19990,N_19942);
nand UO_1920 (O_1920,N_19927,N_19762);
nor UO_1921 (O_1921,N_19972,N_19995);
or UO_1922 (O_1922,N_19990,N_19972);
xor UO_1923 (O_1923,N_19820,N_19965);
xor UO_1924 (O_1924,N_19867,N_19986);
xor UO_1925 (O_1925,N_19755,N_19806);
nor UO_1926 (O_1926,N_19768,N_19847);
nor UO_1927 (O_1927,N_19930,N_19783);
nor UO_1928 (O_1928,N_19776,N_19995);
or UO_1929 (O_1929,N_19875,N_19899);
and UO_1930 (O_1930,N_19776,N_19792);
xor UO_1931 (O_1931,N_19799,N_19931);
nand UO_1932 (O_1932,N_19960,N_19924);
or UO_1933 (O_1933,N_19890,N_19919);
nor UO_1934 (O_1934,N_19886,N_19763);
and UO_1935 (O_1935,N_19914,N_19944);
xor UO_1936 (O_1936,N_19914,N_19979);
nor UO_1937 (O_1937,N_19944,N_19974);
nand UO_1938 (O_1938,N_19882,N_19941);
nand UO_1939 (O_1939,N_19883,N_19832);
or UO_1940 (O_1940,N_19777,N_19885);
xor UO_1941 (O_1941,N_19792,N_19805);
or UO_1942 (O_1942,N_19834,N_19772);
nand UO_1943 (O_1943,N_19984,N_19889);
nor UO_1944 (O_1944,N_19797,N_19936);
nor UO_1945 (O_1945,N_19770,N_19883);
xnor UO_1946 (O_1946,N_19895,N_19831);
or UO_1947 (O_1947,N_19951,N_19778);
nand UO_1948 (O_1948,N_19789,N_19858);
xor UO_1949 (O_1949,N_19963,N_19760);
xnor UO_1950 (O_1950,N_19971,N_19801);
nor UO_1951 (O_1951,N_19899,N_19860);
and UO_1952 (O_1952,N_19994,N_19993);
nand UO_1953 (O_1953,N_19949,N_19757);
xnor UO_1954 (O_1954,N_19986,N_19898);
xnor UO_1955 (O_1955,N_19978,N_19911);
xnor UO_1956 (O_1956,N_19956,N_19853);
and UO_1957 (O_1957,N_19943,N_19941);
xnor UO_1958 (O_1958,N_19921,N_19898);
and UO_1959 (O_1959,N_19989,N_19973);
nor UO_1960 (O_1960,N_19867,N_19974);
nand UO_1961 (O_1961,N_19907,N_19864);
and UO_1962 (O_1962,N_19864,N_19928);
or UO_1963 (O_1963,N_19867,N_19795);
nand UO_1964 (O_1964,N_19835,N_19940);
nand UO_1965 (O_1965,N_19884,N_19767);
nor UO_1966 (O_1966,N_19879,N_19972);
xnor UO_1967 (O_1967,N_19995,N_19992);
or UO_1968 (O_1968,N_19826,N_19890);
nand UO_1969 (O_1969,N_19805,N_19924);
nand UO_1970 (O_1970,N_19809,N_19868);
or UO_1971 (O_1971,N_19931,N_19878);
and UO_1972 (O_1972,N_19756,N_19968);
nand UO_1973 (O_1973,N_19841,N_19855);
nand UO_1974 (O_1974,N_19904,N_19802);
and UO_1975 (O_1975,N_19860,N_19797);
and UO_1976 (O_1976,N_19755,N_19926);
xnor UO_1977 (O_1977,N_19942,N_19987);
and UO_1978 (O_1978,N_19880,N_19793);
and UO_1979 (O_1979,N_19870,N_19895);
and UO_1980 (O_1980,N_19783,N_19906);
xnor UO_1981 (O_1981,N_19935,N_19896);
and UO_1982 (O_1982,N_19924,N_19771);
nor UO_1983 (O_1983,N_19951,N_19767);
nor UO_1984 (O_1984,N_19949,N_19791);
nand UO_1985 (O_1985,N_19902,N_19877);
nand UO_1986 (O_1986,N_19928,N_19848);
nand UO_1987 (O_1987,N_19998,N_19844);
and UO_1988 (O_1988,N_19880,N_19829);
nand UO_1989 (O_1989,N_19850,N_19981);
nand UO_1990 (O_1990,N_19953,N_19763);
nor UO_1991 (O_1991,N_19776,N_19766);
nor UO_1992 (O_1992,N_19976,N_19840);
or UO_1993 (O_1993,N_19987,N_19894);
nand UO_1994 (O_1994,N_19888,N_19977);
xor UO_1995 (O_1995,N_19913,N_19992);
nor UO_1996 (O_1996,N_19784,N_19752);
nand UO_1997 (O_1997,N_19751,N_19930);
and UO_1998 (O_1998,N_19889,N_19755);
xnor UO_1999 (O_1999,N_19812,N_19805);
nand UO_2000 (O_2000,N_19902,N_19797);
nand UO_2001 (O_2001,N_19751,N_19981);
and UO_2002 (O_2002,N_19879,N_19906);
and UO_2003 (O_2003,N_19920,N_19941);
nand UO_2004 (O_2004,N_19885,N_19771);
or UO_2005 (O_2005,N_19907,N_19771);
nand UO_2006 (O_2006,N_19936,N_19877);
or UO_2007 (O_2007,N_19781,N_19916);
nand UO_2008 (O_2008,N_19988,N_19780);
xnor UO_2009 (O_2009,N_19850,N_19777);
nand UO_2010 (O_2010,N_19911,N_19977);
and UO_2011 (O_2011,N_19962,N_19985);
or UO_2012 (O_2012,N_19942,N_19880);
or UO_2013 (O_2013,N_19843,N_19775);
and UO_2014 (O_2014,N_19974,N_19873);
xor UO_2015 (O_2015,N_19885,N_19914);
xor UO_2016 (O_2016,N_19876,N_19796);
or UO_2017 (O_2017,N_19779,N_19930);
or UO_2018 (O_2018,N_19770,N_19988);
nand UO_2019 (O_2019,N_19842,N_19918);
nand UO_2020 (O_2020,N_19968,N_19978);
nand UO_2021 (O_2021,N_19885,N_19811);
or UO_2022 (O_2022,N_19826,N_19993);
nand UO_2023 (O_2023,N_19829,N_19978);
xnor UO_2024 (O_2024,N_19919,N_19958);
xnor UO_2025 (O_2025,N_19939,N_19792);
nand UO_2026 (O_2026,N_19991,N_19907);
or UO_2027 (O_2027,N_19872,N_19963);
and UO_2028 (O_2028,N_19982,N_19950);
nor UO_2029 (O_2029,N_19871,N_19912);
nand UO_2030 (O_2030,N_19865,N_19924);
or UO_2031 (O_2031,N_19884,N_19785);
and UO_2032 (O_2032,N_19864,N_19935);
nor UO_2033 (O_2033,N_19789,N_19798);
and UO_2034 (O_2034,N_19980,N_19961);
nor UO_2035 (O_2035,N_19891,N_19999);
and UO_2036 (O_2036,N_19926,N_19899);
nand UO_2037 (O_2037,N_19817,N_19825);
nor UO_2038 (O_2038,N_19822,N_19867);
nand UO_2039 (O_2039,N_19825,N_19820);
nand UO_2040 (O_2040,N_19999,N_19765);
and UO_2041 (O_2041,N_19870,N_19924);
or UO_2042 (O_2042,N_19855,N_19962);
xnor UO_2043 (O_2043,N_19934,N_19876);
or UO_2044 (O_2044,N_19943,N_19889);
nor UO_2045 (O_2045,N_19900,N_19877);
or UO_2046 (O_2046,N_19760,N_19811);
and UO_2047 (O_2047,N_19876,N_19857);
nor UO_2048 (O_2048,N_19909,N_19943);
nand UO_2049 (O_2049,N_19819,N_19968);
xnor UO_2050 (O_2050,N_19969,N_19975);
xnor UO_2051 (O_2051,N_19954,N_19996);
xnor UO_2052 (O_2052,N_19885,N_19765);
nand UO_2053 (O_2053,N_19866,N_19894);
or UO_2054 (O_2054,N_19751,N_19946);
nand UO_2055 (O_2055,N_19974,N_19764);
nor UO_2056 (O_2056,N_19980,N_19981);
nand UO_2057 (O_2057,N_19816,N_19770);
and UO_2058 (O_2058,N_19772,N_19908);
or UO_2059 (O_2059,N_19986,N_19984);
or UO_2060 (O_2060,N_19772,N_19759);
nor UO_2061 (O_2061,N_19957,N_19838);
nor UO_2062 (O_2062,N_19756,N_19927);
or UO_2063 (O_2063,N_19978,N_19874);
and UO_2064 (O_2064,N_19807,N_19921);
xnor UO_2065 (O_2065,N_19999,N_19961);
xnor UO_2066 (O_2066,N_19979,N_19929);
nor UO_2067 (O_2067,N_19853,N_19858);
xor UO_2068 (O_2068,N_19868,N_19837);
and UO_2069 (O_2069,N_19806,N_19889);
xor UO_2070 (O_2070,N_19846,N_19878);
xor UO_2071 (O_2071,N_19875,N_19972);
xor UO_2072 (O_2072,N_19852,N_19891);
nor UO_2073 (O_2073,N_19974,N_19883);
or UO_2074 (O_2074,N_19791,N_19812);
and UO_2075 (O_2075,N_19764,N_19860);
nor UO_2076 (O_2076,N_19977,N_19779);
and UO_2077 (O_2077,N_19958,N_19799);
nand UO_2078 (O_2078,N_19804,N_19893);
nand UO_2079 (O_2079,N_19877,N_19982);
nor UO_2080 (O_2080,N_19904,N_19785);
and UO_2081 (O_2081,N_19948,N_19857);
nand UO_2082 (O_2082,N_19897,N_19879);
nand UO_2083 (O_2083,N_19750,N_19827);
nor UO_2084 (O_2084,N_19780,N_19928);
nand UO_2085 (O_2085,N_19922,N_19928);
xor UO_2086 (O_2086,N_19900,N_19768);
nand UO_2087 (O_2087,N_19756,N_19929);
and UO_2088 (O_2088,N_19965,N_19880);
or UO_2089 (O_2089,N_19841,N_19754);
xnor UO_2090 (O_2090,N_19859,N_19897);
and UO_2091 (O_2091,N_19872,N_19863);
nand UO_2092 (O_2092,N_19825,N_19863);
or UO_2093 (O_2093,N_19782,N_19971);
nand UO_2094 (O_2094,N_19888,N_19774);
and UO_2095 (O_2095,N_19871,N_19961);
xor UO_2096 (O_2096,N_19854,N_19941);
xnor UO_2097 (O_2097,N_19757,N_19809);
and UO_2098 (O_2098,N_19779,N_19872);
nand UO_2099 (O_2099,N_19977,N_19819);
nor UO_2100 (O_2100,N_19891,N_19830);
nor UO_2101 (O_2101,N_19827,N_19894);
or UO_2102 (O_2102,N_19806,N_19952);
nand UO_2103 (O_2103,N_19960,N_19765);
nand UO_2104 (O_2104,N_19947,N_19804);
nor UO_2105 (O_2105,N_19880,N_19809);
nand UO_2106 (O_2106,N_19826,N_19768);
or UO_2107 (O_2107,N_19760,N_19751);
nor UO_2108 (O_2108,N_19773,N_19793);
and UO_2109 (O_2109,N_19926,N_19979);
and UO_2110 (O_2110,N_19959,N_19832);
nor UO_2111 (O_2111,N_19812,N_19776);
nand UO_2112 (O_2112,N_19878,N_19954);
nand UO_2113 (O_2113,N_19935,N_19930);
xnor UO_2114 (O_2114,N_19846,N_19998);
or UO_2115 (O_2115,N_19769,N_19931);
nand UO_2116 (O_2116,N_19867,N_19790);
nand UO_2117 (O_2117,N_19925,N_19761);
and UO_2118 (O_2118,N_19800,N_19772);
xor UO_2119 (O_2119,N_19862,N_19828);
and UO_2120 (O_2120,N_19866,N_19835);
nand UO_2121 (O_2121,N_19878,N_19922);
xnor UO_2122 (O_2122,N_19840,N_19765);
nor UO_2123 (O_2123,N_19773,N_19854);
nand UO_2124 (O_2124,N_19783,N_19865);
xor UO_2125 (O_2125,N_19827,N_19829);
nand UO_2126 (O_2126,N_19973,N_19809);
nand UO_2127 (O_2127,N_19939,N_19966);
nand UO_2128 (O_2128,N_19985,N_19774);
nand UO_2129 (O_2129,N_19775,N_19877);
nand UO_2130 (O_2130,N_19847,N_19957);
and UO_2131 (O_2131,N_19984,N_19897);
and UO_2132 (O_2132,N_19973,N_19791);
nor UO_2133 (O_2133,N_19867,N_19983);
xnor UO_2134 (O_2134,N_19888,N_19874);
and UO_2135 (O_2135,N_19846,N_19873);
nand UO_2136 (O_2136,N_19911,N_19980);
nand UO_2137 (O_2137,N_19944,N_19830);
or UO_2138 (O_2138,N_19868,N_19920);
or UO_2139 (O_2139,N_19908,N_19878);
nor UO_2140 (O_2140,N_19925,N_19904);
nand UO_2141 (O_2141,N_19915,N_19978);
xnor UO_2142 (O_2142,N_19874,N_19847);
or UO_2143 (O_2143,N_19968,N_19905);
nand UO_2144 (O_2144,N_19787,N_19963);
nor UO_2145 (O_2145,N_19846,N_19895);
xnor UO_2146 (O_2146,N_19841,N_19933);
or UO_2147 (O_2147,N_19947,N_19993);
and UO_2148 (O_2148,N_19757,N_19868);
nor UO_2149 (O_2149,N_19981,N_19975);
nand UO_2150 (O_2150,N_19832,N_19892);
nand UO_2151 (O_2151,N_19860,N_19965);
nand UO_2152 (O_2152,N_19875,N_19903);
nor UO_2153 (O_2153,N_19777,N_19864);
and UO_2154 (O_2154,N_19797,N_19892);
xnor UO_2155 (O_2155,N_19911,N_19912);
nor UO_2156 (O_2156,N_19935,N_19757);
nor UO_2157 (O_2157,N_19876,N_19783);
xor UO_2158 (O_2158,N_19891,N_19919);
nand UO_2159 (O_2159,N_19853,N_19849);
or UO_2160 (O_2160,N_19818,N_19939);
or UO_2161 (O_2161,N_19916,N_19960);
nor UO_2162 (O_2162,N_19796,N_19802);
and UO_2163 (O_2163,N_19825,N_19846);
nand UO_2164 (O_2164,N_19929,N_19950);
nand UO_2165 (O_2165,N_19891,N_19917);
xnor UO_2166 (O_2166,N_19766,N_19996);
or UO_2167 (O_2167,N_19968,N_19951);
nor UO_2168 (O_2168,N_19963,N_19770);
xor UO_2169 (O_2169,N_19921,N_19877);
nand UO_2170 (O_2170,N_19881,N_19956);
nand UO_2171 (O_2171,N_19933,N_19992);
or UO_2172 (O_2172,N_19911,N_19828);
and UO_2173 (O_2173,N_19937,N_19903);
nor UO_2174 (O_2174,N_19900,N_19875);
and UO_2175 (O_2175,N_19761,N_19942);
and UO_2176 (O_2176,N_19793,N_19947);
nor UO_2177 (O_2177,N_19886,N_19839);
nor UO_2178 (O_2178,N_19905,N_19894);
and UO_2179 (O_2179,N_19775,N_19959);
or UO_2180 (O_2180,N_19831,N_19955);
or UO_2181 (O_2181,N_19851,N_19786);
nand UO_2182 (O_2182,N_19980,N_19904);
or UO_2183 (O_2183,N_19786,N_19825);
xor UO_2184 (O_2184,N_19866,N_19750);
and UO_2185 (O_2185,N_19947,N_19753);
xnor UO_2186 (O_2186,N_19942,N_19931);
nand UO_2187 (O_2187,N_19815,N_19932);
nor UO_2188 (O_2188,N_19917,N_19990);
or UO_2189 (O_2189,N_19832,N_19786);
xnor UO_2190 (O_2190,N_19965,N_19757);
nor UO_2191 (O_2191,N_19972,N_19957);
nand UO_2192 (O_2192,N_19936,N_19776);
nand UO_2193 (O_2193,N_19992,N_19890);
nor UO_2194 (O_2194,N_19955,N_19752);
or UO_2195 (O_2195,N_19820,N_19787);
xnor UO_2196 (O_2196,N_19801,N_19788);
nand UO_2197 (O_2197,N_19868,N_19858);
and UO_2198 (O_2198,N_19817,N_19750);
or UO_2199 (O_2199,N_19805,N_19776);
and UO_2200 (O_2200,N_19905,N_19967);
nand UO_2201 (O_2201,N_19983,N_19949);
or UO_2202 (O_2202,N_19787,N_19802);
nand UO_2203 (O_2203,N_19924,N_19910);
and UO_2204 (O_2204,N_19809,N_19793);
nor UO_2205 (O_2205,N_19905,N_19921);
and UO_2206 (O_2206,N_19757,N_19892);
nor UO_2207 (O_2207,N_19761,N_19884);
or UO_2208 (O_2208,N_19853,N_19930);
and UO_2209 (O_2209,N_19925,N_19833);
nand UO_2210 (O_2210,N_19954,N_19992);
or UO_2211 (O_2211,N_19944,N_19780);
nor UO_2212 (O_2212,N_19970,N_19991);
nand UO_2213 (O_2213,N_19870,N_19898);
nor UO_2214 (O_2214,N_19873,N_19889);
xor UO_2215 (O_2215,N_19933,N_19858);
xor UO_2216 (O_2216,N_19963,N_19883);
nor UO_2217 (O_2217,N_19798,N_19942);
or UO_2218 (O_2218,N_19819,N_19937);
or UO_2219 (O_2219,N_19816,N_19781);
nor UO_2220 (O_2220,N_19903,N_19884);
nand UO_2221 (O_2221,N_19924,N_19761);
nand UO_2222 (O_2222,N_19890,N_19976);
and UO_2223 (O_2223,N_19803,N_19906);
xnor UO_2224 (O_2224,N_19951,N_19935);
nor UO_2225 (O_2225,N_19762,N_19953);
or UO_2226 (O_2226,N_19892,N_19913);
nand UO_2227 (O_2227,N_19898,N_19893);
nand UO_2228 (O_2228,N_19774,N_19760);
xor UO_2229 (O_2229,N_19887,N_19974);
xnor UO_2230 (O_2230,N_19860,N_19985);
xnor UO_2231 (O_2231,N_19962,N_19933);
or UO_2232 (O_2232,N_19889,N_19825);
xnor UO_2233 (O_2233,N_19906,N_19837);
or UO_2234 (O_2234,N_19841,N_19843);
xnor UO_2235 (O_2235,N_19993,N_19864);
nand UO_2236 (O_2236,N_19804,N_19856);
or UO_2237 (O_2237,N_19777,N_19883);
xnor UO_2238 (O_2238,N_19842,N_19955);
nor UO_2239 (O_2239,N_19797,N_19925);
xor UO_2240 (O_2240,N_19946,N_19864);
nand UO_2241 (O_2241,N_19967,N_19942);
or UO_2242 (O_2242,N_19838,N_19978);
and UO_2243 (O_2243,N_19892,N_19851);
and UO_2244 (O_2244,N_19839,N_19949);
xnor UO_2245 (O_2245,N_19900,N_19902);
nand UO_2246 (O_2246,N_19990,N_19899);
xnor UO_2247 (O_2247,N_19843,N_19861);
xor UO_2248 (O_2248,N_19872,N_19941);
xor UO_2249 (O_2249,N_19819,N_19780);
nor UO_2250 (O_2250,N_19791,N_19846);
xnor UO_2251 (O_2251,N_19785,N_19834);
and UO_2252 (O_2252,N_19982,N_19899);
and UO_2253 (O_2253,N_19956,N_19893);
nor UO_2254 (O_2254,N_19866,N_19862);
and UO_2255 (O_2255,N_19866,N_19983);
nand UO_2256 (O_2256,N_19939,N_19873);
nand UO_2257 (O_2257,N_19929,N_19889);
nand UO_2258 (O_2258,N_19845,N_19788);
or UO_2259 (O_2259,N_19930,N_19820);
or UO_2260 (O_2260,N_19886,N_19912);
xnor UO_2261 (O_2261,N_19761,N_19829);
xor UO_2262 (O_2262,N_19922,N_19991);
and UO_2263 (O_2263,N_19945,N_19864);
nor UO_2264 (O_2264,N_19754,N_19984);
nand UO_2265 (O_2265,N_19908,N_19989);
nand UO_2266 (O_2266,N_19986,N_19958);
nor UO_2267 (O_2267,N_19859,N_19978);
and UO_2268 (O_2268,N_19961,N_19854);
nand UO_2269 (O_2269,N_19906,N_19960);
xor UO_2270 (O_2270,N_19838,N_19861);
xnor UO_2271 (O_2271,N_19943,N_19786);
nor UO_2272 (O_2272,N_19831,N_19962);
nor UO_2273 (O_2273,N_19991,N_19920);
or UO_2274 (O_2274,N_19810,N_19921);
and UO_2275 (O_2275,N_19780,N_19998);
xnor UO_2276 (O_2276,N_19995,N_19797);
nand UO_2277 (O_2277,N_19846,N_19861);
nor UO_2278 (O_2278,N_19761,N_19982);
nor UO_2279 (O_2279,N_19983,N_19830);
nor UO_2280 (O_2280,N_19954,N_19786);
or UO_2281 (O_2281,N_19964,N_19981);
nand UO_2282 (O_2282,N_19905,N_19964);
or UO_2283 (O_2283,N_19985,N_19987);
xnor UO_2284 (O_2284,N_19885,N_19838);
or UO_2285 (O_2285,N_19861,N_19903);
xnor UO_2286 (O_2286,N_19957,N_19946);
nand UO_2287 (O_2287,N_19945,N_19950);
nand UO_2288 (O_2288,N_19901,N_19885);
or UO_2289 (O_2289,N_19992,N_19751);
nand UO_2290 (O_2290,N_19914,N_19863);
nand UO_2291 (O_2291,N_19812,N_19779);
nand UO_2292 (O_2292,N_19754,N_19824);
nor UO_2293 (O_2293,N_19958,N_19761);
xor UO_2294 (O_2294,N_19886,N_19870);
nand UO_2295 (O_2295,N_19795,N_19869);
nand UO_2296 (O_2296,N_19860,N_19997);
xor UO_2297 (O_2297,N_19796,N_19885);
nand UO_2298 (O_2298,N_19937,N_19859);
nand UO_2299 (O_2299,N_19798,N_19922);
or UO_2300 (O_2300,N_19856,N_19980);
xnor UO_2301 (O_2301,N_19806,N_19919);
and UO_2302 (O_2302,N_19985,N_19761);
nand UO_2303 (O_2303,N_19819,N_19935);
nand UO_2304 (O_2304,N_19865,N_19958);
nor UO_2305 (O_2305,N_19770,N_19904);
or UO_2306 (O_2306,N_19773,N_19977);
nor UO_2307 (O_2307,N_19791,N_19752);
and UO_2308 (O_2308,N_19778,N_19770);
xor UO_2309 (O_2309,N_19957,N_19931);
and UO_2310 (O_2310,N_19857,N_19962);
xor UO_2311 (O_2311,N_19908,N_19807);
or UO_2312 (O_2312,N_19989,N_19780);
nor UO_2313 (O_2313,N_19777,N_19948);
and UO_2314 (O_2314,N_19861,N_19971);
or UO_2315 (O_2315,N_19918,N_19924);
and UO_2316 (O_2316,N_19933,N_19838);
nand UO_2317 (O_2317,N_19971,N_19985);
xnor UO_2318 (O_2318,N_19832,N_19951);
xnor UO_2319 (O_2319,N_19951,N_19809);
nor UO_2320 (O_2320,N_19954,N_19910);
and UO_2321 (O_2321,N_19904,N_19952);
and UO_2322 (O_2322,N_19942,N_19787);
or UO_2323 (O_2323,N_19930,N_19829);
and UO_2324 (O_2324,N_19788,N_19775);
or UO_2325 (O_2325,N_19865,N_19878);
or UO_2326 (O_2326,N_19966,N_19992);
or UO_2327 (O_2327,N_19824,N_19866);
or UO_2328 (O_2328,N_19800,N_19912);
xnor UO_2329 (O_2329,N_19841,N_19840);
nor UO_2330 (O_2330,N_19882,N_19860);
nor UO_2331 (O_2331,N_19883,N_19856);
nand UO_2332 (O_2332,N_19990,N_19995);
or UO_2333 (O_2333,N_19769,N_19927);
and UO_2334 (O_2334,N_19843,N_19877);
or UO_2335 (O_2335,N_19841,N_19857);
xnor UO_2336 (O_2336,N_19910,N_19877);
nand UO_2337 (O_2337,N_19910,N_19942);
nor UO_2338 (O_2338,N_19798,N_19752);
xor UO_2339 (O_2339,N_19895,N_19992);
or UO_2340 (O_2340,N_19939,N_19782);
nor UO_2341 (O_2341,N_19900,N_19762);
xor UO_2342 (O_2342,N_19952,N_19948);
xor UO_2343 (O_2343,N_19919,N_19980);
and UO_2344 (O_2344,N_19969,N_19775);
nor UO_2345 (O_2345,N_19829,N_19811);
nand UO_2346 (O_2346,N_19876,N_19832);
and UO_2347 (O_2347,N_19807,N_19757);
nor UO_2348 (O_2348,N_19982,N_19789);
xor UO_2349 (O_2349,N_19774,N_19989);
xor UO_2350 (O_2350,N_19935,N_19929);
or UO_2351 (O_2351,N_19971,N_19819);
or UO_2352 (O_2352,N_19919,N_19935);
nor UO_2353 (O_2353,N_19917,N_19833);
and UO_2354 (O_2354,N_19868,N_19828);
xnor UO_2355 (O_2355,N_19892,N_19810);
nor UO_2356 (O_2356,N_19759,N_19946);
or UO_2357 (O_2357,N_19909,N_19847);
nand UO_2358 (O_2358,N_19882,N_19769);
nor UO_2359 (O_2359,N_19924,N_19952);
and UO_2360 (O_2360,N_19925,N_19921);
nand UO_2361 (O_2361,N_19982,N_19764);
nand UO_2362 (O_2362,N_19834,N_19751);
xnor UO_2363 (O_2363,N_19857,N_19837);
nand UO_2364 (O_2364,N_19835,N_19855);
and UO_2365 (O_2365,N_19872,N_19822);
nand UO_2366 (O_2366,N_19900,N_19763);
and UO_2367 (O_2367,N_19887,N_19877);
nor UO_2368 (O_2368,N_19994,N_19888);
or UO_2369 (O_2369,N_19895,N_19851);
and UO_2370 (O_2370,N_19944,N_19957);
and UO_2371 (O_2371,N_19984,N_19852);
xor UO_2372 (O_2372,N_19923,N_19874);
and UO_2373 (O_2373,N_19821,N_19931);
nor UO_2374 (O_2374,N_19951,N_19888);
or UO_2375 (O_2375,N_19947,N_19909);
nor UO_2376 (O_2376,N_19755,N_19952);
nand UO_2377 (O_2377,N_19843,N_19911);
or UO_2378 (O_2378,N_19844,N_19786);
xor UO_2379 (O_2379,N_19961,N_19939);
nor UO_2380 (O_2380,N_19957,N_19948);
or UO_2381 (O_2381,N_19832,N_19826);
nor UO_2382 (O_2382,N_19907,N_19954);
nand UO_2383 (O_2383,N_19958,N_19908);
xnor UO_2384 (O_2384,N_19943,N_19940);
nand UO_2385 (O_2385,N_19862,N_19948);
nor UO_2386 (O_2386,N_19911,N_19793);
nand UO_2387 (O_2387,N_19802,N_19970);
nor UO_2388 (O_2388,N_19879,N_19789);
nor UO_2389 (O_2389,N_19757,N_19990);
and UO_2390 (O_2390,N_19825,N_19768);
nor UO_2391 (O_2391,N_19838,N_19871);
xnor UO_2392 (O_2392,N_19987,N_19772);
nand UO_2393 (O_2393,N_19870,N_19855);
nor UO_2394 (O_2394,N_19894,N_19891);
nand UO_2395 (O_2395,N_19869,N_19990);
nor UO_2396 (O_2396,N_19839,N_19823);
and UO_2397 (O_2397,N_19789,N_19969);
xor UO_2398 (O_2398,N_19818,N_19784);
or UO_2399 (O_2399,N_19962,N_19793);
nand UO_2400 (O_2400,N_19797,N_19821);
nand UO_2401 (O_2401,N_19913,N_19884);
or UO_2402 (O_2402,N_19865,N_19957);
nor UO_2403 (O_2403,N_19865,N_19810);
xor UO_2404 (O_2404,N_19805,N_19957);
or UO_2405 (O_2405,N_19933,N_19968);
nand UO_2406 (O_2406,N_19757,N_19846);
nor UO_2407 (O_2407,N_19810,N_19988);
xnor UO_2408 (O_2408,N_19876,N_19885);
or UO_2409 (O_2409,N_19771,N_19872);
or UO_2410 (O_2410,N_19878,N_19972);
and UO_2411 (O_2411,N_19825,N_19975);
nor UO_2412 (O_2412,N_19803,N_19944);
and UO_2413 (O_2413,N_19966,N_19844);
or UO_2414 (O_2414,N_19865,N_19797);
xnor UO_2415 (O_2415,N_19962,N_19907);
nand UO_2416 (O_2416,N_19839,N_19920);
nand UO_2417 (O_2417,N_19805,N_19775);
nor UO_2418 (O_2418,N_19844,N_19793);
xnor UO_2419 (O_2419,N_19829,N_19839);
or UO_2420 (O_2420,N_19762,N_19852);
nor UO_2421 (O_2421,N_19866,N_19925);
or UO_2422 (O_2422,N_19961,N_19997);
nor UO_2423 (O_2423,N_19767,N_19959);
xnor UO_2424 (O_2424,N_19792,N_19809);
or UO_2425 (O_2425,N_19998,N_19797);
nand UO_2426 (O_2426,N_19790,N_19991);
and UO_2427 (O_2427,N_19842,N_19865);
and UO_2428 (O_2428,N_19770,N_19761);
xor UO_2429 (O_2429,N_19998,N_19874);
nand UO_2430 (O_2430,N_19956,N_19844);
nor UO_2431 (O_2431,N_19924,N_19968);
nand UO_2432 (O_2432,N_19776,N_19949);
nand UO_2433 (O_2433,N_19812,N_19817);
nand UO_2434 (O_2434,N_19931,N_19991);
nand UO_2435 (O_2435,N_19900,N_19977);
nor UO_2436 (O_2436,N_19765,N_19846);
nor UO_2437 (O_2437,N_19984,N_19811);
nand UO_2438 (O_2438,N_19850,N_19987);
nand UO_2439 (O_2439,N_19817,N_19800);
nor UO_2440 (O_2440,N_19993,N_19765);
and UO_2441 (O_2441,N_19780,N_19763);
or UO_2442 (O_2442,N_19831,N_19786);
or UO_2443 (O_2443,N_19942,N_19979);
nor UO_2444 (O_2444,N_19764,N_19877);
and UO_2445 (O_2445,N_19856,N_19782);
or UO_2446 (O_2446,N_19930,N_19792);
xnor UO_2447 (O_2447,N_19982,N_19892);
or UO_2448 (O_2448,N_19817,N_19821);
or UO_2449 (O_2449,N_19992,N_19980);
nor UO_2450 (O_2450,N_19873,N_19841);
nand UO_2451 (O_2451,N_19985,N_19981);
and UO_2452 (O_2452,N_19782,N_19857);
xor UO_2453 (O_2453,N_19854,N_19768);
or UO_2454 (O_2454,N_19848,N_19992);
nor UO_2455 (O_2455,N_19918,N_19996);
xor UO_2456 (O_2456,N_19974,N_19965);
xnor UO_2457 (O_2457,N_19767,N_19848);
and UO_2458 (O_2458,N_19949,N_19821);
xor UO_2459 (O_2459,N_19842,N_19946);
nor UO_2460 (O_2460,N_19908,N_19787);
xnor UO_2461 (O_2461,N_19901,N_19861);
or UO_2462 (O_2462,N_19902,N_19879);
xnor UO_2463 (O_2463,N_19951,N_19750);
and UO_2464 (O_2464,N_19864,N_19811);
nand UO_2465 (O_2465,N_19887,N_19892);
nor UO_2466 (O_2466,N_19911,N_19851);
nand UO_2467 (O_2467,N_19981,N_19831);
nor UO_2468 (O_2468,N_19812,N_19866);
xor UO_2469 (O_2469,N_19771,N_19956);
xor UO_2470 (O_2470,N_19925,N_19827);
nand UO_2471 (O_2471,N_19902,N_19969);
and UO_2472 (O_2472,N_19853,N_19861);
and UO_2473 (O_2473,N_19982,N_19874);
nor UO_2474 (O_2474,N_19975,N_19764);
and UO_2475 (O_2475,N_19752,N_19779);
or UO_2476 (O_2476,N_19756,N_19878);
nor UO_2477 (O_2477,N_19920,N_19838);
xnor UO_2478 (O_2478,N_19893,N_19836);
nand UO_2479 (O_2479,N_19892,N_19973);
xor UO_2480 (O_2480,N_19891,N_19790);
or UO_2481 (O_2481,N_19956,N_19872);
and UO_2482 (O_2482,N_19970,N_19984);
nand UO_2483 (O_2483,N_19797,N_19926);
xnor UO_2484 (O_2484,N_19907,N_19841);
nand UO_2485 (O_2485,N_19950,N_19874);
nand UO_2486 (O_2486,N_19844,N_19987);
xor UO_2487 (O_2487,N_19894,N_19974);
nor UO_2488 (O_2488,N_19934,N_19868);
nand UO_2489 (O_2489,N_19929,N_19981);
xnor UO_2490 (O_2490,N_19913,N_19943);
nor UO_2491 (O_2491,N_19862,N_19880);
nor UO_2492 (O_2492,N_19956,N_19988);
nor UO_2493 (O_2493,N_19754,N_19790);
nor UO_2494 (O_2494,N_19888,N_19964);
xnor UO_2495 (O_2495,N_19809,N_19992);
or UO_2496 (O_2496,N_19782,N_19771);
and UO_2497 (O_2497,N_19999,N_19934);
xnor UO_2498 (O_2498,N_19905,N_19970);
nor UO_2499 (O_2499,N_19820,N_19850);
endmodule