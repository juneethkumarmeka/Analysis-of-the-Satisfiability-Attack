module basic_1500_15000_2000_3_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10004,N_10005,N_10006,N_10007,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10035,N_10036,N_10037,N_10043,N_10044,N_10045,N_10046,N_10047,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10059,N_10060,N_10061,N_10062,N_10065,N_10067,N_10068,N_10070,N_10071,N_10072,N_10074,N_10075,N_10076,N_10079,N_10080,N_10082,N_10084,N_10085,N_10086,N_10087,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10097,N_10098,N_10099,N_10100,N_10102,N_10103,N_10104,N_10105,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10116,N_10117,N_10118,N_10120,N_10121,N_10122,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10146,N_10147,N_10148,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10159,N_10160,N_10162,N_10163,N_10164,N_10166,N_10167,N_10168,N_10171,N_10172,N_10173,N_10174,N_10175,N_10177,N_10178,N_10180,N_10182,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10193,N_10194,N_10196,N_10197,N_10198,N_10199,N_10201,N_10202,N_10204,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10231,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10242,N_10243,N_10244,N_10245,N_10246,N_10248,N_10249,N_10250,N_10251,N_10252,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10277,N_10279,N_10280,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10291,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10301,N_10302,N_10304,N_10305,N_10306,N_10308,N_10309,N_10310,N_10311,N_10313,N_10314,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10332,N_10333,N_10334,N_10335,N_10337,N_10338,N_10339,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10360,N_10362,N_10364,N_10365,N_10366,N_10367,N_10368,N_10370,N_10372,N_10374,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10394,N_10395,N_10396,N_10397,N_10399,N_10400,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10423,N_10424,N_10425,N_10426,N_10427,N_10429,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10438,N_10439,N_10441,N_10442,N_10443,N_10444,N_10446,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10460,N_10462,N_10463,N_10465,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10478,N_10479,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10502,N_10503,N_10506,N_10507,N_10508,N_10509,N_10512,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10617,N_10619,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10634,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10654,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10669,N_10670,N_10671,N_10672,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10697,N_10698,N_10699,N_10700,N_10702,N_10703,N_10704,N_10705,N_10706,N_10708,N_10709,N_10710,N_10711,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10749,N_10750,N_10751,N_10752,N_10754,N_10756,N_10758,N_10759,N_10760,N_10761,N_10762,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10773,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10785,N_10786,N_10788,N_10789,N_10790,N_10791,N_10792,N_10795,N_10796,N_10798,N_10799,N_10801,N_10802,N_10803,N_10805,N_10806,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10819,N_10821,N_10822,N_10824,N_10825,N_10826,N_10827,N_10828,N_10831,N_10832,N_10833,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10869,N_10873,N_10874,N_10875,N_10876,N_10877,N_10880,N_10881,N_10882,N_10884,N_10885,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10899,N_10900,N_10902,N_10903,N_10904,N_10905,N_10907,N_10909,N_10910,N_10911,N_10913,N_10914,N_10915,N_10917,N_10918,N_10919,N_10920,N_10921,N_10924,N_10925,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10935,N_10937,N_10938,N_10939,N_10940,N_10941,N_10944,N_10946,N_10948,N_10950,N_10951,N_10952,N_10954,N_10955,N_10956,N_10957,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10976,N_10977,N_10978,N_10979,N_10980,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10990,N_10991,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11009,N_11011,N_11013,N_11014,N_11015,N_11016,N_11018,N_11019,N_11022,N_11023,N_11024,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11033,N_11035,N_11036,N_11037,N_11038,N_11040,N_11041,N_11044,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11068,N_11069,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11095,N_11096,N_11097,N_11098,N_11099,N_11101,N_11102,N_11103,N_11105,N_11106,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11118,N_11119,N_11120,N_11121,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11150,N_11151,N_11152,N_11153,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11162,N_11163,N_11164,N_11165,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11175,N_11176,N_11178,N_11179,N_11180,N_11181,N_11182,N_11184,N_11185,N_11186,N_11187,N_11188,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11212,N_11213,N_11214,N_11215,N_11216,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11245,N_11247,N_11248,N_11250,N_11253,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11265,N_11266,N_11267,N_11269,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11288,N_11289,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11321,N_11323,N_11324,N_11325,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11362,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11388,N_11389,N_11390,N_11391,N_11392,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11401,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11434,N_11435,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11456,N_11457,N_11459,N_11460,N_11461,N_11462,N_11464,N_11465,N_11466,N_11467,N_11469,N_11470,N_11471,N_11472,N_11473,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11484,N_11485,N_11488,N_11492,N_11493,N_11494,N_11496,N_11497,N_11498,N_11500,N_11501,N_11502,N_11503,N_11504,N_11506,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11521,N_11523,N_11524,N_11526,N_11527,N_11528,N_11529,N_11530,N_11532,N_11533,N_11534,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11545,N_11546,N_11547,N_11548,N_11549,N_11551,N_11554,N_11556,N_11557,N_11558,N_11559,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11579,N_11580,N_11581,N_11583,N_11584,N_11585,N_11587,N_11588,N_11590,N_11591,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11635,N_11636,N_11637,N_11638,N_11639,N_11641,N_11642,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11656,N_11657,N_11659,N_11660,N_11661,N_11663,N_11664,N_11666,N_11667,N_11668,N_11669,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11689,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11708,N_11710,N_11711,N_11712,N_11714,N_11716,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11734,N_11735,N_11736,N_11737,N_11738,N_11741,N_11742,N_11743,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11758,N_11759,N_11760,N_11761,N_11763,N_11764,N_11767,N_11768,N_11769,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11807,N_11808,N_11811,N_11812,N_11813,N_11815,N_11816,N_11817,N_11820,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11854,N_11855,N_11857,N_11858,N_11861,N_11862,N_11863,N_11864,N_11865,N_11867,N_11870,N_11872,N_11873,N_11874,N_11875,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11907,N_11909,N_11911,N_11912,N_11914,N_11915,N_11917,N_11919,N_11922,N_11923,N_11924,N_11925,N_11926,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11938,N_11939,N_11940,N_11942,N_11943,N_11944,N_11945,N_11946,N_11948,N_11949,N_11950,N_11952,N_11953,N_11954,N_11956,N_11957,N_11959,N_11961,N_11962,N_11963,N_11964,N_11966,N_11967,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11976,N_11977,N_11978,N_11979,N_11981,N_11983,N_11984,N_11985,N_11986,N_11988,N_11989,N_11990,N_11991,N_11993,N_11994,N_11995,N_11997,N_11998,N_11999,N_12000,N_12002,N_12003,N_12004,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12015,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12037,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12073,N_12074,N_12075,N_12076,N_12077,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12092,N_12093,N_12094,N_12096,N_12097,N_12098,N_12099,N_12101,N_12102,N_12103,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12122,N_12123,N_12124,N_12127,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12144,N_12145,N_12148,N_12149,N_12151,N_12153,N_12154,N_12155,N_12156,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12168,N_12169,N_12170,N_12172,N_12173,N_12174,N_12176,N_12177,N_12180,N_12181,N_12183,N_12184,N_12185,N_12186,N_12188,N_12189,N_12190,N_12191,N_12192,N_12194,N_12195,N_12196,N_12197,N_12198,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12210,N_12211,N_12212,N_12213,N_12214,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12228,N_12229,N_12230,N_12231,N_12233,N_12234,N_12235,N_12238,N_12239,N_12240,N_12243,N_12244,N_12245,N_12247,N_12248,N_12249,N_12250,N_12252,N_12253,N_12255,N_12257,N_12258,N_12259,N_12260,N_12262,N_12263,N_12265,N_12267,N_12268,N_12269,N_12271,N_12272,N_12275,N_12276,N_12278,N_12279,N_12281,N_12283,N_12284,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12293,N_12294,N_12295,N_12298,N_12299,N_12300,N_12301,N_12302,N_12305,N_12306,N_12307,N_12308,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12317,N_12318,N_12319,N_12320,N_12321,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12364,N_12365,N_12366,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12377,N_12378,N_12379,N_12380,N_12381,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12391,N_12392,N_12394,N_12395,N_12396,N_12397,N_12399,N_12400,N_12402,N_12404,N_12405,N_12406,N_12407,N_12409,N_12410,N_12411,N_12412,N_12413,N_12415,N_12419,N_12421,N_12422,N_12423,N_12424,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12449,N_12450,N_12451,N_12452,N_12453,N_12455,N_12456,N_12457,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12481,N_12482,N_12483,N_12484,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12494,N_12495,N_12496,N_12498,N_12499,N_12500,N_12502,N_12503,N_12504,N_12506,N_12507,N_12510,N_12511,N_12512,N_12513,N_12514,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12536,N_12537,N_12538,N_12539,N_12540,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12550,N_12551,N_12552,N_12554,N_12555,N_12556,N_12557,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12568,N_12569,N_12570,N_12572,N_12573,N_12574,N_12575,N_12577,N_12578,N_12579,N_12583,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12594,N_12595,N_12596,N_12598,N_12599,N_12603,N_12604,N_12605,N_12606,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12638,N_12639,N_12641,N_12643,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12656,N_12657,N_12658,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12668,N_12669,N_12670,N_12671,N_12672,N_12674,N_12675,N_12676,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12693,N_12694,N_12695,N_12696,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12706,N_12707,N_12708,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12737,N_12738,N_12739,N_12740,N_12741,N_12744,N_12745,N_12746,N_12747,N_12748,N_12750,N_12751,N_12752,N_12755,N_12756,N_12758,N_12760,N_12761,N_12762,N_12764,N_12765,N_12767,N_12768,N_12769,N_12771,N_12772,N_12773,N_12774,N_12777,N_12778,N_12779,N_12781,N_12782,N_12783,N_12784,N_12786,N_12787,N_12788,N_12789,N_12790,N_12792,N_12793,N_12794,N_12795,N_12796,N_12800,N_12801,N_12803,N_12804,N_12805,N_12806,N_12808,N_12809,N_12811,N_12812,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12822,N_12823,N_12824,N_12827,N_12828,N_12829,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12861,N_12862,N_12863,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12897,N_12898,N_12901,N_12902,N_12903,N_12904,N_12906,N_12907,N_12909,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12918,N_12920,N_12921,N_12922,N_12924,N_12926,N_12927,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12940,N_12941,N_12942,N_12944,N_12946,N_12947,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12987,N_12988,N_12989,N_12992,N_12993,N_12995,N_12997,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13023,N_13024,N_13025,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13047,N_13048,N_13049,N_13050,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13062,N_13063,N_13064,N_13068,N_13069,N_13070,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13084,N_13085,N_13086,N_13088,N_13090,N_13091,N_13093,N_13094,N_13095,N_13097,N_13098,N_13099,N_13100,N_13101,N_13104,N_13105,N_13106,N_13107,N_13109,N_13110,N_13111,N_13113,N_13114,N_13115,N_13116,N_13119,N_13120,N_13122,N_13123,N_13124,N_13125,N_13127,N_13128,N_13129,N_13130,N_13131,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13141,N_13142,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13165,N_13166,N_13168,N_13169,N_13170,N_13172,N_13173,N_13175,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13227,N_13228,N_13229,N_13230,N_13232,N_13233,N_13234,N_13235,N_13236,N_13238,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13269,N_13271,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13284,N_13286,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13298,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13311,N_13314,N_13315,N_13319,N_13320,N_13322,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13332,N_13333,N_13335,N_13336,N_13337,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13347,N_13348,N_13349,N_13350,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13372,N_13373,N_13374,N_13375,N_13377,N_13378,N_13379,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13401,N_13402,N_13403,N_13406,N_13407,N_13409,N_13410,N_13411,N_13412,N_13414,N_13416,N_13417,N_13418,N_13419,N_13420,N_13422,N_13423,N_13425,N_13426,N_13427,N_13428,N_13430,N_13431,N_13432,N_13434,N_13436,N_13438,N_13439,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13457,N_13458,N_13459,N_13460,N_13461,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13476,N_13477,N_13478,N_13479,N_13481,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13490,N_13492,N_13494,N_13496,N_13498,N_13500,N_13501,N_13503,N_13504,N_13505,N_13507,N_13508,N_13511,N_13513,N_13514,N_13515,N_13518,N_13519,N_13520,N_13521,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13535,N_13536,N_13537,N_13538,N_13540,N_13541,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13552,N_13553,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13600,N_13601,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13612,N_13613,N_13614,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13623,N_13624,N_13626,N_13627,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13637,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13648,N_13651,N_13652,N_13653,N_13654,N_13655,N_13657,N_13658,N_13659,N_13660,N_13662,N_13663,N_13665,N_13666,N_13667,N_13669,N_13670,N_13671,N_13672,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13684,N_13685,N_13686,N_13687,N_13688,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13711,N_13712,N_13714,N_13715,N_13717,N_13720,N_13722,N_13723,N_13724,N_13726,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13735,N_13736,N_13737,N_13738,N_13739,N_13741,N_13742,N_13743,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13760,N_13761,N_13764,N_13768,N_13770,N_13771,N_13772,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13813,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13831,N_13832,N_13833,N_13834,N_13836,N_13837,N_13838,N_13839,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13848,N_13849,N_13851,N_13852,N_13853,N_13854,N_13856,N_13857,N_13858,N_13859,N_13860,N_13862,N_13863,N_13865,N_13866,N_13867,N_13870,N_13871,N_13873,N_13874,N_13875,N_13876,N_13877,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13889,N_13890,N_13891,N_13892,N_13894,N_13895,N_13896,N_13897,N_13898,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13921,N_13922,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13931,N_13934,N_13935,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13953,N_13954,N_13956,N_13957,N_13958,N_13959,N_13961,N_13963,N_13964,N_13966,N_13967,N_13968,N_13969,N_13971,N_13972,N_13974,N_13975,N_13976,N_13979,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13990,N_13991,N_13993,N_13994,N_13995,N_13996,N_13998,N_14001,N_14003,N_14004,N_14005,N_14006,N_14008,N_14009,N_14011,N_14013,N_14014,N_14015,N_14016,N_14017,N_14021,N_14022,N_14023,N_14024,N_14026,N_14027,N_14028,N_14031,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14049,N_14050,N_14051,N_14052,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14066,N_14067,N_14068,N_14069,N_14070,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14082,N_14083,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14107,N_14108,N_14109,N_14110,N_14112,N_14113,N_14114,N_14115,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14134,N_14135,N_14136,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14153,N_14154,N_14155,N_14156,N_14158,N_14159,N_14160,N_14161,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14192,N_14193,N_14194,N_14195,N_14196,N_14198,N_14199,N_14200,N_14202,N_14204,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14213,N_14214,N_14216,N_14217,N_14219,N_14220,N_14221,N_14222,N_14224,N_14226,N_14229,N_14230,N_14231,N_14232,N_14233,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14248,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14271,N_14272,N_14273,N_14274,N_14277,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14301,N_14302,N_14303,N_14304,N_14307,N_14308,N_14309,N_14310,N_14311,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14328,N_14329,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14353,N_14354,N_14356,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14371,N_14372,N_14373,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14383,N_14384,N_14387,N_14388,N_14389,N_14390,N_14392,N_14393,N_14394,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14406,N_14407,N_14408,N_14409,N_14411,N_14412,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14423,N_14425,N_14426,N_14429,N_14432,N_14433,N_14435,N_14436,N_14437,N_14438,N_14439,N_14441,N_14442,N_14443,N_14445,N_14446,N_14447,N_14448,N_14449,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14481,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14501,N_14502,N_14503,N_14504,N_14505,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14518,N_14519,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14545,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14557,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14578,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14591,N_14592,N_14593,N_14595,N_14596,N_14597,N_14598,N_14599,N_14601,N_14603,N_14604,N_14605,N_14606,N_14608,N_14609,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14627,N_14628,N_14630,N_14635,N_14636,N_14637,N_14638,N_14639,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14650,N_14652,N_14653,N_14654,N_14656,N_14657,N_14658,N_14659,N_14661,N_14662,N_14663,N_14664,N_14665,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14683,N_14684,N_14685,N_14687,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14696,N_14697,N_14698,N_14699,N_14700,N_14702,N_14703,N_14704,N_14705,N_14706,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14716,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14731,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14744,N_14745,N_14746,N_14749,N_14750,N_14754,N_14755,N_14756,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14776,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14789,N_14790,N_14797,N_14799,N_14800,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14816,N_14819,N_14820,N_14821,N_14822,N_14823,N_14825,N_14826,N_14827,N_14828,N_14830,N_14832,N_14833,N_14835,N_14836,N_14838,N_14839,N_14840,N_14841,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14853,N_14856,N_14858,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14872,N_14873,N_14874,N_14876,N_14877,N_14879,N_14880,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14917,N_14918,N_14919,N_14920,N_14922,N_14923,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14949,N_14950,N_14951,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14961,N_14962,N_14963,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14982,N_14983,N_14984,N_14987,N_14988,N_14989,N_14990,N_14993,N_14994,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_688,In_463);
nand U1 (N_1,In_482,In_848);
or U2 (N_2,In_424,In_669);
and U3 (N_3,In_1099,In_361);
nor U4 (N_4,In_1457,In_157);
nand U5 (N_5,In_770,In_1230);
nand U6 (N_6,In_1136,In_614);
nand U7 (N_7,In_694,In_931);
or U8 (N_8,In_1021,In_494);
and U9 (N_9,In_351,In_252);
nand U10 (N_10,In_970,In_550);
xor U11 (N_11,In_1226,In_263);
nor U12 (N_12,In_775,In_955);
nor U13 (N_13,In_484,In_1450);
or U14 (N_14,In_210,In_603);
nor U15 (N_15,In_1065,In_345);
nand U16 (N_16,In_1435,In_1075);
or U17 (N_17,In_872,In_947);
and U18 (N_18,In_328,In_212);
or U19 (N_19,In_1484,In_979);
nand U20 (N_20,In_428,In_734);
nand U21 (N_21,In_1453,In_867);
nor U22 (N_22,In_711,In_740);
xor U23 (N_23,In_1031,In_259);
xnor U24 (N_24,In_1024,In_1413);
xnor U25 (N_25,In_1258,In_1018);
xnor U26 (N_26,In_780,In_619);
or U27 (N_27,In_673,In_1236);
or U28 (N_28,In_1216,In_1157);
or U29 (N_29,In_445,In_1418);
and U30 (N_30,In_1164,In_1235);
and U31 (N_31,In_975,In_765);
nor U32 (N_32,In_1110,In_1320);
nor U33 (N_33,In_1125,In_1473);
and U34 (N_34,In_981,In_792);
and U35 (N_35,In_1370,In_1172);
and U36 (N_36,In_1141,In_919);
or U37 (N_37,In_826,In_1485);
and U38 (N_38,In_1026,In_1053);
and U39 (N_39,In_1385,In_1);
or U40 (N_40,In_962,In_1354);
nand U41 (N_41,In_670,In_1410);
or U42 (N_42,In_626,In_211);
or U43 (N_43,In_1249,In_987);
or U44 (N_44,In_1460,In_932);
nand U45 (N_45,In_1089,In_429);
nand U46 (N_46,In_983,In_108);
nor U47 (N_47,In_1198,In_870);
nand U48 (N_48,In_243,In_431);
or U49 (N_49,In_203,In_313);
or U50 (N_50,In_965,In_865);
and U51 (N_51,In_235,In_398);
nor U52 (N_52,In_0,In_73);
nor U53 (N_53,In_1306,In_337);
or U54 (N_54,In_1359,In_747);
nand U55 (N_55,In_578,In_1241);
nor U56 (N_56,In_258,In_391);
nor U57 (N_57,In_816,In_1002);
and U58 (N_58,In_717,In_541);
and U59 (N_59,In_735,In_974);
nor U60 (N_60,In_415,In_331);
nor U61 (N_61,In_908,In_878);
or U62 (N_62,In_94,In_293);
or U63 (N_63,In_547,In_1308);
and U64 (N_64,In_98,In_1000);
and U65 (N_65,In_1455,In_275);
or U66 (N_66,In_1232,In_3);
nand U67 (N_67,In_27,In_15);
nand U68 (N_68,In_394,In_527);
nand U69 (N_69,In_715,In_503);
and U70 (N_70,In_774,In_1068);
and U71 (N_71,In_1301,In_411);
nor U72 (N_72,In_265,In_404);
and U73 (N_73,In_399,In_922);
nor U74 (N_74,In_400,In_490);
nor U75 (N_75,In_612,In_1420);
and U76 (N_76,In_950,In_447);
nor U77 (N_77,In_1471,In_1046);
xor U78 (N_78,In_850,In_209);
nor U79 (N_79,In_1076,In_1293);
nand U80 (N_80,In_1206,In_403);
or U81 (N_81,In_1212,In_1185);
or U82 (N_82,In_1144,In_602);
or U83 (N_83,In_942,In_841);
nand U84 (N_84,In_315,In_558);
or U85 (N_85,In_165,In_880);
nor U86 (N_86,In_1456,In_727);
and U87 (N_87,In_902,In_710);
nor U88 (N_88,In_376,In_1154);
and U89 (N_89,In_1339,In_1478);
nand U90 (N_90,In_723,In_167);
nor U91 (N_91,In_191,In_894);
nand U92 (N_92,In_1085,In_1279);
xor U93 (N_93,In_640,In_661);
xnor U94 (N_94,In_1131,In_250);
and U95 (N_95,In_1280,In_998);
or U96 (N_96,In_758,In_319);
or U97 (N_97,In_982,In_247);
or U98 (N_98,In_1094,In_589);
nor U99 (N_99,In_1446,In_750);
xnor U100 (N_100,In_722,In_481);
or U101 (N_101,In_59,In_956);
or U102 (N_102,In_425,In_888);
or U103 (N_103,In_468,In_1174);
nor U104 (N_104,In_889,In_192);
xnor U105 (N_105,In_664,In_104);
or U106 (N_106,In_1401,In_512);
nor U107 (N_107,In_299,In_131);
nand U108 (N_108,In_1093,In_134);
and U109 (N_109,In_1461,In_1404);
xor U110 (N_110,In_1299,In_639);
xnor U111 (N_111,In_1133,In_976);
and U112 (N_112,In_628,In_56);
nand U113 (N_113,In_289,In_837);
nor U114 (N_114,In_1043,In_926);
nor U115 (N_115,In_1439,In_146);
and U116 (N_116,In_312,In_741);
nand U117 (N_117,In_1468,In_1272);
and U118 (N_118,In_1459,In_476);
or U119 (N_119,In_135,In_1149);
nand U120 (N_120,In_545,In_1440);
and U121 (N_121,In_1380,In_782);
nand U122 (N_122,In_1044,In_1143);
or U123 (N_123,In_433,In_129);
or U124 (N_124,In_559,In_799);
or U125 (N_125,In_137,In_563);
and U126 (N_126,In_1493,In_1487);
and U127 (N_127,In_480,In_1324);
nor U128 (N_128,In_968,In_552);
nor U129 (N_129,In_949,In_163);
or U130 (N_130,In_451,In_198);
or U131 (N_131,In_777,In_142);
nand U132 (N_132,In_95,In_1406);
nand U133 (N_133,In_1160,In_1016);
nor U134 (N_134,In_1346,In_1479);
nand U135 (N_135,In_18,In_1292);
xnor U136 (N_136,In_1195,In_276);
nor U137 (N_137,In_830,In_127);
and U138 (N_138,In_86,In_1186);
nor U139 (N_139,In_767,In_405);
or U140 (N_140,In_651,In_1445);
nand U141 (N_141,In_757,In_600);
or U142 (N_142,In_893,In_1289);
nand U143 (N_143,In_1282,In_158);
or U144 (N_144,In_102,In_491);
xor U145 (N_145,In_764,In_1390);
and U146 (N_146,In_455,In_829);
and U147 (N_147,In_1358,In_174);
nor U148 (N_148,In_254,In_1102);
and U149 (N_149,In_763,In_1426);
or U150 (N_150,In_730,In_787);
and U151 (N_151,In_1454,In_665);
nor U152 (N_152,In_1070,In_437);
xor U153 (N_153,In_492,In_1407);
or U154 (N_154,In_1134,In_1351);
nor U155 (N_155,In_631,In_803);
or U156 (N_156,In_1343,In_483);
and U157 (N_157,In_812,In_1364);
or U158 (N_158,In_154,In_1337);
and U159 (N_159,In_242,In_416);
nand U160 (N_160,In_720,In_918);
nand U161 (N_161,In_549,In_301);
or U162 (N_162,In_1317,In_150);
or U163 (N_163,In_1107,In_5);
nand U164 (N_164,In_946,In_1465);
or U165 (N_165,In_377,In_1111);
nor U166 (N_166,In_461,In_1414);
nor U167 (N_167,In_251,In_690);
nand U168 (N_168,In_151,In_283);
nor U169 (N_169,In_114,In_595);
nand U170 (N_170,In_566,In_1266);
nand U171 (N_171,In_1443,In_662);
and U172 (N_172,In_183,In_820);
or U173 (N_173,In_1312,In_540);
and U174 (N_174,In_1431,In_126);
nor U175 (N_175,In_85,In_897);
or U176 (N_176,In_180,In_284);
or U177 (N_177,In_393,In_1108);
nor U178 (N_178,In_853,In_100);
nor U179 (N_179,In_387,In_335);
and U180 (N_180,In_1088,In_362);
nand U181 (N_181,In_389,In_168);
nor U182 (N_182,In_1137,In_223);
and U183 (N_183,In_175,In_1492);
nand U184 (N_184,In_1051,In_65);
nor U185 (N_185,In_1348,In_267);
nand U186 (N_186,In_349,In_326);
nand U187 (N_187,In_10,In_1040);
and U188 (N_188,In_363,In_660);
nor U189 (N_189,In_34,In_995);
xor U190 (N_190,In_769,In_1234);
and U191 (N_191,In_1054,In_232);
nor U192 (N_192,In_33,In_1360);
or U193 (N_193,In_707,In_1091);
and U194 (N_194,In_920,In_1032);
nand U195 (N_195,In_683,In_218);
xnor U196 (N_196,In_1025,In_115);
xnor U197 (N_197,In_802,In_674);
and U198 (N_198,In_1036,In_610);
nand U199 (N_199,In_1434,In_1237);
xor U200 (N_200,In_253,In_1490);
xor U201 (N_201,In_1207,In_72);
nand U202 (N_202,In_493,In_702);
or U203 (N_203,In_588,In_1177);
nor U204 (N_204,In_324,In_1129);
or U205 (N_205,In_1081,In_1012);
nor U206 (N_206,In_350,In_147);
nor U207 (N_207,In_19,In_1098);
or U208 (N_208,In_295,In_1050);
or U209 (N_209,In_996,In_1260);
or U210 (N_210,In_698,In_1117);
nor U211 (N_211,In_1074,In_1495);
and U212 (N_212,In_910,In_9);
nand U213 (N_213,In_364,In_487);
nand U214 (N_214,In_497,In_439);
nor U215 (N_215,In_352,In_721);
nor U216 (N_216,In_675,In_518);
nor U217 (N_217,In_840,In_567);
nor U218 (N_218,In_1336,In_1329);
xnor U219 (N_219,In_1325,In_835);
nand U220 (N_220,In_945,In_1152);
or U221 (N_221,In_273,In_1092);
nand U222 (N_222,In_1436,In_1028);
or U223 (N_223,In_1486,In_347);
and U224 (N_224,In_1083,In_1256);
and U225 (N_225,In_231,In_1225);
nand U226 (N_226,In_66,In_1462);
or U227 (N_227,In_1061,In_1041);
nand U228 (N_228,In_48,In_1394);
or U229 (N_229,In_268,In_355);
nor U230 (N_230,In_245,In_96);
or U231 (N_231,In_1347,In_176);
or U232 (N_232,In_1427,In_169);
nor U233 (N_233,In_796,In_883);
or U234 (N_234,In_1417,In_781);
nor U235 (N_235,In_1135,In_1344);
or U236 (N_236,In_984,In_875);
or U237 (N_237,In_1449,In_903);
nand U238 (N_238,In_857,In_718);
and U239 (N_239,In_1295,In_1373);
nor U240 (N_240,In_386,In_729);
or U241 (N_241,In_544,In_440);
xor U242 (N_242,In_379,In_230);
nor U243 (N_243,In_1077,In_504);
and U244 (N_244,In_611,In_1384);
and U245 (N_245,In_1214,In_937);
or U246 (N_246,In_434,In_458);
nand U247 (N_247,In_1371,In_1227);
or U248 (N_248,In_1388,In_1464);
nor U249 (N_249,In_703,In_257);
nand U250 (N_250,In_580,In_1178);
nand U251 (N_251,In_555,In_456);
and U252 (N_252,In_112,In_1252);
xor U253 (N_253,In_1202,In_1333);
nand U254 (N_254,In_229,In_316);
or U255 (N_255,In_1156,In_1458);
nand U256 (N_256,In_83,In_553);
and U257 (N_257,In_1318,In_847);
nor U258 (N_258,In_291,In_473);
nor U259 (N_259,In_815,In_705);
or U260 (N_260,In_1381,In_973);
and U261 (N_261,In_496,In_153);
or U262 (N_262,In_739,In_264);
and U263 (N_263,In_1165,In_35);
nand U264 (N_264,In_606,In_219);
nand U265 (N_265,In_1416,In_761);
and U266 (N_266,In_145,In_82);
nand U267 (N_267,In_396,In_261);
or U268 (N_268,In_1176,In_392);
and U269 (N_269,In_625,In_475);
nand U270 (N_270,In_1375,In_1196);
nor U271 (N_271,In_599,In_332);
nor U272 (N_272,In_1356,In_113);
and U273 (N_273,In_986,In_296);
or U274 (N_274,In_938,In_725);
or U275 (N_275,In_24,In_686);
or U276 (N_276,In_712,In_262);
or U277 (N_277,In_583,In_372);
nand U278 (N_278,In_1047,In_1132);
xnor U279 (N_279,In_742,In_521);
nor U280 (N_280,In_709,In_28);
nand U281 (N_281,In_530,In_213);
and U282 (N_282,In_1030,In_861);
nand U283 (N_283,In_561,In_162);
nor U284 (N_284,In_408,In_1376);
or U285 (N_285,In_806,In_385);
and U286 (N_286,In_282,In_1438);
and U287 (N_287,In_568,In_322);
nand U288 (N_288,In_292,In_1275);
and U289 (N_289,In_980,In_409);
nor U290 (N_290,In_1319,In_724);
nand U291 (N_291,In_2,In_930);
or U292 (N_292,In_647,In_116);
or U293 (N_293,In_29,In_270);
nor U294 (N_294,In_557,In_240);
nor U295 (N_295,In_430,In_1367);
and U296 (N_296,In_911,In_474);
and U297 (N_297,In_333,In_106);
nor U298 (N_298,In_1153,In_401);
and U299 (N_299,In_498,In_1120);
or U300 (N_300,In_586,In_1330);
or U301 (N_301,In_1447,In_486);
nor U302 (N_302,In_336,In_1345);
or U303 (N_303,In_1210,In_832);
and U304 (N_304,In_676,In_423);
and U305 (N_305,In_277,In_1338);
and U306 (N_306,In_1498,In_943);
nor U307 (N_307,In_344,In_874);
nand U308 (N_308,In_810,In_8);
or U309 (N_309,In_1035,In_1341);
nor U310 (N_310,In_1173,In_141);
nor U311 (N_311,In_768,In_177);
xor U312 (N_312,In_1328,In_1130);
nand U313 (N_313,In_951,In_238);
and U314 (N_314,In_187,In_929);
or U315 (N_315,In_125,In_4);
or U316 (N_316,In_941,In_682);
and U317 (N_317,In_197,In_1208);
xor U318 (N_318,In_749,In_609);
or U319 (N_319,In_139,In_845);
nor U320 (N_320,In_1181,In_587);
or U321 (N_321,In_269,In_1281);
and U322 (N_322,In_1017,In_1073);
nand U323 (N_323,In_144,In_887);
and U324 (N_324,In_1205,In_1494);
or U325 (N_325,In_952,In_1403);
and U326 (N_326,In_1415,In_1169);
nor U327 (N_327,In_788,In_1184);
or U328 (N_328,In_744,In_1062);
or U329 (N_329,In_650,In_1190);
and U330 (N_330,In_890,In_1452);
nor U331 (N_331,In_77,In_924);
or U332 (N_332,In_1221,In_1441);
nor U333 (N_333,In_825,In_620);
xor U334 (N_334,In_824,In_1259);
or U335 (N_335,In_1162,In_1296);
nor U336 (N_336,In_1105,In_1386);
and U337 (N_337,In_68,In_321);
nand U338 (N_338,In_1362,In_828);
and U339 (N_339,In_26,In_1288);
or U340 (N_340,In_1103,In_1127);
nand U341 (N_341,In_1201,In_166);
nor U342 (N_342,In_1271,In_327);
nand U343 (N_343,In_833,In_38);
xnor U344 (N_344,In_330,In_260);
nor U345 (N_345,In_868,In_630);
nor U346 (N_346,In_1071,In_1145);
and U347 (N_347,In_1059,In_689);
xor U348 (N_348,In_1298,In_50);
or U349 (N_349,In_25,In_384);
nor U350 (N_350,In_1267,In_1264);
xor U351 (N_351,In_128,In_1104);
nand U352 (N_352,In_1211,In_813);
nor U353 (N_353,In_789,In_616);
or U354 (N_354,In_248,In_556);
nor U355 (N_355,In_1466,In_149);
xnor U356 (N_356,In_1392,In_1378);
nor U357 (N_357,In_907,In_186);
and U358 (N_358,In_161,In_576);
or U359 (N_359,In_1372,In_641);
nor U360 (N_360,In_452,In_879);
and U361 (N_361,In_20,In_1109);
xor U362 (N_362,In_1250,In_200);
nor U363 (N_363,In_708,In_1368);
nand U364 (N_364,In_236,In_1283);
nor U365 (N_365,In_933,In_1020);
and U366 (N_366,In_348,In_638);
nor U367 (N_367,In_613,In_726);
or U368 (N_368,In_1055,In_1286);
xnor U369 (N_369,In_234,In_52);
nand U370 (N_370,In_1049,In_648);
or U371 (N_371,In_237,In_790);
nor U372 (N_372,In_993,In_713);
and U373 (N_373,In_464,In_569);
nand U374 (N_374,In_807,In_1197);
and U375 (N_375,In_1161,In_778);
and U376 (N_376,In_1228,In_536);
or U377 (N_377,In_369,In_959);
and U378 (N_378,In_659,In_944);
and U379 (N_379,In_17,In_534);
or U380 (N_380,In_953,In_1090);
nand U381 (N_381,In_990,In_846);
and U382 (N_382,In_838,In_657);
nand U383 (N_383,In_16,In_821);
xor U384 (N_384,In_1331,In_1219);
nor U385 (N_385,In_1470,In_23);
and U386 (N_386,In_574,In_1095);
or U387 (N_387,In_743,In_290);
or U388 (N_388,In_671,In_368);
or U389 (N_389,In_1244,In_1251);
nand U390 (N_390,In_1008,In_71);
xor U391 (N_391,In_1277,In_784);
or U392 (N_392,In_804,In_90);
or U393 (N_393,In_1001,In_1009);
or U394 (N_394,In_1496,In_1480);
or U395 (N_395,In_143,In_654);
and U396 (N_396,In_577,In_1423);
nor U397 (N_397,In_560,In_967);
and U398 (N_398,In_1408,In_1019);
nand U399 (N_399,In_1126,In_1353);
nor U400 (N_400,In_539,In_1326);
and U401 (N_401,In_1223,In_877);
or U402 (N_402,In_40,In_817);
nor U403 (N_403,In_1419,In_1387);
or U404 (N_404,In_470,In_43);
nand U405 (N_405,In_999,In_1097);
or U406 (N_406,In_1276,In_642);
nand U407 (N_407,In_1316,In_760);
nor U408 (N_408,In_1138,In_1179);
nor U409 (N_409,In_1409,In_199);
nand U410 (N_410,In_1311,In_1263);
xnor U411 (N_411,In_658,In_905);
or U412 (N_412,In_1124,In_184);
and U413 (N_413,In_488,In_75);
and U414 (N_414,In_912,In_202);
and U415 (N_415,In_1285,In_1374);
nor U416 (N_416,In_548,In_1327);
xnor U417 (N_417,In_380,In_308);
or U418 (N_418,In_55,In_346);
nor U419 (N_419,In_1042,In_178);
nand U420 (N_420,In_225,In_1166);
or U421 (N_421,In_1082,In_340);
xor U422 (N_422,In_1483,In_1304);
nor U423 (N_423,In_341,In_1482);
xor U424 (N_424,In_594,In_582);
nor U425 (N_425,In_1233,In_214);
or U426 (N_426,In_573,In_914);
and U427 (N_427,In_1323,In_138);
xnor U428 (N_428,In_988,In_542);
nand U429 (N_429,In_382,In_649);
or U430 (N_430,In_1167,In_693);
or U431 (N_431,In_1163,In_805);
nand U432 (N_432,In_1052,In_605);
nand U433 (N_433,In_1060,In_762);
or U434 (N_434,In_367,In_1389);
xnor U435 (N_435,In_604,In_1158);
or U436 (N_436,In_511,In_1477);
nor U437 (N_437,In_448,In_1411);
and U438 (N_438,In_1332,In_418);
and U439 (N_439,In_14,In_1314);
nor U440 (N_440,In_844,In_593);
and U441 (N_441,In_274,In_1284);
nand U442 (N_442,In_338,In_966);
or U443 (N_443,In_691,In_656);
xnor U444 (N_444,In_1128,In_477);
or U445 (N_445,In_412,In_1302);
or U446 (N_446,In_280,In_304);
and U447 (N_447,In_895,In_1430);
nor U448 (N_448,In_1335,In_124);
or U449 (N_449,In_1412,In_195);
or U450 (N_450,In_132,In_695);
nand U451 (N_451,In_420,In_1405);
nor U452 (N_452,In_1334,In_343);
or U453 (N_453,In_543,In_701);
nand U454 (N_454,In_522,In_306);
nand U455 (N_455,In_1369,In_495);
nand U456 (N_456,In_1139,In_700);
or U457 (N_457,In_1361,In_501);
and U458 (N_458,In_255,In_1444);
nand U459 (N_459,In_61,In_1193);
nor U460 (N_460,In_901,In_836);
and U461 (N_461,In_92,In_533);
nor U462 (N_462,In_939,In_173);
nor U463 (N_463,In_519,In_748);
and U464 (N_464,In_1004,In_570);
nor U465 (N_465,In_467,In_672);
or U466 (N_466,In_913,In_731);
nand U467 (N_467,In_278,In_371);
and U468 (N_468,In_1180,In_45);
and U469 (N_469,In_1242,In_1116);
or U470 (N_470,In_320,In_1357);
nor U471 (N_471,In_581,In_852);
and U472 (N_472,In_1489,In_1432);
nor U473 (N_473,In_13,In_182);
and U474 (N_474,In_297,In_653);
and U475 (N_475,In_858,In_466);
nor U476 (N_476,In_964,In_514);
nand U477 (N_477,In_1122,In_1397);
or U478 (N_478,In_164,In_99);
or U479 (N_479,In_989,In_766);
and U480 (N_480,In_601,In_357);
and U481 (N_481,In_314,In_1194);
or U482 (N_482,In_866,In_130);
or U483 (N_483,In_892,In_1274);
xor U484 (N_484,In_752,In_1086);
nor U485 (N_485,In_507,In_1310);
and U486 (N_486,In_1476,In_39);
nand U487 (N_487,In_1290,In_562);
xor U488 (N_488,In_1048,In_224);
nor U489 (N_489,In_121,In_107);
or U490 (N_490,In_51,In_873);
xnor U491 (N_491,In_190,In_1248);
and U492 (N_492,In_655,In_37);
or U493 (N_493,In_118,In_886);
nor U494 (N_494,In_472,In_607);
or U495 (N_495,In_793,In_524);
nand U496 (N_496,In_454,In_963);
and U497 (N_497,In_1366,In_442);
and U498 (N_498,In_681,In_1005);
nor U499 (N_499,In_1350,In_948);
nand U500 (N_500,In_148,In_909);
or U501 (N_501,In_302,In_772);
nand U502 (N_502,In_1213,In_1084);
nor U503 (N_503,In_697,In_916);
or U504 (N_504,In_728,In_1087);
and U505 (N_505,In_822,In_860);
nor U506 (N_506,In_869,In_426);
nand U507 (N_507,In_1261,In_215);
nor U508 (N_508,In_422,In_117);
xnor U509 (N_509,In_756,In_171);
nand U510 (N_510,In_921,In_1014);
xor U511 (N_511,In_809,In_310);
nor U512 (N_512,In_11,In_239);
or U513 (N_513,In_678,In_1402);
or U514 (N_514,In_786,In_485);
xor U515 (N_515,In_1015,In_307);
nand U516 (N_516,In_1203,In_1399);
or U517 (N_517,In_531,In_1396);
or U518 (N_518,In_771,In_57);
nand U519 (N_519,In_1475,In_621);
or U520 (N_520,In_1421,In_864);
nor U521 (N_521,In_1146,In_839);
and U522 (N_522,In_871,In_1113);
or U523 (N_523,In_551,In_823);
and U524 (N_524,In_1159,In_111);
or U525 (N_525,In_479,In_358);
nor U526 (N_526,In_1474,In_221);
and U527 (N_527,In_366,In_854);
or U528 (N_528,In_645,In_1270);
and U529 (N_529,In_21,In_70);
nor U530 (N_530,In_719,In_617);
and U531 (N_531,In_42,In_1428);
nand U532 (N_532,In_436,In_294);
nor U533 (N_533,In_204,In_1262);
nand U534 (N_534,In_1463,In_193);
nor U535 (N_535,In_733,In_413);
or U536 (N_536,In_46,In_891);
or U537 (N_537,In_91,In_155);
and U538 (N_538,In_978,In_375);
or U539 (N_539,In_1321,In_585);
xnor U540 (N_540,In_1151,In_1119);
nor U541 (N_541,In_1303,In_502);
nand U542 (N_542,In_1171,In_1497);
nand U543 (N_543,In_365,In_755);
or U544 (N_544,In_1045,In_1499);
and U545 (N_545,In_590,In_592);
or U546 (N_546,In_1010,In_885);
or U547 (N_547,In_1100,In_81);
and U548 (N_548,In_666,In_677);
and U549 (N_549,In_1246,In_1437);
or U550 (N_550,In_58,In_571);
nor U551 (N_551,In_1297,In_615);
nor U552 (N_552,In_1287,In_1123);
nand U553 (N_553,In_863,In_31);
and U554 (N_554,In_935,In_1322);
nand U555 (N_555,In_751,In_505);
or U556 (N_556,In_370,In_529);
xnor U557 (N_557,In_882,In_881);
or U558 (N_558,In_220,In_62);
nand U559 (N_559,In_706,In_181);
nand U560 (N_560,In_795,In_309);
or U561 (N_561,In_643,In_1217);
nand U562 (N_562,In_1039,In_994);
xnor U563 (N_563,In_633,In_776);
nor U564 (N_564,In_407,In_714);
xnor U565 (N_565,In_1467,In_1175);
and U566 (N_566,In_281,In_856);
nand U567 (N_567,In_110,In_194);
nor U568 (N_568,In_644,In_1058);
and U569 (N_569,In_584,In_1269);
and U570 (N_570,In_859,In_272);
or U571 (N_571,In_754,In_287);
nand U572 (N_572,In_1142,In_1222);
nand U573 (N_573,In_597,In_940);
nor U574 (N_574,In_699,In_12);
or U575 (N_575,In_342,In_1307);
nor U576 (N_576,In_119,In_1429);
or U577 (N_577,In_1355,In_736);
nand U578 (N_578,In_624,In_936);
nor U579 (N_579,In_546,In_323);
or U580 (N_580,In_508,In_1300);
and U581 (N_581,In_876,In_1022);
nand U582 (N_582,In_1315,In_381);
nand U583 (N_583,In_915,In_54);
or U584 (N_584,In_1191,In_564);
xor U585 (N_585,In_1121,In_47);
and U586 (N_586,In_318,In_53);
and U587 (N_587,In_843,In_152);
and U588 (N_588,In_185,In_1140);
xor U589 (N_589,In_378,In_667);
or U590 (N_590,In_441,In_450);
nor U591 (N_591,In_244,In_233);
xor U592 (N_592,In_1273,In_923);
or U593 (N_593,In_985,In_1192);
nor U594 (N_594,In_1189,In_1265);
and U595 (N_595,In_421,In_1182);
or U596 (N_596,In_1200,In_460);
nor U597 (N_597,In_207,In_972);
and U598 (N_598,In_598,In_1379);
or U599 (N_599,In_1448,In_1029);
and U600 (N_600,In_596,In_1033);
nand U601 (N_601,In_123,In_329);
nand U602 (N_602,In_1398,In_453);
or U603 (N_603,In_419,In_1106);
and U604 (N_604,In_800,In_286);
xor U605 (N_605,In_1363,In_692);
and U606 (N_606,In_977,In_1188);
or U607 (N_607,In_1342,In_1255);
nand U608 (N_608,In_773,In_69);
nand U609 (N_609,In_216,In_256);
xnor U610 (N_610,In_627,In_1247);
and U611 (N_611,In_925,In_1215);
nand U612 (N_612,In_36,In_438);
xor U613 (N_613,In_759,In_1101);
nor U614 (N_614,In_1425,In_489);
or U615 (N_615,In_78,In_1257);
nand U616 (N_616,In_136,In_851);
xor U617 (N_617,In_74,In_303);
nor U618 (N_618,In_779,In_1003);
and U619 (N_619,In_811,In_285);
nor U620 (N_620,In_60,In_1078);
xor U621 (N_621,In_298,In_1023);
nor U622 (N_622,In_500,In_1383);
or U623 (N_623,In_928,In_904);
or U624 (N_624,In_160,In_575);
or U625 (N_625,In_814,In_591);
xnor U626 (N_626,In_737,In_305);
xnor U627 (N_627,In_1294,In_359);
or U628 (N_628,In_87,In_971);
and U629 (N_629,In_652,In_696);
nor U630 (N_630,In_1067,In_1170);
nand U631 (N_631,In_1240,In_1063);
or U632 (N_632,In_30,In_510);
xor U633 (N_633,In_961,In_785);
or U634 (N_634,In_1155,In_196);
nor U635 (N_635,In_1291,In_927);
nand U636 (N_636,In_89,In_63);
and U637 (N_637,In_834,In_535);
nor U638 (N_638,In_226,In_334);
nor U639 (N_639,In_172,In_1072);
xor U640 (N_640,In_515,In_266);
and U641 (N_641,In_1209,In_1218);
nand U642 (N_642,In_1278,In_862);
nand U643 (N_643,In_105,In_646);
nand U644 (N_644,In_906,In_797);
or U645 (N_645,In_311,In_373);
nor U646 (N_646,In_738,In_808);
and U647 (N_647,In_509,In_156);
or U648 (N_648,In_801,In_1253);
xnor U649 (N_649,In_478,In_133);
nor U650 (N_650,In_954,In_960);
nor U651 (N_651,In_249,In_417);
xnor U652 (N_652,In_992,In_208);
or U653 (N_653,In_1118,In_1442);
and U654 (N_654,In_22,In_406);
xnor U655 (N_655,In_201,In_1006);
nor U656 (N_656,In_317,In_958);
xnor U657 (N_657,In_241,In_471);
xnor U658 (N_658,In_432,In_934);
nand U659 (N_659,In_1395,In_1056);
xor U660 (N_660,In_271,In_855);
and U661 (N_661,In_1268,In_791);
nor U662 (N_662,In_93,In_608);
or U663 (N_663,In_79,In_410);
nand U664 (N_664,In_88,In_680);
nand U665 (N_665,In_618,In_1433);
nand U666 (N_666,In_279,In_554);
and U667 (N_667,In_444,In_462);
nand U668 (N_668,In_1114,In_449);
and U669 (N_669,In_222,In_896);
nor U670 (N_670,In_339,In_537);
and U671 (N_671,In_1147,In_459);
nand U672 (N_672,In_1243,In_831);
nor U673 (N_673,In_991,In_374);
or U674 (N_674,In_189,In_179);
nor U675 (N_675,In_122,In_753);
or U676 (N_676,In_525,In_1340);
and U677 (N_677,In_506,In_1224);
or U678 (N_678,In_120,In_663);
nor U679 (N_679,In_383,In_1066);
or U680 (N_680,In_1382,In_1150);
nor U681 (N_681,In_360,In_44);
and U682 (N_682,In_746,In_1481);
and U683 (N_683,In_1013,In_1377);
xnor U684 (N_684,In_849,In_101);
and U685 (N_685,In_1365,In_356);
or U686 (N_686,In_395,In_109);
or U687 (N_687,In_1034,In_1027);
or U688 (N_688,In_1187,In_1011);
or U689 (N_689,In_103,In_1424);
nor U690 (N_690,In_67,In_1231);
nor U691 (N_691,In_1057,In_579);
nor U692 (N_692,In_41,In_469);
nand U693 (N_693,In_1391,In_353);
nor U694 (N_694,In_679,In_206);
nand U695 (N_695,In_1229,In_526);
or U696 (N_696,In_532,In_900);
or U697 (N_697,In_1096,In_499);
nor U698 (N_698,In_435,In_632);
nand U699 (N_699,In_623,In_1400);
nor U700 (N_700,In_32,In_513);
or U701 (N_701,In_159,In_217);
or U702 (N_702,In_898,In_629);
or U703 (N_703,In_300,In_1393);
and U704 (N_704,In_1422,In_246);
nand U705 (N_705,In_140,In_443);
nor U706 (N_706,In_1472,In_1168);
nand U707 (N_707,In_354,In_1309);
nor U708 (N_708,In_228,In_1112);
nand U709 (N_709,In_899,In_517);
nor U710 (N_710,In_1079,In_465);
nor U711 (N_711,In_637,In_80);
xor U712 (N_712,In_520,In_1469);
or U713 (N_713,In_97,In_1491);
and U714 (N_714,In_1220,In_538);
nand U715 (N_715,In_6,In_402);
and U716 (N_716,In_1254,In_818);
or U717 (N_717,In_997,In_798);
and U718 (N_718,In_1204,In_1183);
and U719 (N_719,In_783,In_957);
nand U720 (N_720,In_684,In_397);
nor U721 (N_721,In_1305,In_516);
or U722 (N_722,In_704,In_572);
or U723 (N_723,In_7,In_227);
and U724 (N_724,In_1245,In_49);
nand U725 (N_725,In_716,In_1080);
nor U726 (N_726,In_745,In_1069);
and U727 (N_727,In_1115,In_732);
xnor U728 (N_728,In_685,In_634);
nor U729 (N_729,In_668,In_687);
nand U730 (N_730,In_1037,In_1488);
or U731 (N_731,In_917,In_827);
nor U732 (N_732,In_288,In_1451);
or U733 (N_733,In_1239,In_427);
or U734 (N_734,In_622,In_842);
nor U735 (N_735,In_1313,In_794);
nor U736 (N_736,In_170,In_205);
xor U737 (N_737,In_1352,In_884);
nor U738 (N_738,In_523,In_388);
and U739 (N_739,In_1007,In_325);
and U740 (N_740,In_1199,In_84);
xnor U741 (N_741,In_414,In_390);
nor U742 (N_742,In_1038,In_635);
xnor U743 (N_743,In_457,In_636);
nand U744 (N_744,In_528,In_969);
and U745 (N_745,In_1238,In_64);
nor U746 (N_746,In_1349,In_1064);
and U747 (N_747,In_1148,In_76);
and U748 (N_748,In_819,In_565);
or U749 (N_749,In_446,In_188);
nand U750 (N_750,In_366,In_39);
and U751 (N_751,In_487,In_1355);
and U752 (N_752,In_860,In_1297);
nor U753 (N_753,In_1363,In_365);
and U754 (N_754,In_1245,In_1347);
xor U755 (N_755,In_1468,In_886);
or U756 (N_756,In_1352,In_577);
xor U757 (N_757,In_502,In_352);
nor U758 (N_758,In_500,In_752);
nor U759 (N_759,In_606,In_1152);
nor U760 (N_760,In_864,In_1473);
nor U761 (N_761,In_63,In_37);
and U762 (N_762,In_1405,In_1170);
or U763 (N_763,In_358,In_1283);
nand U764 (N_764,In_424,In_661);
xnor U765 (N_765,In_937,In_1204);
nand U766 (N_766,In_2,In_654);
or U767 (N_767,In_362,In_760);
xor U768 (N_768,In_1450,In_197);
and U769 (N_769,In_378,In_313);
nor U770 (N_770,In_344,In_502);
xnor U771 (N_771,In_1345,In_1);
and U772 (N_772,In_1151,In_968);
and U773 (N_773,In_127,In_194);
or U774 (N_774,In_224,In_244);
nor U775 (N_775,In_1295,In_420);
and U776 (N_776,In_155,In_766);
nor U777 (N_777,In_235,In_310);
nand U778 (N_778,In_1045,In_1037);
nor U779 (N_779,In_408,In_1496);
nand U780 (N_780,In_82,In_388);
or U781 (N_781,In_621,In_1296);
or U782 (N_782,In_178,In_497);
and U783 (N_783,In_217,In_418);
and U784 (N_784,In_1136,In_966);
nor U785 (N_785,In_707,In_335);
and U786 (N_786,In_888,In_909);
or U787 (N_787,In_20,In_317);
or U788 (N_788,In_853,In_956);
or U789 (N_789,In_525,In_544);
and U790 (N_790,In_483,In_804);
and U791 (N_791,In_816,In_1100);
nor U792 (N_792,In_63,In_250);
nand U793 (N_793,In_703,In_698);
xor U794 (N_794,In_681,In_84);
nor U795 (N_795,In_1210,In_753);
nand U796 (N_796,In_494,In_873);
nor U797 (N_797,In_733,In_1250);
nand U798 (N_798,In_1389,In_500);
nor U799 (N_799,In_129,In_201);
nor U800 (N_800,In_579,In_518);
nand U801 (N_801,In_899,In_1332);
and U802 (N_802,In_1002,In_90);
nand U803 (N_803,In_608,In_903);
nor U804 (N_804,In_539,In_1417);
and U805 (N_805,In_931,In_116);
nor U806 (N_806,In_1481,In_1053);
nor U807 (N_807,In_744,In_461);
nor U808 (N_808,In_746,In_1155);
and U809 (N_809,In_901,In_1119);
nor U810 (N_810,In_164,In_644);
nor U811 (N_811,In_390,In_1272);
nand U812 (N_812,In_1380,In_150);
nor U813 (N_813,In_1108,In_1067);
and U814 (N_814,In_1488,In_536);
and U815 (N_815,In_960,In_558);
and U816 (N_816,In_306,In_439);
and U817 (N_817,In_1408,In_83);
nand U818 (N_818,In_723,In_1215);
or U819 (N_819,In_810,In_1274);
nand U820 (N_820,In_751,In_259);
and U821 (N_821,In_753,In_1165);
and U822 (N_822,In_1229,In_284);
xnor U823 (N_823,In_501,In_403);
or U824 (N_824,In_535,In_1258);
and U825 (N_825,In_1262,In_1460);
nand U826 (N_826,In_209,In_1270);
nor U827 (N_827,In_881,In_1027);
nor U828 (N_828,In_669,In_195);
nor U829 (N_829,In_20,In_696);
or U830 (N_830,In_446,In_594);
nor U831 (N_831,In_620,In_109);
or U832 (N_832,In_175,In_1162);
nor U833 (N_833,In_500,In_1399);
nand U834 (N_834,In_360,In_1177);
or U835 (N_835,In_1410,In_953);
or U836 (N_836,In_873,In_1328);
nand U837 (N_837,In_592,In_1261);
xnor U838 (N_838,In_1447,In_699);
nor U839 (N_839,In_160,In_1232);
nand U840 (N_840,In_481,In_378);
and U841 (N_841,In_259,In_1064);
nor U842 (N_842,In_1053,In_16);
nor U843 (N_843,In_800,In_498);
nand U844 (N_844,In_478,In_349);
nor U845 (N_845,In_1315,In_504);
or U846 (N_846,In_839,In_493);
nor U847 (N_847,In_63,In_497);
nor U848 (N_848,In_1421,In_1335);
nand U849 (N_849,In_1119,In_173);
xnor U850 (N_850,In_715,In_280);
nor U851 (N_851,In_385,In_1303);
xor U852 (N_852,In_455,In_621);
and U853 (N_853,In_1022,In_1065);
nand U854 (N_854,In_423,In_935);
nor U855 (N_855,In_90,In_1007);
or U856 (N_856,In_637,In_1278);
nor U857 (N_857,In_883,In_912);
or U858 (N_858,In_1271,In_958);
nor U859 (N_859,In_170,In_126);
nand U860 (N_860,In_567,In_429);
nand U861 (N_861,In_1444,In_737);
xnor U862 (N_862,In_678,In_1025);
or U863 (N_863,In_1068,In_368);
and U864 (N_864,In_302,In_964);
nand U865 (N_865,In_1140,In_659);
nand U866 (N_866,In_1336,In_1104);
nand U867 (N_867,In_1386,In_1003);
xor U868 (N_868,In_917,In_841);
nor U869 (N_869,In_226,In_341);
and U870 (N_870,In_200,In_993);
nand U871 (N_871,In_257,In_1113);
nand U872 (N_872,In_274,In_1404);
and U873 (N_873,In_846,In_5);
nand U874 (N_874,In_933,In_788);
nand U875 (N_875,In_733,In_943);
nor U876 (N_876,In_960,In_1267);
nor U877 (N_877,In_511,In_935);
and U878 (N_878,In_1005,In_223);
or U879 (N_879,In_1371,In_1470);
nand U880 (N_880,In_1364,In_874);
and U881 (N_881,In_750,In_870);
nand U882 (N_882,In_1424,In_1206);
xor U883 (N_883,In_123,In_330);
nand U884 (N_884,In_883,In_475);
nand U885 (N_885,In_284,In_1334);
nor U886 (N_886,In_1140,In_1425);
nor U887 (N_887,In_1139,In_396);
nand U888 (N_888,In_830,In_733);
xor U889 (N_889,In_937,In_1173);
or U890 (N_890,In_511,In_759);
and U891 (N_891,In_50,In_828);
nor U892 (N_892,In_277,In_1108);
or U893 (N_893,In_298,In_735);
and U894 (N_894,In_287,In_111);
or U895 (N_895,In_1422,In_282);
nor U896 (N_896,In_382,In_592);
nor U897 (N_897,In_536,In_883);
and U898 (N_898,In_202,In_805);
or U899 (N_899,In_399,In_1036);
nor U900 (N_900,In_336,In_949);
or U901 (N_901,In_681,In_1304);
or U902 (N_902,In_624,In_455);
nor U903 (N_903,In_1443,In_1277);
or U904 (N_904,In_584,In_348);
nor U905 (N_905,In_618,In_1402);
xnor U906 (N_906,In_1149,In_1390);
nor U907 (N_907,In_1145,In_1297);
nand U908 (N_908,In_1441,In_442);
nor U909 (N_909,In_596,In_1289);
nor U910 (N_910,In_1441,In_1438);
nand U911 (N_911,In_338,In_1449);
and U912 (N_912,In_905,In_862);
and U913 (N_913,In_1186,In_196);
nor U914 (N_914,In_714,In_1335);
or U915 (N_915,In_15,In_838);
xor U916 (N_916,In_1031,In_174);
nand U917 (N_917,In_631,In_1370);
nor U918 (N_918,In_1070,In_78);
xor U919 (N_919,In_1257,In_1137);
and U920 (N_920,In_1415,In_1212);
nand U921 (N_921,In_957,In_1058);
nor U922 (N_922,In_920,In_1318);
nand U923 (N_923,In_784,In_92);
and U924 (N_924,In_427,In_1395);
nand U925 (N_925,In_1152,In_1146);
nand U926 (N_926,In_461,In_1044);
or U927 (N_927,In_686,In_825);
or U928 (N_928,In_1283,In_387);
nand U929 (N_929,In_155,In_682);
or U930 (N_930,In_702,In_358);
nor U931 (N_931,In_424,In_1196);
nor U932 (N_932,In_16,In_901);
and U933 (N_933,In_189,In_660);
nor U934 (N_934,In_509,In_1257);
and U935 (N_935,In_1148,In_858);
or U936 (N_936,In_8,In_986);
and U937 (N_937,In_1149,In_1214);
or U938 (N_938,In_1093,In_195);
or U939 (N_939,In_1439,In_504);
and U940 (N_940,In_1297,In_241);
nand U941 (N_941,In_42,In_1348);
and U942 (N_942,In_1403,In_1422);
xor U943 (N_943,In_117,In_390);
and U944 (N_944,In_300,In_1073);
and U945 (N_945,In_437,In_1126);
and U946 (N_946,In_742,In_1380);
nand U947 (N_947,In_65,In_919);
nand U948 (N_948,In_1001,In_547);
or U949 (N_949,In_1495,In_44);
xnor U950 (N_950,In_1189,In_1014);
nor U951 (N_951,In_495,In_1100);
nand U952 (N_952,In_1272,In_1343);
xnor U953 (N_953,In_27,In_762);
or U954 (N_954,In_600,In_1173);
xor U955 (N_955,In_4,In_333);
nand U956 (N_956,In_1045,In_260);
and U957 (N_957,In_172,In_648);
or U958 (N_958,In_1256,In_206);
or U959 (N_959,In_1139,In_332);
or U960 (N_960,In_249,In_797);
nor U961 (N_961,In_850,In_1414);
or U962 (N_962,In_948,In_819);
nand U963 (N_963,In_989,In_916);
or U964 (N_964,In_627,In_923);
and U965 (N_965,In_54,In_210);
and U966 (N_966,In_472,In_170);
nand U967 (N_967,In_93,In_1484);
nand U968 (N_968,In_1110,In_44);
nor U969 (N_969,In_761,In_211);
or U970 (N_970,In_1233,In_834);
nor U971 (N_971,In_39,In_876);
xor U972 (N_972,In_667,In_1170);
xor U973 (N_973,In_1034,In_1024);
nor U974 (N_974,In_471,In_732);
nor U975 (N_975,In_954,In_870);
nand U976 (N_976,In_993,In_622);
or U977 (N_977,In_766,In_1187);
or U978 (N_978,In_1400,In_202);
or U979 (N_979,In_833,In_1465);
nand U980 (N_980,In_1174,In_492);
or U981 (N_981,In_1254,In_159);
or U982 (N_982,In_93,In_722);
nor U983 (N_983,In_1293,In_389);
nand U984 (N_984,In_1085,In_171);
nor U985 (N_985,In_427,In_582);
and U986 (N_986,In_659,In_433);
and U987 (N_987,In_473,In_30);
nand U988 (N_988,In_645,In_609);
nand U989 (N_989,In_60,In_1063);
xor U990 (N_990,In_1177,In_422);
nor U991 (N_991,In_1210,In_809);
nor U992 (N_992,In_266,In_313);
or U993 (N_993,In_1291,In_449);
nor U994 (N_994,In_1176,In_629);
nand U995 (N_995,In_509,In_423);
nand U996 (N_996,In_384,In_1127);
nor U997 (N_997,In_95,In_1083);
nand U998 (N_998,In_558,In_830);
and U999 (N_999,In_1247,In_1360);
nor U1000 (N_1000,In_1170,In_1090);
nand U1001 (N_1001,In_500,In_160);
nor U1002 (N_1002,In_1181,In_803);
and U1003 (N_1003,In_1369,In_190);
xor U1004 (N_1004,In_572,In_934);
nor U1005 (N_1005,In_357,In_533);
nor U1006 (N_1006,In_85,In_236);
nor U1007 (N_1007,In_168,In_394);
nand U1008 (N_1008,In_333,In_1334);
nand U1009 (N_1009,In_1064,In_977);
and U1010 (N_1010,In_560,In_962);
and U1011 (N_1011,In_606,In_1208);
nand U1012 (N_1012,In_917,In_938);
nand U1013 (N_1013,In_1163,In_729);
or U1014 (N_1014,In_73,In_237);
or U1015 (N_1015,In_623,In_1121);
and U1016 (N_1016,In_1011,In_1208);
and U1017 (N_1017,In_1432,In_325);
nand U1018 (N_1018,In_667,In_1134);
or U1019 (N_1019,In_176,In_1418);
and U1020 (N_1020,In_1180,In_1144);
xor U1021 (N_1021,In_1438,In_399);
and U1022 (N_1022,In_481,In_173);
nor U1023 (N_1023,In_104,In_1220);
or U1024 (N_1024,In_143,In_560);
nand U1025 (N_1025,In_1102,In_126);
and U1026 (N_1026,In_863,In_1353);
nand U1027 (N_1027,In_674,In_522);
nor U1028 (N_1028,In_338,In_1138);
nand U1029 (N_1029,In_505,In_429);
and U1030 (N_1030,In_1164,In_718);
or U1031 (N_1031,In_20,In_1473);
or U1032 (N_1032,In_1428,In_150);
and U1033 (N_1033,In_1450,In_436);
and U1034 (N_1034,In_952,In_715);
and U1035 (N_1035,In_1276,In_1451);
nor U1036 (N_1036,In_1127,In_371);
and U1037 (N_1037,In_1053,In_1471);
or U1038 (N_1038,In_714,In_1192);
or U1039 (N_1039,In_1366,In_1323);
and U1040 (N_1040,In_190,In_944);
nor U1041 (N_1041,In_1172,In_1280);
xnor U1042 (N_1042,In_170,In_425);
nand U1043 (N_1043,In_1308,In_718);
nand U1044 (N_1044,In_485,In_179);
and U1045 (N_1045,In_881,In_279);
nand U1046 (N_1046,In_1214,In_565);
nor U1047 (N_1047,In_293,In_1401);
xor U1048 (N_1048,In_1075,In_459);
nor U1049 (N_1049,In_214,In_712);
or U1050 (N_1050,In_618,In_619);
or U1051 (N_1051,In_900,In_1245);
or U1052 (N_1052,In_880,In_1298);
nor U1053 (N_1053,In_800,In_1117);
nor U1054 (N_1054,In_700,In_1066);
nor U1055 (N_1055,In_364,In_500);
or U1056 (N_1056,In_870,In_483);
nand U1057 (N_1057,In_488,In_801);
and U1058 (N_1058,In_267,In_527);
nor U1059 (N_1059,In_1416,In_449);
nor U1060 (N_1060,In_1382,In_674);
and U1061 (N_1061,In_821,In_1349);
xnor U1062 (N_1062,In_283,In_26);
nor U1063 (N_1063,In_951,In_435);
nand U1064 (N_1064,In_651,In_1193);
or U1065 (N_1065,In_971,In_393);
or U1066 (N_1066,In_1336,In_1273);
xor U1067 (N_1067,In_1278,In_951);
nand U1068 (N_1068,In_526,In_533);
xnor U1069 (N_1069,In_926,In_1467);
or U1070 (N_1070,In_1368,In_106);
or U1071 (N_1071,In_874,In_237);
nand U1072 (N_1072,In_462,In_1224);
nand U1073 (N_1073,In_1126,In_319);
and U1074 (N_1074,In_795,In_391);
xor U1075 (N_1075,In_783,In_866);
nor U1076 (N_1076,In_301,In_916);
xor U1077 (N_1077,In_837,In_1202);
nor U1078 (N_1078,In_1348,In_1256);
or U1079 (N_1079,In_1479,In_1078);
and U1080 (N_1080,In_1458,In_888);
nand U1081 (N_1081,In_819,In_348);
nand U1082 (N_1082,In_199,In_937);
and U1083 (N_1083,In_592,In_828);
and U1084 (N_1084,In_907,In_989);
or U1085 (N_1085,In_566,In_1026);
and U1086 (N_1086,In_1325,In_883);
and U1087 (N_1087,In_217,In_1373);
nor U1088 (N_1088,In_913,In_1149);
or U1089 (N_1089,In_867,In_1372);
nor U1090 (N_1090,In_606,In_438);
or U1091 (N_1091,In_747,In_1067);
nand U1092 (N_1092,In_1233,In_1347);
xnor U1093 (N_1093,In_817,In_845);
nand U1094 (N_1094,In_1392,In_1152);
xnor U1095 (N_1095,In_968,In_449);
nor U1096 (N_1096,In_1292,In_236);
nand U1097 (N_1097,In_1318,In_1130);
or U1098 (N_1098,In_414,In_1239);
nor U1099 (N_1099,In_673,In_363);
or U1100 (N_1100,In_518,In_212);
and U1101 (N_1101,In_236,In_883);
nor U1102 (N_1102,In_363,In_1093);
or U1103 (N_1103,In_1143,In_1328);
nor U1104 (N_1104,In_1287,In_254);
xnor U1105 (N_1105,In_1096,In_885);
nand U1106 (N_1106,In_436,In_843);
xor U1107 (N_1107,In_827,In_100);
and U1108 (N_1108,In_98,In_1268);
or U1109 (N_1109,In_549,In_1351);
or U1110 (N_1110,In_390,In_1475);
nand U1111 (N_1111,In_732,In_413);
and U1112 (N_1112,In_146,In_840);
nor U1113 (N_1113,In_1198,In_331);
or U1114 (N_1114,In_1449,In_543);
or U1115 (N_1115,In_990,In_1224);
nand U1116 (N_1116,In_438,In_1217);
or U1117 (N_1117,In_111,In_1413);
and U1118 (N_1118,In_698,In_633);
and U1119 (N_1119,In_620,In_22);
or U1120 (N_1120,In_221,In_782);
xnor U1121 (N_1121,In_1130,In_272);
nor U1122 (N_1122,In_521,In_334);
xor U1123 (N_1123,In_585,In_46);
nand U1124 (N_1124,In_296,In_112);
or U1125 (N_1125,In_1234,In_851);
nand U1126 (N_1126,In_164,In_1321);
nor U1127 (N_1127,In_970,In_866);
nor U1128 (N_1128,In_947,In_409);
and U1129 (N_1129,In_1123,In_1331);
and U1130 (N_1130,In_499,In_1001);
nand U1131 (N_1131,In_360,In_167);
or U1132 (N_1132,In_867,In_1427);
nand U1133 (N_1133,In_783,In_725);
and U1134 (N_1134,In_1251,In_689);
nand U1135 (N_1135,In_912,In_376);
and U1136 (N_1136,In_674,In_6);
or U1137 (N_1137,In_1324,In_18);
nor U1138 (N_1138,In_1327,In_247);
or U1139 (N_1139,In_1087,In_210);
nor U1140 (N_1140,In_889,In_773);
nand U1141 (N_1141,In_1197,In_429);
nor U1142 (N_1142,In_945,In_769);
nand U1143 (N_1143,In_798,In_912);
nor U1144 (N_1144,In_307,In_921);
nand U1145 (N_1145,In_700,In_992);
xnor U1146 (N_1146,In_967,In_670);
nor U1147 (N_1147,In_458,In_702);
nand U1148 (N_1148,In_357,In_369);
nor U1149 (N_1149,In_1149,In_127);
nand U1150 (N_1150,In_586,In_104);
nor U1151 (N_1151,In_1349,In_472);
and U1152 (N_1152,In_604,In_136);
nand U1153 (N_1153,In_1291,In_503);
nand U1154 (N_1154,In_481,In_753);
or U1155 (N_1155,In_1405,In_883);
and U1156 (N_1156,In_1219,In_1482);
nor U1157 (N_1157,In_953,In_539);
and U1158 (N_1158,In_1048,In_340);
or U1159 (N_1159,In_847,In_18);
nor U1160 (N_1160,In_764,In_24);
nor U1161 (N_1161,In_358,In_1133);
nand U1162 (N_1162,In_1267,In_1303);
and U1163 (N_1163,In_1449,In_880);
and U1164 (N_1164,In_950,In_405);
or U1165 (N_1165,In_1065,In_777);
and U1166 (N_1166,In_469,In_1184);
and U1167 (N_1167,In_906,In_1317);
or U1168 (N_1168,In_236,In_446);
or U1169 (N_1169,In_345,In_182);
nor U1170 (N_1170,In_1124,In_84);
or U1171 (N_1171,In_1039,In_243);
or U1172 (N_1172,In_238,In_1083);
and U1173 (N_1173,In_1252,In_194);
and U1174 (N_1174,In_886,In_1491);
or U1175 (N_1175,In_709,In_258);
nor U1176 (N_1176,In_344,In_1486);
nor U1177 (N_1177,In_704,In_806);
nor U1178 (N_1178,In_306,In_753);
or U1179 (N_1179,In_1195,In_539);
xor U1180 (N_1180,In_277,In_482);
or U1181 (N_1181,In_1144,In_0);
and U1182 (N_1182,In_1103,In_1099);
nand U1183 (N_1183,In_1118,In_969);
nor U1184 (N_1184,In_614,In_278);
and U1185 (N_1185,In_1126,In_396);
and U1186 (N_1186,In_239,In_1239);
nand U1187 (N_1187,In_1381,In_643);
and U1188 (N_1188,In_571,In_334);
and U1189 (N_1189,In_254,In_173);
nor U1190 (N_1190,In_984,In_1423);
and U1191 (N_1191,In_746,In_1275);
and U1192 (N_1192,In_481,In_1098);
and U1193 (N_1193,In_363,In_119);
or U1194 (N_1194,In_836,In_72);
nand U1195 (N_1195,In_700,In_735);
or U1196 (N_1196,In_677,In_534);
nor U1197 (N_1197,In_810,In_706);
or U1198 (N_1198,In_798,In_882);
and U1199 (N_1199,In_318,In_1072);
or U1200 (N_1200,In_883,In_288);
nor U1201 (N_1201,In_272,In_1204);
or U1202 (N_1202,In_1358,In_736);
or U1203 (N_1203,In_734,In_402);
nand U1204 (N_1204,In_153,In_373);
or U1205 (N_1205,In_451,In_1198);
xor U1206 (N_1206,In_724,In_1178);
nand U1207 (N_1207,In_1022,In_960);
or U1208 (N_1208,In_955,In_1384);
and U1209 (N_1209,In_1121,In_644);
nor U1210 (N_1210,In_261,In_114);
and U1211 (N_1211,In_1398,In_211);
or U1212 (N_1212,In_75,In_1149);
nor U1213 (N_1213,In_1327,In_1237);
and U1214 (N_1214,In_306,In_732);
nor U1215 (N_1215,In_262,In_591);
nor U1216 (N_1216,In_200,In_448);
xnor U1217 (N_1217,In_895,In_1280);
nor U1218 (N_1218,In_1207,In_1204);
nand U1219 (N_1219,In_1045,In_140);
nand U1220 (N_1220,In_685,In_709);
nor U1221 (N_1221,In_998,In_206);
nand U1222 (N_1222,In_865,In_584);
and U1223 (N_1223,In_499,In_1235);
xor U1224 (N_1224,In_1436,In_830);
nand U1225 (N_1225,In_731,In_1313);
and U1226 (N_1226,In_114,In_561);
xnor U1227 (N_1227,In_1351,In_1414);
nand U1228 (N_1228,In_509,In_185);
nand U1229 (N_1229,In_1438,In_326);
or U1230 (N_1230,In_500,In_588);
or U1231 (N_1231,In_1316,In_225);
and U1232 (N_1232,In_1358,In_563);
or U1233 (N_1233,In_106,In_1386);
or U1234 (N_1234,In_441,In_864);
and U1235 (N_1235,In_1063,In_333);
or U1236 (N_1236,In_1440,In_38);
xnor U1237 (N_1237,In_1099,In_541);
or U1238 (N_1238,In_217,In_381);
nand U1239 (N_1239,In_818,In_93);
nand U1240 (N_1240,In_970,In_6);
nand U1241 (N_1241,In_643,In_1013);
nand U1242 (N_1242,In_241,In_529);
and U1243 (N_1243,In_476,In_577);
xor U1244 (N_1244,In_1494,In_1361);
and U1245 (N_1245,In_362,In_383);
or U1246 (N_1246,In_1225,In_1247);
nand U1247 (N_1247,In_344,In_1073);
nor U1248 (N_1248,In_1133,In_662);
and U1249 (N_1249,In_1481,In_1352);
nor U1250 (N_1250,In_1322,In_267);
nor U1251 (N_1251,In_896,In_406);
or U1252 (N_1252,In_116,In_295);
nor U1253 (N_1253,In_831,In_1403);
or U1254 (N_1254,In_13,In_242);
or U1255 (N_1255,In_282,In_253);
and U1256 (N_1256,In_1090,In_506);
nand U1257 (N_1257,In_307,In_546);
or U1258 (N_1258,In_149,In_1419);
or U1259 (N_1259,In_634,In_30);
or U1260 (N_1260,In_15,In_114);
xor U1261 (N_1261,In_54,In_438);
or U1262 (N_1262,In_432,In_1292);
nand U1263 (N_1263,In_402,In_1215);
or U1264 (N_1264,In_1439,In_883);
nand U1265 (N_1265,In_859,In_923);
xor U1266 (N_1266,In_532,In_383);
and U1267 (N_1267,In_311,In_1302);
and U1268 (N_1268,In_1195,In_1455);
and U1269 (N_1269,In_151,In_694);
nand U1270 (N_1270,In_1198,In_1429);
and U1271 (N_1271,In_893,In_806);
and U1272 (N_1272,In_435,In_1105);
nor U1273 (N_1273,In_1282,In_887);
and U1274 (N_1274,In_885,In_863);
and U1275 (N_1275,In_1369,In_1405);
nor U1276 (N_1276,In_1045,In_1177);
nor U1277 (N_1277,In_485,In_1351);
nand U1278 (N_1278,In_71,In_1128);
nand U1279 (N_1279,In_93,In_1256);
and U1280 (N_1280,In_1485,In_1275);
and U1281 (N_1281,In_168,In_1332);
nor U1282 (N_1282,In_42,In_1435);
or U1283 (N_1283,In_78,In_1301);
nor U1284 (N_1284,In_1319,In_1233);
and U1285 (N_1285,In_608,In_1041);
xnor U1286 (N_1286,In_767,In_858);
nor U1287 (N_1287,In_1424,In_1052);
or U1288 (N_1288,In_799,In_117);
and U1289 (N_1289,In_537,In_1350);
nor U1290 (N_1290,In_670,In_970);
nand U1291 (N_1291,In_628,In_845);
xnor U1292 (N_1292,In_1125,In_813);
xor U1293 (N_1293,In_279,In_918);
nand U1294 (N_1294,In_1099,In_1379);
or U1295 (N_1295,In_144,In_1092);
nor U1296 (N_1296,In_688,In_853);
nand U1297 (N_1297,In_1033,In_747);
nor U1298 (N_1298,In_401,In_61);
nand U1299 (N_1299,In_170,In_121);
nand U1300 (N_1300,In_102,In_218);
and U1301 (N_1301,In_223,In_1435);
xor U1302 (N_1302,In_912,In_1215);
nor U1303 (N_1303,In_1462,In_824);
or U1304 (N_1304,In_861,In_329);
nand U1305 (N_1305,In_1300,In_1224);
nor U1306 (N_1306,In_637,In_1427);
nand U1307 (N_1307,In_370,In_1011);
or U1308 (N_1308,In_360,In_560);
or U1309 (N_1309,In_870,In_1422);
xnor U1310 (N_1310,In_93,In_1057);
nand U1311 (N_1311,In_862,In_1423);
nand U1312 (N_1312,In_578,In_1345);
or U1313 (N_1313,In_1159,In_791);
xnor U1314 (N_1314,In_288,In_926);
xnor U1315 (N_1315,In_239,In_1161);
and U1316 (N_1316,In_1105,In_141);
or U1317 (N_1317,In_1335,In_543);
and U1318 (N_1318,In_153,In_95);
xor U1319 (N_1319,In_491,In_646);
and U1320 (N_1320,In_837,In_196);
nor U1321 (N_1321,In_497,In_740);
or U1322 (N_1322,In_863,In_567);
or U1323 (N_1323,In_996,In_1395);
nand U1324 (N_1324,In_201,In_1312);
or U1325 (N_1325,In_771,In_753);
nand U1326 (N_1326,In_792,In_183);
nand U1327 (N_1327,In_608,In_459);
nand U1328 (N_1328,In_327,In_461);
xnor U1329 (N_1329,In_207,In_626);
or U1330 (N_1330,In_829,In_70);
nand U1331 (N_1331,In_1153,In_348);
nor U1332 (N_1332,In_298,In_1385);
or U1333 (N_1333,In_625,In_1156);
or U1334 (N_1334,In_99,In_376);
and U1335 (N_1335,In_1330,In_817);
and U1336 (N_1336,In_1108,In_449);
nand U1337 (N_1337,In_727,In_55);
or U1338 (N_1338,In_1404,In_1266);
xnor U1339 (N_1339,In_653,In_1229);
nor U1340 (N_1340,In_1229,In_424);
or U1341 (N_1341,In_807,In_914);
or U1342 (N_1342,In_363,In_25);
nor U1343 (N_1343,In_477,In_189);
and U1344 (N_1344,In_1372,In_312);
nand U1345 (N_1345,In_497,In_111);
nor U1346 (N_1346,In_14,In_410);
nor U1347 (N_1347,In_254,In_236);
nor U1348 (N_1348,In_304,In_466);
nand U1349 (N_1349,In_564,In_188);
and U1350 (N_1350,In_1403,In_15);
nor U1351 (N_1351,In_491,In_424);
and U1352 (N_1352,In_1073,In_270);
nor U1353 (N_1353,In_803,In_1425);
nand U1354 (N_1354,In_1191,In_76);
nor U1355 (N_1355,In_499,In_513);
xor U1356 (N_1356,In_456,In_719);
and U1357 (N_1357,In_401,In_1068);
xor U1358 (N_1358,In_1256,In_694);
xnor U1359 (N_1359,In_792,In_27);
or U1360 (N_1360,In_936,In_1327);
and U1361 (N_1361,In_629,In_686);
or U1362 (N_1362,In_489,In_743);
nand U1363 (N_1363,In_1243,In_753);
nor U1364 (N_1364,In_1453,In_99);
xnor U1365 (N_1365,In_1356,In_315);
or U1366 (N_1366,In_61,In_1055);
nand U1367 (N_1367,In_1364,In_420);
or U1368 (N_1368,In_568,In_914);
or U1369 (N_1369,In_415,In_714);
nor U1370 (N_1370,In_351,In_622);
or U1371 (N_1371,In_18,In_944);
nand U1372 (N_1372,In_27,In_797);
nand U1373 (N_1373,In_1168,In_1311);
xor U1374 (N_1374,In_921,In_296);
xnor U1375 (N_1375,In_212,In_496);
nand U1376 (N_1376,In_34,In_1070);
or U1377 (N_1377,In_107,In_311);
or U1378 (N_1378,In_18,In_1143);
nand U1379 (N_1379,In_464,In_1189);
nor U1380 (N_1380,In_720,In_1285);
or U1381 (N_1381,In_582,In_1370);
and U1382 (N_1382,In_321,In_397);
nand U1383 (N_1383,In_878,In_97);
or U1384 (N_1384,In_456,In_60);
nor U1385 (N_1385,In_580,In_317);
or U1386 (N_1386,In_1203,In_668);
and U1387 (N_1387,In_1434,In_1206);
and U1388 (N_1388,In_64,In_353);
xor U1389 (N_1389,In_165,In_524);
or U1390 (N_1390,In_882,In_855);
nand U1391 (N_1391,In_1260,In_999);
xnor U1392 (N_1392,In_725,In_1108);
xnor U1393 (N_1393,In_1348,In_99);
nor U1394 (N_1394,In_1169,In_189);
or U1395 (N_1395,In_625,In_379);
nor U1396 (N_1396,In_1098,In_542);
and U1397 (N_1397,In_820,In_416);
nand U1398 (N_1398,In_671,In_1282);
and U1399 (N_1399,In_1268,In_620);
or U1400 (N_1400,In_1045,In_636);
and U1401 (N_1401,In_840,In_848);
nand U1402 (N_1402,In_602,In_1307);
or U1403 (N_1403,In_250,In_1164);
and U1404 (N_1404,In_289,In_312);
nand U1405 (N_1405,In_633,In_418);
and U1406 (N_1406,In_562,In_1233);
nor U1407 (N_1407,In_1343,In_238);
and U1408 (N_1408,In_234,In_1349);
xnor U1409 (N_1409,In_22,In_391);
nand U1410 (N_1410,In_796,In_974);
nand U1411 (N_1411,In_15,In_1107);
and U1412 (N_1412,In_1270,In_1483);
and U1413 (N_1413,In_1293,In_977);
nand U1414 (N_1414,In_1003,In_62);
and U1415 (N_1415,In_704,In_750);
nor U1416 (N_1416,In_444,In_227);
or U1417 (N_1417,In_0,In_1427);
and U1418 (N_1418,In_774,In_677);
xor U1419 (N_1419,In_1421,In_1351);
or U1420 (N_1420,In_585,In_649);
nor U1421 (N_1421,In_1413,In_885);
nor U1422 (N_1422,In_1305,In_1095);
nand U1423 (N_1423,In_1327,In_41);
and U1424 (N_1424,In_496,In_385);
or U1425 (N_1425,In_695,In_255);
nand U1426 (N_1426,In_1253,In_1238);
nand U1427 (N_1427,In_1247,In_895);
nand U1428 (N_1428,In_338,In_1204);
or U1429 (N_1429,In_1439,In_455);
or U1430 (N_1430,In_1482,In_1119);
and U1431 (N_1431,In_468,In_985);
and U1432 (N_1432,In_1317,In_1212);
xnor U1433 (N_1433,In_657,In_1375);
or U1434 (N_1434,In_1141,In_614);
nand U1435 (N_1435,In_281,In_826);
or U1436 (N_1436,In_1488,In_836);
xnor U1437 (N_1437,In_604,In_968);
or U1438 (N_1438,In_1240,In_766);
nand U1439 (N_1439,In_1340,In_1148);
nor U1440 (N_1440,In_1050,In_1313);
or U1441 (N_1441,In_244,In_680);
nand U1442 (N_1442,In_860,In_940);
nor U1443 (N_1443,In_12,In_1153);
and U1444 (N_1444,In_222,In_817);
nand U1445 (N_1445,In_992,In_655);
and U1446 (N_1446,In_364,In_661);
nor U1447 (N_1447,In_1390,In_672);
nor U1448 (N_1448,In_478,In_1340);
nand U1449 (N_1449,In_1178,In_571);
nand U1450 (N_1450,In_1070,In_648);
and U1451 (N_1451,In_331,In_277);
or U1452 (N_1452,In_957,In_525);
or U1453 (N_1453,In_435,In_471);
xnor U1454 (N_1454,In_1420,In_436);
nand U1455 (N_1455,In_1455,In_152);
nor U1456 (N_1456,In_25,In_1225);
xnor U1457 (N_1457,In_53,In_935);
or U1458 (N_1458,In_1320,In_832);
and U1459 (N_1459,In_1130,In_715);
or U1460 (N_1460,In_724,In_1487);
nor U1461 (N_1461,In_857,In_751);
and U1462 (N_1462,In_799,In_372);
or U1463 (N_1463,In_459,In_1477);
xnor U1464 (N_1464,In_436,In_272);
or U1465 (N_1465,In_118,In_13);
or U1466 (N_1466,In_441,In_118);
and U1467 (N_1467,In_1321,In_1390);
xor U1468 (N_1468,In_149,In_1222);
or U1469 (N_1469,In_1292,In_1458);
nand U1470 (N_1470,In_722,In_261);
nand U1471 (N_1471,In_235,In_206);
and U1472 (N_1472,In_217,In_1139);
or U1473 (N_1473,In_383,In_93);
xor U1474 (N_1474,In_1284,In_682);
or U1475 (N_1475,In_760,In_603);
nand U1476 (N_1476,In_1095,In_757);
and U1477 (N_1477,In_843,In_179);
nand U1478 (N_1478,In_108,In_763);
nand U1479 (N_1479,In_829,In_649);
and U1480 (N_1480,In_779,In_617);
nand U1481 (N_1481,In_934,In_634);
and U1482 (N_1482,In_746,In_731);
or U1483 (N_1483,In_766,In_399);
or U1484 (N_1484,In_1146,In_1140);
and U1485 (N_1485,In_1370,In_118);
and U1486 (N_1486,In_1148,In_1315);
nand U1487 (N_1487,In_919,In_985);
nor U1488 (N_1488,In_1190,In_359);
or U1489 (N_1489,In_963,In_86);
nand U1490 (N_1490,In_219,In_238);
or U1491 (N_1491,In_1057,In_1446);
nor U1492 (N_1492,In_1329,In_1373);
and U1493 (N_1493,In_476,In_421);
or U1494 (N_1494,In_164,In_328);
or U1495 (N_1495,In_290,In_1338);
xnor U1496 (N_1496,In_1460,In_457);
nand U1497 (N_1497,In_1427,In_868);
nor U1498 (N_1498,In_886,In_739);
nand U1499 (N_1499,In_200,In_170);
or U1500 (N_1500,In_970,In_1477);
nand U1501 (N_1501,In_649,In_876);
nand U1502 (N_1502,In_789,In_335);
and U1503 (N_1503,In_1249,In_1379);
nor U1504 (N_1504,In_1096,In_665);
and U1505 (N_1505,In_564,In_1392);
xnor U1506 (N_1506,In_205,In_1317);
or U1507 (N_1507,In_585,In_1196);
xnor U1508 (N_1508,In_171,In_778);
nor U1509 (N_1509,In_128,In_1377);
xor U1510 (N_1510,In_334,In_1028);
or U1511 (N_1511,In_959,In_87);
and U1512 (N_1512,In_37,In_309);
or U1513 (N_1513,In_1208,In_963);
or U1514 (N_1514,In_734,In_848);
and U1515 (N_1515,In_536,In_200);
xnor U1516 (N_1516,In_27,In_1430);
nand U1517 (N_1517,In_450,In_962);
nor U1518 (N_1518,In_194,In_1366);
and U1519 (N_1519,In_1007,In_89);
or U1520 (N_1520,In_157,In_1491);
and U1521 (N_1521,In_76,In_365);
nor U1522 (N_1522,In_815,In_987);
xor U1523 (N_1523,In_1335,In_785);
nand U1524 (N_1524,In_417,In_847);
or U1525 (N_1525,In_183,In_1171);
xor U1526 (N_1526,In_997,In_795);
nor U1527 (N_1527,In_1022,In_582);
nand U1528 (N_1528,In_395,In_877);
xor U1529 (N_1529,In_303,In_1490);
or U1530 (N_1530,In_226,In_1234);
and U1531 (N_1531,In_945,In_351);
and U1532 (N_1532,In_1272,In_1479);
nand U1533 (N_1533,In_218,In_1385);
nand U1534 (N_1534,In_903,In_1209);
and U1535 (N_1535,In_187,In_1108);
or U1536 (N_1536,In_256,In_53);
or U1537 (N_1537,In_1159,In_838);
nor U1538 (N_1538,In_1291,In_744);
nor U1539 (N_1539,In_1355,In_1422);
nor U1540 (N_1540,In_70,In_925);
xnor U1541 (N_1541,In_283,In_1074);
or U1542 (N_1542,In_474,In_952);
nand U1543 (N_1543,In_1415,In_62);
xor U1544 (N_1544,In_412,In_471);
nand U1545 (N_1545,In_1068,In_1192);
and U1546 (N_1546,In_1059,In_952);
nor U1547 (N_1547,In_1376,In_739);
or U1548 (N_1548,In_1242,In_1102);
nor U1549 (N_1549,In_149,In_929);
or U1550 (N_1550,In_1379,In_481);
nor U1551 (N_1551,In_854,In_1273);
or U1552 (N_1552,In_1454,In_76);
nor U1553 (N_1553,In_519,In_129);
xnor U1554 (N_1554,In_554,In_321);
or U1555 (N_1555,In_934,In_615);
nand U1556 (N_1556,In_1345,In_1466);
nor U1557 (N_1557,In_543,In_1239);
nor U1558 (N_1558,In_755,In_634);
nand U1559 (N_1559,In_983,In_888);
or U1560 (N_1560,In_356,In_1003);
and U1561 (N_1561,In_724,In_1254);
nand U1562 (N_1562,In_726,In_1455);
or U1563 (N_1563,In_1225,In_626);
nor U1564 (N_1564,In_422,In_1033);
or U1565 (N_1565,In_934,In_1494);
or U1566 (N_1566,In_768,In_353);
or U1567 (N_1567,In_1203,In_893);
nand U1568 (N_1568,In_568,In_1272);
and U1569 (N_1569,In_1147,In_871);
or U1570 (N_1570,In_33,In_662);
and U1571 (N_1571,In_342,In_595);
nand U1572 (N_1572,In_388,In_175);
and U1573 (N_1573,In_499,In_620);
nand U1574 (N_1574,In_754,In_1065);
and U1575 (N_1575,In_827,In_138);
nand U1576 (N_1576,In_399,In_243);
or U1577 (N_1577,In_760,In_722);
and U1578 (N_1578,In_1071,In_255);
nand U1579 (N_1579,In_432,In_213);
and U1580 (N_1580,In_232,In_1128);
nor U1581 (N_1581,In_1494,In_248);
nor U1582 (N_1582,In_63,In_638);
and U1583 (N_1583,In_665,In_1118);
and U1584 (N_1584,In_415,In_25);
and U1585 (N_1585,In_1475,In_133);
xor U1586 (N_1586,In_804,In_1067);
and U1587 (N_1587,In_696,In_332);
and U1588 (N_1588,In_402,In_1200);
and U1589 (N_1589,In_927,In_676);
and U1590 (N_1590,In_1252,In_209);
nor U1591 (N_1591,In_599,In_1115);
and U1592 (N_1592,In_1058,In_1060);
nor U1593 (N_1593,In_501,In_789);
or U1594 (N_1594,In_1055,In_30);
xnor U1595 (N_1595,In_1028,In_1132);
xnor U1596 (N_1596,In_1440,In_343);
or U1597 (N_1597,In_1311,In_275);
nand U1598 (N_1598,In_850,In_721);
and U1599 (N_1599,In_463,In_1471);
nor U1600 (N_1600,In_1449,In_1147);
and U1601 (N_1601,In_217,In_1049);
or U1602 (N_1602,In_1097,In_1163);
nor U1603 (N_1603,In_567,In_1081);
nor U1604 (N_1604,In_709,In_327);
nor U1605 (N_1605,In_512,In_83);
or U1606 (N_1606,In_346,In_752);
or U1607 (N_1607,In_1284,In_1090);
nor U1608 (N_1608,In_246,In_95);
and U1609 (N_1609,In_766,In_812);
nor U1610 (N_1610,In_1053,In_1359);
nand U1611 (N_1611,In_1118,In_1325);
nand U1612 (N_1612,In_161,In_633);
nor U1613 (N_1613,In_1362,In_1167);
nor U1614 (N_1614,In_471,In_437);
nor U1615 (N_1615,In_928,In_298);
nor U1616 (N_1616,In_352,In_1268);
nand U1617 (N_1617,In_910,In_425);
or U1618 (N_1618,In_999,In_1026);
and U1619 (N_1619,In_1381,In_457);
nand U1620 (N_1620,In_1415,In_40);
nand U1621 (N_1621,In_141,In_132);
xor U1622 (N_1622,In_1498,In_575);
nor U1623 (N_1623,In_647,In_699);
and U1624 (N_1624,In_1488,In_196);
xor U1625 (N_1625,In_1474,In_339);
and U1626 (N_1626,In_764,In_556);
nand U1627 (N_1627,In_1149,In_1041);
and U1628 (N_1628,In_239,In_296);
and U1629 (N_1629,In_700,In_398);
or U1630 (N_1630,In_934,In_1234);
nor U1631 (N_1631,In_733,In_1105);
nor U1632 (N_1632,In_1371,In_1167);
nor U1633 (N_1633,In_1096,In_1065);
or U1634 (N_1634,In_648,In_828);
nor U1635 (N_1635,In_141,In_1314);
or U1636 (N_1636,In_560,In_62);
and U1637 (N_1637,In_545,In_1303);
or U1638 (N_1638,In_1474,In_686);
and U1639 (N_1639,In_370,In_366);
xnor U1640 (N_1640,In_267,In_426);
nor U1641 (N_1641,In_1292,In_688);
or U1642 (N_1642,In_238,In_929);
and U1643 (N_1643,In_46,In_1368);
or U1644 (N_1644,In_1351,In_906);
or U1645 (N_1645,In_10,In_400);
or U1646 (N_1646,In_810,In_828);
and U1647 (N_1647,In_843,In_1244);
or U1648 (N_1648,In_495,In_1285);
nor U1649 (N_1649,In_1321,In_284);
nor U1650 (N_1650,In_240,In_835);
and U1651 (N_1651,In_1384,In_1277);
or U1652 (N_1652,In_1158,In_1274);
nand U1653 (N_1653,In_742,In_905);
nor U1654 (N_1654,In_885,In_192);
and U1655 (N_1655,In_1179,In_1337);
and U1656 (N_1656,In_306,In_923);
nand U1657 (N_1657,In_702,In_861);
nor U1658 (N_1658,In_1092,In_1213);
or U1659 (N_1659,In_369,In_1318);
and U1660 (N_1660,In_372,In_1114);
or U1661 (N_1661,In_671,In_692);
or U1662 (N_1662,In_492,In_485);
and U1663 (N_1663,In_572,In_649);
xor U1664 (N_1664,In_535,In_1429);
nor U1665 (N_1665,In_256,In_1231);
and U1666 (N_1666,In_723,In_198);
or U1667 (N_1667,In_371,In_109);
nor U1668 (N_1668,In_602,In_1206);
nand U1669 (N_1669,In_921,In_385);
and U1670 (N_1670,In_1252,In_678);
nor U1671 (N_1671,In_785,In_193);
nor U1672 (N_1672,In_1063,In_181);
nor U1673 (N_1673,In_256,In_1093);
and U1674 (N_1674,In_1132,In_733);
nor U1675 (N_1675,In_642,In_1114);
xnor U1676 (N_1676,In_391,In_1259);
nand U1677 (N_1677,In_45,In_1493);
and U1678 (N_1678,In_202,In_1475);
xnor U1679 (N_1679,In_219,In_1227);
nor U1680 (N_1680,In_91,In_904);
and U1681 (N_1681,In_1188,In_475);
or U1682 (N_1682,In_927,In_1088);
nor U1683 (N_1683,In_589,In_1197);
or U1684 (N_1684,In_352,In_65);
nor U1685 (N_1685,In_1024,In_817);
or U1686 (N_1686,In_1000,In_1244);
nor U1687 (N_1687,In_439,In_1425);
nor U1688 (N_1688,In_594,In_212);
nor U1689 (N_1689,In_920,In_527);
nand U1690 (N_1690,In_1156,In_263);
or U1691 (N_1691,In_378,In_1262);
and U1692 (N_1692,In_1196,In_842);
or U1693 (N_1693,In_78,In_104);
nand U1694 (N_1694,In_568,In_1053);
or U1695 (N_1695,In_380,In_359);
and U1696 (N_1696,In_504,In_49);
and U1697 (N_1697,In_662,In_1228);
or U1698 (N_1698,In_271,In_244);
xor U1699 (N_1699,In_819,In_710);
or U1700 (N_1700,In_1043,In_800);
and U1701 (N_1701,In_1204,In_1085);
and U1702 (N_1702,In_763,In_1080);
nand U1703 (N_1703,In_1310,In_852);
nand U1704 (N_1704,In_259,In_295);
or U1705 (N_1705,In_1273,In_489);
nor U1706 (N_1706,In_378,In_948);
nor U1707 (N_1707,In_650,In_63);
and U1708 (N_1708,In_910,In_278);
nand U1709 (N_1709,In_455,In_54);
xnor U1710 (N_1710,In_951,In_1193);
nand U1711 (N_1711,In_71,In_641);
nor U1712 (N_1712,In_139,In_269);
nand U1713 (N_1713,In_185,In_1173);
nor U1714 (N_1714,In_1328,In_1290);
nand U1715 (N_1715,In_670,In_1238);
or U1716 (N_1716,In_176,In_862);
and U1717 (N_1717,In_349,In_1495);
and U1718 (N_1718,In_634,In_14);
or U1719 (N_1719,In_489,In_89);
nor U1720 (N_1720,In_1256,In_747);
xor U1721 (N_1721,In_96,In_105);
and U1722 (N_1722,In_725,In_326);
xor U1723 (N_1723,In_1329,In_1350);
and U1724 (N_1724,In_842,In_982);
xnor U1725 (N_1725,In_930,In_1075);
and U1726 (N_1726,In_345,In_1102);
nand U1727 (N_1727,In_1128,In_1318);
and U1728 (N_1728,In_197,In_621);
and U1729 (N_1729,In_1095,In_265);
and U1730 (N_1730,In_1106,In_493);
nor U1731 (N_1731,In_236,In_76);
or U1732 (N_1732,In_195,In_1068);
or U1733 (N_1733,In_856,In_993);
nor U1734 (N_1734,In_978,In_1388);
or U1735 (N_1735,In_480,In_345);
and U1736 (N_1736,In_167,In_288);
nor U1737 (N_1737,In_1481,In_36);
nor U1738 (N_1738,In_1479,In_884);
nor U1739 (N_1739,In_484,In_320);
and U1740 (N_1740,In_1310,In_173);
and U1741 (N_1741,In_1345,In_24);
nor U1742 (N_1742,In_81,In_839);
or U1743 (N_1743,In_201,In_1137);
or U1744 (N_1744,In_1060,In_175);
xor U1745 (N_1745,In_956,In_809);
nor U1746 (N_1746,In_380,In_565);
and U1747 (N_1747,In_443,In_611);
or U1748 (N_1748,In_725,In_1001);
nor U1749 (N_1749,In_168,In_675);
nand U1750 (N_1750,In_1423,In_1198);
xor U1751 (N_1751,In_1225,In_365);
and U1752 (N_1752,In_1305,In_1114);
xor U1753 (N_1753,In_1171,In_783);
nor U1754 (N_1754,In_171,In_1109);
nand U1755 (N_1755,In_1347,In_849);
and U1756 (N_1756,In_179,In_870);
nand U1757 (N_1757,In_254,In_188);
nand U1758 (N_1758,In_362,In_77);
nor U1759 (N_1759,In_1382,In_506);
nor U1760 (N_1760,In_859,In_503);
nand U1761 (N_1761,In_662,In_1490);
and U1762 (N_1762,In_582,In_1009);
or U1763 (N_1763,In_1095,In_72);
nand U1764 (N_1764,In_1110,In_1141);
or U1765 (N_1765,In_1278,In_768);
nor U1766 (N_1766,In_181,In_1465);
nor U1767 (N_1767,In_1251,In_1398);
nor U1768 (N_1768,In_1138,In_1007);
nor U1769 (N_1769,In_454,In_1209);
and U1770 (N_1770,In_459,In_1307);
or U1771 (N_1771,In_613,In_466);
or U1772 (N_1772,In_153,In_1390);
xnor U1773 (N_1773,In_298,In_173);
and U1774 (N_1774,In_1271,In_1426);
nor U1775 (N_1775,In_658,In_35);
nor U1776 (N_1776,In_1308,In_382);
nor U1777 (N_1777,In_571,In_1317);
nor U1778 (N_1778,In_448,In_680);
nand U1779 (N_1779,In_165,In_832);
nand U1780 (N_1780,In_660,In_206);
and U1781 (N_1781,In_1307,In_720);
xnor U1782 (N_1782,In_360,In_1080);
nor U1783 (N_1783,In_579,In_871);
nand U1784 (N_1784,In_426,In_1109);
nor U1785 (N_1785,In_1367,In_802);
nand U1786 (N_1786,In_1462,In_96);
nor U1787 (N_1787,In_178,In_85);
nand U1788 (N_1788,In_343,In_1152);
nand U1789 (N_1789,In_304,In_1298);
nand U1790 (N_1790,In_1257,In_759);
nor U1791 (N_1791,In_794,In_724);
and U1792 (N_1792,In_710,In_644);
nor U1793 (N_1793,In_1020,In_853);
or U1794 (N_1794,In_1386,In_594);
and U1795 (N_1795,In_310,In_1147);
nor U1796 (N_1796,In_1002,In_474);
nor U1797 (N_1797,In_369,In_224);
nor U1798 (N_1798,In_1427,In_1214);
xor U1799 (N_1799,In_387,In_56);
nand U1800 (N_1800,In_615,In_428);
nand U1801 (N_1801,In_312,In_1111);
and U1802 (N_1802,In_131,In_269);
nand U1803 (N_1803,In_385,In_664);
or U1804 (N_1804,In_1381,In_401);
nand U1805 (N_1805,In_175,In_527);
nand U1806 (N_1806,In_1485,In_584);
and U1807 (N_1807,In_968,In_897);
nand U1808 (N_1808,In_903,In_174);
and U1809 (N_1809,In_659,In_627);
nand U1810 (N_1810,In_201,In_284);
xnor U1811 (N_1811,In_1380,In_946);
xor U1812 (N_1812,In_939,In_1023);
or U1813 (N_1813,In_1145,In_690);
or U1814 (N_1814,In_1461,In_413);
and U1815 (N_1815,In_147,In_34);
nand U1816 (N_1816,In_95,In_1486);
nor U1817 (N_1817,In_1014,In_533);
or U1818 (N_1818,In_170,In_995);
or U1819 (N_1819,In_1462,In_334);
or U1820 (N_1820,In_1364,In_752);
nand U1821 (N_1821,In_256,In_1099);
nor U1822 (N_1822,In_521,In_952);
or U1823 (N_1823,In_937,In_1304);
or U1824 (N_1824,In_558,In_815);
and U1825 (N_1825,In_1162,In_1245);
nor U1826 (N_1826,In_733,In_844);
or U1827 (N_1827,In_481,In_1288);
and U1828 (N_1828,In_360,In_1056);
nor U1829 (N_1829,In_470,In_1375);
or U1830 (N_1830,In_478,In_176);
and U1831 (N_1831,In_342,In_1474);
and U1832 (N_1832,In_922,In_121);
nand U1833 (N_1833,In_127,In_569);
or U1834 (N_1834,In_629,In_81);
nand U1835 (N_1835,In_1159,In_1165);
and U1836 (N_1836,In_1030,In_701);
and U1837 (N_1837,In_1376,In_634);
xnor U1838 (N_1838,In_1473,In_199);
and U1839 (N_1839,In_629,In_1361);
nand U1840 (N_1840,In_1177,In_824);
nor U1841 (N_1841,In_629,In_698);
and U1842 (N_1842,In_1118,In_905);
or U1843 (N_1843,In_219,In_588);
nand U1844 (N_1844,In_1368,In_342);
nor U1845 (N_1845,In_363,In_31);
nor U1846 (N_1846,In_532,In_255);
and U1847 (N_1847,In_268,In_290);
or U1848 (N_1848,In_957,In_438);
xnor U1849 (N_1849,In_811,In_978);
and U1850 (N_1850,In_1096,In_756);
nand U1851 (N_1851,In_661,In_710);
nor U1852 (N_1852,In_1492,In_383);
and U1853 (N_1853,In_870,In_507);
nand U1854 (N_1854,In_1478,In_865);
nand U1855 (N_1855,In_522,In_362);
and U1856 (N_1856,In_337,In_1260);
or U1857 (N_1857,In_304,In_934);
and U1858 (N_1858,In_26,In_1399);
xor U1859 (N_1859,In_698,In_884);
xnor U1860 (N_1860,In_884,In_430);
nor U1861 (N_1861,In_1475,In_151);
or U1862 (N_1862,In_831,In_149);
or U1863 (N_1863,In_265,In_240);
or U1864 (N_1864,In_1423,In_694);
or U1865 (N_1865,In_1264,In_870);
or U1866 (N_1866,In_340,In_419);
nand U1867 (N_1867,In_951,In_133);
and U1868 (N_1868,In_1124,In_58);
nor U1869 (N_1869,In_15,In_1390);
or U1870 (N_1870,In_1499,In_704);
or U1871 (N_1871,In_455,In_1365);
nand U1872 (N_1872,In_147,In_873);
nand U1873 (N_1873,In_109,In_632);
and U1874 (N_1874,In_119,In_108);
nor U1875 (N_1875,In_1222,In_316);
xor U1876 (N_1876,In_1353,In_704);
or U1877 (N_1877,In_782,In_918);
nor U1878 (N_1878,In_125,In_1332);
nor U1879 (N_1879,In_751,In_94);
or U1880 (N_1880,In_1487,In_350);
nand U1881 (N_1881,In_1161,In_292);
xor U1882 (N_1882,In_430,In_835);
and U1883 (N_1883,In_380,In_48);
and U1884 (N_1884,In_324,In_947);
nor U1885 (N_1885,In_337,In_537);
nand U1886 (N_1886,In_274,In_118);
xnor U1887 (N_1887,In_1132,In_1304);
nand U1888 (N_1888,In_600,In_1301);
nand U1889 (N_1889,In_1492,In_1384);
and U1890 (N_1890,In_894,In_1259);
nor U1891 (N_1891,In_352,In_62);
and U1892 (N_1892,In_204,In_493);
and U1893 (N_1893,In_976,In_169);
nand U1894 (N_1894,In_1105,In_360);
and U1895 (N_1895,In_1053,In_932);
and U1896 (N_1896,In_1385,In_582);
nor U1897 (N_1897,In_814,In_1346);
nor U1898 (N_1898,In_1496,In_821);
xor U1899 (N_1899,In_217,In_486);
or U1900 (N_1900,In_1429,In_376);
nand U1901 (N_1901,In_1181,In_473);
and U1902 (N_1902,In_1442,In_377);
nor U1903 (N_1903,In_809,In_1247);
nor U1904 (N_1904,In_1246,In_526);
xor U1905 (N_1905,In_1163,In_757);
nor U1906 (N_1906,In_1493,In_876);
xnor U1907 (N_1907,In_6,In_1186);
and U1908 (N_1908,In_1096,In_1203);
and U1909 (N_1909,In_96,In_1109);
xnor U1910 (N_1910,In_918,In_510);
or U1911 (N_1911,In_1234,In_415);
or U1912 (N_1912,In_733,In_1429);
nor U1913 (N_1913,In_1247,In_953);
and U1914 (N_1914,In_371,In_719);
nand U1915 (N_1915,In_1262,In_629);
xnor U1916 (N_1916,In_617,In_201);
and U1917 (N_1917,In_971,In_1013);
nand U1918 (N_1918,In_1333,In_413);
nand U1919 (N_1919,In_888,In_6);
nor U1920 (N_1920,In_1003,In_1476);
nand U1921 (N_1921,In_202,In_830);
xnor U1922 (N_1922,In_596,In_670);
nor U1923 (N_1923,In_1261,In_831);
or U1924 (N_1924,In_1409,In_378);
nand U1925 (N_1925,In_974,In_575);
nor U1926 (N_1926,In_385,In_1036);
nand U1927 (N_1927,In_776,In_590);
nor U1928 (N_1928,In_261,In_1483);
and U1929 (N_1929,In_951,In_423);
and U1930 (N_1930,In_877,In_893);
or U1931 (N_1931,In_61,In_849);
or U1932 (N_1932,In_259,In_322);
nor U1933 (N_1933,In_366,In_1184);
and U1934 (N_1934,In_362,In_410);
nand U1935 (N_1935,In_375,In_17);
and U1936 (N_1936,In_1273,In_317);
or U1937 (N_1937,In_957,In_68);
or U1938 (N_1938,In_1091,In_1018);
nor U1939 (N_1939,In_1360,In_982);
and U1940 (N_1940,In_516,In_539);
xnor U1941 (N_1941,In_270,In_198);
nand U1942 (N_1942,In_1320,In_233);
nor U1943 (N_1943,In_1312,In_343);
nor U1944 (N_1944,In_122,In_1169);
or U1945 (N_1945,In_605,In_742);
nor U1946 (N_1946,In_196,In_548);
nand U1947 (N_1947,In_155,In_1421);
nor U1948 (N_1948,In_424,In_787);
xor U1949 (N_1949,In_685,In_965);
and U1950 (N_1950,In_1197,In_104);
nor U1951 (N_1951,In_604,In_429);
and U1952 (N_1952,In_1345,In_1241);
and U1953 (N_1953,In_465,In_381);
or U1954 (N_1954,In_1221,In_648);
and U1955 (N_1955,In_795,In_698);
or U1956 (N_1956,In_529,In_328);
nor U1957 (N_1957,In_646,In_536);
nand U1958 (N_1958,In_906,In_76);
or U1959 (N_1959,In_563,In_1272);
or U1960 (N_1960,In_1347,In_156);
nand U1961 (N_1961,In_431,In_1109);
or U1962 (N_1962,In_1087,In_1275);
and U1963 (N_1963,In_280,In_1297);
or U1964 (N_1964,In_563,In_160);
and U1965 (N_1965,In_458,In_517);
nand U1966 (N_1966,In_796,In_539);
and U1967 (N_1967,In_262,In_1006);
nor U1968 (N_1968,In_759,In_145);
or U1969 (N_1969,In_1104,In_607);
nand U1970 (N_1970,In_26,In_586);
and U1971 (N_1971,In_79,In_353);
nor U1972 (N_1972,In_1182,In_1214);
or U1973 (N_1973,In_366,In_439);
nor U1974 (N_1974,In_884,In_334);
or U1975 (N_1975,In_1418,In_392);
nor U1976 (N_1976,In_363,In_871);
and U1977 (N_1977,In_1391,In_736);
nor U1978 (N_1978,In_1061,In_1232);
nor U1979 (N_1979,In_863,In_777);
or U1980 (N_1980,In_589,In_1217);
and U1981 (N_1981,In_258,In_831);
and U1982 (N_1982,In_943,In_905);
nand U1983 (N_1983,In_31,In_1164);
and U1984 (N_1984,In_29,In_530);
or U1985 (N_1985,In_415,In_980);
xnor U1986 (N_1986,In_944,In_356);
nor U1987 (N_1987,In_140,In_723);
nor U1988 (N_1988,In_999,In_569);
nand U1989 (N_1989,In_570,In_43);
and U1990 (N_1990,In_851,In_128);
or U1991 (N_1991,In_1256,In_1303);
nor U1992 (N_1992,In_1010,In_252);
nor U1993 (N_1993,In_1285,In_337);
and U1994 (N_1994,In_956,In_689);
nand U1995 (N_1995,In_1233,In_51);
nand U1996 (N_1996,In_1348,In_404);
and U1997 (N_1997,In_390,In_1239);
nand U1998 (N_1998,In_137,In_674);
nor U1999 (N_1999,In_234,In_353);
and U2000 (N_2000,In_675,In_652);
or U2001 (N_2001,In_94,In_77);
and U2002 (N_2002,In_209,In_1126);
and U2003 (N_2003,In_487,In_327);
or U2004 (N_2004,In_532,In_67);
nand U2005 (N_2005,In_862,In_509);
nand U2006 (N_2006,In_1204,In_1089);
and U2007 (N_2007,In_1335,In_1069);
and U2008 (N_2008,In_852,In_208);
nand U2009 (N_2009,In_1162,In_717);
nor U2010 (N_2010,In_673,In_734);
nor U2011 (N_2011,In_839,In_1319);
nand U2012 (N_2012,In_149,In_1324);
nand U2013 (N_2013,In_475,In_146);
xor U2014 (N_2014,In_979,In_1068);
nand U2015 (N_2015,In_1,In_46);
and U2016 (N_2016,In_116,In_1221);
nand U2017 (N_2017,In_977,In_1245);
or U2018 (N_2018,In_536,In_66);
or U2019 (N_2019,In_343,In_1290);
or U2020 (N_2020,In_247,In_948);
and U2021 (N_2021,In_1226,In_892);
and U2022 (N_2022,In_198,In_829);
and U2023 (N_2023,In_811,In_1107);
or U2024 (N_2024,In_592,In_1461);
or U2025 (N_2025,In_70,In_366);
or U2026 (N_2026,In_1335,In_1448);
xor U2027 (N_2027,In_951,In_843);
or U2028 (N_2028,In_720,In_1086);
nor U2029 (N_2029,In_1178,In_173);
and U2030 (N_2030,In_308,In_1401);
or U2031 (N_2031,In_1129,In_594);
xnor U2032 (N_2032,In_1126,In_642);
xnor U2033 (N_2033,In_1237,In_1465);
nor U2034 (N_2034,In_1010,In_361);
and U2035 (N_2035,In_249,In_845);
nand U2036 (N_2036,In_1161,In_255);
or U2037 (N_2037,In_840,In_712);
xnor U2038 (N_2038,In_999,In_1246);
and U2039 (N_2039,In_755,In_618);
nor U2040 (N_2040,In_446,In_1068);
nand U2041 (N_2041,In_744,In_283);
xnor U2042 (N_2042,In_883,In_618);
xor U2043 (N_2043,In_1003,In_612);
nand U2044 (N_2044,In_412,In_362);
nand U2045 (N_2045,In_1387,In_788);
nor U2046 (N_2046,In_487,In_696);
nand U2047 (N_2047,In_1322,In_1218);
xor U2048 (N_2048,In_778,In_172);
and U2049 (N_2049,In_102,In_1196);
and U2050 (N_2050,In_86,In_1427);
and U2051 (N_2051,In_1282,In_188);
nor U2052 (N_2052,In_433,In_1159);
and U2053 (N_2053,In_365,In_92);
and U2054 (N_2054,In_517,In_1376);
nor U2055 (N_2055,In_564,In_1235);
nand U2056 (N_2056,In_842,In_945);
nand U2057 (N_2057,In_28,In_392);
nand U2058 (N_2058,In_673,In_1029);
nor U2059 (N_2059,In_423,In_1226);
nand U2060 (N_2060,In_207,In_1083);
nor U2061 (N_2061,In_595,In_111);
or U2062 (N_2062,In_576,In_371);
nand U2063 (N_2063,In_1196,In_713);
and U2064 (N_2064,In_1284,In_781);
nor U2065 (N_2065,In_1442,In_444);
nand U2066 (N_2066,In_217,In_534);
or U2067 (N_2067,In_1244,In_978);
and U2068 (N_2068,In_835,In_1040);
or U2069 (N_2069,In_319,In_1121);
xor U2070 (N_2070,In_534,In_1204);
or U2071 (N_2071,In_258,In_906);
or U2072 (N_2072,In_935,In_324);
nor U2073 (N_2073,In_146,In_204);
nor U2074 (N_2074,In_379,In_181);
nand U2075 (N_2075,In_730,In_1039);
and U2076 (N_2076,In_1214,In_1212);
nand U2077 (N_2077,In_260,In_1112);
and U2078 (N_2078,In_11,In_799);
and U2079 (N_2079,In_252,In_829);
nand U2080 (N_2080,In_1299,In_820);
xnor U2081 (N_2081,In_1482,In_108);
nand U2082 (N_2082,In_668,In_361);
nand U2083 (N_2083,In_732,In_153);
and U2084 (N_2084,In_1367,In_503);
or U2085 (N_2085,In_676,In_723);
or U2086 (N_2086,In_708,In_377);
nand U2087 (N_2087,In_429,In_1466);
nor U2088 (N_2088,In_967,In_829);
or U2089 (N_2089,In_306,In_553);
nor U2090 (N_2090,In_1047,In_164);
and U2091 (N_2091,In_799,In_611);
nand U2092 (N_2092,In_157,In_793);
nand U2093 (N_2093,In_405,In_1008);
and U2094 (N_2094,In_944,In_1354);
and U2095 (N_2095,In_1331,In_565);
or U2096 (N_2096,In_719,In_276);
nor U2097 (N_2097,In_566,In_1233);
and U2098 (N_2098,In_81,In_366);
or U2099 (N_2099,In_723,In_909);
nor U2100 (N_2100,In_461,In_494);
nand U2101 (N_2101,In_1468,In_900);
or U2102 (N_2102,In_1055,In_213);
nand U2103 (N_2103,In_787,In_355);
and U2104 (N_2104,In_432,In_1459);
nor U2105 (N_2105,In_968,In_1142);
or U2106 (N_2106,In_977,In_122);
and U2107 (N_2107,In_733,In_970);
or U2108 (N_2108,In_142,In_1327);
or U2109 (N_2109,In_1001,In_610);
nor U2110 (N_2110,In_624,In_190);
or U2111 (N_2111,In_244,In_900);
nor U2112 (N_2112,In_882,In_1359);
nor U2113 (N_2113,In_366,In_294);
or U2114 (N_2114,In_372,In_740);
and U2115 (N_2115,In_548,In_1169);
nor U2116 (N_2116,In_841,In_1269);
or U2117 (N_2117,In_668,In_1347);
nor U2118 (N_2118,In_1324,In_1237);
or U2119 (N_2119,In_966,In_532);
xnor U2120 (N_2120,In_981,In_1358);
xor U2121 (N_2121,In_1419,In_1146);
nand U2122 (N_2122,In_1185,In_265);
or U2123 (N_2123,In_474,In_1137);
nand U2124 (N_2124,In_376,In_1271);
xor U2125 (N_2125,In_1316,In_773);
or U2126 (N_2126,In_79,In_173);
and U2127 (N_2127,In_1404,In_674);
xnor U2128 (N_2128,In_801,In_1419);
and U2129 (N_2129,In_1441,In_914);
and U2130 (N_2130,In_1402,In_1301);
or U2131 (N_2131,In_793,In_405);
or U2132 (N_2132,In_621,In_24);
and U2133 (N_2133,In_424,In_1395);
or U2134 (N_2134,In_900,In_890);
or U2135 (N_2135,In_1356,In_134);
and U2136 (N_2136,In_720,In_734);
and U2137 (N_2137,In_720,In_1093);
nor U2138 (N_2138,In_1444,In_1028);
nand U2139 (N_2139,In_426,In_1256);
nand U2140 (N_2140,In_870,In_736);
or U2141 (N_2141,In_1141,In_449);
nor U2142 (N_2142,In_375,In_388);
nor U2143 (N_2143,In_96,In_1354);
and U2144 (N_2144,In_256,In_1011);
nand U2145 (N_2145,In_1368,In_914);
or U2146 (N_2146,In_656,In_1266);
nor U2147 (N_2147,In_637,In_1340);
nor U2148 (N_2148,In_451,In_375);
or U2149 (N_2149,In_95,In_1462);
nand U2150 (N_2150,In_83,In_701);
nor U2151 (N_2151,In_1301,In_309);
nor U2152 (N_2152,In_283,In_18);
or U2153 (N_2153,In_1139,In_87);
or U2154 (N_2154,In_769,In_873);
xnor U2155 (N_2155,In_691,In_1149);
or U2156 (N_2156,In_221,In_337);
or U2157 (N_2157,In_197,In_872);
and U2158 (N_2158,In_1495,In_514);
nand U2159 (N_2159,In_1408,In_1010);
nor U2160 (N_2160,In_1067,In_1410);
or U2161 (N_2161,In_1329,In_354);
nand U2162 (N_2162,In_856,In_672);
nor U2163 (N_2163,In_799,In_599);
or U2164 (N_2164,In_1216,In_915);
and U2165 (N_2165,In_270,In_346);
nand U2166 (N_2166,In_1328,In_78);
or U2167 (N_2167,In_268,In_593);
or U2168 (N_2168,In_815,In_179);
or U2169 (N_2169,In_29,In_899);
nor U2170 (N_2170,In_384,In_1066);
nand U2171 (N_2171,In_900,In_1035);
nand U2172 (N_2172,In_1006,In_132);
nor U2173 (N_2173,In_1176,In_393);
and U2174 (N_2174,In_684,In_1086);
nand U2175 (N_2175,In_564,In_1229);
or U2176 (N_2176,In_1135,In_514);
or U2177 (N_2177,In_1018,In_466);
nand U2178 (N_2178,In_251,In_68);
and U2179 (N_2179,In_599,In_1094);
and U2180 (N_2180,In_936,In_940);
nand U2181 (N_2181,In_1089,In_676);
and U2182 (N_2182,In_201,In_312);
nand U2183 (N_2183,In_775,In_1271);
nor U2184 (N_2184,In_301,In_1494);
or U2185 (N_2185,In_417,In_378);
and U2186 (N_2186,In_792,In_222);
and U2187 (N_2187,In_530,In_1157);
xor U2188 (N_2188,In_1103,In_326);
or U2189 (N_2189,In_827,In_604);
nor U2190 (N_2190,In_1406,In_1395);
xor U2191 (N_2191,In_29,In_1320);
and U2192 (N_2192,In_326,In_1436);
nor U2193 (N_2193,In_694,In_604);
or U2194 (N_2194,In_1288,In_281);
or U2195 (N_2195,In_878,In_38);
nor U2196 (N_2196,In_1353,In_1498);
nand U2197 (N_2197,In_335,In_598);
xor U2198 (N_2198,In_1153,In_1297);
and U2199 (N_2199,In_901,In_1075);
nor U2200 (N_2200,In_1492,In_1220);
nor U2201 (N_2201,In_948,In_807);
nand U2202 (N_2202,In_961,In_772);
xnor U2203 (N_2203,In_988,In_1170);
and U2204 (N_2204,In_5,In_101);
nor U2205 (N_2205,In_986,In_958);
xor U2206 (N_2206,In_1389,In_1084);
or U2207 (N_2207,In_1343,In_1328);
or U2208 (N_2208,In_662,In_1019);
nor U2209 (N_2209,In_350,In_987);
or U2210 (N_2210,In_639,In_67);
nor U2211 (N_2211,In_819,In_1);
and U2212 (N_2212,In_847,In_1478);
nor U2213 (N_2213,In_1116,In_1405);
nor U2214 (N_2214,In_704,In_761);
nor U2215 (N_2215,In_159,In_469);
xor U2216 (N_2216,In_628,In_713);
nor U2217 (N_2217,In_176,In_355);
nand U2218 (N_2218,In_41,In_1458);
nor U2219 (N_2219,In_378,In_371);
nor U2220 (N_2220,In_1001,In_603);
or U2221 (N_2221,In_414,In_963);
or U2222 (N_2222,In_967,In_844);
and U2223 (N_2223,In_329,In_231);
nor U2224 (N_2224,In_1451,In_938);
nor U2225 (N_2225,In_1148,In_431);
nand U2226 (N_2226,In_1172,In_1364);
and U2227 (N_2227,In_580,In_45);
nand U2228 (N_2228,In_1264,In_417);
and U2229 (N_2229,In_483,In_614);
and U2230 (N_2230,In_34,In_93);
and U2231 (N_2231,In_1300,In_1158);
nand U2232 (N_2232,In_750,In_1290);
nand U2233 (N_2233,In_878,In_636);
or U2234 (N_2234,In_1403,In_1363);
nor U2235 (N_2235,In_1044,In_384);
nand U2236 (N_2236,In_15,In_333);
and U2237 (N_2237,In_631,In_1129);
or U2238 (N_2238,In_1000,In_1330);
nor U2239 (N_2239,In_284,In_960);
and U2240 (N_2240,In_231,In_530);
xor U2241 (N_2241,In_148,In_407);
nand U2242 (N_2242,In_10,In_947);
nand U2243 (N_2243,In_532,In_21);
nor U2244 (N_2244,In_51,In_1055);
or U2245 (N_2245,In_606,In_1147);
nand U2246 (N_2246,In_803,In_515);
and U2247 (N_2247,In_793,In_531);
nor U2248 (N_2248,In_1243,In_434);
nor U2249 (N_2249,In_584,In_171);
nand U2250 (N_2250,In_853,In_580);
nand U2251 (N_2251,In_94,In_1120);
and U2252 (N_2252,In_777,In_438);
or U2253 (N_2253,In_9,In_1355);
or U2254 (N_2254,In_504,In_584);
nand U2255 (N_2255,In_696,In_109);
nor U2256 (N_2256,In_896,In_1099);
nand U2257 (N_2257,In_1350,In_455);
xnor U2258 (N_2258,In_443,In_261);
nor U2259 (N_2259,In_1296,In_540);
nor U2260 (N_2260,In_107,In_1458);
nor U2261 (N_2261,In_1370,In_868);
xor U2262 (N_2262,In_213,In_593);
or U2263 (N_2263,In_870,In_730);
nand U2264 (N_2264,In_1128,In_222);
or U2265 (N_2265,In_781,In_431);
and U2266 (N_2266,In_732,In_1178);
and U2267 (N_2267,In_1414,In_387);
nand U2268 (N_2268,In_11,In_988);
or U2269 (N_2269,In_84,In_1260);
or U2270 (N_2270,In_250,In_1453);
or U2271 (N_2271,In_632,In_1163);
xnor U2272 (N_2272,In_39,In_1359);
nor U2273 (N_2273,In_443,In_1458);
nand U2274 (N_2274,In_26,In_1263);
or U2275 (N_2275,In_959,In_1111);
or U2276 (N_2276,In_1366,In_211);
xor U2277 (N_2277,In_1307,In_1248);
nand U2278 (N_2278,In_908,In_988);
nor U2279 (N_2279,In_126,In_1265);
and U2280 (N_2280,In_1360,In_702);
nor U2281 (N_2281,In_729,In_940);
and U2282 (N_2282,In_768,In_392);
and U2283 (N_2283,In_1436,In_1038);
and U2284 (N_2284,In_351,In_1191);
nor U2285 (N_2285,In_1251,In_588);
and U2286 (N_2286,In_1435,In_227);
or U2287 (N_2287,In_777,In_212);
xnor U2288 (N_2288,In_1427,In_390);
xor U2289 (N_2289,In_1441,In_950);
or U2290 (N_2290,In_427,In_1491);
xnor U2291 (N_2291,In_1420,In_1312);
nor U2292 (N_2292,In_1123,In_922);
nand U2293 (N_2293,In_77,In_736);
xnor U2294 (N_2294,In_708,In_1281);
or U2295 (N_2295,In_615,In_1431);
or U2296 (N_2296,In_1195,In_867);
nor U2297 (N_2297,In_393,In_1267);
nand U2298 (N_2298,In_1147,In_261);
nor U2299 (N_2299,In_538,In_302);
nor U2300 (N_2300,In_213,In_84);
nand U2301 (N_2301,In_8,In_1146);
nor U2302 (N_2302,In_195,In_265);
nor U2303 (N_2303,In_1219,In_337);
and U2304 (N_2304,In_1014,In_855);
nor U2305 (N_2305,In_1173,In_706);
or U2306 (N_2306,In_1059,In_1459);
or U2307 (N_2307,In_1448,In_1217);
nor U2308 (N_2308,In_820,In_1127);
nor U2309 (N_2309,In_941,In_1264);
nand U2310 (N_2310,In_390,In_751);
xnor U2311 (N_2311,In_639,In_238);
nand U2312 (N_2312,In_15,In_37);
nand U2313 (N_2313,In_1351,In_720);
or U2314 (N_2314,In_1077,In_135);
nor U2315 (N_2315,In_400,In_899);
nand U2316 (N_2316,In_296,In_507);
and U2317 (N_2317,In_133,In_1109);
and U2318 (N_2318,In_1004,In_1375);
and U2319 (N_2319,In_568,In_476);
nor U2320 (N_2320,In_1251,In_1289);
nor U2321 (N_2321,In_54,In_1247);
or U2322 (N_2322,In_486,In_1295);
nor U2323 (N_2323,In_547,In_996);
nor U2324 (N_2324,In_1140,In_1136);
or U2325 (N_2325,In_613,In_52);
nand U2326 (N_2326,In_1076,In_216);
or U2327 (N_2327,In_660,In_400);
nor U2328 (N_2328,In_688,In_391);
nor U2329 (N_2329,In_1429,In_635);
nand U2330 (N_2330,In_1212,In_555);
or U2331 (N_2331,In_1273,In_710);
and U2332 (N_2332,In_1085,In_26);
nand U2333 (N_2333,In_1320,In_151);
xnor U2334 (N_2334,In_1479,In_1107);
or U2335 (N_2335,In_977,In_1421);
nor U2336 (N_2336,In_20,In_1452);
nand U2337 (N_2337,In_1476,In_1407);
nand U2338 (N_2338,In_515,In_1149);
or U2339 (N_2339,In_452,In_891);
xor U2340 (N_2340,In_10,In_402);
and U2341 (N_2341,In_602,In_1374);
and U2342 (N_2342,In_393,In_256);
or U2343 (N_2343,In_717,In_1134);
xor U2344 (N_2344,In_294,In_493);
and U2345 (N_2345,In_1192,In_312);
nor U2346 (N_2346,In_866,In_775);
or U2347 (N_2347,In_251,In_1194);
nor U2348 (N_2348,In_1342,In_1486);
or U2349 (N_2349,In_1299,In_1128);
nor U2350 (N_2350,In_154,In_1027);
or U2351 (N_2351,In_514,In_30);
nor U2352 (N_2352,In_1011,In_27);
or U2353 (N_2353,In_37,In_52);
nand U2354 (N_2354,In_947,In_239);
xor U2355 (N_2355,In_862,In_640);
nand U2356 (N_2356,In_386,In_202);
nor U2357 (N_2357,In_1039,In_708);
nor U2358 (N_2358,In_804,In_42);
xor U2359 (N_2359,In_105,In_372);
nand U2360 (N_2360,In_1170,In_999);
nor U2361 (N_2361,In_1351,In_1060);
nor U2362 (N_2362,In_610,In_484);
or U2363 (N_2363,In_947,In_419);
nor U2364 (N_2364,In_159,In_174);
xnor U2365 (N_2365,In_646,In_953);
nor U2366 (N_2366,In_717,In_606);
nand U2367 (N_2367,In_1443,In_449);
and U2368 (N_2368,In_441,In_1336);
nand U2369 (N_2369,In_1068,In_510);
or U2370 (N_2370,In_499,In_384);
or U2371 (N_2371,In_1041,In_272);
xor U2372 (N_2372,In_284,In_735);
nor U2373 (N_2373,In_294,In_1351);
nor U2374 (N_2374,In_406,In_1268);
xnor U2375 (N_2375,In_311,In_553);
nor U2376 (N_2376,In_68,In_1343);
nor U2377 (N_2377,In_965,In_1123);
nor U2378 (N_2378,In_965,In_573);
and U2379 (N_2379,In_980,In_1207);
and U2380 (N_2380,In_1436,In_1043);
nand U2381 (N_2381,In_244,In_1037);
nand U2382 (N_2382,In_1194,In_301);
nor U2383 (N_2383,In_240,In_643);
or U2384 (N_2384,In_1271,In_648);
nor U2385 (N_2385,In_480,In_858);
and U2386 (N_2386,In_541,In_1272);
and U2387 (N_2387,In_602,In_463);
or U2388 (N_2388,In_320,In_450);
nor U2389 (N_2389,In_0,In_1392);
nand U2390 (N_2390,In_1158,In_670);
nor U2391 (N_2391,In_126,In_827);
nor U2392 (N_2392,In_91,In_1162);
nand U2393 (N_2393,In_426,In_665);
or U2394 (N_2394,In_678,In_17);
nand U2395 (N_2395,In_939,In_1316);
and U2396 (N_2396,In_1246,In_1451);
nand U2397 (N_2397,In_1164,In_1390);
and U2398 (N_2398,In_1081,In_69);
or U2399 (N_2399,In_522,In_1331);
nand U2400 (N_2400,In_201,In_1460);
nor U2401 (N_2401,In_145,In_1258);
nor U2402 (N_2402,In_1333,In_1272);
nor U2403 (N_2403,In_1032,In_70);
and U2404 (N_2404,In_1226,In_473);
and U2405 (N_2405,In_1460,In_1393);
nor U2406 (N_2406,In_1133,In_180);
and U2407 (N_2407,In_429,In_466);
and U2408 (N_2408,In_1007,In_1258);
or U2409 (N_2409,In_1296,In_1360);
nor U2410 (N_2410,In_377,In_1356);
nor U2411 (N_2411,In_810,In_773);
nand U2412 (N_2412,In_691,In_965);
or U2413 (N_2413,In_1310,In_835);
nor U2414 (N_2414,In_895,In_806);
or U2415 (N_2415,In_532,In_582);
nand U2416 (N_2416,In_455,In_928);
and U2417 (N_2417,In_871,In_420);
nand U2418 (N_2418,In_182,In_493);
nor U2419 (N_2419,In_1207,In_81);
or U2420 (N_2420,In_10,In_1033);
nor U2421 (N_2421,In_412,In_953);
nand U2422 (N_2422,In_589,In_1456);
and U2423 (N_2423,In_836,In_1190);
and U2424 (N_2424,In_176,In_130);
and U2425 (N_2425,In_156,In_17);
xor U2426 (N_2426,In_104,In_1094);
and U2427 (N_2427,In_175,In_1414);
or U2428 (N_2428,In_962,In_221);
nor U2429 (N_2429,In_1395,In_1191);
nand U2430 (N_2430,In_684,In_36);
or U2431 (N_2431,In_1039,In_343);
and U2432 (N_2432,In_1040,In_1081);
or U2433 (N_2433,In_505,In_1339);
nand U2434 (N_2434,In_1054,In_155);
xor U2435 (N_2435,In_577,In_735);
nand U2436 (N_2436,In_340,In_271);
nor U2437 (N_2437,In_110,In_364);
or U2438 (N_2438,In_1161,In_544);
or U2439 (N_2439,In_244,In_661);
xor U2440 (N_2440,In_437,In_821);
and U2441 (N_2441,In_753,In_191);
or U2442 (N_2442,In_1421,In_636);
xnor U2443 (N_2443,In_505,In_768);
and U2444 (N_2444,In_1468,In_432);
nand U2445 (N_2445,In_159,In_1286);
and U2446 (N_2446,In_1083,In_427);
nor U2447 (N_2447,In_704,In_1433);
nand U2448 (N_2448,In_96,In_1196);
nor U2449 (N_2449,In_1196,In_671);
and U2450 (N_2450,In_1430,In_1139);
nand U2451 (N_2451,In_1375,In_1328);
nor U2452 (N_2452,In_816,In_393);
or U2453 (N_2453,In_37,In_1399);
nor U2454 (N_2454,In_225,In_593);
xor U2455 (N_2455,In_718,In_260);
or U2456 (N_2456,In_71,In_564);
nor U2457 (N_2457,In_726,In_1203);
nand U2458 (N_2458,In_940,In_318);
nand U2459 (N_2459,In_1411,In_788);
nand U2460 (N_2460,In_252,In_241);
and U2461 (N_2461,In_1102,In_1211);
and U2462 (N_2462,In_915,In_364);
and U2463 (N_2463,In_770,In_476);
nand U2464 (N_2464,In_1359,In_142);
nor U2465 (N_2465,In_1249,In_1179);
nor U2466 (N_2466,In_452,In_1004);
or U2467 (N_2467,In_856,In_590);
or U2468 (N_2468,In_173,In_220);
nor U2469 (N_2469,In_172,In_970);
and U2470 (N_2470,In_858,In_446);
xnor U2471 (N_2471,In_1355,In_67);
or U2472 (N_2472,In_309,In_1186);
and U2473 (N_2473,In_654,In_1373);
or U2474 (N_2474,In_23,In_576);
xnor U2475 (N_2475,In_341,In_46);
nor U2476 (N_2476,In_1380,In_695);
and U2477 (N_2477,In_1328,In_968);
and U2478 (N_2478,In_1078,In_657);
nand U2479 (N_2479,In_690,In_917);
or U2480 (N_2480,In_887,In_422);
and U2481 (N_2481,In_1371,In_335);
and U2482 (N_2482,In_586,In_1486);
nand U2483 (N_2483,In_30,In_1471);
or U2484 (N_2484,In_394,In_212);
and U2485 (N_2485,In_1447,In_599);
or U2486 (N_2486,In_460,In_714);
or U2487 (N_2487,In_1248,In_208);
or U2488 (N_2488,In_878,In_817);
nand U2489 (N_2489,In_464,In_737);
nand U2490 (N_2490,In_953,In_800);
nor U2491 (N_2491,In_1011,In_247);
and U2492 (N_2492,In_1045,In_222);
nor U2493 (N_2493,In_189,In_246);
xor U2494 (N_2494,In_848,In_1019);
xnor U2495 (N_2495,In_673,In_17);
nor U2496 (N_2496,In_1041,In_70);
nor U2497 (N_2497,In_265,In_1083);
and U2498 (N_2498,In_935,In_993);
nand U2499 (N_2499,In_84,In_46);
or U2500 (N_2500,In_248,In_1001);
xnor U2501 (N_2501,In_433,In_751);
nand U2502 (N_2502,In_818,In_442);
or U2503 (N_2503,In_1437,In_214);
and U2504 (N_2504,In_160,In_977);
nand U2505 (N_2505,In_498,In_1380);
and U2506 (N_2506,In_181,In_749);
or U2507 (N_2507,In_1045,In_236);
and U2508 (N_2508,In_581,In_776);
or U2509 (N_2509,In_1366,In_352);
nand U2510 (N_2510,In_1031,In_873);
nand U2511 (N_2511,In_1043,In_638);
and U2512 (N_2512,In_1414,In_903);
and U2513 (N_2513,In_244,In_1272);
or U2514 (N_2514,In_391,In_1107);
xnor U2515 (N_2515,In_1284,In_1123);
nor U2516 (N_2516,In_1342,In_1212);
xor U2517 (N_2517,In_1009,In_1047);
and U2518 (N_2518,In_356,In_327);
nor U2519 (N_2519,In_405,In_1224);
or U2520 (N_2520,In_926,In_1417);
or U2521 (N_2521,In_409,In_600);
and U2522 (N_2522,In_1453,In_138);
and U2523 (N_2523,In_1333,In_1064);
nand U2524 (N_2524,In_1400,In_26);
nand U2525 (N_2525,In_89,In_88);
or U2526 (N_2526,In_1003,In_586);
or U2527 (N_2527,In_599,In_735);
or U2528 (N_2528,In_1170,In_62);
nor U2529 (N_2529,In_1184,In_641);
or U2530 (N_2530,In_791,In_1059);
and U2531 (N_2531,In_1059,In_825);
xor U2532 (N_2532,In_767,In_1486);
and U2533 (N_2533,In_1199,In_1361);
nand U2534 (N_2534,In_1082,In_1328);
nand U2535 (N_2535,In_1194,In_851);
or U2536 (N_2536,In_688,In_846);
and U2537 (N_2537,In_1117,In_740);
or U2538 (N_2538,In_91,In_1207);
nand U2539 (N_2539,In_890,In_1208);
or U2540 (N_2540,In_149,In_933);
nor U2541 (N_2541,In_1061,In_910);
nand U2542 (N_2542,In_1047,In_44);
and U2543 (N_2543,In_1136,In_402);
nor U2544 (N_2544,In_341,In_1364);
nand U2545 (N_2545,In_844,In_880);
xnor U2546 (N_2546,In_1351,In_124);
and U2547 (N_2547,In_778,In_602);
nand U2548 (N_2548,In_1053,In_691);
nor U2549 (N_2549,In_1158,In_546);
or U2550 (N_2550,In_975,In_788);
nand U2551 (N_2551,In_537,In_618);
nor U2552 (N_2552,In_666,In_1155);
nor U2553 (N_2553,In_713,In_1038);
nor U2554 (N_2554,In_48,In_160);
nor U2555 (N_2555,In_749,In_674);
nor U2556 (N_2556,In_1066,In_682);
nand U2557 (N_2557,In_639,In_519);
nand U2558 (N_2558,In_991,In_128);
nor U2559 (N_2559,In_659,In_623);
and U2560 (N_2560,In_669,In_796);
nor U2561 (N_2561,In_1310,In_566);
or U2562 (N_2562,In_503,In_134);
xor U2563 (N_2563,In_1056,In_661);
xor U2564 (N_2564,In_754,In_1297);
and U2565 (N_2565,In_1008,In_638);
and U2566 (N_2566,In_1468,In_30);
nor U2567 (N_2567,In_48,In_1061);
nor U2568 (N_2568,In_1267,In_915);
or U2569 (N_2569,In_588,In_244);
or U2570 (N_2570,In_1373,In_411);
nor U2571 (N_2571,In_790,In_879);
nand U2572 (N_2572,In_466,In_376);
and U2573 (N_2573,In_960,In_1000);
xor U2574 (N_2574,In_195,In_1473);
nor U2575 (N_2575,In_950,In_539);
nand U2576 (N_2576,In_427,In_302);
xor U2577 (N_2577,In_303,In_1004);
and U2578 (N_2578,In_362,In_253);
nor U2579 (N_2579,In_666,In_795);
or U2580 (N_2580,In_887,In_931);
or U2581 (N_2581,In_444,In_926);
or U2582 (N_2582,In_58,In_325);
and U2583 (N_2583,In_1047,In_1289);
nor U2584 (N_2584,In_923,In_1182);
and U2585 (N_2585,In_1353,In_779);
and U2586 (N_2586,In_397,In_1230);
or U2587 (N_2587,In_205,In_1363);
nor U2588 (N_2588,In_764,In_225);
or U2589 (N_2589,In_551,In_1394);
nand U2590 (N_2590,In_780,In_616);
nor U2591 (N_2591,In_917,In_651);
nand U2592 (N_2592,In_855,In_1051);
or U2593 (N_2593,In_783,In_850);
nor U2594 (N_2594,In_258,In_1380);
xnor U2595 (N_2595,In_742,In_252);
and U2596 (N_2596,In_654,In_408);
and U2597 (N_2597,In_1388,In_969);
nor U2598 (N_2598,In_1498,In_35);
nand U2599 (N_2599,In_1338,In_1001);
nor U2600 (N_2600,In_313,In_250);
nor U2601 (N_2601,In_1244,In_468);
or U2602 (N_2602,In_631,In_1163);
xnor U2603 (N_2603,In_941,In_1024);
xnor U2604 (N_2604,In_1027,In_802);
and U2605 (N_2605,In_1498,In_1409);
nor U2606 (N_2606,In_529,In_530);
nor U2607 (N_2607,In_575,In_86);
nor U2608 (N_2608,In_1380,In_1496);
nand U2609 (N_2609,In_732,In_1318);
nand U2610 (N_2610,In_3,In_581);
and U2611 (N_2611,In_461,In_1053);
or U2612 (N_2612,In_1059,In_311);
or U2613 (N_2613,In_737,In_729);
nand U2614 (N_2614,In_107,In_903);
or U2615 (N_2615,In_1054,In_174);
and U2616 (N_2616,In_733,In_606);
nand U2617 (N_2617,In_857,In_1266);
or U2618 (N_2618,In_235,In_256);
nor U2619 (N_2619,In_576,In_241);
and U2620 (N_2620,In_1218,In_189);
and U2621 (N_2621,In_380,In_475);
nand U2622 (N_2622,In_894,In_1113);
nor U2623 (N_2623,In_446,In_1067);
or U2624 (N_2624,In_1140,In_449);
xor U2625 (N_2625,In_270,In_1425);
xnor U2626 (N_2626,In_1317,In_1447);
or U2627 (N_2627,In_1213,In_954);
and U2628 (N_2628,In_451,In_570);
and U2629 (N_2629,In_1072,In_1268);
nor U2630 (N_2630,In_587,In_624);
or U2631 (N_2631,In_462,In_1439);
or U2632 (N_2632,In_8,In_338);
or U2633 (N_2633,In_435,In_475);
or U2634 (N_2634,In_962,In_314);
or U2635 (N_2635,In_1468,In_1489);
nand U2636 (N_2636,In_1070,In_62);
and U2637 (N_2637,In_113,In_486);
nor U2638 (N_2638,In_1469,In_1033);
or U2639 (N_2639,In_39,In_595);
nor U2640 (N_2640,In_47,In_1039);
nand U2641 (N_2641,In_619,In_12);
nor U2642 (N_2642,In_127,In_221);
nand U2643 (N_2643,In_355,In_855);
or U2644 (N_2644,In_1149,In_588);
nand U2645 (N_2645,In_1092,In_978);
and U2646 (N_2646,In_1153,In_929);
or U2647 (N_2647,In_1476,In_649);
or U2648 (N_2648,In_1378,In_1105);
xor U2649 (N_2649,In_1020,In_713);
or U2650 (N_2650,In_395,In_1234);
or U2651 (N_2651,In_609,In_372);
or U2652 (N_2652,In_232,In_116);
nor U2653 (N_2653,In_1415,In_390);
or U2654 (N_2654,In_788,In_1134);
nor U2655 (N_2655,In_665,In_618);
and U2656 (N_2656,In_209,In_30);
and U2657 (N_2657,In_384,In_1294);
or U2658 (N_2658,In_290,In_548);
nor U2659 (N_2659,In_1372,In_564);
and U2660 (N_2660,In_1372,In_216);
and U2661 (N_2661,In_1155,In_966);
and U2662 (N_2662,In_450,In_352);
or U2663 (N_2663,In_213,In_1381);
nand U2664 (N_2664,In_73,In_21);
nor U2665 (N_2665,In_172,In_57);
and U2666 (N_2666,In_220,In_74);
and U2667 (N_2667,In_1051,In_527);
xor U2668 (N_2668,In_349,In_188);
nor U2669 (N_2669,In_36,In_874);
or U2670 (N_2670,In_948,In_1099);
or U2671 (N_2671,In_679,In_1330);
and U2672 (N_2672,In_1479,In_680);
nand U2673 (N_2673,In_1383,In_1288);
nor U2674 (N_2674,In_313,In_1338);
and U2675 (N_2675,In_958,In_72);
nand U2676 (N_2676,In_1007,In_663);
or U2677 (N_2677,In_52,In_1401);
or U2678 (N_2678,In_191,In_1288);
nor U2679 (N_2679,In_1482,In_605);
nor U2680 (N_2680,In_377,In_75);
and U2681 (N_2681,In_863,In_1422);
nor U2682 (N_2682,In_14,In_788);
nor U2683 (N_2683,In_799,In_686);
xnor U2684 (N_2684,In_1271,In_290);
xnor U2685 (N_2685,In_407,In_1333);
and U2686 (N_2686,In_1363,In_1356);
nor U2687 (N_2687,In_1479,In_753);
and U2688 (N_2688,In_928,In_509);
nor U2689 (N_2689,In_1032,In_333);
nor U2690 (N_2690,In_778,In_264);
or U2691 (N_2691,In_973,In_1245);
nor U2692 (N_2692,In_1016,In_1381);
or U2693 (N_2693,In_558,In_1380);
nand U2694 (N_2694,In_186,In_835);
nand U2695 (N_2695,In_3,In_1323);
and U2696 (N_2696,In_1490,In_432);
or U2697 (N_2697,In_810,In_800);
xor U2698 (N_2698,In_924,In_963);
or U2699 (N_2699,In_1078,In_959);
or U2700 (N_2700,In_690,In_797);
nand U2701 (N_2701,In_1098,In_44);
xor U2702 (N_2702,In_946,In_638);
nand U2703 (N_2703,In_913,In_142);
xor U2704 (N_2704,In_168,In_1269);
xnor U2705 (N_2705,In_664,In_1423);
nor U2706 (N_2706,In_13,In_158);
and U2707 (N_2707,In_978,In_976);
nor U2708 (N_2708,In_211,In_582);
nor U2709 (N_2709,In_1075,In_1116);
or U2710 (N_2710,In_791,In_77);
and U2711 (N_2711,In_197,In_1329);
and U2712 (N_2712,In_1105,In_1376);
nand U2713 (N_2713,In_1120,In_1474);
and U2714 (N_2714,In_784,In_181);
or U2715 (N_2715,In_1317,In_1082);
or U2716 (N_2716,In_563,In_1258);
or U2717 (N_2717,In_682,In_1423);
nand U2718 (N_2718,In_1425,In_792);
and U2719 (N_2719,In_951,In_1309);
and U2720 (N_2720,In_1259,In_1449);
or U2721 (N_2721,In_1039,In_1264);
nor U2722 (N_2722,In_1182,In_1054);
and U2723 (N_2723,In_623,In_872);
or U2724 (N_2724,In_583,In_839);
nor U2725 (N_2725,In_854,In_892);
and U2726 (N_2726,In_491,In_234);
and U2727 (N_2727,In_481,In_1230);
or U2728 (N_2728,In_448,In_686);
nand U2729 (N_2729,In_1152,In_402);
or U2730 (N_2730,In_1412,In_275);
or U2731 (N_2731,In_710,In_1343);
nand U2732 (N_2732,In_377,In_364);
and U2733 (N_2733,In_241,In_1083);
nand U2734 (N_2734,In_688,In_1201);
nand U2735 (N_2735,In_981,In_1406);
nand U2736 (N_2736,In_1414,In_602);
and U2737 (N_2737,In_531,In_1310);
nor U2738 (N_2738,In_515,In_1249);
nor U2739 (N_2739,In_710,In_622);
or U2740 (N_2740,In_430,In_1480);
and U2741 (N_2741,In_144,In_1036);
and U2742 (N_2742,In_1047,In_204);
nand U2743 (N_2743,In_1351,In_1287);
nor U2744 (N_2744,In_1439,In_341);
nor U2745 (N_2745,In_1070,In_397);
and U2746 (N_2746,In_538,In_831);
and U2747 (N_2747,In_228,In_729);
nand U2748 (N_2748,In_968,In_1258);
or U2749 (N_2749,In_1308,In_578);
or U2750 (N_2750,In_917,In_471);
or U2751 (N_2751,In_35,In_1205);
and U2752 (N_2752,In_113,In_1028);
nor U2753 (N_2753,In_734,In_502);
and U2754 (N_2754,In_840,In_143);
nor U2755 (N_2755,In_1325,In_1007);
and U2756 (N_2756,In_887,In_893);
nor U2757 (N_2757,In_168,In_1420);
and U2758 (N_2758,In_1411,In_1478);
nor U2759 (N_2759,In_1067,In_101);
nor U2760 (N_2760,In_700,In_929);
nor U2761 (N_2761,In_516,In_465);
and U2762 (N_2762,In_101,In_1226);
or U2763 (N_2763,In_373,In_321);
nor U2764 (N_2764,In_1184,In_1261);
nor U2765 (N_2765,In_627,In_635);
nor U2766 (N_2766,In_998,In_393);
and U2767 (N_2767,In_644,In_1460);
or U2768 (N_2768,In_819,In_1326);
nand U2769 (N_2769,In_499,In_874);
or U2770 (N_2770,In_357,In_430);
nor U2771 (N_2771,In_569,In_546);
nand U2772 (N_2772,In_135,In_312);
and U2773 (N_2773,In_617,In_413);
or U2774 (N_2774,In_76,In_1053);
xor U2775 (N_2775,In_220,In_392);
nor U2776 (N_2776,In_891,In_515);
xnor U2777 (N_2777,In_748,In_1365);
and U2778 (N_2778,In_1123,In_1062);
nand U2779 (N_2779,In_928,In_903);
nand U2780 (N_2780,In_1250,In_812);
and U2781 (N_2781,In_141,In_126);
and U2782 (N_2782,In_1275,In_1040);
xnor U2783 (N_2783,In_84,In_584);
nand U2784 (N_2784,In_1403,In_1228);
or U2785 (N_2785,In_519,In_110);
or U2786 (N_2786,In_143,In_20);
nand U2787 (N_2787,In_779,In_1068);
and U2788 (N_2788,In_47,In_640);
and U2789 (N_2789,In_545,In_125);
or U2790 (N_2790,In_759,In_599);
nand U2791 (N_2791,In_676,In_547);
nor U2792 (N_2792,In_1028,In_1204);
or U2793 (N_2793,In_698,In_353);
nand U2794 (N_2794,In_692,In_1495);
nor U2795 (N_2795,In_1150,In_71);
nand U2796 (N_2796,In_816,In_1189);
xor U2797 (N_2797,In_600,In_507);
nand U2798 (N_2798,In_303,In_9);
nand U2799 (N_2799,In_329,In_198);
or U2800 (N_2800,In_198,In_648);
or U2801 (N_2801,In_1390,In_1230);
nand U2802 (N_2802,In_132,In_1024);
or U2803 (N_2803,In_160,In_784);
nand U2804 (N_2804,In_361,In_900);
nor U2805 (N_2805,In_389,In_736);
nand U2806 (N_2806,In_109,In_190);
and U2807 (N_2807,In_1201,In_664);
nand U2808 (N_2808,In_223,In_626);
or U2809 (N_2809,In_1414,In_104);
or U2810 (N_2810,In_727,In_763);
nand U2811 (N_2811,In_1192,In_177);
nor U2812 (N_2812,In_1145,In_940);
or U2813 (N_2813,In_1262,In_186);
or U2814 (N_2814,In_1344,In_1413);
and U2815 (N_2815,In_717,In_1060);
and U2816 (N_2816,In_289,In_957);
nand U2817 (N_2817,In_525,In_599);
xor U2818 (N_2818,In_600,In_1265);
or U2819 (N_2819,In_1044,In_896);
or U2820 (N_2820,In_454,In_707);
nand U2821 (N_2821,In_962,In_383);
nand U2822 (N_2822,In_399,In_340);
nor U2823 (N_2823,In_646,In_124);
and U2824 (N_2824,In_1037,In_627);
xor U2825 (N_2825,In_1279,In_1048);
xor U2826 (N_2826,In_1126,In_1437);
nand U2827 (N_2827,In_951,In_973);
nor U2828 (N_2828,In_947,In_1344);
nand U2829 (N_2829,In_214,In_264);
xor U2830 (N_2830,In_1196,In_754);
or U2831 (N_2831,In_1106,In_15);
and U2832 (N_2832,In_265,In_979);
and U2833 (N_2833,In_1348,In_1020);
and U2834 (N_2834,In_288,In_256);
and U2835 (N_2835,In_1382,In_685);
xor U2836 (N_2836,In_995,In_179);
and U2837 (N_2837,In_1272,In_52);
nor U2838 (N_2838,In_902,In_1039);
or U2839 (N_2839,In_439,In_1369);
and U2840 (N_2840,In_1150,In_173);
xnor U2841 (N_2841,In_969,In_1208);
and U2842 (N_2842,In_333,In_981);
nand U2843 (N_2843,In_888,In_501);
and U2844 (N_2844,In_545,In_166);
and U2845 (N_2845,In_1056,In_806);
or U2846 (N_2846,In_121,In_443);
or U2847 (N_2847,In_1341,In_1162);
nand U2848 (N_2848,In_37,In_566);
nand U2849 (N_2849,In_135,In_1140);
and U2850 (N_2850,In_653,In_127);
nor U2851 (N_2851,In_405,In_568);
and U2852 (N_2852,In_859,In_1495);
xor U2853 (N_2853,In_444,In_167);
or U2854 (N_2854,In_1373,In_811);
xor U2855 (N_2855,In_939,In_91);
nor U2856 (N_2856,In_786,In_1127);
xor U2857 (N_2857,In_1048,In_142);
nand U2858 (N_2858,In_707,In_864);
nor U2859 (N_2859,In_930,In_34);
nand U2860 (N_2860,In_742,In_802);
xor U2861 (N_2861,In_1126,In_530);
xnor U2862 (N_2862,In_1162,In_1096);
nand U2863 (N_2863,In_648,In_1270);
nor U2864 (N_2864,In_91,In_768);
xnor U2865 (N_2865,In_949,In_1434);
or U2866 (N_2866,In_1292,In_754);
nor U2867 (N_2867,In_841,In_934);
and U2868 (N_2868,In_491,In_141);
xor U2869 (N_2869,In_1037,In_614);
nor U2870 (N_2870,In_984,In_1428);
or U2871 (N_2871,In_82,In_676);
nand U2872 (N_2872,In_816,In_1066);
nand U2873 (N_2873,In_63,In_1050);
and U2874 (N_2874,In_1490,In_1005);
or U2875 (N_2875,In_26,In_1096);
and U2876 (N_2876,In_192,In_1390);
or U2877 (N_2877,In_1328,In_875);
nor U2878 (N_2878,In_998,In_881);
xnor U2879 (N_2879,In_1166,In_180);
nand U2880 (N_2880,In_1194,In_95);
or U2881 (N_2881,In_4,In_89);
nand U2882 (N_2882,In_1114,In_253);
xnor U2883 (N_2883,In_852,In_1412);
nand U2884 (N_2884,In_1199,In_513);
nor U2885 (N_2885,In_399,In_384);
nor U2886 (N_2886,In_1208,In_105);
nor U2887 (N_2887,In_1378,In_518);
nor U2888 (N_2888,In_345,In_1092);
or U2889 (N_2889,In_1341,In_912);
and U2890 (N_2890,In_354,In_518);
and U2891 (N_2891,In_345,In_1349);
and U2892 (N_2892,In_60,In_1068);
and U2893 (N_2893,In_486,In_206);
and U2894 (N_2894,In_13,In_1403);
xnor U2895 (N_2895,In_1002,In_1492);
nand U2896 (N_2896,In_1126,In_611);
nand U2897 (N_2897,In_1183,In_1171);
or U2898 (N_2898,In_690,In_939);
and U2899 (N_2899,In_324,In_318);
and U2900 (N_2900,In_217,In_785);
and U2901 (N_2901,In_259,In_780);
nand U2902 (N_2902,In_1347,In_1176);
nand U2903 (N_2903,In_1305,In_102);
and U2904 (N_2904,In_934,In_1065);
or U2905 (N_2905,In_1249,In_628);
nand U2906 (N_2906,In_924,In_1383);
nand U2907 (N_2907,In_28,In_579);
and U2908 (N_2908,In_1033,In_300);
or U2909 (N_2909,In_975,In_656);
nor U2910 (N_2910,In_89,In_442);
nand U2911 (N_2911,In_1334,In_1038);
and U2912 (N_2912,In_1079,In_187);
nor U2913 (N_2913,In_779,In_842);
and U2914 (N_2914,In_808,In_448);
and U2915 (N_2915,In_230,In_262);
nor U2916 (N_2916,In_1198,In_1024);
nor U2917 (N_2917,In_365,In_950);
nand U2918 (N_2918,In_737,In_1357);
nor U2919 (N_2919,In_1394,In_315);
and U2920 (N_2920,In_1330,In_1413);
nand U2921 (N_2921,In_273,In_784);
nand U2922 (N_2922,In_1418,In_622);
nand U2923 (N_2923,In_1299,In_728);
nor U2924 (N_2924,In_80,In_1131);
and U2925 (N_2925,In_1477,In_1101);
nor U2926 (N_2926,In_1426,In_1359);
and U2927 (N_2927,In_382,In_1259);
and U2928 (N_2928,In_1073,In_631);
or U2929 (N_2929,In_654,In_147);
or U2930 (N_2930,In_1434,In_1169);
nand U2931 (N_2931,In_553,In_448);
nand U2932 (N_2932,In_549,In_1236);
and U2933 (N_2933,In_806,In_1026);
and U2934 (N_2934,In_234,In_572);
nor U2935 (N_2935,In_254,In_85);
and U2936 (N_2936,In_389,In_582);
nand U2937 (N_2937,In_1001,In_431);
nor U2938 (N_2938,In_8,In_1492);
or U2939 (N_2939,In_1436,In_885);
or U2940 (N_2940,In_255,In_1345);
or U2941 (N_2941,In_929,In_1078);
nand U2942 (N_2942,In_832,In_113);
or U2943 (N_2943,In_334,In_400);
nand U2944 (N_2944,In_1396,In_1454);
nor U2945 (N_2945,In_983,In_1356);
and U2946 (N_2946,In_976,In_614);
or U2947 (N_2947,In_912,In_658);
nand U2948 (N_2948,In_143,In_118);
or U2949 (N_2949,In_70,In_374);
or U2950 (N_2950,In_1274,In_60);
and U2951 (N_2951,In_1203,In_104);
or U2952 (N_2952,In_954,In_1227);
nand U2953 (N_2953,In_676,In_703);
and U2954 (N_2954,In_10,In_656);
nand U2955 (N_2955,In_153,In_347);
and U2956 (N_2956,In_1490,In_612);
or U2957 (N_2957,In_952,In_396);
nand U2958 (N_2958,In_709,In_1170);
xnor U2959 (N_2959,In_1028,In_1224);
and U2960 (N_2960,In_1226,In_1123);
or U2961 (N_2961,In_1000,In_1047);
xnor U2962 (N_2962,In_1216,In_264);
or U2963 (N_2963,In_666,In_1434);
xor U2964 (N_2964,In_821,In_1417);
nor U2965 (N_2965,In_998,In_807);
and U2966 (N_2966,In_901,In_489);
or U2967 (N_2967,In_1108,In_222);
nor U2968 (N_2968,In_237,In_1339);
nand U2969 (N_2969,In_161,In_695);
or U2970 (N_2970,In_563,In_950);
and U2971 (N_2971,In_362,In_255);
nor U2972 (N_2972,In_1212,In_69);
nand U2973 (N_2973,In_1415,In_186);
xor U2974 (N_2974,In_1166,In_364);
xnor U2975 (N_2975,In_24,In_1367);
nand U2976 (N_2976,In_171,In_1149);
xor U2977 (N_2977,In_644,In_414);
xnor U2978 (N_2978,In_1285,In_310);
nand U2979 (N_2979,In_126,In_1488);
and U2980 (N_2980,In_205,In_729);
nor U2981 (N_2981,In_1420,In_1268);
nor U2982 (N_2982,In_311,In_1385);
or U2983 (N_2983,In_1152,In_901);
or U2984 (N_2984,In_1239,In_447);
nor U2985 (N_2985,In_1075,In_238);
and U2986 (N_2986,In_733,In_1492);
and U2987 (N_2987,In_285,In_368);
or U2988 (N_2988,In_1287,In_607);
and U2989 (N_2989,In_396,In_63);
nand U2990 (N_2990,In_359,In_1487);
xor U2991 (N_2991,In_116,In_1140);
nand U2992 (N_2992,In_927,In_453);
nor U2993 (N_2993,In_754,In_1431);
nor U2994 (N_2994,In_277,In_1398);
and U2995 (N_2995,In_943,In_1170);
or U2996 (N_2996,In_789,In_1094);
nor U2997 (N_2997,In_532,In_950);
and U2998 (N_2998,In_776,In_1053);
nand U2999 (N_2999,In_482,In_631);
nand U3000 (N_3000,In_1411,In_643);
xnor U3001 (N_3001,In_1448,In_97);
and U3002 (N_3002,In_600,In_920);
nand U3003 (N_3003,In_286,In_1219);
nor U3004 (N_3004,In_772,In_362);
xor U3005 (N_3005,In_445,In_991);
and U3006 (N_3006,In_350,In_508);
and U3007 (N_3007,In_1088,In_980);
or U3008 (N_3008,In_1449,In_387);
nor U3009 (N_3009,In_590,In_799);
nor U3010 (N_3010,In_202,In_1195);
nor U3011 (N_3011,In_963,In_216);
nor U3012 (N_3012,In_521,In_286);
nand U3013 (N_3013,In_1469,In_636);
nor U3014 (N_3014,In_488,In_15);
and U3015 (N_3015,In_654,In_469);
and U3016 (N_3016,In_942,In_1026);
nand U3017 (N_3017,In_945,In_836);
and U3018 (N_3018,In_734,In_703);
nor U3019 (N_3019,In_1159,In_79);
nor U3020 (N_3020,In_615,In_450);
nand U3021 (N_3021,In_654,In_594);
nand U3022 (N_3022,In_1034,In_917);
or U3023 (N_3023,In_1425,In_598);
nand U3024 (N_3024,In_1141,In_799);
or U3025 (N_3025,In_193,In_819);
nand U3026 (N_3026,In_84,In_782);
and U3027 (N_3027,In_463,In_437);
nand U3028 (N_3028,In_423,In_752);
nor U3029 (N_3029,In_1298,In_1386);
nand U3030 (N_3030,In_645,In_302);
or U3031 (N_3031,In_1176,In_764);
nand U3032 (N_3032,In_784,In_374);
xnor U3033 (N_3033,In_388,In_307);
nor U3034 (N_3034,In_563,In_432);
nand U3035 (N_3035,In_1469,In_238);
or U3036 (N_3036,In_630,In_854);
and U3037 (N_3037,In_523,In_1093);
or U3038 (N_3038,In_966,In_895);
and U3039 (N_3039,In_890,In_750);
nand U3040 (N_3040,In_1187,In_1157);
and U3041 (N_3041,In_1462,In_1027);
nand U3042 (N_3042,In_194,In_857);
nor U3043 (N_3043,In_1413,In_827);
nor U3044 (N_3044,In_392,In_1261);
nand U3045 (N_3045,In_887,In_1214);
and U3046 (N_3046,In_1254,In_954);
xnor U3047 (N_3047,In_823,In_226);
and U3048 (N_3048,In_1186,In_677);
xnor U3049 (N_3049,In_239,In_594);
or U3050 (N_3050,In_1255,In_1412);
and U3051 (N_3051,In_1070,In_144);
and U3052 (N_3052,In_441,In_847);
nor U3053 (N_3053,In_657,In_1158);
or U3054 (N_3054,In_868,In_540);
nand U3055 (N_3055,In_1320,In_1301);
xor U3056 (N_3056,In_1207,In_9);
nor U3057 (N_3057,In_455,In_650);
nand U3058 (N_3058,In_1274,In_1001);
nor U3059 (N_3059,In_256,In_601);
nor U3060 (N_3060,In_646,In_587);
or U3061 (N_3061,In_710,In_873);
nor U3062 (N_3062,In_596,In_727);
and U3063 (N_3063,In_527,In_348);
xor U3064 (N_3064,In_1383,In_496);
nand U3065 (N_3065,In_57,In_719);
and U3066 (N_3066,In_980,In_1043);
nor U3067 (N_3067,In_1321,In_891);
nand U3068 (N_3068,In_486,In_1027);
nor U3069 (N_3069,In_1422,In_1146);
and U3070 (N_3070,In_1149,In_1049);
xnor U3071 (N_3071,In_1300,In_565);
xor U3072 (N_3072,In_1237,In_1004);
and U3073 (N_3073,In_656,In_373);
or U3074 (N_3074,In_1005,In_530);
xor U3075 (N_3075,In_767,In_589);
and U3076 (N_3076,In_138,In_361);
and U3077 (N_3077,In_947,In_1291);
nand U3078 (N_3078,In_1073,In_696);
nor U3079 (N_3079,In_1104,In_382);
and U3080 (N_3080,In_659,In_1029);
nand U3081 (N_3081,In_1392,In_1390);
nor U3082 (N_3082,In_588,In_1465);
nor U3083 (N_3083,In_1030,In_207);
or U3084 (N_3084,In_839,In_577);
nor U3085 (N_3085,In_285,In_816);
or U3086 (N_3086,In_1465,In_569);
nand U3087 (N_3087,In_353,In_1291);
nand U3088 (N_3088,In_190,In_799);
or U3089 (N_3089,In_919,In_1493);
xor U3090 (N_3090,In_698,In_369);
or U3091 (N_3091,In_1069,In_1177);
and U3092 (N_3092,In_197,In_478);
nor U3093 (N_3093,In_1388,In_1479);
nor U3094 (N_3094,In_329,In_1271);
xor U3095 (N_3095,In_905,In_175);
and U3096 (N_3096,In_727,In_1224);
and U3097 (N_3097,In_1383,In_85);
xnor U3098 (N_3098,In_1463,In_337);
and U3099 (N_3099,In_668,In_1192);
xnor U3100 (N_3100,In_1048,In_293);
and U3101 (N_3101,In_400,In_907);
and U3102 (N_3102,In_923,In_340);
nand U3103 (N_3103,In_1027,In_811);
and U3104 (N_3104,In_1233,In_170);
nand U3105 (N_3105,In_278,In_1352);
or U3106 (N_3106,In_210,In_710);
and U3107 (N_3107,In_316,In_541);
xor U3108 (N_3108,In_161,In_1345);
nand U3109 (N_3109,In_123,In_607);
xnor U3110 (N_3110,In_1408,In_1158);
and U3111 (N_3111,In_127,In_87);
and U3112 (N_3112,In_5,In_1325);
nor U3113 (N_3113,In_1305,In_891);
nor U3114 (N_3114,In_255,In_1065);
or U3115 (N_3115,In_1272,In_197);
and U3116 (N_3116,In_1178,In_1099);
and U3117 (N_3117,In_1478,In_1249);
nor U3118 (N_3118,In_751,In_575);
xnor U3119 (N_3119,In_35,In_608);
or U3120 (N_3120,In_206,In_1311);
or U3121 (N_3121,In_760,In_1142);
xnor U3122 (N_3122,In_158,In_233);
nor U3123 (N_3123,In_771,In_761);
and U3124 (N_3124,In_958,In_259);
nor U3125 (N_3125,In_351,In_456);
and U3126 (N_3126,In_1391,In_495);
nor U3127 (N_3127,In_141,In_241);
nand U3128 (N_3128,In_163,In_1455);
nor U3129 (N_3129,In_1264,In_1358);
and U3130 (N_3130,In_334,In_183);
nor U3131 (N_3131,In_819,In_828);
or U3132 (N_3132,In_1453,In_481);
nand U3133 (N_3133,In_930,In_719);
or U3134 (N_3134,In_1345,In_1492);
nor U3135 (N_3135,In_1312,In_1304);
and U3136 (N_3136,In_1140,In_935);
or U3137 (N_3137,In_1238,In_713);
and U3138 (N_3138,In_1121,In_147);
and U3139 (N_3139,In_114,In_1298);
nor U3140 (N_3140,In_796,In_801);
nand U3141 (N_3141,In_323,In_610);
and U3142 (N_3142,In_109,In_1300);
or U3143 (N_3143,In_771,In_362);
nor U3144 (N_3144,In_856,In_726);
nand U3145 (N_3145,In_114,In_1443);
nor U3146 (N_3146,In_31,In_85);
and U3147 (N_3147,In_1436,In_1497);
xor U3148 (N_3148,In_163,In_372);
xor U3149 (N_3149,In_623,In_962);
xor U3150 (N_3150,In_365,In_727);
and U3151 (N_3151,In_278,In_199);
and U3152 (N_3152,In_1260,In_440);
or U3153 (N_3153,In_466,In_449);
nand U3154 (N_3154,In_786,In_1205);
nand U3155 (N_3155,In_990,In_1440);
nand U3156 (N_3156,In_408,In_170);
or U3157 (N_3157,In_1153,In_1318);
or U3158 (N_3158,In_1117,In_88);
xnor U3159 (N_3159,In_285,In_1241);
or U3160 (N_3160,In_372,In_1157);
and U3161 (N_3161,In_783,In_1117);
nor U3162 (N_3162,In_1289,In_483);
and U3163 (N_3163,In_471,In_143);
and U3164 (N_3164,In_479,In_95);
and U3165 (N_3165,In_744,In_1139);
or U3166 (N_3166,In_474,In_1402);
or U3167 (N_3167,In_115,In_102);
or U3168 (N_3168,In_1120,In_404);
nor U3169 (N_3169,In_1276,In_799);
or U3170 (N_3170,In_1465,In_898);
nor U3171 (N_3171,In_1365,In_211);
xor U3172 (N_3172,In_334,In_105);
nand U3173 (N_3173,In_336,In_1101);
nand U3174 (N_3174,In_928,In_705);
nor U3175 (N_3175,In_1050,In_917);
xor U3176 (N_3176,In_1467,In_381);
or U3177 (N_3177,In_22,In_8);
nor U3178 (N_3178,In_504,In_125);
nor U3179 (N_3179,In_1421,In_363);
xnor U3180 (N_3180,In_213,In_81);
and U3181 (N_3181,In_1011,In_10);
or U3182 (N_3182,In_859,In_341);
and U3183 (N_3183,In_60,In_914);
or U3184 (N_3184,In_1103,In_798);
nor U3185 (N_3185,In_362,In_1033);
and U3186 (N_3186,In_604,In_748);
and U3187 (N_3187,In_370,In_1441);
and U3188 (N_3188,In_746,In_74);
nand U3189 (N_3189,In_622,In_1264);
or U3190 (N_3190,In_854,In_1386);
nand U3191 (N_3191,In_1415,In_1469);
nand U3192 (N_3192,In_956,In_346);
nand U3193 (N_3193,In_1211,In_1354);
or U3194 (N_3194,In_1282,In_614);
nor U3195 (N_3195,In_707,In_384);
and U3196 (N_3196,In_13,In_1094);
nand U3197 (N_3197,In_480,In_1117);
nor U3198 (N_3198,In_298,In_293);
and U3199 (N_3199,In_167,In_827);
or U3200 (N_3200,In_1221,In_514);
nor U3201 (N_3201,In_747,In_779);
or U3202 (N_3202,In_980,In_74);
nor U3203 (N_3203,In_879,In_700);
nand U3204 (N_3204,In_1156,In_220);
nor U3205 (N_3205,In_553,In_95);
and U3206 (N_3206,In_437,In_65);
nand U3207 (N_3207,In_1090,In_1193);
and U3208 (N_3208,In_1485,In_1382);
and U3209 (N_3209,In_1283,In_1247);
nand U3210 (N_3210,In_839,In_133);
nor U3211 (N_3211,In_1084,In_1498);
nor U3212 (N_3212,In_378,In_1366);
or U3213 (N_3213,In_134,In_1041);
nor U3214 (N_3214,In_889,In_157);
or U3215 (N_3215,In_149,In_537);
nand U3216 (N_3216,In_444,In_1062);
xor U3217 (N_3217,In_863,In_707);
or U3218 (N_3218,In_1473,In_603);
nor U3219 (N_3219,In_1442,In_1408);
or U3220 (N_3220,In_1416,In_93);
nor U3221 (N_3221,In_857,In_615);
xnor U3222 (N_3222,In_263,In_1083);
and U3223 (N_3223,In_832,In_638);
xnor U3224 (N_3224,In_813,In_1079);
and U3225 (N_3225,In_1340,In_632);
nand U3226 (N_3226,In_634,In_905);
nor U3227 (N_3227,In_487,In_1137);
nor U3228 (N_3228,In_1124,In_458);
and U3229 (N_3229,In_1114,In_1076);
nor U3230 (N_3230,In_435,In_136);
nand U3231 (N_3231,In_1199,In_910);
nor U3232 (N_3232,In_136,In_1163);
and U3233 (N_3233,In_1222,In_1124);
nand U3234 (N_3234,In_6,In_1262);
and U3235 (N_3235,In_1295,In_599);
and U3236 (N_3236,In_1080,In_431);
nand U3237 (N_3237,In_119,In_1280);
nand U3238 (N_3238,In_1472,In_1249);
and U3239 (N_3239,In_659,In_1096);
nor U3240 (N_3240,In_1073,In_1277);
nand U3241 (N_3241,In_1103,In_1124);
nor U3242 (N_3242,In_563,In_712);
and U3243 (N_3243,In_888,In_350);
nand U3244 (N_3244,In_759,In_429);
or U3245 (N_3245,In_575,In_1312);
or U3246 (N_3246,In_1359,In_1186);
nand U3247 (N_3247,In_1136,In_113);
and U3248 (N_3248,In_967,In_314);
or U3249 (N_3249,In_372,In_1116);
and U3250 (N_3250,In_814,In_396);
and U3251 (N_3251,In_828,In_1116);
xor U3252 (N_3252,In_1376,In_315);
nor U3253 (N_3253,In_147,In_363);
nor U3254 (N_3254,In_666,In_658);
nand U3255 (N_3255,In_21,In_341);
nor U3256 (N_3256,In_951,In_957);
or U3257 (N_3257,In_72,In_46);
nand U3258 (N_3258,In_1479,In_1400);
nand U3259 (N_3259,In_1257,In_230);
and U3260 (N_3260,In_1099,In_1239);
and U3261 (N_3261,In_1034,In_459);
or U3262 (N_3262,In_43,In_1245);
nor U3263 (N_3263,In_300,In_602);
nor U3264 (N_3264,In_195,In_642);
nand U3265 (N_3265,In_1288,In_1326);
nor U3266 (N_3266,In_845,In_626);
and U3267 (N_3267,In_390,In_1123);
or U3268 (N_3268,In_385,In_1322);
and U3269 (N_3269,In_1047,In_572);
or U3270 (N_3270,In_1066,In_851);
or U3271 (N_3271,In_1417,In_1149);
and U3272 (N_3272,In_75,In_823);
xor U3273 (N_3273,In_438,In_1330);
nand U3274 (N_3274,In_924,In_939);
nor U3275 (N_3275,In_395,In_938);
nor U3276 (N_3276,In_43,In_1045);
xnor U3277 (N_3277,In_276,In_1462);
nand U3278 (N_3278,In_1034,In_643);
nor U3279 (N_3279,In_373,In_1059);
nand U3280 (N_3280,In_13,In_711);
nor U3281 (N_3281,In_1287,In_568);
nand U3282 (N_3282,In_721,In_92);
or U3283 (N_3283,In_241,In_1227);
xor U3284 (N_3284,In_861,In_970);
or U3285 (N_3285,In_420,In_1256);
and U3286 (N_3286,In_959,In_790);
nor U3287 (N_3287,In_881,In_1167);
or U3288 (N_3288,In_1372,In_1059);
or U3289 (N_3289,In_802,In_1153);
or U3290 (N_3290,In_643,In_262);
nor U3291 (N_3291,In_938,In_1339);
xnor U3292 (N_3292,In_1442,In_672);
and U3293 (N_3293,In_251,In_1169);
or U3294 (N_3294,In_1023,In_1196);
or U3295 (N_3295,In_1324,In_120);
nand U3296 (N_3296,In_36,In_685);
nand U3297 (N_3297,In_1204,In_497);
or U3298 (N_3298,In_539,In_653);
and U3299 (N_3299,In_722,In_571);
nor U3300 (N_3300,In_1339,In_225);
nand U3301 (N_3301,In_692,In_1132);
or U3302 (N_3302,In_290,In_1267);
nand U3303 (N_3303,In_238,In_213);
or U3304 (N_3304,In_1405,In_1179);
and U3305 (N_3305,In_106,In_450);
or U3306 (N_3306,In_1231,In_571);
and U3307 (N_3307,In_1372,In_570);
and U3308 (N_3308,In_1338,In_269);
nand U3309 (N_3309,In_162,In_413);
nand U3310 (N_3310,In_215,In_96);
or U3311 (N_3311,In_1433,In_605);
or U3312 (N_3312,In_964,In_1455);
nand U3313 (N_3313,In_592,In_1090);
or U3314 (N_3314,In_340,In_307);
nand U3315 (N_3315,In_681,In_749);
and U3316 (N_3316,In_377,In_925);
or U3317 (N_3317,In_402,In_363);
nor U3318 (N_3318,In_89,In_1370);
nand U3319 (N_3319,In_398,In_1448);
nand U3320 (N_3320,In_722,In_901);
or U3321 (N_3321,In_343,In_723);
nor U3322 (N_3322,In_1324,In_1142);
nor U3323 (N_3323,In_262,In_1260);
nor U3324 (N_3324,In_1013,In_1414);
nand U3325 (N_3325,In_601,In_432);
and U3326 (N_3326,In_1471,In_1081);
and U3327 (N_3327,In_201,In_370);
and U3328 (N_3328,In_94,In_1314);
or U3329 (N_3329,In_716,In_1306);
or U3330 (N_3330,In_768,In_1485);
nand U3331 (N_3331,In_1169,In_404);
and U3332 (N_3332,In_420,In_774);
nor U3333 (N_3333,In_599,In_1329);
xnor U3334 (N_3334,In_45,In_665);
and U3335 (N_3335,In_867,In_1180);
nor U3336 (N_3336,In_278,In_1254);
or U3337 (N_3337,In_1401,In_76);
xor U3338 (N_3338,In_1469,In_1342);
nor U3339 (N_3339,In_1425,In_1204);
nand U3340 (N_3340,In_72,In_580);
nor U3341 (N_3341,In_315,In_1157);
nand U3342 (N_3342,In_1449,In_245);
xnor U3343 (N_3343,In_117,In_1073);
nor U3344 (N_3344,In_980,In_1357);
xor U3345 (N_3345,In_1454,In_1482);
nor U3346 (N_3346,In_855,In_648);
or U3347 (N_3347,In_1496,In_383);
and U3348 (N_3348,In_560,In_1489);
and U3349 (N_3349,In_1120,In_205);
and U3350 (N_3350,In_1418,In_21);
or U3351 (N_3351,In_482,In_541);
nand U3352 (N_3352,In_430,In_701);
or U3353 (N_3353,In_490,In_5);
or U3354 (N_3354,In_1398,In_120);
nor U3355 (N_3355,In_326,In_636);
nor U3356 (N_3356,In_265,In_345);
nand U3357 (N_3357,In_128,In_882);
or U3358 (N_3358,In_219,In_742);
or U3359 (N_3359,In_277,In_132);
and U3360 (N_3360,In_942,In_1062);
nor U3361 (N_3361,In_553,In_350);
and U3362 (N_3362,In_350,In_163);
or U3363 (N_3363,In_946,In_955);
and U3364 (N_3364,In_1005,In_350);
and U3365 (N_3365,In_1138,In_18);
or U3366 (N_3366,In_970,In_465);
nand U3367 (N_3367,In_294,In_202);
and U3368 (N_3368,In_580,In_811);
and U3369 (N_3369,In_1044,In_322);
xnor U3370 (N_3370,In_453,In_804);
nor U3371 (N_3371,In_341,In_1189);
or U3372 (N_3372,In_1341,In_1402);
or U3373 (N_3373,In_1228,In_614);
nor U3374 (N_3374,In_671,In_775);
nor U3375 (N_3375,In_628,In_560);
nor U3376 (N_3376,In_506,In_1347);
or U3377 (N_3377,In_864,In_616);
nand U3378 (N_3378,In_1043,In_1051);
nand U3379 (N_3379,In_939,In_8);
nor U3380 (N_3380,In_1158,In_608);
nand U3381 (N_3381,In_917,In_339);
nand U3382 (N_3382,In_935,In_1342);
nand U3383 (N_3383,In_722,In_664);
nand U3384 (N_3384,In_818,In_1028);
or U3385 (N_3385,In_896,In_1140);
nor U3386 (N_3386,In_894,In_195);
xor U3387 (N_3387,In_944,In_371);
nor U3388 (N_3388,In_1032,In_1298);
or U3389 (N_3389,In_1336,In_67);
nor U3390 (N_3390,In_1431,In_772);
and U3391 (N_3391,In_1456,In_1264);
nor U3392 (N_3392,In_1035,In_419);
nor U3393 (N_3393,In_1087,In_1016);
or U3394 (N_3394,In_600,In_237);
nand U3395 (N_3395,In_914,In_894);
nor U3396 (N_3396,In_403,In_268);
nand U3397 (N_3397,In_556,In_8);
nor U3398 (N_3398,In_310,In_375);
nor U3399 (N_3399,In_1396,In_117);
and U3400 (N_3400,In_497,In_938);
or U3401 (N_3401,In_367,In_946);
nand U3402 (N_3402,In_841,In_1065);
or U3403 (N_3403,In_1048,In_903);
nand U3404 (N_3404,In_896,In_1283);
and U3405 (N_3405,In_754,In_208);
nor U3406 (N_3406,In_1476,In_642);
nand U3407 (N_3407,In_118,In_1239);
nor U3408 (N_3408,In_670,In_1309);
nor U3409 (N_3409,In_964,In_282);
nor U3410 (N_3410,In_437,In_1036);
nor U3411 (N_3411,In_998,In_790);
or U3412 (N_3412,In_1086,In_237);
or U3413 (N_3413,In_228,In_368);
nor U3414 (N_3414,In_514,In_1223);
and U3415 (N_3415,In_1013,In_271);
nand U3416 (N_3416,In_1051,In_248);
and U3417 (N_3417,In_1445,In_879);
nand U3418 (N_3418,In_46,In_259);
or U3419 (N_3419,In_942,In_753);
nand U3420 (N_3420,In_805,In_20);
nor U3421 (N_3421,In_349,In_748);
nor U3422 (N_3422,In_386,In_1388);
or U3423 (N_3423,In_274,In_374);
and U3424 (N_3424,In_1349,In_278);
or U3425 (N_3425,In_761,In_1163);
nor U3426 (N_3426,In_416,In_716);
xnor U3427 (N_3427,In_675,In_899);
and U3428 (N_3428,In_984,In_663);
and U3429 (N_3429,In_1285,In_698);
nand U3430 (N_3430,In_287,In_739);
nand U3431 (N_3431,In_515,In_787);
or U3432 (N_3432,In_663,In_836);
xnor U3433 (N_3433,In_631,In_687);
or U3434 (N_3434,In_683,In_535);
and U3435 (N_3435,In_1294,In_472);
or U3436 (N_3436,In_334,In_1008);
and U3437 (N_3437,In_863,In_429);
nand U3438 (N_3438,In_1007,In_1360);
and U3439 (N_3439,In_901,In_271);
and U3440 (N_3440,In_1076,In_732);
or U3441 (N_3441,In_27,In_774);
xnor U3442 (N_3442,In_1080,In_265);
nor U3443 (N_3443,In_86,In_1330);
xor U3444 (N_3444,In_361,In_273);
and U3445 (N_3445,In_152,In_1226);
nor U3446 (N_3446,In_1266,In_845);
or U3447 (N_3447,In_1233,In_532);
and U3448 (N_3448,In_1345,In_1388);
nand U3449 (N_3449,In_1161,In_176);
and U3450 (N_3450,In_1292,In_966);
and U3451 (N_3451,In_642,In_0);
and U3452 (N_3452,In_1439,In_162);
nor U3453 (N_3453,In_319,In_328);
nor U3454 (N_3454,In_1228,In_837);
and U3455 (N_3455,In_1327,In_1136);
or U3456 (N_3456,In_866,In_753);
or U3457 (N_3457,In_945,In_1354);
and U3458 (N_3458,In_111,In_606);
or U3459 (N_3459,In_925,In_1220);
xnor U3460 (N_3460,In_667,In_630);
nor U3461 (N_3461,In_1474,In_218);
nor U3462 (N_3462,In_934,In_625);
xnor U3463 (N_3463,In_444,In_487);
or U3464 (N_3464,In_36,In_498);
or U3465 (N_3465,In_81,In_797);
or U3466 (N_3466,In_1349,In_1088);
or U3467 (N_3467,In_282,In_410);
nor U3468 (N_3468,In_1167,In_1044);
or U3469 (N_3469,In_1077,In_575);
xor U3470 (N_3470,In_795,In_640);
nor U3471 (N_3471,In_1458,In_1247);
nor U3472 (N_3472,In_574,In_1275);
or U3473 (N_3473,In_1293,In_829);
and U3474 (N_3474,In_79,In_342);
xnor U3475 (N_3475,In_1085,In_1407);
or U3476 (N_3476,In_1359,In_296);
or U3477 (N_3477,In_28,In_506);
nor U3478 (N_3478,In_349,In_1334);
nand U3479 (N_3479,In_29,In_94);
and U3480 (N_3480,In_776,In_719);
and U3481 (N_3481,In_603,In_823);
nor U3482 (N_3482,In_663,In_153);
or U3483 (N_3483,In_969,In_55);
xnor U3484 (N_3484,In_768,In_43);
or U3485 (N_3485,In_464,In_1273);
nand U3486 (N_3486,In_993,In_15);
nand U3487 (N_3487,In_1337,In_749);
xor U3488 (N_3488,In_388,In_646);
nor U3489 (N_3489,In_133,In_869);
nand U3490 (N_3490,In_326,In_128);
or U3491 (N_3491,In_116,In_528);
or U3492 (N_3492,In_1396,In_1423);
nor U3493 (N_3493,In_200,In_1171);
nand U3494 (N_3494,In_403,In_354);
and U3495 (N_3495,In_195,In_1414);
and U3496 (N_3496,In_1176,In_1092);
nor U3497 (N_3497,In_424,In_924);
nand U3498 (N_3498,In_268,In_1189);
nor U3499 (N_3499,In_989,In_1226);
nand U3500 (N_3500,In_723,In_945);
and U3501 (N_3501,In_372,In_1492);
nand U3502 (N_3502,In_1303,In_1262);
and U3503 (N_3503,In_675,In_1327);
nor U3504 (N_3504,In_1048,In_250);
or U3505 (N_3505,In_12,In_216);
and U3506 (N_3506,In_1169,In_1139);
or U3507 (N_3507,In_1414,In_193);
nor U3508 (N_3508,In_1341,In_533);
and U3509 (N_3509,In_622,In_623);
or U3510 (N_3510,In_521,In_6);
nor U3511 (N_3511,In_1486,In_1094);
nand U3512 (N_3512,In_1017,In_172);
or U3513 (N_3513,In_1182,In_767);
or U3514 (N_3514,In_130,In_1283);
nor U3515 (N_3515,In_264,In_407);
nand U3516 (N_3516,In_443,In_955);
nand U3517 (N_3517,In_558,In_150);
and U3518 (N_3518,In_1400,In_395);
and U3519 (N_3519,In_1427,In_665);
or U3520 (N_3520,In_1317,In_1283);
or U3521 (N_3521,In_207,In_1392);
nor U3522 (N_3522,In_325,In_301);
or U3523 (N_3523,In_852,In_98);
nor U3524 (N_3524,In_1437,In_842);
and U3525 (N_3525,In_978,In_410);
or U3526 (N_3526,In_410,In_992);
nand U3527 (N_3527,In_545,In_564);
or U3528 (N_3528,In_557,In_513);
nor U3529 (N_3529,In_1196,In_441);
xor U3530 (N_3530,In_922,In_677);
nand U3531 (N_3531,In_878,In_885);
nand U3532 (N_3532,In_210,In_115);
or U3533 (N_3533,In_534,In_430);
nand U3534 (N_3534,In_1162,In_1155);
or U3535 (N_3535,In_460,In_717);
nor U3536 (N_3536,In_809,In_1145);
xnor U3537 (N_3537,In_810,In_958);
or U3538 (N_3538,In_158,In_1057);
or U3539 (N_3539,In_1087,In_813);
and U3540 (N_3540,In_258,In_727);
nor U3541 (N_3541,In_1307,In_1076);
or U3542 (N_3542,In_800,In_860);
xnor U3543 (N_3543,In_1283,In_618);
and U3544 (N_3544,In_1067,In_774);
or U3545 (N_3545,In_1039,In_1335);
nor U3546 (N_3546,In_99,In_869);
or U3547 (N_3547,In_494,In_1074);
and U3548 (N_3548,In_1311,In_1130);
and U3549 (N_3549,In_599,In_1);
and U3550 (N_3550,In_1289,In_619);
and U3551 (N_3551,In_1421,In_685);
and U3552 (N_3552,In_1302,In_1442);
and U3553 (N_3553,In_220,In_275);
and U3554 (N_3554,In_39,In_609);
and U3555 (N_3555,In_1364,In_864);
nand U3556 (N_3556,In_684,In_1153);
nor U3557 (N_3557,In_913,In_1427);
or U3558 (N_3558,In_286,In_1158);
and U3559 (N_3559,In_172,In_1000);
nand U3560 (N_3560,In_1224,In_224);
and U3561 (N_3561,In_307,In_1408);
xor U3562 (N_3562,In_536,In_946);
nor U3563 (N_3563,In_1207,In_377);
or U3564 (N_3564,In_120,In_500);
or U3565 (N_3565,In_1130,In_1284);
and U3566 (N_3566,In_587,In_820);
and U3567 (N_3567,In_1058,In_457);
nor U3568 (N_3568,In_281,In_928);
nor U3569 (N_3569,In_741,In_1155);
nor U3570 (N_3570,In_1115,In_1204);
nor U3571 (N_3571,In_690,In_35);
or U3572 (N_3572,In_93,In_1348);
or U3573 (N_3573,In_333,In_1439);
and U3574 (N_3574,In_626,In_101);
or U3575 (N_3575,In_1052,In_642);
nand U3576 (N_3576,In_45,In_33);
and U3577 (N_3577,In_1348,In_306);
nor U3578 (N_3578,In_330,In_1412);
nand U3579 (N_3579,In_792,In_1182);
or U3580 (N_3580,In_939,In_1413);
or U3581 (N_3581,In_413,In_303);
nand U3582 (N_3582,In_73,In_599);
nand U3583 (N_3583,In_1028,In_675);
and U3584 (N_3584,In_1324,In_30);
and U3585 (N_3585,In_551,In_1204);
nand U3586 (N_3586,In_1456,In_1402);
or U3587 (N_3587,In_387,In_361);
or U3588 (N_3588,In_209,In_49);
xor U3589 (N_3589,In_632,In_767);
or U3590 (N_3590,In_883,In_594);
and U3591 (N_3591,In_1282,In_1099);
nor U3592 (N_3592,In_1231,In_361);
nor U3593 (N_3593,In_18,In_829);
and U3594 (N_3594,In_1429,In_69);
nor U3595 (N_3595,In_1018,In_856);
xor U3596 (N_3596,In_1357,In_357);
and U3597 (N_3597,In_236,In_449);
or U3598 (N_3598,In_79,In_1187);
nor U3599 (N_3599,In_637,In_967);
nand U3600 (N_3600,In_1357,In_363);
or U3601 (N_3601,In_880,In_510);
nand U3602 (N_3602,In_780,In_934);
xnor U3603 (N_3603,In_826,In_1256);
or U3604 (N_3604,In_1383,In_723);
or U3605 (N_3605,In_248,In_1288);
or U3606 (N_3606,In_305,In_292);
xor U3607 (N_3607,In_736,In_958);
nor U3608 (N_3608,In_1321,In_1156);
or U3609 (N_3609,In_1028,In_46);
nand U3610 (N_3610,In_89,In_850);
and U3611 (N_3611,In_1468,In_658);
or U3612 (N_3612,In_39,In_888);
or U3613 (N_3613,In_1261,In_267);
and U3614 (N_3614,In_560,In_582);
nand U3615 (N_3615,In_622,In_291);
and U3616 (N_3616,In_1353,In_465);
or U3617 (N_3617,In_1343,In_475);
or U3618 (N_3618,In_1268,In_1188);
nand U3619 (N_3619,In_311,In_838);
or U3620 (N_3620,In_627,In_1382);
and U3621 (N_3621,In_888,In_399);
nand U3622 (N_3622,In_1437,In_453);
nand U3623 (N_3623,In_575,In_944);
or U3624 (N_3624,In_1059,In_1334);
nor U3625 (N_3625,In_1043,In_781);
or U3626 (N_3626,In_532,In_23);
nand U3627 (N_3627,In_474,In_945);
or U3628 (N_3628,In_1178,In_451);
xnor U3629 (N_3629,In_682,In_1005);
nand U3630 (N_3630,In_888,In_1264);
xnor U3631 (N_3631,In_57,In_380);
or U3632 (N_3632,In_1104,In_1429);
nor U3633 (N_3633,In_391,In_952);
nand U3634 (N_3634,In_800,In_648);
nand U3635 (N_3635,In_1427,In_561);
xnor U3636 (N_3636,In_623,In_140);
and U3637 (N_3637,In_12,In_0);
nand U3638 (N_3638,In_1195,In_312);
or U3639 (N_3639,In_972,In_1129);
nor U3640 (N_3640,In_327,In_1216);
nor U3641 (N_3641,In_615,In_1490);
and U3642 (N_3642,In_216,In_1222);
and U3643 (N_3643,In_1064,In_203);
nor U3644 (N_3644,In_25,In_1279);
nand U3645 (N_3645,In_365,In_1272);
xnor U3646 (N_3646,In_216,In_1377);
xor U3647 (N_3647,In_788,In_1471);
or U3648 (N_3648,In_1336,In_1120);
and U3649 (N_3649,In_152,In_190);
nand U3650 (N_3650,In_1290,In_1423);
nor U3651 (N_3651,In_653,In_962);
nor U3652 (N_3652,In_1095,In_673);
and U3653 (N_3653,In_63,In_1395);
and U3654 (N_3654,In_1131,In_1235);
or U3655 (N_3655,In_453,In_344);
nor U3656 (N_3656,In_493,In_94);
xor U3657 (N_3657,In_24,In_1480);
xnor U3658 (N_3658,In_1373,In_275);
nand U3659 (N_3659,In_789,In_575);
or U3660 (N_3660,In_1085,In_498);
nor U3661 (N_3661,In_728,In_1060);
nor U3662 (N_3662,In_1165,In_682);
nor U3663 (N_3663,In_1205,In_1476);
or U3664 (N_3664,In_1214,In_1110);
nand U3665 (N_3665,In_526,In_428);
and U3666 (N_3666,In_745,In_558);
nand U3667 (N_3667,In_1005,In_210);
nor U3668 (N_3668,In_421,In_611);
nor U3669 (N_3669,In_1455,In_1250);
nand U3670 (N_3670,In_49,In_329);
or U3671 (N_3671,In_678,In_336);
and U3672 (N_3672,In_188,In_626);
and U3673 (N_3673,In_1002,In_346);
nor U3674 (N_3674,In_338,In_433);
nand U3675 (N_3675,In_1310,In_419);
or U3676 (N_3676,In_1310,In_814);
nor U3677 (N_3677,In_1317,In_1225);
or U3678 (N_3678,In_21,In_1257);
nand U3679 (N_3679,In_488,In_1285);
nand U3680 (N_3680,In_264,In_800);
nand U3681 (N_3681,In_1150,In_1066);
nor U3682 (N_3682,In_172,In_351);
and U3683 (N_3683,In_225,In_328);
nand U3684 (N_3684,In_554,In_601);
xor U3685 (N_3685,In_1481,In_1408);
nand U3686 (N_3686,In_1140,In_1389);
or U3687 (N_3687,In_823,In_30);
and U3688 (N_3688,In_127,In_724);
nand U3689 (N_3689,In_1019,In_838);
nor U3690 (N_3690,In_1088,In_1242);
nor U3691 (N_3691,In_746,In_490);
or U3692 (N_3692,In_351,In_1427);
nor U3693 (N_3693,In_1491,In_1465);
nand U3694 (N_3694,In_148,In_1472);
nor U3695 (N_3695,In_403,In_708);
or U3696 (N_3696,In_1496,In_29);
and U3697 (N_3697,In_357,In_893);
nand U3698 (N_3698,In_886,In_68);
xnor U3699 (N_3699,In_707,In_1202);
nand U3700 (N_3700,In_1195,In_445);
or U3701 (N_3701,In_1030,In_379);
nand U3702 (N_3702,In_1138,In_1081);
nand U3703 (N_3703,In_646,In_809);
or U3704 (N_3704,In_649,In_632);
nor U3705 (N_3705,In_687,In_1151);
nor U3706 (N_3706,In_1015,In_865);
xor U3707 (N_3707,In_59,In_154);
and U3708 (N_3708,In_711,In_489);
nor U3709 (N_3709,In_1216,In_1282);
and U3710 (N_3710,In_765,In_970);
or U3711 (N_3711,In_1009,In_879);
xnor U3712 (N_3712,In_1276,In_207);
xor U3713 (N_3713,In_662,In_126);
nand U3714 (N_3714,In_178,In_1300);
xnor U3715 (N_3715,In_901,In_644);
and U3716 (N_3716,In_1066,In_1030);
or U3717 (N_3717,In_262,In_971);
nor U3718 (N_3718,In_167,In_1416);
or U3719 (N_3719,In_112,In_934);
and U3720 (N_3720,In_977,In_297);
and U3721 (N_3721,In_910,In_1149);
and U3722 (N_3722,In_353,In_982);
or U3723 (N_3723,In_753,In_1475);
or U3724 (N_3724,In_690,In_680);
and U3725 (N_3725,In_905,In_366);
or U3726 (N_3726,In_95,In_810);
or U3727 (N_3727,In_436,In_818);
xnor U3728 (N_3728,In_1323,In_366);
or U3729 (N_3729,In_992,In_425);
nor U3730 (N_3730,In_999,In_363);
nor U3731 (N_3731,In_547,In_953);
or U3732 (N_3732,In_451,In_1170);
or U3733 (N_3733,In_801,In_450);
nand U3734 (N_3734,In_783,In_464);
nand U3735 (N_3735,In_376,In_969);
nand U3736 (N_3736,In_1394,In_1313);
or U3737 (N_3737,In_1122,In_5);
nor U3738 (N_3738,In_925,In_759);
and U3739 (N_3739,In_1023,In_547);
nor U3740 (N_3740,In_802,In_893);
and U3741 (N_3741,In_1429,In_400);
or U3742 (N_3742,In_158,In_1033);
nor U3743 (N_3743,In_1301,In_343);
nand U3744 (N_3744,In_1478,In_1298);
and U3745 (N_3745,In_448,In_936);
nand U3746 (N_3746,In_1188,In_317);
and U3747 (N_3747,In_889,In_1169);
nor U3748 (N_3748,In_796,In_211);
and U3749 (N_3749,In_383,In_738);
or U3750 (N_3750,In_428,In_353);
nor U3751 (N_3751,In_423,In_643);
nand U3752 (N_3752,In_236,In_891);
or U3753 (N_3753,In_1011,In_1093);
or U3754 (N_3754,In_413,In_1076);
nor U3755 (N_3755,In_1249,In_351);
nand U3756 (N_3756,In_81,In_183);
or U3757 (N_3757,In_997,In_835);
nand U3758 (N_3758,In_1071,In_1452);
nand U3759 (N_3759,In_98,In_608);
and U3760 (N_3760,In_726,In_1162);
nand U3761 (N_3761,In_958,In_225);
or U3762 (N_3762,In_1383,In_1041);
and U3763 (N_3763,In_1052,In_444);
or U3764 (N_3764,In_1337,In_807);
nand U3765 (N_3765,In_121,In_166);
nand U3766 (N_3766,In_730,In_1395);
or U3767 (N_3767,In_18,In_183);
nand U3768 (N_3768,In_51,In_1077);
nand U3769 (N_3769,In_77,In_52);
nor U3770 (N_3770,In_223,In_1007);
and U3771 (N_3771,In_156,In_1204);
and U3772 (N_3772,In_1212,In_641);
nor U3773 (N_3773,In_817,In_1454);
and U3774 (N_3774,In_1149,In_5);
and U3775 (N_3775,In_349,In_744);
nor U3776 (N_3776,In_984,In_1240);
and U3777 (N_3777,In_266,In_292);
or U3778 (N_3778,In_689,In_274);
nor U3779 (N_3779,In_790,In_266);
and U3780 (N_3780,In_955,In_1122);
and U3781 (N_3781,In_762,In_1143);
and U3782 (N_3782,In_1240,In_264);
and U3783 (N_3783,In_1210,In_1203);
and U3784 (N_3784,In_1366,In_570);
nand U3785 (N_3785,In_162,In_781);
nor U3786 (N_3786,In_1251,In_66);
and U3787 (N_3787,In_451,In_155);
nand U3788 (N_3788,In_1066,In_688);
nand U3789 (N_3789,In_929,In_1193);
xor U3790 (N_3790,In_662,In_833);
or U3791 (N_3791,In_1413,In_823);
nand U3792 (N_3792,In_686,In_888);
and U3793 (N_3793,In_1497,In_695);
nor U3794 (N_3794,In_303,In_1442);
or U3795 (N_3795,In_255,In_176);
or U3796 (N_3796,In_592,In_1460);
xnor U3797 (N_3797,In_1327,In_722);
nor U3798 (N_3798,In_534,In_999);
nor U3799 (N_3799,In_87,In_52);
nor U3800 (N_3800,In_240,In_951);
nand U3801 (N_3801,In_662,In_235);
nand U3802 (N_3802,In_420,In_1234);
nand U3803 (N_3803,In_561,In_232);
or U3804 (N_3804,In_274,In_743);
or U3805 (N_3805,In_869,In_450);
nand U3806 (N_3806,In_648,In_1113);
nand U3807 (N_3807,In_1393,In_1007);
nand U3808 (N_3808,In_716,In_260);
nor U3809 (N_3809,In_62,In_1462);
or U3810 (N_3810,In_602,In_434);
nand U3811 (N_3811,In_1486,In_289);
or U3812 (N_3812,In_1087,In_1337);
and U3813 (N_3813,In_1378,In_604);
nand U3814 (N_3814,In_471,In_635);
nor U3815 (N_3815,In_975,In_755);
nor U3816 (N_3816,In_195,In_1204);
nand U3817 (N_3817,In_1448,In_456);
xnor U3818 (N_3818,In_75,In_12);
nor U3819 (N_3819,In_951,In_1462);
nor U3820 (N_3820,In_610,In_100);
or U3821 (N_3821,In_561,In_871);
and U3822 (N_3822,In_913,In_1339);
nor U3823 (N_3823,In_223,In_905);
and U3824 (N_3824,In_540,In_3);
nand U3825 (N_3825,In_1045,In_126);
nand U3826 (N_3826,In_212,In_189);
and U3827 (N_3827,In_135,In_682);
nor U3828 (N_3828,In_652,In_553);
and U3829 (N_3829,In_864,In_161);
xnor U3830 (N_3830,In_247,In_137);
xnor U3831 (N_3831,In_949,In_369);
and U3832 (N_3832,In_1089,In_1020);
and U3833 (N_3833,In_456,In_465);
and U3834 (N_3834,In_969,In_247);
and U3835 (N_3835,In_699,In_1163);
and U3836 (N_3836,In_1457,In_1485);
nor U3837 (N_3837,In_657,In_673);
nand U3838 (N_3838,In_1308,In_1237);
and U3839 (N_3839,In_178,In_1441);
nand U3840 (N_3840,In_694,In_587);
nor U3841 (N_3841,In_1016,In_673);
or U3842 (N_3842,In_995,In_577);
nand U3843 (N_3843,In_760,In_37);
nor U3844 (N_3844,In_133,In_352);
and U3845 (N_3845,In_836,In_371);
and U3846 (N_3846,In_355,In_41);
and U3847 (N_3847,In_1380,In_1478);
xnor U3848 (N_3848,In_1195,In_1433);
nand U3849 (N_3849,In_1264,In_158);
xnor U3850 (N_3850,In_261,In_906);
nor U3851 (N_3851,In_843,In_1331);
xnor U3852 (N_3852,In_544,In_1329);
or U3853 (N_3853,In_24,In_564);
or U3854 (N_3854,In_295,In_1029);
or U3855 (N_3855,In_1431,In_875);
nand U3856 (N_3856,In_279,In_584);
or U3857 (N_3857,In_515,In_1122);
nor U3858 (N_3858,In_1117,In_158);
nor U3859 (N_3859,In_712,In_1402);
nand U3860 (N_3860,In_713,In_1031);
xnor U3861 (N_3861,In_174,In_1462);
nor U3862 (N_3862,In_1025,In_725);
and U3863 (N_3863,In_1136,In_1336);
nand U3864 (N_3864,In_384,In_378);
nor U3865 (N_3865,In_907,In_94);
nand U3866 (N_3866,In_1464,In_1366);
nor U3867 (N_3867,In_1498,In_196);
or U3868 (N_3868,In_25,In_1413);
nor U3869 (N_3869,In_66,In_1113);
nand U3870 (N_3870,In_210,In_688);
or U3871 (N_3871,In_884,In_402);
nor U3872 (N_3872,In_289,In_1477);
xnor U3873 (N_3873,In_493,In_1052);
or U3874 (N_3874,In_603,In_1495);
nor U3875 (N_3875,In_1311,In_893);
and U3876 (N_3876,In_776,In_364);
or U3877 (N_3877,In_1075,In_704);
nor U3878 (N_3878,In_1468,In_127);
xnor U3879 (N_3879,In_1033,In_735);
xor U3880 (N_3880,In_607,In_1496);
or U3881 (N_3881,In_1041,In_642);
or U3882 (N_3882,In_1324,In_1113);
nor U3883 (N_3883,In_660,In_243);
and U3884 (N_3884,In_354,In_565);
nor U3885 (N_3885,In_1486,In_980);
nor U3886 (N_3886,In_711,In_1251);
xnor U3887 (N_3887,In_1352,In_457);
xnor U3888 (N_3888,In_1111,In_29);
and U3889 (N_3889,In_1009,In_1471);
or U3890 (N_3890,In_1177,In_1432);
and U3891 (N_3891,In_1146,In_568);
or U3892 (N_3892,In_1136,In_301);
and U3893 (N_3893,In_341,In_469);
nor U3894 (N_3894,In_922,In_1408);
and U3895 (N_3895,In_400,In_1298);
xor U3896 (N_3896,In_1434,In_1141);
or U3897 (N_3897,In_992,In_1196);
nor U3898 (N_3898,In_1209,In_612);
or U3899 (N_3899,In_1369,In_104);
nand U3900 (N_3900,In_1404,In_302);
nand U3901 (N_3901,In_392,In_939);
and U3902 (N_3902,In_849,In_183);
nand U3903 (N_3903,In_340,In_976);
nand U3904 (N_3904,In_438,In_772);
nor U3905 (N_3905,In_665,In_564);
and U3906 (N_3906,In_1007,In_319);
nand U3907 (N_3907,In_576,In_40);
nand U3908 (N_3908,In_642,In_128);
nor U3909 (N_3909,In_657,In_721);
nand U3910 (N_3910,In_29,In_417);
and U3911 (N_3911,In_1344,In_1118);
nand U3912 (N_3912,In_172,In_478);
and U3913 (N_3913,In_1252,In_182);
and U3914 (N_3914,In_332,In_192);
xor U3915 (N_3915,In_632,In_389);
nor U3916 (N_3916,In_606,In_400);
nand U3917 (N_3917,In_83,In_257);
nor U3918 (N_3918,In_235,In_528);
nor U3919 (N_3919,In_535,In_1420);
or U3920 (N_3920,In_707,In_630);
or U3921 (N_3921,In_1270,In_1432);
nor U3922 (N_3922,In_876,In_286);
nor U3923 (N_3923,In_657,In_656);
or U3924 (N_3924,In_166,In_922);
or U3925 (N_3925,In_1150,In_578);
xnor U3926 (N_3926,In_879,In_480);
and U3927 (N_3927,In_487,In_673);
nor U3928 (N_3928,In_1368,In_474);
or U3929 (N_3929,In_1383,In_1302);
nand U3930 (N_3930,In_1287,In_18);
nor U3931 (N_3931,In_218,In_1280);
nor U3932 (N_3932,In_78,In_1494);
nand U3933 (N_3933,In_29,In_737);
and U3934 (N_3934,In_53,In_155);
nor U3935 (N_3935,In_1276,In_344);
or U3936 (N_3936,In_1001,In_1467);
xnor U3937 (N_3937,In_1283,In_317);
nand U3938 (N_3938,In_383,In_204);
or U3939 (N_3939,In_445,In_78);
or U3940 (N_3940,In_1390,In_1375);
or U3941 (N_3941,In_998,In_786);
or U3942 (N_3942,In_914,In_1012);
nor U3943 (N_3943,In_325,In_291);
xor U3944 (N_3944,In_430,In_891);
and U3945 (N_3945,In_285,In_561);
nor U3946 (N_3946,In_909,In_387);
or U3947 (N_3947,In_1101,In_769);
and U3948 (N_3948,In_673,In_65);
nand U3949 (N_3949,In_305,In_1025);
and U3950 (N_3950,In_972,In_1228);
xor U3951 (N_3951,In_1358,In_596);
or U3952 (N_3952,In_754,In_113);
and U3953 (N_3953,In_663,In_268);
and U3954 (N_3954,In_1050,In_1341);
or U3955 (N_3955,In_1456,In_1008);
nor U3956 (N_3956,In_239,In_827);
nor U3957 (N_3957,In_509,In_1481);
or U3958 (N_3958,In_1328,In_1412);
xnor U3959 (N_3959,In_125,In_1429);
and U3960 (N_3960,In_734,In_432);
nand U3961 (N_3961,In_1384,In_785);
and U3962 (N_3962,In_611,In_556);
nand U3963 (N_3963,In_637,In_941);
nand U3964 (N_3964,In_571,In_252);
nor U3965 (N_3965,In_72,In_44);
nor U3966 (N_3966,In_869,In_578);
or U3967 (N_3967,In_421,In_1);
nand U3968 (N_3968,In_283,In_1404);
nor U3969 (N_3969,In_1213,In_515);
nor U3970 (N_3970,In_843,In_1099);
and U3971 (N_3971,In_197,In_1419);
nand U3972 (N_3972,In_267,In_996);
nor U3973 (N_3973,In_243,In_1287);
or U3974 (N_3974,In_61,In_1353);
xnor U3975 (N_3975,In_292,In_516);
xor U3976 (N_3976,In_67,In_607);
and U3977 (N_3977,In_1386,In_695);
or U3978 (N_3978,In_770,In_650);
nand U3979 (N_3979,In_988,In_778);
and U3980 (N_3980,In_23,In_1078);
and U3981 (N_3981,In_640,In_1330);
xor U3982 (N_3982,In_991,In_55);
nand U3983 (N_3983,In_1450,In_301);
xnor U3984 (N_3984,In_688,In_1232);
or U3985 (N_3985,In_290,In_992);
or U3986 (N_3986,In_538,In_996);
or U3987 (N_3987,In_296,In_129);
nor U3988 (N_3988,In_866,In_976);
and U3989 (N_3989,In_639,In_1241);
xnor U3990 (N_3990,In_476,In_289);
and U3991 (N_3991,In_545,In_450);
or U3992 (N_3992,In_68,In_478);
xor U3993 (N_3993,In_452,In_1117);
nand U3994 (N_3994,In_336,In_38);
and U3995 (N_3995,In_993,In_243);
or U3996 (N_3996,In_660,In_913);
or U3997 (N_3997,In_646,In_618);
or U3998 (N_3998,In_1423,In_1157);
and U3999 (N_3999,In_130,In_1449);
or U4000 (N_4000,In_509,In_1372);
nand U4001 (N_4001,In_1406,In_629);
or U4002 (N_4002,In_803,In_757);
nand U4003 (N_4003,In_373,In_124);
and U4004 (N_4004,In_216,In_744);
nand U4005 (N_4005,In_1445,In_490);
nand U4006 (N_4006,In_591,In_337);
nand U4007 (N_4007,In_868,In_414);
and U4008 (N_4008,In_332,In_654);
or U4009 (N_4009,In_1267,In_1141);
xnor U4010 (N_4010,In_15,In_134);
or U4011 (N_4011,In_249,In_729);
and U4012 (N_4012,In_511,In_1387);
and U4013 (N_4013,In_275,In_355);
and U4014 (N_4014,In_1299,In_970);
nand U4015 (N_4015,In_923,In_1101);
nand U4016 (N_4016,In_277,In_850);
and U4017 (N_4017,In_122,In_218);
nand U4018 (N_4018,In_1483,In_65);
and U4019 (N_4019,In_1004,In_533);
xnor U4020 (N_4020,In_1103,In_888);
nor U4021 (N_4021,In_415,In_631);
or U4022 (N_4022,In_289,In_576);
nor U4023 (N_4023,In_271,In_503);
nand U4024 (N_4024,In_655,In_371);
or U4025 (N_4025,In_890,In_508);
and U4026 (N_4026,In_176,In_495);
or U4027 (N_4027,In_1394,In_568);
and U4028 (N_4028,In_1382,In_79);
or U4029 (N_4029,In_290,In_1395);
or U4030 (N_4030,In_124,In_859);
nand U4031 (N_4031,In_528,In_536);
nand U4032 (N_4032,In_1136,In_535);
or U4033 (N_4033,In_426,In_852);
xor U4034 (N_4034,In_291,In_923);
nor U4035 (N_4035,In_491,In_1355);
nand U4036 (N_4036,In_529,In_916);
and U4037 (N_4037,In_869,In_271);
or U4038 (N_4038,In_1283,In_1477);
or U4039 (N_4039,In_909,In_465);
nand U4040 (N_4040,In_888,In_14);
and U4041 (N_4041,In_885,In_1118);
and U4042 (N_4042,In_1243,In_928);
or U4043 (N_4043,In_459,In_745);
nand U4044 (N_4044,In_33,In_5);
nand U4045 (N_4045,In_1410,In_774);
and U4046 (N_4046,In_1228,In_711);
nand U4047 (N_4047,In_138,In_724);
or U4048 (N_4048,In_442,In_23);
or U4049 (N_4049,In_1209,In_1101);
and U4050 (N_4050,In_355,In_890);
or U4051 (N_4051,In_1240,In_1143);
and U4052 (N_4052,In_980,In_336);
nor U4053 (N_4053,In_224,In_337);
and U4054 (N_4054,In_945,In_646);
nand U4055 (N_4055,In_614,In_517);
and U4056 (N_4056,In_106,In_545);
nand U4057 (N_4057,In_48,In_473);
and U4058 (N_4058,In_884,In_901);
or U4059 (N_4059,In_265,In_151);
nand U4060 (N_4060,In_1274,In_1106);
nor U4061 (N_4061,In_224,In_1011);
nand U4062 (N_4062,In_766,In_1168);
nor U4063 (N_4063,In_89,In_1176);
and U4064 (N_4064,In_572,In_1191);
or U4065 (N_4065,In_129,In_331);
or U4066 (N_4066,In_914,In_1065);
nand U4067 (N_4067,In_13,In_288);
nor U4068 (N_4068,In_126,In_69);
or U4069 (N_4069,In_269,In_37);
xor U4070 (N_4070,In_1066,In_976);
nor U4071 (N_4071,In_973,In_73);
nand U4072 (N_4072,In_1269,In_665);
or U4073 (N_4073,In_686,In_514);
xnor U4074 (N_4074,In_1280,In_550);
or U4075 (N_4075,In_478,In_486);
or U4076 (N_4076,In_415,In_1039);
and U4077 (N_4077,In_1272,In_610);
or U4078 (N_4078,In_785,In_1300);
or U4079 (N_4079,In_225,In_127);
xnor U4080 (N_4080,In_440,In_218);
or U4081 (N_4081,In_838,In_133);
and U4082 (N_4082,In_1439,In_1399);
nor U4083 (N_4083,In_221,In_364);
nor U4084 (N_4084,In_928,In_1396);
xnor U4085 (N_4085,In_1136,In_160);
and U4086 (N_4086,In_154,In_1250);
or U4087 (N_4087,In_100,In_268);
and U4088 (N_4088,In_191,In_380);
xor U4089 (N_4089,In_1168,In_817);
nor U4090 (N_4090,In_316,In_1141);
nand U4091 (N_4091,In_212,In_783);
and U4092 (N_4092,In_1080,In_151);
nand U4093 (N_4093,In_135,In_192);
and U4094 (N_4094,In_823,In_1122);
nand U4095 (N_4095,In_481,In_471);
and U4096 (N_4096,In_164,In_306);
nor U4097 (N_4097,In_25,In_1428);
or U4098 (N_4098,In_737,In_878);
nand U4099 (N_4099,In_175,In_1225);
or U4100 (N_4100,In_678,In_634);
xnor U4101 (N_4101,In_710,In_365);
or U4102 (N_4102,In_705,In_1366);
nor U4103 (N_4103,In_1402,In_133);
or U4104 (N_4104,In_661,In_69);
or U4105 (N_4105,In_816,In_418);
xor U4106 (N_4106,In_1137,In_341);
nand U4107 (N_4107,In_856,In_311);
nand U4108 (N_4108,In_1463,In_13);
or U4109 (N_4109,In_111,In_1156);
xor U4110 (N_4110,In_1005,In_1068);
nor U4111 (N_4111,In_1311,In_925);
and U4112 (N_4112,In_1044,In_155);
nand U4113 (N_4113,In_1275,In_317);
nor U4114 (N_4114,In_1283,In_1416);
nor U4115 (N_4115,In_1478,In_14);
and U4116 (N_4116,In_999,In_907);
nor U4117 (N_4117,In_956,In_30);
and U4118 (N_4118,In_399,In_1396);
or U4119 (N_4119,In_1415,In_128);
nor U4120 (N_4120,In_1074,In_308);
nor U4121 (N_4121,In_802,In_75);
xor U4122 (N_4122,In_903,In_90);
nor U4123 (N_4123,In_39,In_661);
nand U4124 (N_4124,In_303,In_906);
nor U4125 (N_4125,In_114,In_1492);
nand U4126 (N_4126,In_728,In_409);
or U4127 (N_4127,In_1056,In_381);
nor U4128 (N_4128,In_1458,In_1442);
and U4129 (N_4129,In_561,In_1385);
or U4130 (N_4130,In_223,In_932);
nor U4131 (N_4131,In_356,In_1225);
and U4132 (N_4132,In_10,In_229);
or U4133 (N_4133,In_265,In_1173);
nand U4134 (N_4134,In_426,In_596);
nor U4135 (N_4135,In_977,In_755);
nand U4136 (N_4136,In_24,In_497);
nor U4137 (N_4137,In_171,In_795);
nand U4138 (N_4138,In_847,In_1366);
and U4139 (N_4139,In_1354,In_1485);
and U4140 (N_4140,In_815,In_165);
and U4141 (N_4141,In_676,In_818);
and U4142 (N_4142,In_769,In_622);
nand U4143 (N_4143,In_490,In_123);
xor U4144 (N_4144,In_473,In_1247);
or U4145 (N_4145,In_522,In_9);
or U4146 (N_4146,In_808,In_113);
nor U4147 (N_4147,In_821,In_628);
nor U4148 (N_4148,In_1377,In_815);
nand U4149 (N_4149,In_1498,In_178);
and U4150 (N_4150,In_1213,In_1411);
nor U4151 (N_4151,In_567,In_906);
or U4152 (N_4152,In_318,In_885);
nand U4153 (N_4153,In_70,In_895);
xor U4154 (N_4154,In_1353,In_46);
nor U4155 (N_4155,In_454,In_183);
nand U4156 (N_4156,In_790,In_616);
or U4157 (N_4157,In_146,In_344);
and U4158 (N_4158,In_1170,In_960);
or U4159 (N_4159,In_404,In_1273);
and U4160 (N_4160,In_1294,In_528);
nor U4161 (N_4161,In_291,In_352);
nor U4162 (N_4162,In_1189,In_1159);
and U4163 (N_4163,In_970,In_1400);
or U4164 (N_4164,In_515,In_649);
nor U4165 (N_4165,In_801,In_633);
and U4166 (N_4166,In_318,In_1275);
or U4167 (N_4167,In_1453,In_905);
nor U4168 (N_4168,In_270,In_484);
nand U4169 (N_4169,In_943,In_1264);
nor U4170 (N_4170,In_653,In_774);
nand U4171 (N_4171,In_1025,In_1207);
nand U4172 (N_4172,In_798,In_1078);
nor U4173 (N_4173,In_323,In_595);
xor U4174 (N_4174,In_728,In_1454);
and U4175 (N_4175,In_1419,In_51);
and U4176 (N_4176,In_670,In_470);
or U4177 (N_4177,In_768,In_670);
or U4178 (N_4178,In_67,In_352);
nor U4179 (N_4179,In_1473,In_495);
nand U4180 (N_4180,In_1186,In_1035);
nand U4181 (N_4181,In_1379,In_82);
and U4182 (N_4182,In_1123,In_1324);
or U4183 (N_4183,In_581,In_1408);
nor U4184 (N_4184,In_284,In_878);
nor U4185 (N_4185,In_1187,In_714);
xor U4186 (N_4186,In_93,In_1265);
or U4187 (N_4187,In_703,In_1159);
xor U4188 (N_4188,In_1065,In_1113);
or U4189 (N_4189,In_314,In_106);
or U4190 (N_4190,In_598,In_1292);
nand U4191 (N_4191,In_1482,In_26);
and U4192 (N_4192,In_276,In_1308);
nand U4193 (N_4193,In_1101,In_850);
and U4194 (N_4194,In_278,In_1258);
or U4195 (N_4195,In_1271,In_583);
nand U4196 (N_4196,In_1427,In_877);
and U4197 (N_4197,In_1480,In_886);
nand U4198 (N_4198,In_1348,In_1220);
nand U4199 (N_4199,In_316,In_468);
xor U4200 (N_4200,In_1362,In_462);
nand U4201 (N_4201,In_1345,In_964);
nor U4202 (N_4202,In_679,In_672);
nand U4203 (N_4203,In_614,In_158);
nor U4204 (N_4204,In_461,In_1332);
nor U4205 (N_4205,In_881,In_526);
or U4206 (N_4206,In_1321,In_795);
nand U4207 (N_4207,In_1250,In_682);
nor U4208 (N_4208,In_1212,In_799);
nand U4209 (N_4209,In_844,In_1208);
nand U4210 (N_4210,In_516,In_707);
xor U4211 (N_4211,In_1017,In_173);
or U4212 (N_4212,In_514,In_408);
nor U4213 (N_4213,In_1004,In_1209);
nand U4214 (N_4214,In_672,In_542);
nand U4215 (N_4215,In_1158,In_856);
and U4216 (N_4216,In_768,In_1219);
xor U4217 (N_4217,In_1449,In_1433);
nor U4218 (N_4218,In_1213,In_546);
and U4219 (N_4219,In_1432,In_1471);
or U4220 (N_4220,In_860,In_311);
nor U4221 (N_4221,In_565,In_836);
nor U4222 (N_4222,In_375,In_271);
and U4223 (N_4223,In_258,In_133);
and U4224 (N_4224,In_422,In_256);
or U4225 (N_4225,In_426,In_35);
nor U4226 (N_4226,In_809,In_133);
or U4227 (N_4227,In_243,In_258);
nor U4228 (N_4228,In_1172,In_960);
and U4229 (N_4229,In_329,In_275);
nor U4230 (N_4230,In_740,In_710);
nor U4231 (N_4231,In_504,In_271);
and U4232 (N_4232,In_755,In_601);
and U4233 (N_4233,In_1471,In_300);
or U4234 (N_4234,In_736,In_210);
or U4235 (N_4235,In_1207,In_394);
nand U4236 (N_4236,In_1313,In_506);
or U4237 (N_4237,In_1287,In_1344);
and U4238 (N_4238,In_639,In_988);
or U4239 (N_4239,In_129,In_839);
or U4240 (N_4240,In_965,In_331);
xnor U4241 (N_4241,In_381,In_1493);
nor U4242 (N_4242,In_663,In_1379);
nor U4243 (N_4243,In_1461,In_1435);
nand U4244 (N_4244,In_735,In_365);
nor U4245 (N_4245,In_461,In_1173);
xor U4246 (N_4246,In_940,In_1155);
and U4247 (N_4247,In_1321,In_1302);
nand U4248 (N_4248,In_994,In_798);
or U4249 (N_4249,In_759,In_253);
and U4250 (N_4250,In_315,In_1019);
nor U4251 (N_4251,In_1308,In_326);
nand U4252 (N_4252,In_11,In_1409);
xor U4253 (N_4253,In_998,In_1123);
nor U4254 (N_4254,In_153,In_622);
nor U4255 (N_4255,In_1073,In_22);
or U4256 (N_4256,In_1429,In_458);
xor U4257 (N_4257,In_200,In_697);
nor U4258 (N_4258,In_1231,In_84);
or U4259 (N_4259,In_219,In_1196);
xor U4260 (N_4260,In_677,In_974);
or U4261 (N_4261,In_1002,In_245);
xnor U4262 (N_4262,In_99,In_978);
nand U4263 (N_4263,In_11,In_535);
nand U4264 (N_4264,In_357,In_630);
nor U4265 (N_4265,In_10,In_1408);
or U4266 (N_4266,In_797,In_1386);
or U4267 (N_4267,In_1320,In_220);
nand U4268 (N_4268,In_1278,In_702);
nor U4269 (N_4269,In_49,In_37);
nand U4270 (N_4270,In_124,In_104);
and U4271 (N_4271,In_33,In_821);
nor U4272 (N_4272,In_154,In_1368);
xnor U4273 (N_4273,In_1248,In_874);
nor U4274 (N_4274,In_1377,In_992);
nand U4275 (N_4275,In_763,In_914);
and U4276 (N_4276,In_1083,In_662);
nand U4277 (N_4277,In_1187,In_805);
or U4278 (N_4278,In_131,In_1464);
or U4279 (N_4279,In_1221,In_422);
or U4280 (N_4280,In_395,In_919);
nor U4281 (N_4281,In_900,In_602);
or U4282 (N_4282,In_1436,In_1072);
and U4283 (N_4283,In_1370,In_969);
or U4284 (N_4284,In_1443,In_917);
or U4285 (N_4285,In_781,In_1439);
or U4286 (N_4286,In_1265,In_504);
nand U4287 (N_4287,In_307,In_80);
nand U4288 (N_4288,In_772,In_640);
and U4289 (N_4289,In_191,In_1227);
or U4290 (N_4290,In_13,In_1350);
xor U4291 (N_4291,In_895,In_1231);
and U4292 (N_4292,In_23,In_51);
or U4293 (N_4293,In_884,In_639);
and U4294 (N_4294,In_1067,In_612);
and U4295 (N_4295,In_807,In_920);
nor U4296 (N_4296,In_1172,In_371);
and U4297 (N_4297,In_1265,In_834);
nand U4298 (N_4298,In_600,In_596);
xor U4299 (N_4299,In_1055,In_786);
and U4300 (N_4300,In_953,In_325);
nor U4301 (N_4301,In_1064,In_114);
nand U4302 (N_4302,In_1461,In_316);
or U4303 (N_4303,In_869,In_1181);
and U4304 (N_4304,In_363,In_708);
or U4305 (N_4305,In_514,In_611);
nor U4306 (N_4306,In_983,In_637);
nor U4307 (N_4307,In_781,In_1476);
or U4308 (N_4308,In_520,In_1061);
and U4309 (N_4309,In_1165,In_1324);
or U4310 (N_4310,In_623,In_527);
and U4311 (N_4311,In_994,In_560);
or U4312 (N_4312,In_1266,In_133);
or U4313 (N_4313,In_378,In_1479);
or U4314 (N_4314,In_971,In_1140);
nor U4315 (N_4315,In_900,In_628);
and U4316 (N_4316,In_23,In_223);
or U4317 (N_4317,In_1464,In_1035);
nor U4318 (N_4318,In_479,In_184);
and U4319 (N_4319,In_897,In_548);
and U4320 (N_4320,In_432,In_1016);
nand U4321 (N_4321,In_857,In_1071);
or U4322 (N_4322,In_1028,In_509);
nand U4323 (N_4323,In_1064,In_107);
or U4324 (N_4324,In_1206,In_727);
nand U4325 (N_4325,In_759,In_191);
and U4326 (N_4326,In_832,In_589);
xnor U4327 (N_4327,In_612,In_1130);
nand U4328 (N_4328,In_1234,In_1375);
nand U4329 (N_4329,In_1236,In_1302);
or U4330 (N_4330,In_407,In_278);
and U4331 (N_4331,In_769,In_803);
nand U4332 (N_4332,In_930,In_19);
and U4333 (N_4333,In_381,In_1455);
or U4334 (N_4334,In_1465,In_1293);
and U4335 (N_4335,In_1150,In_1050);
and U4336 (N_4336,In_1431,In_36);
nor U4337 (N_4337,In_1009,In_1247);
nand U4338 (N_4338,In_512,In_770);
nand U4339 (N_4339,In_1111,In_99);
nor U4340 (N_4340,In_431,In_1273);
nor U4341 (N_4341,In_859,In_917);
nand U4342 (N_4342,In_1059,In_856);
xnor U4343 (N_4343,In_228,In_1214);
xnor U4344 (N_4344,In_156,In_36);
or U4345 (N_4345,In_278,In_466);
or U4346 (N_4346,In_1474,In_349);
nand U4347 (N_4347,In_1003,In_1340);
nand U4348 (N_4348,In_1019,In_515);
nor U4349 (N_4349,In_168,In_717);
nand U4350 (N_4350,In_1432,In_1456);
nor U4351 (N_4351,In_634,In_1191);
or U4352 (N_4352,In_34,In_546);
nor U4353 (N_4353,In_578,In_1439);
nor U4354 (N_4354,In_278,In_330);
xor U4355 (N_4355,In_306,In_1045);
nand U4356 (N_4356,In_316,In_235);
nor U4357 (N_4357,In_790,In_1308);
and U4358 (N_4358,In_836,In_876);
nor U4359 (N_4359,In_300,In_699);
nand U4360 (N_4360,In_1409,In_603);
and U4361 (N_4361,In_793,In_759);
nand U4362 (N_4362,In_327,In_594);
or U4363 (N_4363,In_358,In_396);
nand U4364 (N_4364,In_1091,In_550);
nand U4365 (N_4365,In_1151,In_530);
nor U4366 (N_4366,In_1242,In_515);
or U4367 (N_4367,In_207,In_1445);
nor U4368 (N_4368,In_174,In_388);
xor U4369 (N_4369,In_634,In_149);
nand U4370 (N_4370,In_840,In_1330);
nor U4371 (N_4371,In_897,In_765);
or U4372 (N_4372,In_1128,In_351);
and U4373 (N_4373,In_903,In_1339);
or U4374 (N_4374,In_731,In_1050);
or U4375 (N_4375,In_656,In_315);
nand U4376 (N_4376,In_138,In_807);
and U4377 (N_4377,In_593,In_1486);
and U4378 (N_4378,In_366,In_649);
and U4379 (N_4379,In_163,In_4);
nand U4380 (N_4380,In_1277,In_1221);
nor U4381 (N_4381,In_1411,In_731);
nor U4382 (N_4382,In_1398,In_326);
nand U4383 (N_4383,In_101,In_215);
nor U4384 (N_4384,In_1032,In_1181);
nor U4385 (N_4385,In_1336,In_76);
nand U4386 (N_4386,In_988,In_718);
nor U4387 (N_4387,In_771,In_153);
and U4388 (N_4388,In_1069,In_1317);
nand U4389 (N_4389,In_409,In_1084);
or U4390 (N_4390,In_447,In_384);
nand U4391 (N_4391,In_346,In_241);
nand U4392 (N_4392,In_388,In_1162);
nor U4393 (N_4393,In_1061,In_609);
nor U4394 (N_4394,In_1379,In_212);
xnor U4395 (N_4395,In_68,In_334);
nor U4396 (N_4396,In_1350,In_982);
nand U4397 (N_4397,In_240,In_106);
or U4398 (N_4398,In_1285,In_845);
and U4399 (N_4399,In_440,In_795);
or U4400 (N_4400,In_1176,In_164);
nand U4401 (N_4401,In_5,In_949);
nand U4402 (N_4402,In_1063,In_53);
xnor U4403 (N_4403,In_1088,In_1081);
nand U4404 (N_4404,In_963,In_1224);
nand U4405 (N_4405,In_764,In_1154);
and U4406 (N_4406,In_1271,In_768);
and U4407 (N_4407,In_435,In_479);
or U4408 (N_4408,In_1230,In_585);
or U4409 (N_4409,In_443,In_12);
or U4410 (N_4410,In_14,In_43);
nor U4411 (N_4411,In_1358,In_366);
nor U4412 (N_4412,In_1019,In_916);
or U4413 (N_4413,In_168,In_438);
and U4414 (N_4414,In_791,In_1290);
nor U4415 (N_4415,In_725,In_185);
nand U4416 (N_4416,In_918,In_853);
and U4417 (N_4417,In_27,In_812);
nor U4418 (N_4418,In_1102,In_1275);
nand U4419 (N_4419,In_296,In_10);
nand U4420 (N_4420,In_1040,In_212);
and U4421 (N_4421,In_933,In_243);
and U4422 (N_4422,In_694,In_463);
nand U4423 (N_4423,In_60,In_1009);
nand U4424 (N_4424,In_749,In_495);
and U4425 (N_4425,In_324,In_275);
nand U4426 (N_4426,In_390,In_249);
and U4427 (N_4427,In_1307,In_352);
and U4428 (N_4428,In_861,In_257);
and U4429 (N_4429,In_901,In_1258);
or U4430 (N_4430,In_223,In_479);
xor U4431 (N_4431,In_1100,In_137);
and U4432 (N_4432,In_824,In_1406);
and U4433 (N_4433,In_28,In_620);
and U4434 (N_4434,In_757,In_189);
and U4435 (N_4435,In_1161,In_58);
nand U4436 (N_4436,In_483,In_316);
and U4437 (N_4437,In_1154,In_1243);
and U4438 (N_4438,In_1057,In_1370);
nand U4439 (N_4439,In_257,In_1204);
and U4440 (N_4440,In_332,In_1386);
xnor U4441 (N_4441,In_1217,In_951);
nor U4442 (N_4442,In_31,In_1294);
nand U4443 (N_4443,In_188,In_328);
and U4444 (N_4444,In_784,In_505);
or U4445 (N_4445,In_1242,In_146);
nand U4446 (N_4446,In_980,In_555);
or U4447 (N_4447,In_885,In_458);
or U4448 (N_4448,In_1065,In_1216);
or U4449 (N_4449,In_1244,In_374);
and U4450 (N_4450,In_1184,In_523);
and U4451 (N_4451,In_1460,In_681);
nor U4452 (N_4452,In_561,In_182);
or U4453 (N_4453,In_654,In_900);
and U4454 (N_4454,In_1392,In_838);
or U4455 (N_4455,In_289,In_310);
xor U4456 (N_4456,In_1254,In_842);
and U4457 (N_4457,In_946,In_330);
nor U4458 (N_4458,In_263,In_408);
and U4459 (N_4459,In_0,In_448);
nor U4460 (N_4460,In_777,In_683);
or U4461 (N_4461,In_515,In_432);
xnor U4462 (N_4462,In_1160,In_836);
nand U4463 (N_4463,In_498,In_230);
or U4464 (N_4464,In_1207,In_298);
nand U4465 (N_4465,In_695,In_294);
nor U4466 (N_4466,In_588,In_1115);
and U4467 (N_4467,In_469,In_779);
nand U4468 (N_4468,In_542,In_215);
nand U4469 (N_4469,In_453,In_1289);
and U4470 (N_4470,In_1049,In_987);
and U4471 (N_4471,In_453,In_17);
or U4472 (N_4472,In_777,In_490);
or U4473 (N_4473,In_1473,In_525);
xor U4474 (N_4474,In_888,In_217);
and U4475 (N_4475,In_51,In_343);
nand U4476 (N_4476,In_105,In_1180);
xnor U4477 (N_4477,In_1154,In_731);
nor U4478 (N_4478,In_1248,In_1138);
xnor U4479 (N_4479,In_1466,In_488);
or U4480 (N_4480,In_794,In_1159);
and U4481 (N_4481,In_333,In_572);
nand U4482 (N_4482,In_1270,In_164);
or U4483 (N_4483,In_1179,In_585);
nor U4484 (N_4484,In_1038,In_1435);
nor U4485 (N_4485,In_40,In_1222);
nor U4486 (N_4486,In_1377,In_762);
nand U4487 (N_4487,In_187,In_1296);
nor U4488 (N_4488,In_809,In_519);
nand U4489 (N_4489,In_1369,In_554);
xor U4490 (N_4490,In_1437,In_515);
and U4491 (N_4491,In_551,In_985);
and U4492 (N_4492,In_609,In_716);
nor U4493 (N_4493,In_959,In_293);
and U4494 (N_4494,In_440,In_267);
nor U4495 (N_4495,In_994,In_492);
or U4496 (N_4496,In_624,In_995);
nor U4497 (N_4497,In_327,In_813);
or U4498 (N_4498,In_592,In_260);
nand U4499 (N_4499,In_994,In_300);
or U4500 (N_4500,In_103,In_1183);
nor U4501 (N_4501,In_89,In_1023);
and U4502 (N_4502,In_1302,In_781);
nand U4503 (N_4503,In_965,In_1445);
nor U4504 (N_4504,In_603,In_714);
or U4505 (N_4505,In_1332,In_699);
nor U4506 (N_4506,In_1075,In_1295);
xnor U4507 (N_4507,In_479,In_313);
nand U4508 (N_4508,In_134,In_621);
and U4509 (N_4509,In_475,In_355);
or U4510 (N_4510,In_706,In_1180);
nand U4511 (N_4511,In_449,In_1221);
and U4512 (N_4512,In_477,In_715);
nand U4513 (N_4513,In_661,In_305);
nor U4514 (N_4514,In_802,In_1448);
nand U4515 (N_4515,In_1171,In_1014);
and U4516 (N_4516,In_764,In_769);
nor U4517 (N_4517,In_1451,In_1461);
or U4518 (N_4518,In_1254,In_61);
nor U4519 (N_4519,In_1310,In_912);
nor U4520 (N_4520,In_830,In_1257);
nor U4521 (N_4521,In_834,In_146);
or U4522 (N_4522,In_862,In_770);
nor U4523 (N_4523,In_209,In_166);
nand U4524 (N_4524,In_363,In_577);
nand U4525 (N_4525,In_1358,In_664);
or U4526 (N_4526,In_1039,In_826);
nand U4527 (N_4527,In_1265,In_694);
nor U4528 (N_4528,In_900,In_530);
or U4529 (N_4529,In_127,In_1207);
nor U4530 (N_4530,In_476,In_710);
and U4531 (N_4531,In_1256,In_932);
nor U4532 (N_4532,In_224,In_1078);
nor U4533 (N_4533,In_957,In_160);
and U4534 (N_4534,In_288,In_773);
and U4535 (N_4535,In_944,In_251);
or U4536 (N_4536,In_111,In_322);
and U4537 (N_4537,In_520,In_147);
nand U4538 (N_4538,In_842,In_368);
and U4539 (N_4539,In_432,In_127);
nand U4540 (N_4540,In_608,In_315);
or U4541 (N_4541,In_202,In_762);
xnor U4542 (N_4542,In_293,In_492);
and U4543 (N_4543,In_201,In_26);
nor U4544 (N_4544,In_582,In_658);
and U4545 (N_4545,In_749,In_1010);
nand U4546 (N_4546,In_163,In_734);
nand U4547 (N_4547,In_637,In_896);
nor U4548 (N_4548,In_102,In_951);
nor U4549 (N_4549,In_357,In_312);
and U4550 (N_4550,In_1446,In_1356);
or U4551 (N_4551,In_407,In_211);
nand U4552 (N_4552,In_1086,In_1355);
and U4553 (N_4553,In_309,In_1150);
and U4554 (N_4554,In_442,In_319);
nor U4555 (N_4555,In_374,In_837);
and U4556 (N_4556,In_511,In_825);
nor U4557 (N_4557,In_888,In_275);
nor U4558 (N_4558,In_1343,In_313);
and U4559 (N_4559,In_1293,In_1379);
nor U4560 (N_4560,In_1116,In_747);
or U4561 (N_4561,In_86,In_539);
or U4562 (N_4562,In_634,In_966);
nand U4563 (N_4563,In_590,In_230);
and U4564 (N_4564,In_1247,In_147);
and U4565 (N_4565,In_637,In_741);
nand U4566 (N_4566,In_675,In_48);
and U4567 (N_4567,In_443,In_1002);
and U4568 (N_4568,In_1479,In_24);
nor U4569 (N_4569,In_288,In_998);
nand U4570 (N_4570,In_1024,In_814);
nand U4571 (N_4571,In_152,In_1106);
nor U4572 (N_4572,In_83,In_1249);
or U4573 (N_4573,In_383,In_133);
nand U4574 (N_4574,In_444,In_1387);
nor U4575 (N_4575,In_1492,In_323);
and U4576 (N_4576,In_1466,In_788);
nand U4577 (N_4577,In_208,In_1484);
nor U4578 (N_4578,In_1379,In_696);
nand U4579 (N_4579,In_350,In_611);
or U4580 (N_4580,In_146,In_567);
xor U4581 (N_4581,In_192,In_697);
nand U4582 (N_4582,In_511,In_723);
nor U4583 (N_4583,In_1246,In_1449);
and U4584 (N_4584,In_68,In_652);
nor U4585 (N_4585,In_876,In_1281);
or U4586 (N_4586,In_1106,In_62);
nand U4587 (N_4587,In_1302,In_28);
and U4588 (N_4588,In_1445,In_200);
xnor U4589 (N_4589,In_831,In_1431);
and U4590 (N_4590,In_714,In_1200);
and U4591 (N_4591,In_484,In_713);
nor U4592 (N_4592,In_1383,In_6);
nand U4593 (N_4593,In_49,In_1261);
and U4594 (N_4594,In_416,In_664);
or U4595 (N_4595,In_116,In_1382);
xor U4596 (N_4596,In_153,In_1333);
nand U4597 (N_4597,In_165,In_397);
nor U4598 (N_4598,In_334,In_427);
or U4599 (N_4599,In_424,In_304);
and U4600 (N_4600,In_1204,In_952);
nand U4601 (N_4601,In_51,In_114);
xor U4602 (N_4602,In_943,In_1128);
and U4603 (N_4603,In_1011,In_988);
and U4604 (N_4604,In_80,In_853);
nor U4605 (N_4605,In_538,In_170);
nor U4606 (N_4606,In_1012,In_587);
or U4607 (N_4607,In_626,In_1420);
and U4608 (N_4608,In_133,In_1244);
nor U4609 (N_4609,In_1387,In_943);
nor U4610 (N_4610,In_732,In_173);
nand U4611 (N_4611,In_212,In_847);
and U4612 (N_4612,In_1002,In_639);
nor U4613 (N_4613,In_936,In_883);
nand U4614 (N_4614,In_823,In_480);
nor U4615 (N_4615,In_805,In_1075);
and U4616 (N_4616,In_621,In_454);
and U4617 (N_4617,In_262,In_1128);
or U4618 (N_4618,In_917,In_830);
nor U4619 (N_4619,In_74,In_1418);
and U4620 (N_4620,In_1094,In_1028);
nand U4621 (N_4621,In_1264,In_831);
xnor U4622 (N_4622,In_227,In_1048);
nor U4623 (N_4623,In_279,In_207);
nor U4624 (N_4624,In_294,In_182);
nand U4625 (N_4625,In_1444,In_371);
and U4626 (N_4626,In_1174,In_1056);
nand U4627 (N_4627,In_663,In_790);
nand U4628 (N_4628,In_1379,In_976);
nand U4629 (N_4629,In_1033,In_185);
and U4630 (N_4630,In_1360,In_570);
nor U4631 (N_4631,In_854,In_812);
xnor U4632 (N_4632,In_878,In_862);
nand U4633 (N_4633,In_201,In_830);
xnor U4634 (N_4634,In_789,In_1294);
nor U4635 (N_4635,In_1316,In_1267);
or U4636 (N_4636,In_1357,In_1288);
and U4637 (N_4637,In_1351,In_228);
nor U4638 (N_4638,In_1327,In_623);
and U4639 (N_4639,In_22,In_1469);
or U4640 (N_4640,In_196,In_582);
and U4641 (N_4641,In_258,In_704);
nor U4642 (N_4642,In_1186,In_1314);
or U4643 (N_4643,In_696,In_1415);
nor U4644 (N_4644,In_1197,In_423);
nor U4645 (N_4645,In_86,In_667);
nand U4646 (N_4646,In_501,In_1299);
nor U4647 (N_4647,In_585,In_65);
nand U4648 (N_4648,In_1164,In_962);
nand U4649 (N_4649,In_351,In_1014);
and U4650 (N_4650,In_499,In_1217);
nor U4651 (N_4651,In_735,In_238);
nor U4652 (N_4652,In_1027,In_1263);
and U4653 (N_4653,In_450,In_661);
and U4654 (N_4654,In_571,In_785);
nand U4655 (N_4655,In_1304,In_1431);
nor U4656 (N_4656,In_765,In_1183);
xor U4657 (N_4657,In_851,In_881);
nor U4658 (N_4658,In_1416,In_1392);
nand U4659 (N_4659,In_168,In_204);
and U4660 (N_4660,In_379,In_510);
xnor U4661 (N_4661,In_505,In_983);
nand U4662 (N_4662,In_1022,In_1042);
or U4663 (N_4663,In_122,In_8);
and U4664 (N_4664,In_1073,In_98);
nor U4665 (N_4665,In_1043,In_209);
xor U4666 (N_4666,In_1349,In_1081);
and U4667 (N_4667,In_67,In_390);
and U4668 (N_4668,In_634,In_843);
or U4669 (N_4669,In_794,In_657);
and U4670 (N_4670,In_436,In_985);
or U4671 (N_4671,In_574,In_798);
nor U4672 (N_4672,In_413,In_1183);
or U4673 (N_4673,In_813,In_797);
xnor U4674 (N_4674,In_863,In_472);
nand U4675 (N_4675,In_424,In_206);
and U4676 (N_4676,In_1154,In_310);
nor U4677 (N_4677,In_1033,In_586);
xor U4678 (N_4678,In_459,In_1487);
nor U4679 (N_4679,In_576,In_1200);
nand U4680 (N_4680,In_1424,In_371);
nor U4681 (N_4681,In_951,In_1206);
nor U4682 (N_4682,In_1005,In_1361);
and U4683 (N_4683,In_327,In_407);
nor U4684 (N_4684,In_31,In_1243);
and U4685 (N_4685,In_1353,In_610);
and U4686 (N_4686,In_1047,In_105);
nand U4687 (N_4687,In_716,In_148);
and U4688 (N_4688,In_56,In_759);
xor U4689 (N_4689,In_1251,In_1069);
nand U4690 (N_4690,In_245,In_411);
and U4691 (N_4691,In_1105,In_501);
nand U4692 (N_4692,In_812,In_24);
xor U4693 (N_4693,In_219,In_1182);
or U4694 (N_4694,In_1136,In_1369);
nor U4695 (N_4695,In_762,In_1273);
xor U4696 (N_4696,In_464,In_547);
xnor U4697 (N_4697,In_2,In_1193);
nand U4698 (N_4698,In_856,In_1376);
nand U4699 (N_4699,In_842,In_990);
or U4700 (N_4700,In_181,In_520);
and U4701 (N_4701,In_1036,In_1303);
or U4702 (N_4702,In_381,In_535);
or U4703 (N_4703,In_549,In_880);
or U4704 (N_4704,In_1115,In_563);
and U4705 (N_4705,In_109,In_627);
and U4706 (N_4706,In_46,In_570);
xor U4707 (N_4707,In_1487,In_1473);
xnor U4708 (N_4708,In_144,In_652);
or U4709 (N_4709,In_1115,In_345);
nor U4710 (N_4710,In_640,In_954);
nand U4711 (N_4711,In_1123,In_895);
xor U4712 (N_4712,In_820,In_1363);
nor U4713 (N_4713,In_1195,In_797);
or U4714 (N_4714,In_1135,In_649);
nor U4715 (N_4715,In_23,In_1131);
or U4716 (N_4716,In_554,In_504);
and U4717 (N_4717,In_737,In_424);
or U4718 (N_4718,In_963,In_159);
nor U4719 (N_4719,In_280,In_1479);
nor U4720 (N_4720,In_853,In_902);
nor U4721 (N_4721,In_1011,In_977);
or U4722 (N_4722,In_478,In_967);
nor U4723 (N_4723,In_1228,In_379);
and U4724 (N_4724,In_521,In_1061);
nand U4725 (N_4725,In_1267,In_642);
and U4726 (N_4726,In_1378,In_516);
and U4727 (N_4727,In_1160,In_282);
or U4728 (N_4728,In_594,In_616);
nor U4729 (N_4729,In_392,In_34);
nor U4730 (N_4730,In_802,In_182);
and U4731 (N_4731,In_1320,In_1489);
and U4732 (N_4732,In_843,In_1338);
nor U4733 (N_4733,In_932,In_1491);
nand U4734 (N_4734,In_1077,In_1001);
nand U4735 (N_4735,In_1483,In_1191);
nor U4736 (N_4736,In_26,In_862);
nor U4737 (N_4737,In_879,In_40);
and U4738 (N_4738,In_991,In_45);
and U4739 (N_4739,In_1314,In_275);
and U4740 (N_4740,In_15,In_558);
and U4741 (N_4741,In_838,In_425);
or U4742 (N_4742,In_890,In_229);
and U4743 (N_4743,In_656,In_1092);
nand U4744 (N_4744,In_1199,In_613);
nand U4745 (N_4745,In_644,In_1145);
nor U4746 (N_4746,In_1144,In_1411);
or U4747 (N_4747,In_58,In_123);
and U4748 (N_4748,In_798,In_1434);
nor U4749 (N_4749,In_14,In_461);
nand U4750 (N_4750,In_708,In_1382);
nor U4751 (N_4751,In_625,In_956);
nor U4752 (N_4752,In_764,In_240);
xnor U4753 (N_4753,In_670,In_845);
nor U4754 (N_4754,In_813,In_1139);
and U4755 (N_4755,In_451,In_348);
nor U4756 (N_4756,In_1005,In_1061);
nor U4757 (N_4757,In_1264,In_77);
or U4758 (N_4758,In_340,In_963);
nand U4759 (N_4759,In_1003,In_241);
nand U4760 (N_4760,In_654,In_1377);
nor U4761 (N_4761,In_1013,In_1203);
or U4762 (N_4762,In_1317,In_672);
or U4763 (N_4763,In_1479,In_1320);
or U4764 (N_4764,In_1126,In_1440);
nand U4765 (N_4765,In_932,In_1404);
nor U4766 (N_4766,In_1292,In_95);
nor U4767 (N_4767,In_233,In_153);
and U4768 (N_4768,In_135,In_352);
and U4769 (N_4769,In_781,In_752);
or U4770 (N_4770,In_218,In_415);
nand U4771 (N_4771,In_248,In_247);
and U4772 (N_4772,In_251,In_1362);
or U4773 (N_4773,In_636,In_156);
or U4774 (N_4774,In_192,In_450);
xor U4775 (N_4775,In_719,In_976);
nor U4776 (N_4776,In_126,In_894);
and U4777 (N_4777,In_307,In_770);
or U4778 (N_4778,In_470,In_1036);
or U4779 (N_4779,In_1064,In_721);
and U4780 (N_4780,In_468,In_93);
or U4781 (N_4781,In_1401,In_1270);
xnor U4782 (N_4782,In_988,In_172);
and U4783 (N_4783,In_561,In_645);
nand U4784 (N_4784,In_960,In_1408);
or U4785 (N_4785,In_138,In_1284);
nand U4786 (N_4786,In_954,In_424);
nand U4787 (N_4787,In_744,In_1195);
nand U4788 (N_4788,In_666,In_1276);
nand U4789 (N_4789,In_38,In_1280);
nand U4790 (N_4790,In_1357,In_179);
nor U4791 (N_4791,In_1410,In_1332);
nand U4792 (N_4792,In_262,In_385);
nor U4793 (N_4793,In_450,In_1092);
or U4794 (N_4794,In_15,In_1072);
nand U4795 (N_4795,In_221,In_410);
xor U4796 (N_4796,In_703,In_761);
xor U4797 (N_4797,In_454,In_238);
nor U4798 (N_4798,In_340,In_385);
nor U4799 (N_4799,In_41,In_1206);
and U4800 (N_4800,In_1081,In_257);
and U4801 (N_4801,In_1194,In_687);
or U4802 (N_4802,In_86,In_795);
and U4803 (N_4803,In_39,In_686);
nor U4804 (N_4804,In_688,In_183);
and U4805 (N_4805,In_1256,In_387);
and U4806 (N_4806,In_783,In_105);
or U4807 (N_4807,In_810,In_428);
or U4808 (N_4808,In_174,In_241);
or U4809 (N_4809,In_1340,In_661);
nand U4810 (N_4810,In_1389,In_319);
or U4811 (N_4811,In_292,In_74);
nand U4812 (N_4812,In_965,In_1252);
and U4813 (N_4813,In_801,In_857);
nor U4814 (N_4814,In_175,In_752);
nand U4815 (N_4815,In_325,In_717);
or U4816 (N_4816,In_160,In_1095);
and U4817 (N_4817,In_1485,In_1091);
and U4818 (N_4818,In_740,In_1094);
nor U4819 (N_4819,In_452,In_1034);
nand U4820 (N_4820,In_999,In_253);
and U4821 (N_4821,In_1463,In_792);
or U4822 (N_4822,In_474,In_105);
and U4823 (N_4823,In_25,In_1192);
and U4824 (N_4824,In_947,In_87);
nand U4825 (N_4825,In_187,In_1126);
and U4826 (N_4826,In_756,In_143);
and U4827 (N_4827,In_1398,In_84);
and U4828 (N_4828,In_497,In_1158);
xnor U4829 (N_4829,In_1366,In_899);
or U4830 (N_4830,In_458,In_765);
nand U4831 (N_4831,In_441,In_658);
nor U4832 (N_4832,In_344,In_1205);
nor U4833 (N_4833,In_991,In_1193);
and U4834 (N_4834,In_429,In_652);
nand U4835 (N_4835,In_779,In_712);
nor U4836 (N_4836,In_809,In_907);
nand U4837 (N_4837,In_607,In_1013);
and U4838 (N_4838,In_55,In_1093);
nand U4839 (N_4839,In_483,In_369);
or U4840 (N_4840,In_263,In_330);
and U4841 (N_4841,In_345,In_644);
nand U4842 (N_4842,In_839,In_1125);
and U4843 (N_4843,In_827,In_374);
or U4844 (N_4844,In_1434,In_87);
nor U4845 (N_4845,In_1390,In_818);
or U4846 (N_4846,In_288,In_1256);
xor U4847 (N_4847,In_949,In_528);
nor U4848 (N_4848,In_1484,In_583);
xnor U4849 (N_4849,In_1022,In_1187);
xnor U4850 (N_4850,In_755,In_552);
nor U4851 (N_4851,In_1393,In_314);
xnor U4852 (N_4852,In_223,In_6);
xnor U4853 (N_4853,In_1094,In_1480);
or U4854 (N_4854,In_1374,In_855);
xnor U4855 (N_4855,In_797,In_597);
and U4856 (N_4856,In_865,In_1220);
nand U4857 (N_4857,In_749,In_321);
nand U4858 (N_4858,In_1131,In_343);
or U4859 (N_4859,In_1007,In_286);
or U4860 (N_4860,In_577,In_101);
and U4861 (N_4861,In_91,In_813);
nand U4862 (N_4862,In_250,In_780);
and U4863 (N_4863,In_791,In_226);
and U4864 (N_4864,In_1199,In_739);
and U4865 (N_4865,In_800,In_390);
or U4866 (N_4866,In_60,In_934);
or U4867 (N_4867,In_1087,In_857);
and U4868 (N_4868,In_896,In_1310);
and U4869 (N_4869,In_240,In_568);
and U4870 (N_4870,In_392,In_1219);
or U4871 (N_4871,In_392,In_299);
xnor U4872 (N_4872,In_241,In_313);
nand U4873 (N_4873,In_1357,In_818);
nor U4874 (N_4874,In_265,In_1223);
and U4875 (N_4875,In_1308,In_13);
nand U4876 (N_4876,In_570,In_1484);
nand U4877 (N_4877,In_853,In_30);
or U4878 (N_4878,In_1152,In_738);
and U4879 (N_4879,In_833,In_1024);
nand U4880 (N_4880,In_129,In_752);
and U4881 (N_4881,In_324,In_1323);
nor U4882 (N_4882,In_373,In_1436);
and U4883 (N_4883,In_155,In_417);
or U4884 (N_4884,In_175,In_1218);
xnor U4885 (N_4885,In_1474,In_4);
nand U4886 (N_4886,In_66,In_951);
nand U4887 (N_4887,In_207,In_645);
and U4888 (N_4888,In_110,In_761);
nor U4889 (N_4889,In_785,In_1102);
xor U4890 (N_4890,In_292,In_1199);
and U4891 (N_4891,In_322,In_176);
and U4892 (N_4892,In_633,In_157);
and U4893 (N_4893,In_283,In_1473);
nor U4894 (N_4894,In_328,In_1260);
nand U4895 (N_4895,In_76,In_902);
nor U4896 (N_4896,In_1347,In_29);
nor U4897 (N_4897,In_1279,In_76);
or U4898 (N_4898,In_332,In_178);
nor U4899 (N_4899,In_608,In_6);
nor U4900 (N_4900,In_1060,In_1175);
nand U4901 (N_4901,In_577,In_1372);
and U4902 (N_4902,In_418,In_1115);
nor U4903 (N_4903,In_798,In_52);
or U4904 (N_4904,In_158,In_694);
xor U4905 (N_4905,In_1054,In_539);
or U4906 (N_4906,In_362,In_467);
or U4907 (N_4907,In_1342,In_862);
nand U4908 (N_4908,In_1430,In_642);
nand U4909 (N_4909,In_137,In_799);
nand U4910 (N_4910,In_455,In_315);
and U4911 (N_4911,In_1103,In_1178);
or U4912 (N_4912,In_1480,In_614);
nand U4913 (N_4913,In_937,In_674);
and U4914 (N_4914,In_32,In_688);
nand U4915 (N_4915,In_1009,In_270);
nor U4916 (N_4916,In_1327,In_315);
nand U4917 (N_4917,In_1002,In_1429);
nand U4918 (N_4918,In_453,In_897);
and U4919 (N_4919,In_1227,In_64);
or U4920 (N_4920,In_858,In_766);
xnor U4921 (N_4921,In_709,In_779);
or U4922 (N_4922,In_224,In_339);
or U4923 (N_4923,In_1352,In_412);
or U4924 (N_4924,In_819,In_229);
nand U4925 (N_4925,In_335,In_56);
and U4926 (N_4926,In_1101,In_963);
and U4927 (N_4927,In_1411,In_901);
nand U4928 (N_4928,In_542,In_1045);
and U4929 (N_4929,In_850,In_842);
nand U4930 (N_4930,In_350,In_661);
or U4931 (N_4931,In_1365,In_716);
and U4932 (N_4932,In_775,In_619);
nand U4933 (N_4933,In_1325,In_711);
or U4934 (N_4934,In_164,In_735);
nor U4935 (N_4935,In_568,In_205);
xor U4936 (N_4936,In_242,In_303);
nand U4937 (N_4937,In_1055,In_86);
nor U4938 (N_4938,In_901,In_793);
nand U4939 (N_4939,In_817,In_1142);
nand U4940 (N_4940,In_481,In_1426);
and U4941 (N_4941,In_823,In_1447);
and U4942 (N_4942,In_760,In_783);
nand U4943 (N_4943,In_1162,In_611);
xnor U4944 (N_4944,In_1129,In_1115);
and U4945 (N_4945,In_472,In_223);
or U4946 (N_4946,In_1119,In_244);
or U4947 (N_4947,In_1168,In_1099);
or U4948 (N_4948,In_290,In_395);
and U4949 (N_4949,In_936,In_1078);
xnor U4950 (N_4950,In_277,In_1412);
nor U4951 (N_4951,In_1240,In_824);
nor U4952 (N_4952,In_186,In_1330);
and U4953 (N_4953,In_568,In_1178);
xnor U4954 (N_4954,In_1201,In_14);
and U4955 (N_4955,In_1337,In_508);
nand U4956 (N_4956,In_477,In_1447);
nand U4957 (N_4957,In_1293,In_1129);
or U4958 (N_4958,In_1408,In_1064);
or U4959 (N_4959,In_58,In_474);
nor U4960 (N_4960,In_1199,In_1164);
or U4961 (N_4961,In_371,In_262);
or U4962 (N_4962,In_1226,In_1135);
and U4963 (N_4963,In_1143,In_177);
nand U4964 (N_4964,In_782,In_169);
xor U4965 (N_4965,In_408,In_895);
or U4966 (N_4966,In_445,In_752);
nor U4967 (N_4967,In_764,In_443);
or U4968 (N_4968,In_145,In_1445);
xor U4969 (N_4969,In_497,In_7);
nand U4970 (N_4970,In_247,In_417);
nand U4971 (N_4971,In_1249,In_432);
or U4972 (N_4972,In_410,In_1457);
and U4973 (N_4973,In_1153,In_446);
and U4974 (N_4974,In_1197,In_577);
nor U4975 (N_4975,In_150,In_841);
xnor U4976 (N_4976,In_479,In_987);
or U4977 (N_4977,In_673,In_777);
nand U4978 (N_4978,In_708,In_754);
or U4979 (N_4979,In_1418,In_1442);
xor U4980 (N_4980,In_1293,In_995);
and U4981 (N_4981,In_513,In_742);
and U4982 (N_4982,In_998,In_1063);
or U4983 (N_4983,In_374,In_1313);
xor U4984 (N_4984,In_247,In_244);
nor U4985 (N_4985,In_148,In_1296);
nor U4986 (N_4986,In_619,In_1353);
nor U4987 (N_4987,In_1379,In_273);
nand U4988 (N_4988,In_775,In_573);
or U4989 (N_4989,In_409,In_813);
or U4990 (N_4990,In_193,In_1399);
and U4991 (N_4991,In_577,In_1288);
or U4992 (N_4992,In_282,In_408);
xor U4993 (N_4993,In_1223,In_1312);
nor U4994 (N_4994,In_540,In_995);
nor U4995 (N_4995,In_291,In_1416);
xnor U4996 (N_4996,In_1053,In_552);
or U4997 (N_4997,In_1155,In_1228);
nand U4998 (N_4998,In_1220,In_99);
and U4999 (N_4999,In_125,In_560);
and U5000 (N_5000,N_4065,N_1999);
nand U5001 (N_5001,N_2206,N_3354);
nor U5002 (N_5002,N_4615,N_3935);
nor U5003 (N_5003,N_76,N_2698);
and U5004 (N_5004,N_3641,N_4800);
nor U5005 (N_5005,N_2277,N_650);
or U5006 (N_5006,N_4209,N_2756);
or U5007 (N_5007,N_1245,N_389);
xor U5008 (N_5008,N_1966,N_2487);
nor U5009 (N_5009,N_1791,N_4240);
nor U5010 (N_5010,N_1239,N_2604);
nor U5011 (N_5011,N_968,N_2526);
or U5012 (N_5012,N_1867,N_1337);
and U5013 (N_5013,N_3140,N_3341);
nand U5014 (N_5014,N_711,N_936);
and U5015 (N_5015,N_1428,N_4019);
and U5016 (N_5016,N_926,N_2796);
nor U5017 (N_5017,N_2385,N_511);
or U5018 (N_5018,N_2426,N_1353);
or U5019 (N_5019,N_143,N_64);
or U5020 (N_5020,N_2153,N_243);
nor U5021 (N_5021,N_1134,N_1125);
and U5022 (N_5022,N_544,N_61);
or U5023 (N_5023,N_3145,N_1233);
xnor U5024 (N_5024,N_4702,N_4253);
nor U5025 (N_5025,N_2328,N_669);
and U5026 (N_5026,N_823,N_2427);
and U5027 (N_5027,N_3106,N_3812);
nand U5028 (N_5028,N_1741,N_4134);
or U5029 (N_5029,N_2457,N_4119);
and U5030 (N_5030,N_4136,N_1361);
and U5031 (N_5031,N_3230,N_3207);
nand U5032 (N_5032,N_3380,N_4329);
nand U5033 (N_5033,N_1807,N_1121);
or U5034 (N_5034,N_489,N_2065);
nor U5035 (N_5035,N_578,N_1360);
nor U5036 (N_5036,N_3210,N_861);
nand U5037 (N_5037,N_1745,N_1435);
or U5038 (N_5038,N_1806,N_4631);
and U5039 (N_5039,N_771,N_3218);
and U5040 (N_5040,N_3400,N_1088);
xnor U5041 (N_5041,N_728,N_2629);
nand U5042 (N_5042,N_362,N_3128);
nand U5043 (N_5043,N_268,N_2);
nand U5044 (N_5044,N_3397,N_4250);
and U5045 (N_5045,N_3849,N_3945);
nor U5046 (N_5046,N_2996,N_3531);
and U5047 (N_5047,N_1029,N_2325);
nand U5048 (N_5048,N_2519,N_4137);
nor U5049 (N_5049,N_4741,N_4907);
xnor U5050 (N_5050,N_4767,N_1785);
xor U5051 (N_5051,N_4040,N_553);
or U5052 (N_5052,N_3367,N_2212);
nand U5053 (N_5053,N_4578,N_2908);
nor U5054 (N_5054,N_1303,N_3177);
nor U5055 (N_5055,N_2974,N_39);
or U5056 (N_5056,N_2360,N_2594);
or U5057 (N_5057,N_2407,N_4732);
xnor U5058 (N_5058,N_1605,N_66);
nand U5059 (N_5059,N_1574,N_1795);
and U5060 (N_5060,N_4048,N_121);
nand U5061 (N_5061,N_1302,N_4959);
nand U5062 (N_5062,N_87,N_3676);
nor U5063 (N_5063,N_2632,N_641);
nand U5064 (N_5064,N_164,N_2431);
nor U5065 (N_5065,N_37,N_2187);
xor U5066 (N_5066,N_4200,N_4377);
and U5067 (N_5067,N_481,N_2428);
or U5068 (N_5068,N_73,N_4906);
xnor U5069 (N_5069,N_4050,N_1209);
nor U5070 (N_5070,N_2418,N_4207);
nor U5071 (N_5071,N_4372,N_2762);
or U5072 (N_5072,N_699,N_1097);
or U5073 (N_5073,N_3977,N_4171);
and U5074 (N_5074,N_4326,N_2786);
or U5075 (N_5075,N_287,N_2667);
xor U5076 (N_5076,N_2343,N_2521);
or U5077 (N_5077,N_4052,N_1877);
nor U5078 (N_5078,N_3509,N_910);
nand U5079 (N_5079,N_3956,N_634);
or U5080 (N_5080,N_1194,N_658);
nand U5081 (N_5081,N_2572,N_835);
nor U5082 (N_5082,N_4966,N_3603);
nand U5083 (N_5083,N_4573,N_4391);
and U5084 (N_5084,N_474,N_135);
nand U5085 (N_5085,N_2848,N_2913);
and U5086 (N_5086,N_3768,N_4092);
xor U5087 (N_5087,N_2522,N_1102);
and U5088 (N_5088,N_3348,N_3115);
nand U5089 (N_5089,N_2186,N_2546);
nand U5090 (N_5090,N_4331,N_1611);
or U5091 (N_5091,N_3907,N_3396);
and U5092 (N_5092,N_4911,N_3663);
or U5093 (N_5093,N_3474,N_4368);
nand U5094 (N_5094,N_1851,N_1646);
and U5095 (N_5095,N_2134,N_4104);
nor U5096 (N_5096,N_2250,N_3105);
or U5097 (N_5097,N_809,N_954);
nand U5098 (N_5098,N_333,N_4210);
nand U5099 (N_5099,N_991,N_2367);
nand U5100 (N_5100,N_2997,N_4698);
nor U5101 (N_5101,N_3614,N_2067);
or U5102 (N_5102,N_2718,N_3906);
nor U5103 (N_5103,N_4729,N_2834);
nor U5104 (N_5104,N_3905,N_1398);
nor U5105 (N_5105,N_2649,N_1478);
or U5106 (N_5106,N_985,N_478);
nor U5107 (N_5107,N_1790,N_922);
and U5108 (N_5108,N_849,N_4362);
and U5109 (N_5109,N_888,N_3025);
nand U5110 (N_5110,N_2740,N_3413);
nor U5111 (N_5111,N_515,N_2617);
nor U5112 (N_5112,N_2927,N_2489);
nand U5113 (N_5113,N_3087,N_3781);
nand U5114 (N_5114,N_3858,N_3371);
xnor U5115 (N_5115,N_4298,N_4941);
xnor U5116 (N_5116,N_1828,N_3510);
nor U5117 (N_5117,N_4601,N_295);
or U5118 (N_5118,N_4353,N_3517);
nand U5119 (N_5119,N_1467,N_847);
nand U5120 (N_5120,N_518,N_56);
or U5121 (N_5121,N_2788,N_2413);
xor U5122 (N_5122,N_4416,N_2823);
nand U5123 (N_5123,N_3112,N_562);
nor U5124 (N_5124,N_2851,N_3052);
and U5125 (N_5125,N_3859,N_4289);
and U5126 (N_5126,N_4076,N_3308);
xor U5127 (N_5127,N_907,N_4921);
nor U5128 (N_5128,N_1271,N_4196);
and U5129 (N_5129,N_1408,N_4621);
and U5130 (N_5130,N_4056,N_4726);
nor U5131 (N_5131,N_4228,N_419);
nand U5132 (N_5132,N_2877,N_3469);
and U5133 (N_5133,N_690,N_3164);
xor U5134 (N_5134,N_2540,N_794);
nor U5135 (N_5135,N_2031,N_2085);
nor U5136 (N_5136,N_4697,N_2759);
xor U5137 (N_5137,N_7,N_4044);
nand U5138 (N_5138,N_1046,N_2100);
nand U5139 (N_5139,N_3243,N_3989);
xnor U5140 (N_5140,N_4357,N_1942);
and U5141 (N_5141,N_315,N_2801);
nor U5142 (N_5142,N_2044,N_181);
or U5143 (N_5143,N_3636,N_2636);
or U5144 (N_5144,N_606,N_4806);
nor U5145 (N_5145,N_4748,N_3002);
and U5146 (N_5146,N_3840,N_1368);
or U5147 (N_5147,N_1433,N_1815);
nand U5148 (N_5148,N_852,N_929);
nor U5149 (N_5149,N_1796,N_4672);
nor U5150 (N_5150,N_3537,N_4675);
and U5151 (N_5151,N_318,N_455);
and U5152 (N_5152,N_4097,N_4917);
and U5153 (N_5153,N_2215,N_1734);
and U5154 (N_5154,N_3362,N_1446);
and U5155 (N_5155,N_3000,N_1554);
and U5156 (N_5156,N_4860,N_2993);
and U5157 (N_5157,N_2003,N_322);
or U5158 (N_5158,N_3556,N_2852);
and U5159 (N_5159,N_4833,N_2755);
or U5160 (N_5160,N_134,N_1172);
nor U5161 (N_5161,N_2259,N_241);
or U5162 (N_5162,N_1445,N_2873);
or U5163 (N_5163,N_4643,N_543);
nand U5164 (N_5164,N_3158,N_1567);
or U5165 (N_5165,N_3761,N_574);
nor U5166 (N_5166,N_885,N_356);
nand U5167 (N_5167,N_1104,N_447);
nor U5168 (N_5168,N_3794,N_2822);
and U5169 (N_5169,N_897,N_242);
nand U5170 (N_5170,N_4255,N_2789);
nor U5171 (N_5171,N_4584,N_453);
nor U5172 (N_5172,N_3877,N_948);
or U5173 (N_5173,N_4001,N_2799);
nand U5174 (N_5174,N_3608,N_1719);
nor U5175 (N_5175,N_276,N_1925);
nor U5176 (N_5176,N_1002,N_24);
nand U5177 (N_5177,N_4920,N_984);
or U5178 (N_5178,N_4743,N_1026);
nand U5179 (N_5179,N_4075,N_4905);
and U5180 (N_5180,N_3757,N_3346);
or U5181 (N_5181,N_4246,N_280);
nand U5182 (N_5182,N_4229,N_615);
xor U5183 (N_5183,N_4144,N_2430);
nand U5184 (N_5184,N_1802,N_3003);
nor U5185 (N_5185,N_789,N_3670);
nor U5186 (N_5186,N_2610,N_668);
and U5187 (N_5187,N_4389,N_4722);
nand U5188 (N_5188,N_585,N_2229);
or U5189 (N_5189,N_36,N_4036);
or U5190 (N_5190,N_4664,N_4063);
or U5191 (N_5191,N_696,N_4283);
nand U5192 (N_5192,N_2497,N_2790);
or U5193 (N_5193,N_1938,N_1436);
nor U5194 (N_5194,N_449,N_102);
or U5195 (N_5195,N_4031,N_602);
nand U5196 (N_5196,N_4463,N_1915);
xnor U5197 (N_5197,N_841,N_2271);
nand U5198 (N_5198,N_1346,N_540);
nand U5199 (N_5199,N_4466,N_3828);
nor U5200 (N_5200,N_50,N_4378);
nand U5201 (N_5201,N_3780,N_491);
xor U5202 (N_5202,N_2897,N_1120);
or U5203 (N_5203,N_4205,N_2387);
nand U5204 (N_5204,N_867,N_4013);
or U5205 (N_5205,N_1399,N_586);
and U5206 (N_5206,N_1631,N_695);
xnor U5207 (N_5207,N_3853,N_189);
xnor U5208 (N_5208,N_4891,N_4354);
and U5209 (N_5209,N_4894,N_4296);
and U5210 (N_5210,N_4269,N_2356);
or U5211 (N_5211,N_4842,N_2797);
or U5212 (N_5212,N_2911,N_3523);
nand U5213 (N_5213,N_682,N_3898);
or U5214 (N_5214,N_3173,N_2599);
nand U5215 (N_5215,N_2716,N_4451);
xnor U5216 (N_5216,N_2432,N_2013);
nand U5217 (N_5217,N_1893,N_1821);
and U5218 (N_5218,N_2240,N_4565);
nand U5219 (N_5219,N_4035,N_248);
nor U5220 (N_5220,N_2143,N_1268);
or U5221 (N_5221,N_2712,N_4945);
nor U5222 (N_5222,N_4895,N_381);
nor U5223 (N_5223,N_63,N_2006);
nand U5224 (N_5224,N_1639,N_3999);
nor U5225 (N_5225,N_85,N_2383);
or U5226 (N_5226,N_3805,N_4147);
nor U5227 (N_5227,N_2892,N_440);
nor U5228 (N_5228,N_2750,N_3918);
xnor U5229 (N_5229,N_548,N_3008);
nor U5230 (N_5230,N_636,N_2254);
and U5231 (N_5231,N_4381,N_2009);
and U5232 (N_5232,N_401,N_1941);
nand U5233 (N_5233,N_1697,N_4591);
or U5234 (N_5234,N_3649,N_1038);
nand U5235 (N_5235,N_4193,N_4666);
nand U5236 (N_5236,N_2373,N_1106);
nor U5237 (N_5237,N_2896,N_3508);
nor U5238 (N_5238,N_3719,N_4469);
nand U5239 (N_5239,N_4878,N_2425);
nor U5240 (N_5240,N_4370,N_1524);
or U5241 (N_5241,N_3643,N_1119);
or U5242 (N_5242,N_2630,N_1555);
nand U5243 (N_5243,N_537,N_1873);
nor U5244 (N_5244,N_3047,N_1047);
or U5245 (N_5245,N_2298,N_2995);
and U5246 (N_5246,N_3248,N_3806);
nand U5247 (N_5247,N_1579,N_4956);
or U5248 (N_5248,N_4815,N_818);
and U5249 (N_5249,N_4140,N_4058);
nor U5250 (N_5250,N_2622,N_508);
or U5251 (N_5251,N_4765,N_2050);
nor U5252 (N_5252,N_843,N_4940);
nand U5253 (N_5253,N_3810,N_3921);
or U5254 (N_5254,N_417,N_1378);
and U5255 (N_5255,N_1855,N_408);
and U5256 (N_5256,N_1421,N_1765);
nor U5257 (N_5257,N_4838,N_196);
and U5258 (N_5258,N_750,N_4819);
or U5259 (N_5259,N_277,N_3317);
or U5260 (N_5260,N_2701,N_1927);
nor U5261 (N_5261,N_4768,N_3657);
or U5262 (N_5262,N_448,N_2929);
xnor U5263 (N_5263,N_3707,N_1318);
nand U5264 (N_5264,N_3738,N_3333);
or U5265 (N_5265,N_4008,N_4609);
nand U5266 (N_5266,N_1799,N_424);
xnor U5267 (N_5267,N_3798,N_532);
nand U5268 (N_5268,N_3094,N_721);
nor U5269 (N_5269,N_795,N_330);
nand U5270 (N_5270,N_2722,N_1737);
or U5271 (N_5271,N_3040,N_4996);
or U5272 (N_5272,N_2653,N_1919);
nor U5273 (N_5273,N_785,N_3984);
nand U5274 (N_5274,N_4449,N_3815);
or U5275 (N_5275,N_1978,N_490);
nand U5276 (N_5276,N_1278,N_4101);
nor U5277 (N_5277,N_10,N_3401);
xnor U5278 (N_5278,N_4915,N_1515);
or U5279 (N_5279,N_3571,N_4005);
nand U5280 (N_5280,N_1533,N_4641);
nor U5281 (N_5281,N_4060,N_2481);
xnor U5282 (N_5282,N_140,N_4173);
nor U5283 (N_5283,N_1808,N_2902);
or U5284 (N_5284,N_4902,N_935);
or U5285 (N_5285,N_2160,N_2948);
or U5286 (N_5286,N_3804,N_1382);
or U5287 (N_5287,N_1934,N_2399);
and U5288 (N_5288,N_2598,N_2939);
nand U5289 (N_5289,N_2347,N_2045);
nor U5290 (N_5290,N_2348,N_132);
nand U5291 (N_5291,N_3573,N_3208);
nor U5292 (N_5292,N_640,N_2248);
xnor U5293 (N_5293,N_3829,N_4775);
or U5294 (N_5294,N_4066,N_4841);
nand U5295 (N_5295,N_2607,N_139);
or U5296 (N_5296,N_3240,N_3438);
nand U5297 (N_5297,N_3493,N_297);
xor U5298 (N_5298,N_3152,N_499);
nor U5299 (N_5299,N_1753,N_1);
nand U5300 (N_5300,N_1173,N_1036);
xnor U5301 (N_5301,N_2841,N_321);
or U5302 (N_5302,N_4410,N_3314);
xnor U5303 (N_5303,N_1014,N_2438);
nor U5304 (N_5304,N_270,N_3626);
and U5305 (N_5305,N_4382,N_2221);
nand U5306 (N_5306,N_3419,N_4241);
and U5307 (N_5307,N_2077,N_4829);
or U5308 (N_5308,N_67,N_3514);
nor U5309 (N_5309,N_3272,N_148);
nand U5310 (N_5310,N_514,N_1838);
nor U5311 (N_5311,N_1082,N_4432);
nand U5312 (N_5312,N_1469,N_4394);
or U5313 (N_5313,N_1731,N_4464);
and U5314 (N_5314,N_4476,N_4674);
or U5315 (N_5315,N_2560,N_476);
nand U5316 (N_5316,N_870,N_863);
nor U5317 (N_5317,N_4564,N_1576);
and U5318 (N_5318,N_1261,N_4349);
nand U5319 (N_5319,N_3163,N_4753);
nand U5320 (N_5320,N_3350,N_137);
nor U5321 (N_5321,N_1405,N_1888);
or U5322 (N_5322,N_1908,N_4492);
nor U5323 (N_5323,N_1279,N_388);
and U5324 (N_5324,N_790,N_4976);
and U5325 (N_5325,N_3251,N_479);
nand U5326 (N_5326,N_1336,N_2810);
or U5327 (N_5327,N_3119,N_2439);
nor U5328 (N_5328,N_2916,N_1392);
and U5329 (N_5329,N_2469,N_1006);
nor U5330 (N_5330,N_1073,N_2233);
and U5331 (N_5331,N_4582,N_1115);
nor U5332 (N_5332,N_4541,N_1461);
nand U5333 (N_5333,N_1714,N_4595);
nand U5334 (N_5334,N_2069,N_2331);
and U5335 (N_5335,N_2375,N_933);
or U5336 (N_5336,N_1003,N_2128);
nor U5337 (N_5337,N_2861,N_198);
and U5338 (N_5338,N_3760,N_4855);
and U5339 (N_5339,N_811,N_4236);
xnor U5340 (N_5340,N_4531,N_2976);
nand U5341 (N_5341,N_1845,N_1389);
nor U5342 (N_5342,N_1671,N_990);
nand U5343 (N_5343,N_2696,N_2682);
nor U5344 (N_5344,N_3767,N_384);
nor U5345 (N_5345,N_1441,N_1775);
or U5346 (N_5346,N_2269,N_1198);
nor U5347 (N_5347,N_3961,N_3733);
nand U5348 (N_5348,N_2000,N_956);
nand U5349 (N_5349,N_3518,N_4094);
xnor U5350 (N_5350,N_3561,N_1559);
nand U5351 (N_5351,N_247,N_1191);
or U5352 (N_5352,N_2026,N_724);
nand U5353 (N_5353,N_1219,N_3363);
and U5354 (N_5354,N_1730,N_663);
nand U5355 (N_5355,N_1393,N_3028);
and U5356 (N_5356,N_2666,N_3437);
or U5357 (N_5357,N_188,N_4203);
or U5358 (N_5358,N_291,N_4662);
xnor U5359 (N_5359,N_317,N_1819);
or U5360 (N_5360,N_3309,N_3712);
or U5361 (N_5361,N_3709,N_2391);
xnor U5362 (N_5362,N_15,N_1650);
or U5363 (N_5363,N_3577,N_18);
xnor U5364 (N_5364,N_2954,N_1188);
nand U5365 (N_5365,N_1666,N_2648);
nor U5366 (N_5366,N_2825,N_848);
xnor U5367 (N_5367,N_3644,N_4170);
and U5368 (N_5368,N_71,N_764);
nand U5369 (N_5369,N_3943,N_1606);
nor U5370 (N_5370,N_2595,N_288);
and U5371 (N_5371,N_1301,N_2422);
or U5372 (N_5372,N_3440,N_624);
or U5373 (N_5373,N_454,N_1472);
xor U5374 (N_5374,N_3927,N_1385);
or U5375 (N_5375,N_3963,N_3558);
nand U5376 (N_5376,N_2188,N_2404);
xnor U5377 (N_5377,N_3069,N_752);
nor U5378 (N_5378,N_4846,N_3847);
nor U5379 (N_5379,N_4095,N_4007);
nand U5380 (N_5380,N_1933,N_917);
xnor U5381 (N_5381,N_4716,N_3807);
nor U5382 (N_5382,N_892,N_1911);
and U5383 (N_5383,N_4714,N_4089);
nand U5384 (N_5384,N_2910,N_3058);
xor U5385 (N_5385,N_1876,N_3741);
or U5386 (N_5386,N_2196,N_170);
nor U5387 (N_5387,N_261,N_589);
or U5388 (N_5388,N_1993,N_1707);
and U5389 (N_5389,N_4696,N_531);
or U5390 (N_5390,N_2286,N_2864);
and U5391 (N_5391,N_2219,N_1608);
or U5392 (N_5392,N_1422,N_4887);
nand U5393 (N_5393,N_3347,N_1166);
nor U5394 (N_5394,N_2849,N_1369);
xnor U5395 (N_5395,N_1983,N_2455);
and U5396 (N_5396,N_672,N_1388);
nor U5397 (N_5397,N_4683,N_3234);
or U5398 (N_5398,N_3349,N_186);
or U5399 (N_5399,N_1497,N_3791);
nor U5400 (N_5400,N_1149,N_1871);
nor U5401 (N_5401,N_4169,N_1957);
and U5402 (N_5402,N_2032,N_4736);
nor U5403 (N_5403,N_2859,N_3484);
nor U5404 (N_5404,N_3964,N_2978);
nor U5405 (N_5405,N_231,N_1442);
nand U5406 (N_5406,N_3273,N_3216);
nand U5407 (N_5407,N_1585,N_1503);
nor U5408 (N_5408,N_693,N_41);
and U5409 (N_5409,N_2818,N_3200);
or U5410 (N_5410,N_3778,N_1215);
nand U5411 (N_5411,N_4330,N_1454);
nor U5412 (N_5412,N_705,N_1685);
nand U5413 (N_5413,N_1406,N_3458);
or U5414 (N_5414,N_2541,N_2255);
xor U5415 (N_5415,N_185,N_3465);
and U5416 (N_5416,N_3700,N_4374);
nor U5417 (N_5417,N_4886,N_2287);
nor U5418 (N_5418,N_3129,N_733);
nand U5419 (N_5419,N_4213,N_3045);
and U5420 (N_5420,N_2224,N_3180);
nor U5421 (N_5421,N_1507,N_3749);
or U5422 (N_5422,N_1694,N_2289);
nor U5423 (N_5423,N_4195,N_3973);
nor U5424 (N_5424,N_2544,N_2891);
or U5425 (N_5425,N_4529,N_1327);
and U5426 (N_5426,N_2491,N_3);
nor U5427 (N_5427,N_1858,N_4017);
or U5428 (N_5428,N_503,N_3001);
nor U5429 (N_5429,N_3629,N_1429);
and U5430 (N_5430,N_3311,N_3247);
or U5431 (N_5431,N_4133,N_3376);
nor U5432 (N_5432,N_83,N_1072);
nor U5433 (N_5433,N_1265,N_1904);
nand U5434 (N_5434,N_4681,N_2882);
xor U5435 (N_5435,N_1375,N_4419);
and U5436 (N_5436,N_4212,N_4371);
or U5437 (N_5437,N_2177,N_3364);
nor U5438 (N_5438,N_773,N_4975);
nor U5439 (N_5439,N_2127,N_2819);
and U5440 (N_5440,N_4218,N_4030);
nand U5441 (N_5441,N_3193,N_727);
xnor U5442 (N_5442,N_2965,N_4226);
and U5443 (N_5443,N_390,N_3845);
nand U5444 (N_5444,N_2454,N_1324);
and U5445 (N_5445,N_2461,N_4239);
or U5446 (N_5446,N_498,N_4157);
nor U5447 (N_5447,N_4225,N_1913);
nand U5448 (N_5448,N_2173,N_3773);
xnor U5449 (N_5449,N_172,N_868);
or U5450 (N_5450,N_97,N_168);
and U5451 (N_5451,N_521,N_1623);
and U5452 (N_5452,N_4339,N_127);
and U5453 (N_5453,N_2043,N_4460);
and U5454 (N_5454,N_3107,N_1651);
nor U5455 (N_5455,N_2022,N_2472);
nand U5456 (N_5456,N_2523,N_3992);
nor U5457 (N_5457,N_3222,N_1332);
or U5458 (N_5458,N_678,N_475);
nand U5459 (N_5459,N_599,N_4712);
or U5460 (N_5460,N_3132,N_3278);
nand U5461 (N_5461,N_4158,N_762);
nand U5462 (N_5462,N_1415,N_569);
nor U5463 (N_5463,N_3360,N_1976);
nand U5464 (N_5464,N_3692,N_3904);
nand U5465 (N_5465,N_3383,N_2072);
nor U5466 (N_5466,N_2372,N_2914);
nor U5467 (N_5467,N_3968,N_2014);
or U5468 (N_5468,N_755,N_334);
and U5469 (N_5469,N_3777,N_2366);
and U5470 (N_5470,N_4291,N_660);
or U5471 (N_5471,N_776,N_3550);
nand U5472 (N_5472,N_1460,N_2922);
nor U5473 (N_5473,N_416,N_1669);
nor U5474 (N_5474,N_793,N_4152);
nand U5475 (N_5475,N_4851,N_3135);
and U5476 (N_5476,N_1695,N_3734);
nand U5477 (N_5477,N_30,N_3082);
nor U5478 (N_5478,N_2327,N_1833);
and U5479 (N_5479,N_1617,N_633);
and U5480 (N_5480,N_946,N_1133);
nand U5481 (N_5481,N_4561,N_463);
nor U5482 (N_5482,N_2549,N_4143);
xor U5483 (N_5483,N_3192,N_1284);
and U5484 (N_5484,N_1401,N_4340);
and U5485 (N_5485,N_662,N_2641);
or U5486 (N_5486,N_3451,N_1206);
nor U5487 (N_5487,N_2613,N_3928);
and U5488 (N_5488,N_4079,N_677);
nor U5489 (N_5489,N_4360,N_3224);
nand U5490 (N_5490,N_496,N_1773);
nor U5491 (N_5491,N_1109,N_232);
nor U5492 (N_5492,N_4148,N_2525);
and U5493 (N_5493,N_431,N_4957);
and U5494 (N_5494,N_3096,N_2977);
nand U5495 (N_5495,N_1162,N_1224);
nor U5496 (N_5496,N_2833,N_689);
or U5497 (N_5497,N_2903,N_2563);
xor U5498 (N_5498,N_3519,N_2757);
and U5499 (N_5499,N_1295,N_1456);
nand U5500 (N_5500,N_207,N_3390);
nor U5501 (N_5501,N_1403,N_379);
and U5502 (N_5502,N_1201,N_1420);
nor U5503 (N_5503,N_3103,N_1747);
nor U5504 (N_5504,N_2941,N_4754);
or U5505 (N_5505,N_1766,N_4764);
nand U5506 (N_5506,N_4408,N_1015);
or U5507 (N_5507,N_1080,N_3729);
xnor U5508 (N_5508,N_4475,N_4034);
and U5509 (N_5509,N_301,N_1584);
xor U5510 (N_5510,N_1609,N_4083);
and U5511 (N_5511,N_4918,N_4122);
or U5512 (N_5512,N_4725,N_1214);
nand U5513 (N_5513,N_3885,N_3015);
nor U5514 (N_5514,N_4358,N_4820);
xor U5515 (N_5515,N_2638,N_1672);
nand U5516 (N_5516,N_1792,N_2083);
xor U5517 (N_5517,N_3104,N_1110);
xor U5518 (N_5518,N_3165,N_2424);
nor U5519 (N_5519,N_4575,N_2130);
and U5520 (N_5520,N_2550,N_4088);
and U5521 (N_5521,N_4880,N_2753);
xnor U5522 (N_5522,N_4916,N_3338);
or U5523 (N_5523,N_4870,N_200);
xnor U5524 (N_5524,N_1811,N_2602);
and U5525 (N_5525,N_2267,N_519);
nor U5526 (N_5526,N_4084,N_1306);
and U5527 (N_5527,N_4505,N_1699);
nand U5528 (N_5528,N_3392,N_197);
or U5529 (N_5529,N_3793,N_1857);
xor U5530 (N_5530,N_2213,N_1820);
xnor U5531 (N_5531,N_2062,N_3753);
xnor U5532 (N_5532,N_4086,N_2673);
nand U5533 (N_5533,N_194,N_959);
nand U5534 (N_5534,N_3996,N_3634);
or U5535 (N_5535,N_925,N_736);
nor U5536 (N_5536,N_1391,N_4482);
or U5537 (N_5537,N_1103,N_349);
or U5538 (N_5538,N_95,N_2582);
or U5539 (N_5539,N_2702,N_3985);
nor U5540 (N_5540,N_4055,N_4292);
and U5541 (N_5541,N_4166,N_2732);
and U5542 (N_5542,N_2496,N_3512);
nor U5543 (N_5543,N_1241,N_3220);
nand U5544 (N_5544,N_3095,N_2222);
nor U5545 (N_5545,N_4530,N_4650);
nand U5546 (N_5546,N_212,N_1410);
and U5547 (N_5547,N_942,N_421);
nor U5548 (N_5548,N_1329,N_1298);
and U5549 (N_5549,N_441,N_3442);
or U5550 (N_5550,N_1184,N_1289);
or U5551 (N_5551,N_1553,N_2290);
and U5552 (N_5552,N_2410,N_4993);
or U5553 (N_5553,N_1527,N_3598);
and U5554 (N_5554,N_3244,N_2983);
nand U5555 (N_5555,N_2713,N_3587);
or U5556 (N_5556,N_4572,N_3183);
nand U5557 (N_5557,N_3219,N_461);
xnor U5558 (N_5558,N_4532,N_3126);
or U5559 (N_5559,N_233,N_704);
and U5560 (N_5560,N_1453,N_2088);
nor U5561 (N_5561,N_2104,N_79);
nand U5562 (N_5562,N_1449,N_2202);
nor U5563 (N_5563,N_4642,N_1069);
nor U5564 (N_5564,N_4596,N_3637);
and U5565 (N_5565,N_2476,N_3073);
nor U5566 (N_5566,N_1634,N_4102);
and U5567 (N_5567,N_2835,N_4801);
xor U5568 (N_5568,N_2612,N_4009);
and U5569 (N_5569,N_3576,N_1086);
nor U5570 (N_5570,N_2813,N_4123);
or U5571 (N_5571,N_1678,N_1190);
nor U5572 (N_5572,N_4995,N_193);
nand U5573 (N_5573,N_2775,N_1117);
nor U5574 (N_5574,N_4670,N_4311);
nand U5575 (N_5575,N_1018,N_4398);
nand U5576 (N_5576,N_4570,N_4049);
or U5577 (N_5577,N_1081,N_228);
nand U5578 (N_5578,N_2952,N_989);
nor U5579 (N_5579,N_238,N_2618);
and U5580 (N_5580,N_2087,N_3168);
xnor U5581 (N_5581,N_1540,N_361);
and U5582 (N_5582,N_1179,N_882);
nand U5583 (N_5583,N_4407,N_1762);
or U5584 (N_5584,N_1060,N_4780);
and U5585 (N_5585,N_458,N_1750);
or U5586 (N_5586,N_2693,N_4261);
nand U5587 (N_5587,N_664,N_208);
or U5588 (N_5588,N_3274,N_828);
nand U5589 (N_5589,N_4647,N_3495);
and U5590 (N_5590,N_3099,N_1805);
and U5591 (N_5591,N_3994,N_4189);
or U5592 (N_5592,N_1980,N_2596);
nor U5593 (N_5593,N_3978,N_2398);
or U5594 (N_5594,N_928,N_783);
xor U5595 (N_5595,N_1656,N_3141);
nand U5596 (N_5596,N_2152,N_1593);
nor U5597 (N_5597,N_4904,N_4939);
nor U5598 (N_5598,N_4731,N_4737);
or U5599 (N_5599,N_1023,N_1012);
nor U5600 (N_5600,N_110,N_1708);
nor U5601 (N_5601,N_2225,N_4301);
xor U5602 (N_5602,N_2076,N_2817);
and U5603 (N_5603,N_4843,N_1591);
and U5604 (N_5604,N_4898,N_568);
or U5605 (N_5605,N_4333,N_1087);
and U5606 (N_5606,N_1757,N_3452);
nand U5607 (N_5607,N_3237,N_4925);
or U5608 (N_5608,N_2812,N_3920);
nor U5609 (N_5609,N_1374,N_2646);
or U5610 (N_5610,N_1092,N_2587);
or U5611 (N_5611,N_3620,N_3116);
xnor U5612 (N_5612,N_2265,N_674);
and U5613 (N_5613,N_4438,N_554);
nand U5614 (N_5614,N_2114,N_4411);
or U5615 (N_5615,N_1658,N_2513);
nor U5616 (N_5616,N_2020,N_3701);
and U5617 (N_5617,N_1798,N_4808);
nor U5618 (N_5618,N_1779,N_1160);
or U5619 (N_5619,N_2482,N_3880);
nand U5620 (N_5620,N_1962,N_1287);
and U5621 (N_5621,N_404,N_1655);
nor U5622 (N_5622,N_3619,N_302);
nand U5623 (N_5623,N_4965,N_3085);
nand U5624 (N_5624,N_4400,N_1466);
nand U5625 (N_5625,N_3933,N_2056);
xor U5626 (N_5626,N_1124,N_2095);
nand U5627 (N_5627,N_3894,N_0);
or U5628 (N_5628,N_187,N_3854);
nand U5629 (N_5629,N_14,N_3264);
and U5630 (N_5630,N_1660,N_975);
or U5631 (N_5631,N_1681,N_1434);
or U5632 (N_5632,N_4622,N_3948);
nand U5633 (N_5633,N_1457,N_4569);
and U5634 (N_5634,N_1771,N_4576);
xnor U5635 (N_5635,N_3063,N_2600);
nand U5636 (N_5636,N_960,N_3051);
and U5637 (N_5637,N_4054,N_4625);
or U5638 (N_5638,N_4555,N_3589);
or U5639 (N_5639,N_3211,N_2764);
nor U5640 (N_5640,N_3525,N_1034);
and U5641 (N_5641,N_632,N_3693);
nor U5642 (N_5642,N_4640,N_3627);
or U5643 (N_5643,N_1463,N_1949);
or U5644 (N_5644,N_1939,N_887);
and U5645 (N_5645,N_3271,N_4828);
or U5646 (N_5646,N_829,N_352);
nor U5647 (N_5647,N_3604,N_405);
nor U5648 (N_5648,N_3133,N_1884);
xor U5649 (N_5649,N_3108,N_1339);
and U5650 (N_5650,N_2854,N_4299);
and U5651 (N_5651,N_3954,N_1270);
nand U5652 (N_5652,N_869,N_3542);
or U5653 (N_5653,N_947,N_4837);
nor U5654 (N_5654,N_4869,N_1490);
or U5655 (N_5655,N_1743,N_623);
nand U5656 (N_5656,N_3032,N_227);
nand U5657 (N_5657,N_3752,N_4610);
nand U5658 (N_5658,N_1948,N_4024);
xnor U5659 (N_5659,N_3754,N_857);
and U5660 (N_5660,N_2208,N_2004);
nand U5661 (N_5661,N_4412,N_3249);
or U5662 (N_5662,N_851,N_4623);
or U5663 (N_5663,N_2706,N_2953);
nor U5664 (N_5664,N_2479,N_590);
and U5665 (N_5665,N_2699,N_47);
and U5666 (N_5666,N_2408,N_710);
or U5667 (N_5667,N_1366,N_4443);
or U5668 (N_5668,N_4982,N_307);
nor U5669 (N_5669,N_4871,N_1973);
nor U5670 (N_5670,N_2777,N_2510);
and U5671 (N_5671,N_4946,N_1596);
and U5672 (N_5672,N_4470,N_2297);
or U5673 (N_5673,N_1065,N_2341);
or U5674 (N_5674,N_1735,N_898);
and U5675 (N_5675,N_2495,N_579);
nand U5676 (N_5676,N_3146,N_944);
nor U5677 (N_5677,N_3694,N_2938);
nor U5678 (N_5678,N_4231,N_2162);
nor U5679 (N_5679,N_2266,N_940);
nand U5680 (N_5680,N_1560,N_3316);
and U5681 (N_5681,N_1267,N_673);
xnor U5682 (N_5682,N_3862,N_4720);
nand U5683 (N_5683,N_856,N_4520);
nand U5684 (N_5684,N_2082,N_2520);
or U5685 (N_5685,N_3900,N_2771);
xor U5686 (N_5686,N_3762,N_1290);
and U5687 (N_5687,N_3801,N_1341);
nand U5688 (N_5688,N_1019,N_4659);
xor U5689 (N_5689,N_1041,N_2832);
nor U5690 (N_5690,N_2511,N_4405);
xnor U5691 (N_5691,N_4618,N_4093);
or U5692 (N_5692,N_2316,N_2282);
nor U5693 (N_5693,N_1865,N_2943);
and U5694 (N_5694,N_746,N_4537);
nand U5695 (N_5695,N_82,N_350);
and U5696 (N_5696,N_3288,N_1404);
or U5697 (N_5697,N_81,N_4297);
or U5698 (N_5698,N_1786,N_3870);
xnor U5699 (N_5699,N_2138,N_1661);
nor U5700 (N_5700,N_4445,N_715);
and U5701 (N_5701,N_3846,N_3797);
or U5702 (N_5702,N_4897,N_1968);
nor U5703 (N_5703,N_2611,N_1066);
and U5704 (N_5704,N_1144,N_3705);
nor U5705 (N_5705,N_114,N_3473);
nor U5706 (N_5706,N_3756,N_4461);
nor U5707 (N_5707,N_2165,N_2565);
xnor U5708 (N_5708,N_1071,N_4305);
nor U5709 (N_5709,N_3011,N_1789);
nor U5710 (N_5710,N_1550,N_1520);
or U5711 (N_5711,N_1629,N_1326);
nor U5712 (N_5712,N_3262,N_758);
xor U5713 (N_5713,N_747,N_2656);
nand U5714 (N_5714,N_4688,N_2547);
nand U5715 (N_5715,N_1958,N_2574);
and U5716 (N_5716,N_1253,N_714);
nand U5717 (N_5717,N_3242,N_2011);
nand U5718 (N_5718,N_763,N_1910);
and U5719 (N_5719,N_4175,N_1659);
nor U5720 (N_5720,N_2195,N_1444);
nor U5721 (N_5721,N_768,N_3259);
xor U5722 (N_5722,N_4938,N_655);
and U5723 (N_5723,N_4761,N_3529);
xnor U5724 (N_5724,N_3856,N_860);
and U5725 (N_5725,N_1381,N_1565);
or U5726 (N_5726,N_2691,N_2760);
and U5727 (N_5727,N_4671,N_1485);
or U5728 (N_5728,N_6,N_3776);
nand U5729 (N_5729,N_937,N_3205);
and U5730 (N_5730,N_4450,N_1926);
nand U5731 (N_5731,N_2415,N_730);
nor U5732 (N_5732,N_1242,N_1511);
nor U5733 (N_5733,N_620,N_4522);
xnor U5734 (N_5734,N_3231,N_3787);
and U5735 (N_5735,N_4003,N_1498);
or U5736 (N_5736,N_635,N_1817);
and U5737 (N_5737,N_152,N_3621);
and U5738 (N_5738,N_1847,N_2686);
or U5739 (N_5739,N_4877,N_1592);
and U5740 (N_5740,N_3403,N_1297);
nor U5741 (N_5741,N_2919,N_1068);
or U5742 (N_5742,N_3923,N_3779);
and U5743 (N_5743,N_149,N_1482);
and U5744 (N_5744,N_161,N_3110);
nor U5745 (N_5745,N_3330,N_4217);
nor U5746 (N_5746,N_1698,N_3730);
and U5747 (N_5747,N_131,N_1649);
or U5748 (N_5748,N_2411,N_93);
nor U5749 (N_5749,N_3111,N_3199);
and U5750 (N_5750,N_2785,N_2872);
nand U5751 (N_5751,N_2831,N_3726);
or U5752 (N_5752,N_3328,N_833);
nor U5753 (N_5753,N_4562,N_1447);
or U5754 (N_5754,N_3593,N_3312);
and U5755 (N_5755,N_4,N_4802);
nand U5756 (N_5756,N_343,N_106);
nor U5757 (N_5757,N_2555,N_4864);
nor U5758 (N_5758,N_2326,N_2249);
nor U5759 (N_5759,N_2039,N_314);
nand U5760 (N_5760,N_3492,N_3034);
or U5761 (N_5761,N_4341,N_2449);
nand U5762 (N_5762,N_413,N_1501);
nand U5763 (N_5763,N_311,N_26);
and U5764 (N_5764,N_3824,N_2111);
nor U5765 (N_5765,N_2564,N_1491);
or U5766 (N_5766,N_2767,N_2235);
or U5767 (N_5767,N_2241,N_4180);
nor U5768 (N_5768,N_1342,N_4668);
xor U5769 (N_5769,N_3886,N_1158);
nor U5770 (N_5770,N_4159,N_899);
or U5771 (N_5771,N_683,N_4127);
and U5772 (N_5772,N_2230,N_1922);
nor U5773 (N_5773,N_1351,N_957);
nand U5774 (N_5774,N_485,N_3871);
nand U5775 (N_5775,N_4312,N_4818);
or U5776 (N_5776,N_4513,N_1256);
or U5777 (N_5777,N_1720,N_1972);
and U5778 (N_5778,N_3373,N_3892);
and U5779 (N_5779,N_346,N_4715);
or U5780 (N_5780,N_1519,N_2845);
xor U5781 (N_5781,N_1759,N_3171);
xnor U5782 (N_5782,N_4632,N_1570);
nor U5783 (N_5783,N_1203,N_4694);
nand U5784 (N_5784,N_2371,N_1696);
nand U5785 (N_5785,N_4547,N_4281);
nand U5786 (N_5786,N_3901,N_2689);
nand U5787 (N_5787,N_800,N_4247);
nand U5788 (N_5788,N_2164,N_2828);
and U5789 (N_5789,N_2276,N_371);
nand U5790 (N_5790,N_592,N_3470);
or U5791 (N_5791,N_4201,N_1243);
or U5792 (N_5792,N_1552,N_549);
xnor U5793 (N_5793,N_2416,N_4579);
or U5794 (N_5794,N_3503,N_1989);
nor U5795 (N_5795,N_1504,N_2223);
nand U5796 (N_5796,N_1960,N_4949);
nand U5797 (N_5797,N_3161,N_3021);
or U5798 (N_5798,N_3157,N_2898);
and U5799 (N_5799,N_1169,N_4757);
nand U5800 (N_5800,N_3291,N_117);
nor U5801 (N_5801,N_600,N_3792);
xor U5802 (N_5802,N_1004,N_1680);
nand U5803 (N_5803,N_559,N_1643);
nor U5804 (N_5804,N_2330,N_4107);
nor U5805 (N_5805,N_2967,N_2019);
nand U5806 (N_5806,N_3585,N_274);
nor U5807 (N_5807,N_748,N_1832);
nor U5808 (N_5808,N_3655,N_2211);
or U5809 (N_5809,N_4960,N_1717);
nand U5810 (N_5810,N_4032,N_1357);
nand U5811 (N_5811,N_3671,N_4272);
and U5812 (N_5812,N_512,N_3908);
or U5813 (N_5813,N_3983,N_309);
nand U5814 (N_5814,N_3151,N_2583);
and U5815 (N_5815,N_4216,N_2683);
and U5816 (N_5816,N_1863,N_2106);
and U5817 (N_5817,N_3664,N_3315);
or U5818 (N_5818,N_4186,N_282);
xor U5819 (N_5819,N_4256,N_2321);
and U5820 (N_5820,N_2585,N_741);
nand U5821 (N_5821,N_3102,N_1859);
xnor U5822 (N_5822,N_2216,N_219);
nand U5823 (N_5823,N_3515,N_59);
and U5824 (N_5824,N_337,N_2030);
nand U5825 (N_5825,N_1211,N_433);
and U5826 (N_5826,N_4639,N_1535);
and U5827 (N_5827,N_4727,N_3718);
xor U5828 (N_5828,N_2163,N_222);
or U5829 (N_5829,N_1732,N_488);
and U5830 (N_5830,N_3821,N_826);
and U5831 (N_5831,N_3331,N_3261);
nand U5832 (N_5832,N_3748,N_1848);
xor U5833 (N_5833,N_2783,N_2957);
nor U5834 (N_5834,N_3639,N_2350);
nor U5835 (N_5835,N_2028,N_953);
nand U5836 (N_5836,N_3922,N_3446);
and U5837 (N_5837,N_4483,N_2576);
or U5838 (N_5838,N_1474,N_3681);
nand U5839 (N_5839,N_203,N_1955);
nand U5840 (N_5840,N_46,N_2284);
nand U5841 (N_5841,N_425,N_1338);
and U5842 (N_5842,N_218,N_399);
nor U5843 (N_5843,N_21,N_3372);
xnor U5844 (N_5844,N_179,N_3526);
nor U5845 (N_5845,N_2975,N_84);
nand U5846 (N_5846,N_3318,N_4111);
or U5847 (N_5847,N_3398,N_3266);
xnor U5848 (N_5848,N_1221,N_4593);
nand U5849 (N_5849,N_4057,N_1756);
xnor U5850 (N_5850,N_2097,N_4383);
and U5851 (N_5851,N_4208,N_4627);
or U5852 (N_5852,N_2340,N_3698);
and U5853 (N_5853,N_3030,N_3121);
and U5854 (N_5854,N_3482,N_2745);
and U5855 (N_5855,N_4544,N_4947);
and U5856 (N_5856,N_2963,N_157);
nor U5857 (N_5857,N_972,N_3414);
and U5858 (N_5858,N_2296,N_310);
and U5859 (N_5859,N_380,N_2203);
and U5860 (N_5860,N_1031,N_1137);
nand U5861 (N_5861,N_3969,N_9);
and U5862 (N_5862,N_955,N_2887);
and U5863 (N_5863,N_2894,N_4319);
nor U5864 (N_5864,N_3393,N_2784);
nor U5865 (N_5865,N_1648,N_4192);
nand U5866 (N_5866,N_3091,N_1840);
and U5867 (N_5867,N_3743,N_2466);
nor U5868 (N_5868,N_3277,N_526);
and U5869 (N_5869,N_1924,N_2727);
nor U5870 (N_5870,N_3570,N_4747);
xor U5871 (N_5871,N_1431,N_834);
and U5872 (N_5872,N_921,N_751);
nor U5873 (N_5873,N_2369,N_912);
and U5874 (N_5874,N_3631,N_1834);
nand U5875 (N_5875,N_4577,N_4361);
or U5876 (N_5876,N_130,N_523);
xnor U5877 (N_5877,N_2605,N_1413);
nand U5878 (N_5878,N_4997,N_1304);
nor U5879 (N_5879,N_3374,N_385);
xor U5880 (N_5880,N_3018,N_4974);
nor U5881 (N_5881,N_3123,N_3951);
nor U5882 (N_5882,N_4420,N_1218);
nor U5883 (N_5883,N_2158,N_1350);
and U5884 (N_5884,N_4719,N_169);
and U5885 (N_5885,N_732,N_4708);
nor U5886 (N_5886,N_3428,N_1965);
nor U5887 (N_5887,N_4776,N_891);
and U5888 (N_5888,N_2597,N_210);
and U5889 (N_5889,N_4164,N_3714);
or U5890 (N_5890,N_2590,N_2606);
and U5891 (N_5891,N_2609,N_3717);
nor U5892 (N_5892,N_4271,N_4336);
or U5893 (N_5893,N_1111,N_2795);
or U5894 (N_5894,N_2349,N_821);
xor U5895 (N_5895,N_4937,N_1323);
and U5896 (N_5896,N_2458,N_4634);
nand U5897 (N_5897,N_4585,N_4616);
nand U5898 (N_5898,N_4162,N_3056);
nor U5899 (N_5899,N_2643,N_3687);
and U5900 (N_5900,N_1891,N_3053);
or U5901 (N_5901,N_3539,N_1465);
nor U5902 (N_5902,N_1208,N_266);
xor U5903 (N_5903,N_1776,N_1654);
nand U5904 (N_5904,N_4752,N_2644);
and U5905 (N_5905,N_4850,N_1624);
or U5906 (N_5906,N_1536,N_575);
or U5907 (N_5907,N_2151,N_723);
nand U5908 (N_5908,N_4771,N_3578);
xor U5909 (N_5909,N_3313,N_2124);
and U5910 (N_5910,N_883,N_4633);
nand U5911 (N_5911,N_2561,N_4910);
or U5912 (N_5912,N_725,N_4862);
nor U5913 (N_5913,N_1823,N_698);
and U5914 (N_5914,N_1384,N_2036);
nor U5915 (N_5915,N_2578,N_3050);
nand U5916 (N_5916,N_4991,N_4259);
nor U5917 (N_5917,N_2492,N_4512);
nor U5918 (N_5918,N_576,N_890);
or U5919 (N_5919,N_486,N_259);
or U5920 (N_5920,N_2392,N_550);
nor U5921 (N_5921,N_3062,N_3178);
and U5922 (N_5922,N_2293,N_4417);
nand U5923 (N_5923,N_3737,N_1849);
xnor U5924 (N_5924,N_1630,N_2189);
or U5925 (N_5925,N_3642,N_3149);
or U5926 (N_5926,N_1963,N_4276);
nand U5927 (N_5927,N_4390,N_4981);
and U5928 (N_5928,N_1246,N_1174);
nor U5929 (N_5929,N_3294,N_1322);
and U5930 (N_5930,N_1614,N_2412);
and U5931 (N_5931,N_769,N_23);
and U5932 (N_5932,N_2869,N_3075);
nand U5933 (N_5933,N_294,N_3257);
nor U5934 (N_5934,N_363,N_3214);
and U5935 (N_5935,N_1981,N_3980);
xnor U5936 (N_5936,N_436,N_4508);
nand U5937 (N_5937,N_4499,N_359);
and U5938 (N_5938,N_3618,N_2980);
nor U5939 (N_5939,N_1517,N_4302);
nor U5940 (N_5940,N_1556,N_3638);
or U5941 (N_5941,N_1512,N_3101);
and U5942 (N_5942,N_1744,N_4418);
and U5943 (N_5943,N_1892,N_3131);
and U5944 (N_5944,N_2220,N_1217);
or U5945 (N_5945,N_4258,N_786);
nand U5946 (N_5946,N_465,N_367);
nor U5947 (N_5947,N_3410,N_2738);
nor U5948 (N_5948,N_1027,N_1638);
or U5949 (N_5949,N_3420,N_3065);
xor U5950 (N_5950,N_3324,N_1107);
nor U5951 (N_5951,N_924,N_1618);
or U5952 (N_5952,N_2695,N_2518);
xnor U5953 (N_5953,N_3468,N_2531);
and U5954 (N_5954,N_2456,N_3289);
nor U5955 (N_5955,N_57,N_4242);
or U5956 (N_5956,N_2078,N_3290);
nor U5957 (N_5957,N_2530,N_2192);
nand U5958 (N_5958,N_2661,N_675);
and U5959 (N_5959,N_328,N_4080);
or U5960 (N_5960,N_915,N_3988);
and U5961 (N_5961,N_158,N_4795);
or U5962 (N_5962,N_952,N_3566);
xor U5963 (N_5963,N_1598,N_2793);
nor U5964 (N_5964,N_2467,N_649);
or U5965 (N_5965,N_122,N_1935);
or U5966 (N_5966,N_802,N_1992);
xor U5967 (N_5967,N_8,N_1684);
nand U5968 (N_5968,N_587,N_1514);
nand U5969 (N_5969,N_2051,N_916);
or U5970 (N_5970,N_2782,N_4511);
nand U5971 (N_5971,N_4888,N_3864);
nor U5972 (N_5972,N_4112,N_98);
xnor U5973 (N_5973,N_884,N_2508);
nand U5974 (N_5974,N_4465,N_2826);
nand U5975 (N_5975,N_3148,N_4222);
nor U5976 (N_5976,N_1518,N_4534);
nor U5977 (N_5977,N_1418,N_1044);
xnor U5978 (N_5978,N_4167,N_142);
and U5979 (N_5979,N_4314,N_4777);
xnor U5980 (N_5980,N_2514,N_2537);
nand U5981 (N_5981,N_3565,N_1875);
or U5982 (N_5982,N_3190,N_4379);
nor U5983 (N_5983,N_2023,N_3086);
and U5984 (N_5984,N_3544,N_377);
nor U5985 (N_5985,N_2338,N_1313);
or U5986 (N_5986,N_2988,N_3673);
nand U5987 (N_5987,N_426,N_2113);
nor U5988 (N_5988,N_1602,N_824);
xor U5989 (N_5989,N_495,N_1039);
nor U5990 (N_5990,N_4797,N_3605);
and U5991 (N_5991,N_2318,N_4724);
nor U5992 (N_5992,N_1477,N_450);
nor U5993 (N_5993,N_2365,N_1113);
or U5994 (N_5994,N_101,N_3491);
and U5995 (N_5995,N_378,N_1254);
nand U5996 (N_5996,N_1183,N_4356);
or U5997 (N_5997,N_816,N_3580);
xor U5998 (N_5998,N_3476,N_1930);
or U5999 (N_5999,N_2962,N_3505);
nor U6000 (N_6000,N_1425,N_118);
and U6001 (N_6001,N_2344,N_2261);
or U6002 (N_6002,N_2575,N_4230);
and U6003 (N_6003,N_1645,N_1768);
or U6004 (N_6004,N_3345,N_4868);
or U6005 (N_6005,N_3502,N_1061);
nand U6006 (N_6006,N_837,N_215);
and U6007 (N_6007,N_2109,N_3022);
and U6008 (N_6008,N_1492,N_3203);
nand U6009 (N_6009,N_1663,N_1123);
nand U6010 (N_6010,N_3959,N_49);
and U6011 (N_6011,N_3284,N_1531);
xnor U6012 (N_6012,N_2987,N_3960);
nor U6013 (N_6013,N_1937,N_3607);
and U6014 (N_6014,N_4324,N_4699);
nand U6015 (N_6015,N_1285,N_3506);
and U6016 (N_6016,N_3569,N_3496);
and U6017 (N_6017,N_757,N_1356);
or U6018 (N_6018,N_4424,N_4899);
nor U6019 (N_6019,N_4713,N_3879);
or U6020 (N_6020,N_4594,N_2982);
nand U6021 (N_6021,N_351,N_3130);
nor U6022 (N_6022,N_3990,N_1982);
and U6023 (N_6023,N_1647,N_628);
or U6024 (N_6024,N_3695,N_712);
nor U6025 (N_6025,N_3645,N_2161);
nor U6026 (N_6026,N_2417,N_1986);
nand U6027 (N_6027,N_4433,N_2401);
nor U6028 (N_6028,N_2969,N_971);
and U6029 (N_6029,N_1021,N_994);
nand U6030 (N_6030,N_1255,N_177);
nor U6031 (N_6031,N_2794,N_183);
or U6032 (N_6032,N_4778,N_2568);
nor U6033 (N_6033,N_2867,N_4745);
xor U6034 (N_6034,N_225,N_3747);
or U6035 (N_6035,N_4456,N_2055);
nor U6036 (N_6036,N_697,N_1263);
and U6037 (N_6037,N_4586,N_4929);
nor U6038 (N_6038,N_1542,N_3941);
nor U6039 (N_6039,N_2769,N_459);
nor U6040 (N_6040,N_4637,N_4125);
xor U6041 (N_6041,N_701,N_510);
or U6042 (N_6042,N_1733,N_706);
xnor U6043 (N_6043,N_2294,N_4188);
xor U6044 (N_6044,N_594,N_3568);
nor U6045 (N_6045,N_2930,N_3370);
nand U6046 (N_6046,N_1280,N_889);
and U6047 (N_6047,N_652,N_2463);
and U6048 (N_6048,N_1943,N_3929);
nor U6049 (N_6049,N_1488,N_2506);
nand U6050 (N_6050,N_1262,N_4481);
nor U6051 (N_6051,N_1521,N_4163);
nor U6052 (N_6052,N_407,N_341);
or U6053 (N_6053,N_3986,N_4142);
and U6054 (N_6054,N_1665,N_3699);
nor U6055 (N_6055,N_289,N_604);
nand U6056 (N_6056,N_2724,N_2675);
xnor U6057 (N_6057,N_2419,N_1526);
nor U6058 (N_6058,N_2270,N_3691);
and U6059 (N_6059,N_3682,N_484);
nand U6060 (N_6060,N_3245,N_3464);
and U6061 (N_6061,N_3097,N_973);
nand U6062 (N_6062,N_1705,N_2314);
or U6063 (N_6063,N_292,N_2035);
nand U6064 (N_6064,N_4992,N_1831);
and U6065 (N_6065,N_4085,N_2685);
nor U6066 (N_6066,N_3653,N_2926);
or U6067 (N_6067,N_4490,N_1010);
and U6068 (N_6068,N_3254,N_3223);
nor U6069 (N_6069,N_4145,N_1176);
nor U6070 (N_6070,N_4606,N_2736);
nand U6071 (N_6071,N_4687,N_422);
or U6072 (N_6072,N_1128,N_2105);
or U6073 (N_6073,N_112,N_1161);
nand U6074 (N_6074,N_4150,N_4078);
and U6075 (N_6075,N_3581,N_4901);
nor U6076 (N_6076,N_3339,N_4011);
nor U6077 (N_6077,N_2979,N_2942);
xnor U6078 (N_6078,N_720,N_89);
and U6079 (N_6079,N_2608,N_462);
and U6080 (N_6080,N_932,N_2236);
nand U6081 (N_6081,N_3296,N_1774);
and U6082 (N_6082,N_3395,N_3041);
nor U6083 (N_6083,N_2099,N_2700);
nand U6084 (N_6084,N_1222,N_3453);
nand U6085 (N_6085,N_1070,N_43);
and U6086 (N_6086,N_195,N_464);
and U6087 (N_6087,N_1616,N_3891);
nand U6088 (N_6088,N_665,N_3702);
xor U6089 (N_6089,N_1471,N_1564);
nand U6090 (N_6090,N_2787,N_3287);
and U6091 (N_6091,N_3009,N_2421);
and U6092 (N_6092,N_1583,N_3276);
nor U6093 (N_6093,N_4717,N_1749);
nand U6094 (N_6094,N_2021,N_3735);
nor U6095 (N_6095,N_2498,N_766);
xor U6096 (N_6096,N_530,N_3813);
nor U6097 (N_6097,N_3213,N_2231);
and U6098 (N_6098,N_3613,N_1084);
or U6099 (N_6099,N_1700,N_2405);
nor U6100 (N_6100,N_4983,N_761);
nor U6101 (N_6101,N_2460,N_1971);
nor U6102 (N_6102,N_2384,N_1830);
nand U6103 (N_6103,N_2999,N_685);
nand U6104 (N_6104,N_3808,N_2300);
and U6105 (N_6105,N_4557,N_1387);
and U6106 (N_6106,N_2262,N_442);
nand U6107 (N_6107,N_2772,N_4509);
and U6108 (N_6108,N_3083,N_4498);
nand U6109 (N_6109,N_2601,N_3169);
nand U6110 (N_6110,N_2535,N_3122);
or U6111 (N_6111,N_53,N_4507);
and U6112 (N_6112,N_4010,N_4440);
and U6113 (N_6113,N_629,N_2836);
or U6114 (N_6114,N_2803,N_1881);
nand U6115 (N_6115,N_1909,N_1895);
and U6116 (N_6116,N_3591,N_564);
nor U6117 (N_6117,N_2660,N_4962);
or U6118 (N_6118,N_4603,N_676);
and U6119 (N_6119,N_1670,N_2351);
nor U6120 (N_6120,N_3866,N_1582);
and U6121 (N_6121,N_603,N_4630);
xor U6122 (N_6122,N_1252,N_4288);
or U6123 (N_6123,N_2207,N_108);
xnor U6124 (N_6124,N_383,N_918);
nor U6125 (N_6125,N_1742,N_1826);
or U6126 (N_6126,N_4514,N_819);
or U6127 (N_6127,N_3176,N_3703);
nor U6128 (N_6128,N_1114,N_4961);
and U6129 (N_6129,N_1568,N_756);
nand U6130 (N_6130,N_805,N_374);
nor U6131 (N_6131,N_3255,N_364);
nor U6132 (N_6132,N_4185,N_1918);
nor U6133 (N_6133,N_4914,N_1777);
and U6134 (N_6134,N_1094,N_3770);
xor U6135 (N_6135,N_900,N_3739);
or U6136 (N_6136,N_1170,N_3803);
nor U6137 (N_6137,N_2320,N_263);
and U6138 (N_6138,N_2181,N_107);
nand U6139 (N_6139,N_4493,N_4172);
and U6140 (N_6140,N_3830,N_4220);
nand U6141 (N_6141,N_2332,N_4376);
nor U6142 (N_6142,N_504,N_4091);
or U6143 (N_6143,N_4187,N_3471);
nor U6144 (N_6144,N_3415,N_687);
nand U6145 (N_6145,N_316,N_4146);
nand U6146 (N_6146,N_509,N_607);
nand U6147 (N_6147,N_31,N_3834);
and U6148 (N_6148,N_713,N_4844);
or U6149 (N_6149,N_1500,N_1464);
xor U6150 (N_6150,N_396,N_2830);
nand U6151 (N_6151,N_3449,N_3124);
nand U6152 (N_6152,N_4168,N_1854);
nand U6153 (N_6153,N_516,N_2335);
and U6154 (N_6154,N_4430,N_16);
or U6155 (N_6155,N_4004,N_3426);
nor U6156 (N_6156,N_3895,N_2588);
nor U6157 (N_6157,N_4181,N_2364);
nor U6158 (N_6158,N_1626,N_2345);
nor U6159 (N_6159,N_4474,N_3351);
xor U6160 (N_6160,N_3113,N_4215);
nand U6161 (N_6161,N_3068,N_217);
nand U6162 (N_6162,N_4293,N_657);
or U6163 (N_6163,N_2147,N_3868);
and U6164 (N_6164,N_557,N_4387);
and U6165 (N_6165,N_2707,N_527);
nand U6166 (N_6166,N_1112,N_4267);
and U6167 (N_6167,N_722,N_572);
and U6168 (N_6168,N_3282,N_702);
xnor U6169 (N_6169,N_1688,N_141);
nor U6170 (N_6170,N_3489,N_3723);
or U6171 (N_6171,N_4758,N_3873);
or U6172 (N_6172,N_3049,N_3184);
nand U6173 (N_6173,N_2313,N_2543);
nor U6174 (N_6174,N_4211,N_2503);
nor U6175 (N_6175,N_1721,N_951);
nand U6176 (N_6176,N_1984,N_4571);
xor U6177 (N_6177,N_1824,N_4310);
and U6178 (N_6178,N_2579,N_4069);
nand U6179 (N_6179,N_1769,N_4468);
and U6180 (N_6180,N_4087,N_482);
and U6181 (N_6181,N_2960,N_2317);
or U6182 (N_6182,N_4859,N_4355);
nor U6183 (N_6183,N_375,N_1673);
and U6184 (N_6184,N_1686,N_684);
nand U6185 (N_6185,N_2866,N_3925);
nor U6186 (N_6186,N_4316,N_1186);
nor U6187 (N_6187,N_3722,N_3890);
nor U6188 (N_6188,N_1827,N_830);
nor U6189 (N_6189,N_2781,N_4703);
nand U6190 (N_6190,N_4179,N_1724);
or U6191 (N_6191,N_871,N_1479);
and U6192 (N_6192,N_3301,N_492);
nor U6193 (N_6193,N_4317,N_331);
nand U6194 (N_6194,N_4810,N_3601);
xnor U6195 (N_6195,N_551,N_533);
and U6196 (N_6196,N_3995,N_3382);
nor U6197 (N_6197,N_174,N_4738);
and U6198 (N_6198,N_3109,N_2311);
and U6199 (N_6199,N_2352,N_1380);
nand U6200 (N_6200,N_2742,N_3480);
and U6201 (N_6201,N_3574,N_2734);
or U6202 (N_6202,N_3716,N_1064);
nor U6203 (N_6203,N_4364,N_1604);
nor U6204 (N_6204,N_2167,N_4273);
or U6205 (N_6205,N_3731,N_2169);
nor U6206 (N_6206,N_4835,N_2016);
or U6207 (N_6207,N_4624,N_858);
nand U6208 (N_6208,N_981,N_4178);
and U6209 (N_6209,N_3596,N_927);
xor U6210 (N_6210,N_4989,N_670);
nor U6211 (N_6211,N_497,N_4351);
nor U6212 (N_6212,N_2857,N_2509);
nor U6213 (N_6213,N_4990,N_1682);
xor U6214 (N_6214,N_4588,N_4985);
or U6215 (N_6215,N_2218,N_4113);
and U6216 (N_6216,N_129,N_1846);
or U6217 (N_6217,N_2748,N_3795);
xnor U6218 (N_6218,N_2809,N_2446);
and U6219 (N_6219,N_2934,N_2041);
nor U6220 (N_6220,N_1495,N_2054);
or U6221 (N_6221,N_1229,N_3343);
or U6222 (N_6222,N_2336,N_3012);
or U6223 (N_6223,N_1586,N_4197);
and U6224 (N_6224,N_4656,N_4282);
or U6225 (N_6225,N_875,N_336);
and U6226 (N_6226,N_271,N_262);
nor U6227 (N_6227,N_1899,N_4951);
nand U6228 (N_6228,N_4114,N_3381);
nand U6229 (N_6229,N_1936,N_1800);
or U6230 (N_6230,N_2037,N_4343);
nand U6231 (N_6231,N_3540,N_4964);
or U6232 (N_6232,N_3628,N_3648);
nand U6233 (N_6233,N_4130,N_1580);
nor U6234 (N_6234,N_4038,N_2694);
nor U6235 (N_6235,N_4772,N_258);
nand U6236 (N_6236,N_3533,N_3926);
nand U6237 (N_6237,N_2368,N_3407);
and U6238 (N_6238,N_842,N_737);
and U6239 (N_6239,N_729,N_4836);
or U6240 (N_6240,N_4701,N_2199);
nand U6241 (N_6241,N_400,N_3310);
or U6242 (N_6242,N_11,N_2304);
and U6243 (N_6243,N_2945,N_647);
and U6244 (N_6244,N_392,N_3427);
and U6245 (N_6245,N_2157,N_3883);
xor U6246 (N_6246,N_1637,N_2917);
or U6247 (N_6247,N_1213,N_799);
and U6248 (N_6248,N_3386,N_4110);
and U6249 (N_6249,N_3379,N_4183);
nor U6250 (N_6250,N_230,N_3728);
nand U6251 (N_6251,N_4224,N_4262);
nand U6252 (N_6252,N_3600,N_4309);
nand U6253 (N_6253,N_4980,N_4900);
or U6254 (N_6254,N_4545,N_4458);
or U6255 (N_6255,N_1764,N_4015);
nor U6256 (N_6256,N_524,N_3952);
xor U6257 (N_6257,N_4867,N_4805);
and U6258 (N_6258,N_2403,N_2380);
or U6259 (N_6259,N_1723,N_4592);
and U6260 (N_6260,N_1767,N_4131);
nor U6261 (N_6261,N_1199,N_1007);
or U6262 (N_6262,N_2061,N_1506);
nor U6263 (N_6263,N_3521,N_3946);
and U6264 (N_6264,N_4488,N_2049);
nand U6265 (N_6265,N_3553,N_1946);
and U6266 (N_6266,N_4428,N_4824);
and U6267 (N_6267,N_1083,N_4046);
nor U6268 (N_6268,N_1632,N_236);
nand U6269 (N_6269,N_3162,N_1419);
and U6270 (N_6270,N_609,N_1706);
nand U6271 (N_6271,N_2396,N_2126);
and U6272 (N_6272,N_376,N_3060);
or U6273 (N_6273,N_2363,N_536);
nor U6274 (N_6274,N_2060,N_1228);
or U6275 (N_6275,N_3668,N_224);
xnor U6276 (N_6276,N_1153,N_895);
or U6277 (N_6277,N_2185,N_1979);
and U6278 (N_6278,N_2517,N_2389);
or U6279 (N_6279,N_3019,N_1455);
nor U6280 (N_6280,N_3633,N_3742);
or U6281 (N_6281,N_4873,N_1308);
xor U6282 (N_6282,N_1054,N_4294);
nor U6283 (N_6283,N_176,N_3822);
nand U6284 (N_6284,N_4190,N_1017);
nor U6285 (N_6285,N_2257,N_865);
and U6286 (N_6286,N_651,N_3842);
or U6287 (N_6287,N_2839,N_3377);
nor U6288 (N_6288,N_4135,N_2746);
or U6289 (N_6289,N_4684,N_4814);
nor U6290 (N_6290,N_4550,N_654);
and U6291 (N_6291,N_3966,N_4275);
and U6292 (N_6292,N_4306,N_4711);
and U6293 (N_6293,N_2132,N_2814);
nand U6294 (N_6294,N_1090,N_1940);
nand U6295 (N_6295,N_3005,N_1091);
or U6296 (N_6296,N_4799,N_3835);
nand U6297 (N_6297,N_2704,N_2679);
or U6298 (N_6298,N_2234,N_4548);
and U6299 (N_6299,N_4237,N_1754);
and U6300 (N_6300,N_4709,N_3836);
nand U6301 (N_6301,N_4963,N_545);
nand U6302 (N_6302,N_2058,N_4567);
or U6303 (N_6303,N_2554,N_4278);
and U6304 (N_6304,N_1273,N_4931);
xor U6305 (N_6305,N_1641,N_1078);
nor U6306 (N_6306,N_391,N_4373);
or U6307 (N_6307,N_1781,N_4812);
nand U6308 (N_6308,N_4202,N_1571);
or U6309 (N_6309,N_1257,N_3740);
and U6310 (N_6310,N_4248,N_306);
nand U6311 (N_6311,N_3538,N_296);
nand U6312 (N_6312,N_2299,N_3635);
or U6313 (N_6313,N_3771,N_681);
nand U6314 (N_6314,N_2664,N_2477);
and U6315 (N_6315,N_3524,N_528);
or U6316 (N_6316,N_2878,N_3799);
and U6317 (N_6317,N_305,N_4679);
xnor U6318 (N_6318,N_1152,N_3098);
and U6319 (N_6319,N_3516,N_555);
or U6320 (N_6320,N_2393,N_4067);
nand U6321 (N_6321,N_3972,N_1178);
or U6322 (N_6322,N_1887,N_2672);
or U6323 (N_6323,N_3562,N_2475);
and U6324 (N_6324,N_3147,N_4421);
or U6325 (N_6325,N_4199,N_1296);
nor U6326 (N_6326,N_2655,N_163);
nand U6327 (N_6327,N_541,N_281);
and U6328 (N_6328,N_260,N_192);
and U6329 (N_6329,N_1923,N_3661);
and U6330 (N_6330,N_4636,N_2774);
nand U6331 (N_6331,N_3488,N_1452);
nand U6332 (N_6332,N_3975,N_3647);
nor U6333 (N_6333,N_2815,N_2156);
xnor U6334 (N_6334,N_4177,N_2870);
nand U6335 (N_6335,N_4037,N_1539);
and U6336 (N_6336,N_1543,N_151);
xor U6337 (N_6337,N_1739,N_4626);
and U6338 (N_6338,N_2166,N_1898);
and U6339 (N_6339,N_327,N_3789);
xor U6340 (N_6340,N_3355,N_3564);
nand U6341 (N_6341,N_2098,N_3070);
and U6342 (N_6342,N_3783,N_3297);
nand U6343 (N_6343,N_4414,N_621);
and U6344 (N_6344,N_988,N_2627);
nor U6345 (N_6345,N_645,N_4518);
or U6346 (N_6346,N_4770,N_4315);
nor U6347 (N_6347,N_534,N_3046);
and U6348 (N_6348,N_1325,N_3915);
or U6349 (N_6349,N_1722,N_90);
or U6350 (N_6350,N_738,N_4395);
nor U6351 (N_6351,N_4485,N_2329);
nor U6352 (N_6352,N_2776,N_4264);
nand U6353 (N_6353,N_312,N_2295);
xnor U6354 (N_6354,N_2743,N_1822);
nand U6355 (N_6355,N_4494,N_982);
and U6356 (N_6356,N_949,N_3154);
nand U6357 (N_6357,N_2723,N_1483);
nand U6358 (N_6358,N_251,N_2180);
and U6359 (N_6359,N_962,N_1142);
and U6360 (N_6360,N_731,N_2949);
nand U6361 (N_6361,N_2063,N_4825);
or U6362 (N_6362,N_1397,N_525);
and U6363 (N_6363,N_1067,N_2409);
xnor U6364 (N_6364,N_2681,N_4287);
xor U6365 (N_6365,N_1035,N_1359);
or U6366 (N_6366,N_506,N_1883);
nand U6367 (N_6367,N_214,N_2763);
and U6368 (N_6368,N_1370,N_1165);
or U6369 (N_6369,N_4733,N_945);
or U6370 (N_6370,N_4928,N_1947);
and U6371 (N_6371,N_3079,N_4660);
and U6372 (N_6372,N_3486,N_1997);
nand U6373 (N_6373,N_2005,N_2485);
and U6374 (N_6374,N_4909,N_2017);
or U6375 (N_6375,N_4599,N_529);
nand U6376 (N_6376,N_1192,N_4605);
or U6377 (N_6377,N_133,N_2122);
nand U6378 (N_6378,N_171,N_1704);
nand U6379 (N_6379,N_3599,N_1502);
xor U6380 (N_6380,N_246,N_3195);
nor U6381 (N_6381,N_70,N_806);
nor U6382 (N_6382,N_2322,N_2697);
nor U6383 (N_6383,N_3175,N_2747);
nand U6384 (N_6384,N_2172,N_1510);
nor U6385 (N_6385,N_3555,N_573);
nor U6386 (N_6386,N_4155,N_1077);
nor U6387 (N_6387,N_1878,N_3674);
or U6388 (N_6388,N_4811,N_4973);
nand U6389 (N_6389,N_980,N_2557);
nand U6390 (N_6390,N_4385,N_3466);
nor U6391 (N_6391,N_4071,N_3909);
and U6392 (N_6392,N_1850,N_1236);
nor U6393 (N_6393,N_4471,N_4404);
xnor U6394 (N_6394,N_2944,N_2197);
nand U6395 (N_6395,N_1702,N_1711);
and U6396 (N_6396,N_2863,N_1712);
and U6397 (N_6397,N_2048,N_1277);
nand U6398 (N_6398,N_4380,N_1193);
nand U6399 (N_6399,N_2247,N_854);
nor U6400 (N_6400,N_4695,N_3865);
and U6401 (N_6401,N_4025,N_4536);
or U6402 (N_6402,N_4426,N_1045);
xnor U6403 (N_6403,N_4845,N_1761);
xnor U6404 (N_6404,N_4984,N_54);
or U6405 (N_6405,N_3546,N_27);
nor U6406 (N_6406,N_4366,N_2802);
nor U6407 (N_6407,N_2821,N_2959);
and U6408 (N_6408,N_3286,N_1489);
nand U6409 (N_6409,N_3782,N_3319);
nand U6410 (N_6410,N_3993,N_78);
nor U6411 (N_6411,N_3534,N_4942);
nor U6412 (N_6412,N_4363,N_1001);
nor U6413 (N_6413,N_3750,N_4447);
or U6414 (N_6414,N_3143,N_3875);
nor U6415 (N_6415,N_4848,N_1998);
nor U6416 (N_6416,N_4029,N_2237);
xnor U6417 (N_6417,N_718,N_4872);
or U6418 (N_6418,N_3820,N_3997);
and U6419 (N_6419,N_4375,N_3624);
or U6420 (N_6420,N_3666,N_2007);
xnor U6421 (N_6421,N_303,N_1813);
and U6422 (N_6422,N_4350,N_611);
and U6423 (N_6423,N_1458,N_2145);
or U6424 (N_6424,N_116,N_3825);
or U6425 (N_6425,N_3775,N_881);
xnor U6426 (N_6426,N_2645,N_2715);
or U6427 (N_6427,N_4386,N_964);
and U6428 (N_6428,N_4979,N_3976);
and U6429 (N_6429,N_2933,N_2437);
nor U6430 (N_6430,N_3481,N_2779);
or U6431 (N_6431,N_2174,N_4039);
and U6432 (N_6432,N_796,N_1901);
nand U6433 (N_6433,N_4788,N_3160);
xor U6434 (N_6434,N_3187,N_2303);
or U6435 (N_6435,N_4290,N_3462);
and U6436 (N_6436,N_1880,N_3690);
nand U6437 (N_6437,N_1523,N_434);
nor U6438 (N_6438,N_1266,N_2720);
nand U6439 (N_6439,N_1248,N_1175);
xor U6440 (N_6440,N_4323,N_3329);
nand U6441 (N_6441,N_1394,N_3715);
or U6442 (N_6442,N_1816,N_4462);
and U6443 (N_6443,N_552,N_138);
nand U6444 (N_6444,N_1677,N_1844);
nor U6445 (N_6445,N_500,N_4798);
or U6446 (N_6446,N_1058,N_4721);
and U6447 (N_6447,N_2714,N_4813);
nor U6448 (N_6448,N_4830,N_216);
xor U6449 (N_6449,N_2205,N_427);
or U6450 (N_6450,N_1063,N_4459);
nor U6451 (N_6451,N_803,N_4021);
nand U6452 (N_6452,N_4611,N_313);
nand U6453 (N_6453,N_853,N_709);
nand U6454 (N_6454,N_355,N_3498);
xnor U6455 (N_6455,N_3602,N_1076);
or U6456 (N_6456,N_4081,N_4692);
nand U6457 (N_6457,N_2209,N_1309);
nor U6458 (N_6458,N_3487,N_3852);
nor U6459 (N_6459,N_470,N_4422);
or U6460 (N_6460,N_666,N_269);
xnor U6461 (N_6461,N_2486,N_1331);
and U6462 (N_6462,N_2884,N_4840);
or U6463 (N_6463,N_4042,N_2642);
nand U6464 (N_6464,N_4787,N_692);
and U6465 (N_6465,N_2434,N_2516);
or U6466 (N_6466,N_4614,N_423);
nand U6467 (N_6467,N_1244,N_4401);
nand U6468 (N_6468,N_202,N_618);
nor U6469 (N_6469,N_2118,N_4332);
nor U6470 (N_6470,N_1390,N_970);
and U6471 (N_6471,N_2073,N_4817);
nand U6472 (N_6472,N_556,N_3499);
and U6473 (N_6473,N_4554,N_1025);
nand U6474 (N_6474,N_2141,N_3680);
and U6475 (N_6475,N_2843,N_1928);
nor U6476 (N_6476,N_4165,N_4839);
nor U6477 (N_6477,N_3914,N_4307);
and U6478 (N_6478,N_2778,N_2433);
or U6479 (N_6479,N_3020,N_3204);
nor U6480 (N_6480,N_3685,N_3384);
and U6481 (N_6481,N_680,N_639);
and U6482 (N_6482,N_4415,N_4117);
nor U6483 (N_6483,N_402,N_3406);
nand U6484 (N_6484,N_1987,N_4495);
nor U6485 (N_6485,N_1432,N_1612);
nor U6486 (N_6486,N_4875,N_1085);
and U6487 (N_6487,N_4510,N_2451);
nor U6488 (N_6488,N_3456,N_1177);
nor U6489 (N_6489,N_1760,N_4680);
xor U6490 (N_6490,N_3844,N_3252);
xor U6491 (N_6491,N_2046,N_1451);
or U6492 (N_6492,N_3118,N_4827);
nor U6493 (N_6493,N_787,N_2538);
xor U6494 (N_6494,N_1897,N_3772);
and U6495 (N_6495,N_1288,N_2155);
xor U6496 (N_6496,N_2515,N_4082);
and U6497 (N_6497,N_4478,N_716);
and U6498 (N_6498,N_3155,N_4645);
xnor U6499 (N_6499,N_2394,N_1468);
xnor U6500 (N_6500,N_2961,N_4313);
and U6501 (N_6501,N_4243,N_285);
or U6502 (N_6502,N_1509,N_3831);
xnor U6503 (N_6503,N_255,N_1042);
and U6504 (N_6504,N_1282,N_913);
and U6505 (N_6505,N_4335,N_3306);
or U6506 (N_6506,N_2507,N_2628);
and U6507 (N_6507,N_2092,N_734);
or U6508 (N_6508,N_1496,N_300);
or U6509 (N_6509,N_3725,N_1150);
nand U6510 (N_6510,N_3023,N_4393);
or U6511 (N_6511,N_4334,N_3751);
nor U6512 (N_6512,N_4852,N_4912);
nor U6513 (N_6513,N_3522,N_1020);
and U6514 (N_6514,N_513,N_2268);
or U6515 (N_6515,N_4746,N_3352);
or U6516 (N_6516,N_2024,N_1100);
nand U6517 (N_6517,N_1716,N_4608);
xor U6518 (N_6518,N_3336,N_1348);
or U6519 (N_6519,N_2308,N_2256);
or U6520 (N_6520,N_2868,N_2668);
xor U6521 (N_6521,N_2895,N_2947);
xnor U6522 (N_6522,N_1145,N_272);
xnor U6523 (N_6523,N_115,N_211);
nand U6524 (N_6524,N_1842,N_3368);
nor U6525 (N_6525,N_4099,N_2842);
or U6526 (N_6526,N_3622,N_4751);
and U6527 (N_6527,N_3953,N_3552);
nor U6528 (N_6528,N_3048,N_2820);
and U6529 (N_6529,N_3532,N_166);
nand U6530 (N_6530,N_2733,N_3567);
nor U6531 (N_6531,N_1305,N_1890);
xnor U6532 (N_6532,N_2972,N_1437);
xor U6533 (N_6533,N_1349,N_2623);
and U6534 (N_6534,N_1627,N_4691);
nor U6535 (N_6535,N_1522,N_4762);
nor U6536 (N_6536,N_686,N_2692);
nand U6537 (N_6537,N_3863,N_3093);
or U6538 (N_6538,N_4861,N_4487);
or U6539 (N_6539,N_3860,N_3924);
or U6540 (N_6540,N_2937,N_4160);
nor U6541 (N_6541,N_2765,N_3679);
and U6542 (N_6542,N_4304,N_825);
xor U6543 (N_6543,N_4402,N_267);
nor U6544 (N_6544,N_2154,N_920);
nand U6545 (N_6545,N_3405,N_2402);
nand U6546 (N_6546,N_1127,N_1545);
and U6547 (N_6547,N_2621,N_1674);
xnor U6548 (N_6548,N_4516,N_4014);
and U6549 (N_6549,N_2837,N_4546);
and U6550 (N_6550,N_4635,N_4783);
and U6551 (N_6551,N_412,N_1906);
nand U6552 (N_6552,N_3520,N_3811);
nor U6553 (N_6553,N_4628,N_153);
nand U6554 (N_6554,N_2871,N_3412);
or U6555 (N_6555,N_1264,N_2791);
and U6556 (N_6556,N_4551,N_3678);
or U6557 (N_6557,N_1274,N_1843);
or U6558 (N_6558,N_987,N_4124);
and U6559 (N_6559,N_1758,N_3970);
nor U6560 (N_6560,N_3903,N_4325);
nor U6561 (N_6561,N_4345,N_3745);
nand U6562 (N_6562,N_209,N_4020);
or U6563 (N_6563,N_2631,N_4233);
and U6564 (N_6564,N_1055,N_4045);
and U6565 (N_6565,N_4988,N_4396);
and U6566 (N_6566,N_2010,N_570);
or U6567 (N_6567,N_2614,N_3270);
nor U6568 (N_6568,N_4502,N_2064);
nor U6569 (N_6569,N_1216,N_4539);
nor U6570 (N_6570,N_1856,N_4454);
nor U6571 (N_6571,N_844,N_1148);
nor U6572 (N_6572,N_3485,N_4816);
and U6573 (N_6573,N_3704,N_2619);
and U6574 (N_6574,N_1577,N_961);
xor U6575 (N_6575,N_2091,N_1903);
xnor U6576 (N_6576,N_2855,N_3979);
nand U6577 (N_6577,N_48,N_3855);
nand U6578 (N_6578,N_3375,N_3394);
nand U6579 (N_6579,N_3055,N_3814);
and U6580 (N_6580,N_4455,N_3888);
nand U6581 (N_6581,N_4425,N_2761);
nor U6582 (N_6582,N_1367,N_1736);
nor U6583 (N_6583,N_2901,N_4619);
or U6584 (N_6584,N_249,N_4527);
nand U6585 (N_6585,N_2038,N_4707);
nor U6586 (N_6586,N_2676,N_4232);
nand U6587 (N_6587,N_4506,N_4543);
and U6588 (N_6588,N_1016,N_3014);
and U6589 (N_6589,N_1916,N_1991);
and U6590 (N_6590,N_2505,N_3659);
and U6591 (N_6591,N_2478,N_3232);
nor U6592 (N_6592,N_4286,N_3434);
nand U6593 (N_6593,N_2200,N_477);
or U6594 (N_6594,N_12,N_445);
nor U6595 (N_6595,N_1809,N_3039);
xor U6596 (N_6596,N_1379,N_2397);
nand U6597 (N_6597,N_804,N_4235);
or U6598 (N_6598,N_591,N_120);
nand U6599 (N_6599,N_2150,N_2570);
and U6600 (N_6600,N_2139,N_4033);
and U6601 (N_6601,N_1310,N_967);
nor U6602 (N_6602,N_1156,N_4853);
nor U6603 (N_6603,N_1725,N_1024);
nand U6604 (N_6604,N_1028,N_3586);
nor U6605 (N_6605,N_3432,N_3938);
nand U6606 (N_6606,N_4047,N_3746);
or U6607 (N_6607,N_3226,N_3786);
or U6608 (N_6608,N_1484,N_3281);
nor U6609 (N_6609,N_3292,N_1952);
nand U6610 (N_6610,N_4138,N_745);
nor U6611 (N_6611,N_4392,N_1448);
nor U6612 (N_6612,N_4436,N_4108);
nor U6613 (N_6613,N_4587,N_4194);
nor U6614 (N_6614,N_3940,N_1715);
nand U6615 (N_6615,N_1009,N_320);
xor U6616 (N_6616,N_1691,N_3389);
nor U6617 (N_6617,N_539,N_411);
nor U6618 (N_6618,N_4028,N_4061);
nand U6619 (N_6619,N_3583,N_254);
and U6620 (N_6620,N_304,N_977);
or U6621 (N_6621,N_4322,N_2388);
and U6622 (N_6622,N_3217,N_1837);
nand U6623 (N_6623,N_3139,N_4710);
nor U6624 (N_6624,N_4934,N_4477);
nand U6625 (N_6625,N_4972,N_2474);
or U6626 (N_6626,N_51,N_4265);
nand U6627 (N_6627,N_3688,N_648);
or U6628 (N_6628,N_4359,N_144);
or U6629 (N_6629,N_2123,N_4923);
and U6630 (N_6630,N_2182,N_1653);
or U6631 (N_6631,N_1549,N_2571);
and U6632 (N_6632,N_1226,N_368);
or U6633 (N_6633,N_2658,N_3800);
nand U6634 (N_6634,N_1197,N_3153);
and U6635 (N_6635,N_3818,N_2951);
nor U6636 (N_6636,N_4739,N_4434);
nand U6637 (N_6637,N_4549,N_358);
and U6638 (N_6638,N_4321,N_1563);
or U6639 (N_6639,N_969,N_1227);
nand U6640 (N_6640,N_428,N_2292);
nand U6641 (N_6641,N_4930,N_873);
nand U6642 (N_6642,N_3878,N_703);
nor U6643 (N_6643,N_4971,N_3127);
nand U6644 (N_6644,N_466,N_2958);
nand U6645 (N_6645,N_430,N_4184);
and U6646 (N_6646,N_2377,N_2880);
nor U6647 (N_6647,N_2749,N_2912);
xor U6648 (N_6648,N_612,N_2283);
xnor U6649 (N_6649,N_1335,N_2033);
nand U6650 (N_6650,N_765,N_2556);
xor U6651 (N_6651,N_3268,N_850);
or U6652 (N_6652,N_175,N_1929);
nor U6653 (N_6653,N_345,N_3340);
nand U6654 (N_6654,N_3962,N_2501);
nand U6655 (N_6655,N_2483,N_4006);
and U6656 (N_6656,N_2264,N_2370);
nand U6657 (N_6657,N_357,N_983);
nor U6658 (N_6658,N_707,N_1052);
or U6659 (N_6659,N_1062,N_100);
nand U6660 (N_6660,N_3911,N_2808);
nand U6661 (N_6661,N_3325,N_827);
nor U6662 (N_6662,N_3445,N_1662);
and U6663 (N_6663,N_3594,N_3971);
nand U6664 (N_6664,N_3031,N_2992);
nor U6665 (N_6665,N_2452,N_4927);
nand U6666 (N_6666,N_3931,N_1644);
or U6667 (N_6667,N_3066,N_2101);
or U6668 (N_6668,N_150,N_2909);
and U6669 (N_6669,N_4613,N_2390);
or U6670 (N_6670,N_1964,N_1787);
nand U6671 (N_6671,N_3044,N_3448);
xnor U6672 (N_6672,N_2529,N_409);
nor U6673 (N_6673,N_4590,N_4967);
nand U6674 (N_6674,N_3837,N_1628);
or U6675 (N_6675,N_2214,N_1825);
nor U6676 (N_6676,N_3913,N_2302);
xnor U6677 (N_6677,N_4277,N_2773);
and U6678 (N_6678,N_3337,N_2305);
nand U6679 (N_6679,N_111,N_4244);
or U6680 (N_6680,N_777,N_2149);
or U6681 (N_6681,N_1801,N_3513);
or U6682 (N_6682,N_1151,N_3912);
nand U6683 (N_6683,N_1532,N_2581);
or U6684 (N_6684,N_2275,N_3675);
nor U6685 (N_6685,N_3423,N_2665);
nor U6686 (N_6686,N_2252,N_1159);
nor U6687 (N_6687,N_4924,N_4064);
nand U6688 (N_6688,N_3897,N_744);
and U6689 (N_6689,N_2860,N_4074);
and U6690 (N_6690,N_1056,N_2047);
or U6691 (N_6691,N_2971,N_2981);
and U6692 (N_6692,N_4790,N_4766);
or U6693 (N_6693,N_65,N_420);
nand U6694 (N_6694,N_2770,N_4059);
and U6695 (N_6695,N_3563,N_3447);
nand U6696 (N_6696,N_1620,N_2107);
xnor U6697 (N_6697,N_1932,N_1633);
nor U6698 (N_6698,N_1907,N_256);
or U6699 (N_6699,N_2324,N_3387);
or U6700 (N_6700,N_3958,N_3303);
nand U6701 (N_6701,N_2441,N_1530);
and U6702 (N_6702,N_784,N_5);
or U6703 (N_6703,N_1333,N_4792);
nor U6704 (N_6704,N_3887,N_1607);
nor U6705 (N_6705,N_1202,N_45);
or U6706 (N_6706,N_1613,N_4969);
nand U6707 (N_6707,N_2751,N_726);
xnor U6708 (N_6708,N_4337,N_2245);
and U6709 (N_6709,N_4822,N_4051);
xnor U6710 (N_6710,N_1409,N_1238);
nand U6711 (N_6711,N_2226,N_584);
nand U6712 (N_6712,N_4893,N_1529);
and U6713 (N_6713,N_993,N_273);
or U6714 (N_6714,N_2015,N_2093);
xor U6715 (N_6715,N_1022,N_3632);
nor U6716 (N_6716,N_4338,N_3579);
nand U6717 (N_6717,N_1272,N_4023);
nand U6718 (N_6718,N_3478,N_753);
and U6719 (N_6719,N_1075,N_3179);
and U6720 (N_6720,N_3285,N_3490);
nand U6721 (N_6721,N_4227,N_1364);
nor U6722 (N_6722,N_1402,N_1414);
and U6723 (N_6723,N_1954,N_2447);
and U6724 (N_6724,N_2471,N_2353);
or U6725 (N_6725,N_1718,N_831);
nand U6726 (N_6726,N_1281,N_365);
and U6727 (N_6727,N_909,N_1098);
nor U6728 (N_6728,N_1330,N_2244);
nand U6729 (N_6729,N_2635,N_3560);
or U6730 (N_6730,N_1480,N_2110);
nor U6731 (N_6731,N_614,N_4663);
nor U6732 (N_6732,N_1185,N_3233);
nand U6733 (N_6733,N_4501,N_4234);
and U6734 (N_6734,N_1207,N_2670);
nand U6735 (N_6735,N_616,N_2499);
and U6736 (N_6736,N_2881,N_4807);
or U6737 (N_6737,N_2964,N_501);
xnor U6738 (N_6738,N_1462,N_3080);
nand U6739 (N_6739,N_1135,N_199);
xor U6740 (N_6740,N_4090,N_2709);
or U6741 (N_6741,N_2940,N_4785);
or U6742 (N_6742,N_387,N_1879);
and U6743 (N_6743,N_3597,N_3665);
or U6744 (N_6744,N_2807,N_1862);
and U6745 (N_6745,N_3322,N_2075);
nor U6746 (N_6746,N_840,N_4161);
nand U6747 (N_6747,N_3212,N_3416);
nor U6748 (N_6748,N_1751,N_1829);
nor U6749 (N_6749,N_2440,N_4773);
nor U6750 (N_6750,N_1168,N_1667);
nor U6751 (N_6751,N_20,N_245);
or U6752 (N_6752,N_749,N_68);
or U6753 (N_6753,N_3930,N_644);
or U6754 (N_6754,N_535,N_4077);
nor U6755 (N_6755,N_4574,N_627);
or U6756 (N_6756,N_4018,N_3358);
nor U6757 (N_6757,N_439,N_3227);
or U6758 (N_6758,N_4700,N_3029);
and U6759 (N_6759,N_1096,N_3689);
or U6760 (N_6760,N_4491,N_1138);
and U6761 (N_6761,N_1836,N_901);
or U6762 (N_6762,N_4756,N_2730);
and U6763 (N_6763,N_2567,N_3326);
and U6764 (N_6764,N_3623,N_2480);
nand U6765 (N_6765,N_4750,N_74);
and U6766 (N_6766,N_1230,N_3299);
nor U6767 (N_6767,N_3919,N_2386);
xnor U6768 (N_6768,N_2381,N_3356);
nor U6769 (N_6769,N_3450,N_1050);
and U6770 (N_6770,N_1868,N_52);
or U6771 (N_6771,N_1804,N_1600);
and U6772 (N_6772,N_2309,N_398);
xor U6773 (N_6773,N_3088,N_1676);
nand U6774 (N_6774,N_29,N_659);
and U6775 (N_6775,N_2758,N_4760);
nor U6776 (N_6776,N_1251,N_1108);
or U6777 (N_6777,N_4284,N_1977);
and U6778 (N_6778,N_2991,N_2354);
or U6779 (N_6779,N_1487,N_772);
and U6780 (N_6780,N_996,N_2620);
or U6781 (N_6781,N_1129,N_1300);
nor U6782 (N_6782,N_974,N_4480);
nand U6783 (N_6783,N_3059,N_807);
xor U6784 (N_6784,N_2333,N_1212);
nand U6785 (N_6785,N_4892,N_4658);
and U6786 (N_6786,N_812,N_4174);
nor U6787 (N_6787,N_3893,N_2194);
and U6788 (N_6788,N_2435,N_3454);
or U6789 (N_6789,N_3535,N_2117);
nor U6790 (N_6790,N_4496,N_1118);
nand U6791 (N_6791,N_1473,N_3221);
or U6792 (N_6792,N_740,N_3305);
nand U6793 (N_6793,N_3194,N_1293);
and U6794 (N_6794,N_1595,N_62);
and U6795 (N_6795,N_2310,N_3174);
nor U6796 (N_6796,N_2171,N_339);
or U6797 (N_6797,N_105,N_2890);
and U6798 (N_6798,N_3902,N_1920);
and U6799 (N_6799,N_2086,N_1513);
xnor U6800 (N_6800,N_4597,N_123);
nand U6801 (N_6801,N_2662,N_1727);
or U6802 (N_6802,N_2042,N_2406);
and U6803 (N_6803,N_3991,N_4890);
or U6804 (N_6804,N_2462,N_493);
nand U6805 (N_6805,N_1163,N_4678);
xnor U6806 (N_6806,N_456,N_3429);
and U6807 (N_6807,N_4718,N_4348);
nor U6808 (N_6808,N_3832,N_2616);
or U6809 (N_6809,N_91,N_3074);
xnor U6810 (N_6810,N_397,N_201);
and U6811 (N_6811,N_3857,N_1237);
or U6812 (N_6812,N_4413,N_3876);
nor U6813 (N_6813,N_3280,N_2137);
or U6814 (N_6814,N_414,N_4320);
nand U6815 (N_6815,N_2068,N_4268);
nand U6816 (N_6816,N_2108,N_904);
nand U6817 (N_6817,N_4823,N_1610);
nor U6818 (N_6818,N_653,N_3982);
nor U6819 (N_6819,N_4896,N_147);
or U6820 (N_6820,N_2232,N_3250);
and U6821 (N_6821,N_3937,N_2493);
and U6822 (N_6822,N_583,N_265);
and U6823 (N_6823,N_2968,N_791);
and U6824 (N_6824,N_1316,N_1642);
and U6825 (N_6825,N_938,N_3802);
or U6826 (N_6826,N_1951,N_1588);
nand U6827 (N_6827,N_4693,N_1788);
nand U6828 (N_6828,N_2355,N_3100);
nand U6829 (N_6829,N_3974,N_3483);
or U6830 (N_6830,N_893,N_3279);
nand U6831 (N_6831,N_3035,N_2120);
nor U6832 (N_6832,N_1231,N_1187);
and U6833 (N_6833,N_2102,N_4686);
nand U6834 (N_6834,N_2306,N_104);
or U6835 (N_6835,N_3949,N_2624);
and U6836 (N_6836,N_3609,N_1376);
or U6837 (N_6837,N_1439,N_3076);
or U6838 (N_6838,N_3736,N_3408);
or U6839 (N_6839,N_4791,N_3759);
nor U6840 (N_6840,N_4252,N_2001);
and U6841 (N_6841,N_4856,N_4563);
or U6842 (N_6842,N_4948,N_3125);
nand U6843 (N_6843,N_3796,N_4423);
and U6844 (N_6844,N_4399,N_4388);
nand U6845 (N_6845,N_3441,N_2273);
xor U6846 (N_6846,N_4834,N_2260);
or U6847 (N_6847,N_3201,N_1033);
and U6848 (N_6848,N_124,N_184);
and U6849 (N_6849,N_4149,N_3557);
and U6850 (N_6850,N_4429,N_4043);
nor U6851 (N_6851,N_3430,N_253);
or U6852 (N_6852,N_3630,N_279);
nand U6853 (N_6853,N_373,N_1373);
nand U6854 (N_6854,N_2074,N_3159);
xor U6855 (N_6855,N_3706,N_1141);
nand U6856 (N_6856,N_778,N_1746);
nand U6857 (N_6857,N_1417,N_229);
nor U6858 (N_6858,N_3256,N_444);
nor U6859 (N_6859,N_4540,N_173);
and U6860 (N_6860,N_250,N_2879);
xnor U6861 (N_6861,N_290,N_4796);
and U6862 (N_6862,N_1541,N_2634);
and U6863 (N_6863,N_4318,N_4106);
and U6864 (N_6864,N_2735,N_872);
nor U6865 (N_6865,N_3667,N_3156);
or U6866 (N_6866,N_3293,N_597);
nor U6867 (N_6867,N_3590,N_792);
or U6868 (N_6868,N_719,N_3409);
and U6869 (N_6869,N_661,N_1358);
nor U6870 (N_6870,N_638,N_329);
and U6871 (N_6871,N_3708,N_275);
or U6872 (N_6872,N_443,N_2533);
and U6873 (N_6873,N_3402,N_3120);
nor U6874 (N_6874,N_1095,N_234);
nor U6875 (N_6875,N_348,N_775);
and U6876 (N_6876,N_1544,N_2687);
or U6877 (N_6877,N_1040,N_1200);
or U6878 (N_6878,N_1396,N_3307);
nor U6879 (N_6879,N_4328,N_4120);
nor U6880 (N_6880,N_4704,N_4781);
nand U6881 (N_6881,N_4661,N_667);
or U6882 (N_6882,N_2936,N_1713);
and U6883 (N_6883,N_4854,N_2726);
nand U6884 (N_6884,N_2562,N_4583);
and U6885 (N_6885,N_832,N_2337);
and U6886 (N_6886,N_1793,N_1126);
nor U6887 (N_6887,N_4139,N_4883);
nand U6888 (N_6888,N_4515,N_3298);
or U6889 (N_6889,N_2450,N_1220);
nor U6890 (N_6890,N_3359,N_257);
xor U6891 (N_6891,N_2729,N_1269);
or U6892 (N_6892,N_2659,N_2116);
and U6893 (N_6893,N_3378,N_299);
nand U6894 (N_6894,N_3501,N_4073);
or U6895 (N_6895,N_3239,N_1164);
and U6896 (N_6896,N_4251,N_3027);
or U6897 (N_6897,N_33,N_4204);
nand U6898 (N_6898,N_2827,N_2838);
nor U6899 (N_6899,N_3335,N_4504);
or U6900 (N_6900,N_2135,N_1778);
or U6901 (N_6901,N_2566,N_4153);
or U6902 (N_6902,N_324,N_1689);
and U6903 (N_6903,N_418,N_4121);
and U6904 (N_6904,N_1037,N_1057);
or U6905 (N_6905,N_4849,N_3934);
nor U6906 (N_6906,N_1709,N_1347);
and U6907 (N_6907,N_4740,N_3235);
nand U6908 (N_6908,N_963,N_3010);
nand U6909 (N_6909,N_3683,N_3037);
or U6910 (N_6910,N_4612,N_3114);
nand U6911 (N_6911,N_99,N_2663);
and U6912 (N_6912,N_2008,N_1594);
nor U6913 (N_6913,N_2307,N_3436);
and U6914 (N_6914,N_2928,N_223);
and U6915 (N_6915,N_1470,N_237);
nor U6916 (N_6916,N_2654,N_4874);
nand U6917 (N_6917,N_4598,N_1101);
nor U6918 (N_6918,N_3137,N_4876);
nor U6919 (N_6919,N_468,N_619);
or U6920 (N_6920,N_2752,N_119);
nor U6921 (N_6921,N_3809,N_69);
and U6922 (N_6922,N_4728,N_1443);
or U6923 (N_6923,N_3541,N_3477);
or U6924 (N_6924,N_3790,N_999);
nor U6925 (N_6925,N_4526,N_1294);
and U6926 (N_6926,N_2652,N_3817);
or U6927 (N_6927,N_1557,N_4191);
nand U6928 (N_6928,N_2798,N_1622);
nand U6929 (N_6929,N_4245,N_2805);
or U6930 (N_6930,N_1961,N_4863);
and U6931 (N_6931,N_252,N_2524);
nand U6932 (N_6932,N_502,N_3584);
xnor U6933 (N_6933,N_3344,N_3774);
nand U6934 (N_6934,N_1438,N_1729);
nand U6935 (N_6935,N_846,N_2115);
or U6936 (N_6936,N_2899,N_3007);
or U6937 (N_6937,N_3823,N_4804);
and U6938 (N_6938,N_3625,N_2766);
and U6939 (N_6939,N_2227,N_1223);
nor U6940 (N_6940,N_1240,N_298);
nor U6941 (N_6941,N_2577,N_2768);
and U6942 (N_6942,N_4533,N_4100);
nand U6943 (N_6943,N_1569,N_3422);
nand U6944 (N_6944,N_2025,N_3654);
or U6945 (N_6945,N_3197,N_1597);
and U6946 (N_6946,N_679,N_2414);
or U6947 (N_6947,N_3166,N_3170);
nor U6948 (N_6948,N_3472,N_1234);
xnor U6949 (N_6949,N_278,N_3889);
and U6950 (N_6950,N_930,N_1974);
nor U6951 (N_6951,N_3592,N_1371);
nand U6952 (N_6952,N_4857,N_3755);
nand U6953 (N_6953,N_1395,N_4789);
and U6954 (N_6954,N_1547,N_943);
or U6955 (N_6955,N_1548,N_2906);
or U6956 (N_6956,N_3391,N_128);
or U6957 (N_6957,N_2319,N_1196);
or U6958 (N_6958,N_2719,N_3006);
and U6959 (N_6959,N_1450,N_1426);
and U6960 (N_6960,N_4295,N_4308);
or U6961 (N_6961,N_3896,N_2029);
and U6962 (N_6962,N_2990,N_4068);
nor U6963 (N_6963,N_2639,N_2534);
nand U6964 (N_6964,N_2274,N_3202);
nor U6965 (N_6965,N_35,N_2626);
xnor U6966 (N_6966,N_4352,N_1956);
nand U6967 (N_6967,N_4431,N_522);
nand U6968 (N_6968,N_1546,N_4977);
or U6969 (N_6969,N_3172,N_622);
nor U6970 (N_6970,N_939,N_1870);
and U6971 (N_6971,N_2059,N_2925);
and U6972 (N_6972,N_581,N_1143);
nor U6973 (N_6973,N_1581,N_1763);
nor U6974 (N_6974,N_3851,N_3323);
and U6975 (N_6975,N_1738,N_4943);
nand U6976 (N_6976,N_2027,N_1874);
nand U6977 (N_6977,N_1625,N_1640);
xnor U6978 (N_6978,N_3090,N_191);
nand U6979 (N_6979,N_3861,N_2129);
nor U6980 (N_6980,N_866,N_3548);
nand U6981 (N_6981,N_1841,N_3651);
and U6982 (N_6982,N_1810,N_1755);
nor U6983 (N_6983,N_1818,N_1314);
and U6984 (N_6984,N_4865,N_3206);
and U6985 (N_6985,N_2502,N_813);
nand U6986 (N_6986,N_3658,N_469);
nor U6987 (N_6987,N_3713,N_1516);
nand U6988 (N_6988,N_965,N_1944);
nor U6989 (N_6989,N_1412,N_878);
and U6990 (N_6990,N_4779,N_979);
or U6991 (N_6991,N_1486,N_4589);
or U6992 (N_6992,N_1861,N_1292);
nand U6993 (N_6993,N_3646,N_2935);
nand U6994 (N_6994,N_708,N_774);
or U6995 (N_6995,N_2272,N_1701);
and U6996 (N_6996,N_2242,N_2885);
and U6997 (N_6997,N_1853,N_2553);
or U6998 (N_6998,N_1772,N_3295);
nor U6999 (N_6999,N_3072,N_2312);
or U7000 (N_7000,N_2800,N_2144);
nor U7001 (N_7001,N_1636,N_4774);
and U7002 (N_7002,N_2754,N_42);
or U7003 (N_7003,N_372,N_136);
or U7004 (N_7004,N_1171,N_4954);
nor U7005 (N_7005,N_3057,N_239);
and U7006 (N_7006,N_323,N_2504);
nor U7007 (N_7007,N_3872,N_4198);
nand U7008 (N_7008,N_1247,N_4214);
and U7009 (N_7009,N_4553,N_1258);
nand U7010 (N_7010,N_2362,N_1181);
nand U7011 (N_7011,N_1994,N_1131);
and U7012 (N_7012,N_3744,N_3463);
nand U7013 (N_7013,N_3530,N_1921);
xor U7014 (N_7014,N_3827,N_2217);
or U7015 (N_7015,N_1424,N_4689);
or U7016 (N_7016,N_4367,N_1283);
and U7017 (N_7017,N_4070,N_472);
or U7018 (N_7018,N_2625,N_1286);
nor U7019 (N_7019,N_1852,N_2710);
nor U7020 (N_7020,N_4882,N_2512);
or U7021 (N_7021,N_3188,N_366);
nor U7022 (N_7022,N_2018,N_4479);
nor U7023 (N_7023,N_4676,N_3366);
nand U7024 (N_7024,N_2536,N_3595);
nand U7025 (N_7025,N_178,N_2125);
xnor U7026 (N_7026,N_1657,N_2183);
and U7027 (N_7027,N_2423,N_4903);
and U7028 (N_7028,N_3267,N_864);
nand U7029 (N_7029,N_567,N_3536);
or U7030 (N_7030,N_4617,N_836);
and U7031 (N_7031,N_593,N_386);
and U7032 (N_7032,N_546,N_1959);
nor U7033 (N_7033,N_2900,N_2263);
nand U7034 (N_7034,N_1354,N_3957);
and U7035 (N_7035,N_3241,N_4219);
or U7036 (N_7036,N_3215,N_2739);
and U7037 (N_7037,N_72,N_2744);
nand U7038 (N_7038,N_2931,N_204);
nand U7039 (N_7039,N_4667,N_3265);
nor U7040 (N_7040,N_4096,N_1703);
or U7041 (N_7041,N_220,N_1043);
and U7042 (N_7042,N_3321,N_483);
nor U7043 (N_7043,N_3479,N_3369);
or U7044 (N_7044,N_3732,N_3932);
nor U7045 (N_7045,N_3606,N_1835);
nor U7046 (N_7046,N_3077,N_221);
or U7047 (N_7047,N_1652,N_1315);
nand U7048 (N_7048,N_3662,N_2159);
nor U7049 (N_7049,N_781,N_4484);
or U7050 (N_7050,N_4128,N_3841);
or U7051 (N_7051,N_1635,N_1383);
nand U7052 (N_7052,N_656,N_3572);
or U7053 (N_7053,N_2573,N_3433);
nor U7054 (N_7054,N_3881,N_3320);
xor U7055 (N_7055,N_3327,N_1307);
or U7056 (N_7056,N_3848,N_3043);
nor U7057 (N_7057,N_3839,N_1917);
xnor U7058 (N_7058,N_17,N_3064);
nor U7059 (N_7059,N_2669,N_617);
nand U7060 (N_7060,N_3246,N_2904);
or U7061 (N_7061,N_332,N_1950);
or U7062 (N_7062,N_2131,N_2034);
nor U7063 (N_7063,N_637,N_2918);
or U7064 (N_7064,N_2473,N_2121);
and U7065 (N_7065,N_1566,N_4638);
nor U7066 (N_7066,N_2146,N_457);
nor U7067 (N_7067,N_1675,N_2193);
nand U7068 (N_7068,N_4538,N_4646);
or U7069 (N_7069,N_3987,N_2346);
nor U7070 (N_7070,N_1139,N_547);
or U7071 (N_7071,N_2876,N_4105);
nand U7072 (N_7072,N_3575,N_4809);
nor U7073 (N_7073,N_3652,N_3766);
xnor U7074 (N_7074,N_2168,N_4558);
nor U7075 (N_7075,N_4500,N_1494);
nand U7076 (N_7076,N_2875,N_3819);
nand U7077 (N_7077,N_4176,N_2542);
or U7078 (N_7078,N_2191,N_4803);
or U7079 (N_7079,N_3253,N_2846);
and U7080 (N_7080,N_1990,N_1182);
or U7081 (N_7081,N_4452,N_2633);
nor U7082 (N_7082,N_25,N_4409);
or U7083 (N_7083,N_4129,N_3507);
and U7084 (N_7084,N_145,N_4986);
and U7085 (N_7085,N_902,N_1783);
or U7086 (N_7086,N_3067,N_1601);
nand U7087 (N_7087,N_2444,N_429);
and U7088 (N_7088,N_4620,N_2731);
nor U7089 (N_7089,N_1537,N_2850);
nor U7090 (N_7090,N_1900,N_3365);
nand U7091 (N_7091,N_2112,N_876);
nor U7092 (N_7092,N_3697,N_180);
and U7093 (N_7093,N_4403,N_3142);
nand U7094 (N_7094,N_1573,N_3411);
nor U7095 (N_7095,N_3117,N_1860);
or U7096 (N_7096,N_4936,N_4669);
nand U7097 (N_7097,N_2179,N_3024);
or U7098 (N_7098,N_1132,N_1146);
and U7099 (N_7099,N_2057,N_801);
nor U7100 (N_7100,N_1430,N_360);
and U7101 (N_7101,N_1953,N_146);
xnor U7102 (N_7102,N_1866,N_3724);
xnor U7103 (N_7103,N_505,N_2640);
nor U7104 (N_7104,N_1249,N_4950);
or U7105 (N_7105,N_808,N_1664);
xor U7106 (N_7106,N_997,N_520);
and U7107 (N_7107,N_3763,N_3417);
or U7108 (N_7108,N_4344,N_471);
or U7109 (N_7109,N_2400,N_3884);
xor U7110 (N_7110,N_2889,N_743);
and U7111 (N_7111,N_308,N_460);
or U7112 (N_7112,N_1005,N_4126);
nor U7113 (N_7113,N_4655,N_4525);
nor U7114 (N_7114,N_2442,N_877);
xor U7115 (N_7115,N_3612,N_1499);
nor U7116 (N_7116,N_3357,N_820);
or U7117 (N_7117,N_4027,N_1493);
and U7118 (N_7118,N_1578,N_3461);
xnor U7119 (N_7119,N_2615,N_4690);
nand U7120 (N_7120,N_1988,N_4602);
xnor U7121 (N_7121,N_2545,N_2140);
nor U7122 (N_7122,N_58,N_978);
or U7123 (N_7123,N_1074,N_2650);
nor U7124 (N_7124,N_3838,N_886);
nor U7125 (N_7125,N_4519,N_3185);
nor U7126 (N_7126,N_3078,N_958);
nand U7127 (N_7127,N_1914,N_4652);
and U7128 (N_7128,N_4473,N_3617);
nor U7129 (N_7129,N_3850,N_4919);
or U7130 (N_7130,N_2459,N_2973);
or U7131 (N_7131,N_3942,N_2994);
or U7132 (N_7132,N_3545,N_798);
nor U7133 (N_7133,N_2253,N_4677);
and U7134 (N_7134,N_986,N_3721);
nor U7135 (N_7135,N_1299,N_3081);
nor U7136 (N_7136,N_452,N_4987);
nand U7137 (N_7137,N_1372,N_2552);
nor U7138 (N_7138,N_1794,N_2847);
nand U7139 (N_7139,N_3275,N_1538);
nor U7140 (N_7140,N_1030,N_3867);
and U7141 (N_7141,N_382,N_3435);
and U7142 (N_7142,N_1334,N_1872);
and U7143 (N_7143,N_2559,N_283);
or U7144 (N_7144,N_2728,N_2040);
or U7145 (N_7145,N_473,N_1355);
nand U7146 (N_7146,N_2053,N_992);
or U7147 (N_7147,N_2070,N_340);
and U7148 (N_7148,N_77,N_1276);
nand U7149 (N_7149,N_4369,N_538);
and U7150 (N_7150,N_2239,N_558);
nor U7151 (N_7151,N_2201,N_80);
xor U7152 (N_7152,N_2488,N_1784);
nand U7153 (N_7153,N_767,N_4968);
and U7154 (N_7154,N_1905,N_1340);
or U7155 (N_7155,N_86,N_4581);
and U7156 (N_7156,N_156,N_1475);
or U7157 (N_7157,N_4497,N_4560);
nand U7158 (N_7158,N_507,N_235);
or U7159 (N_7159,N_2657,N_2998);
and U7160 (N_7160,N_3764,N_162);
xnor U7161 (N_7161,N_2558,N_2464);
xor U7162 (N_7162,N_2721,N_4427);
nand U7163 (N_7163,N_2584,N_3554);
xor U7164 (N_7164,N_3225,N_494);
nor U7165 (N_7165,N_2436,N_3660);
nor U7166 (N_7166,N_4734,N_2711);
or U7167 (N_7167,N_4300,N_839);
nor U7168 (N_7168,N_32,N_264);
nand U7169 (N_7169,N_2856,N_2378);
and U7170 (N_7170,N_560,N_4866);
xnor U7171 (N_7171,N_3944,N_4651);
and U7172 (N_7172,N_4604,N_3640);
nand U7173 (N_7173,N_109,N_3967);
or U7174 (N_7174,N_2089,N_4437);
nand U7175 (N_7175,N_3710,N_3981);
nand U7176 (N_7176,N_4397,N_760);
and U7177 (N_7177,N_4782,N_1740);
nor U7178 (N_7178,N_880,N_2923);
and U7179 (N_7179,N_3439,N_4238);
nand U7180 (N_7180,N_2429,N_1967);
nand U7181 (N_7181,N_437,N_2920);
or U7182 (N_7182,N_1770,N_1969);
nor U7183 (N_7183,N_2678,N_438);
nor U7184 (N_7184,N_4384,N_642);
and U7185 (N_7185,N_911,N_631);
nor U7186 (N_7186,N_1423,N_4730);
or U7187 (N_7187,N_1587,N_2228);
or U7188 (N_7188,N_1590,N_2251);
nor U7189 (N_7189,N_3672,N_4257);
or U7190 (N_7190,N_4644,N_1344);
or U7191 (N_7191,N_3588,N_4673);
and U7192 (N_7192,N_4580,N_3785);
nand U7193 (N_7193,N_671,N_3547);
nor U7194 (N_7194,N_2915,N_2084);
or U7195 (N_7195,N_2883,N_2677);
and U7196 (N_7196,N_1416,N_1599);
nor U7197 (N_7197,N_165,N_3017);
nand U7198 (N_7198,N_1589,N_1693);
nor U7199 (N_7199,N_1996,N_4742);
nand U7200 (N_7200,N_3181,N_2853);
xor U7201 (N_7201,N_4303,N_335);
nand U7202 (N_7202,N_2342,N_4744);
xor U7203 (N_7203,N_1400,N_2090);
and U7204 (N_7204,N_1317,N_563);
and U7205 (N_7205,N_2204,N_2970);
and U7206 (N_7206,N_4879,N_1427);
nor U7207 (N_7207,N_923,N_3431);
nor U7208 (N_7208,N_1204,N_2066);
and U7209 (N_7209,N_2175,N_2190);
nand U7210 (N_7210,N_28,N_2291);
nor U7211 (N_7211,N_542,N_2301);
nand U7212 (N_7212,N_517,N_1995);
nand U7213 (N_7213,N_3421,N_4072);
or U7214 (N_7214,N_3084,N_797);
nor U7215 (N_7215,N_906,N_3939);
and U7216 (N_7216,N_451,N_1528);
nor U7217 (N_7217,N_4206,N_2589);
or U7218 (N_7218,N_182,N_2737);
or U7219 (N_7219,N_432,N_2717);
or U7220 (N_7220,N_4648,N_3418);
nand U7221 (N_7221,N_4970,N_3769);
or U7222 (N_7222,N_646,N_2905);
and U7223 (N_7223,N_2490,N_4600);
nor U7224 (N_7224,N_75,N_2445);
nand U7225 (N_7225,N_4523,N_3186);
and U7226 (N_7226,N_914,N_1985);
xor U7227 (N_7227,N_3263,N_1328);
nor U7228 (N_7228,N_4347,N_4270);
or U7229 (N_7229,N_4568,N_4629);
xor U7230 (N_7230,N_2374,N_4556);
and U7231 (N_7231,N_4933,N_1558);
or U7232 (N_7232,N_2528,N_1099);
and U7233 (N_7233,N_4346,N_4908);
xnor U7234 (N_7234,N_2453,N_4831);
nor U7235 (N_7235,N_1945,N_845);
nor U7236 (N_7236,N_4524,N_4221);
and U7237 (N_7237,N_3686,N_2985);
or U7238 (N_7238,N_1210,N_2198);
and U7239 (N_7239,N_780,N_1726);
nand U7240 (N_7240,N_1812,N_919);
or U7241 (N_7241,N_3826,N_4657);
xor U7242 (N_7242,N_2647,N_353);
or U7243 (N_7243,N_2280,N_2448);
or U7244 (N_7244,N_4542,N_38);
nand U7245 (N_7245,N_1748,N_284);
nand U7246 (N_7246,N_1896,N_903);
or U7247 (N_7247,N_4953,N_3198);
or U7248 (N_7248,N_4249,N_4266);
nor U7249 (N_7249,N_4999,N_4735);
nor U7250 (N_7250,N_60,N_4439);
nor U7251 (N_7251,N_4472,N_3677);
nand U7252 (N_7252,N_598,N_1136);
nand U7253 (N_7253,N_2603,N_393);
xnor U7254 (N_7254,N_2500,N_19);
or U7255 (N_7255,N_613,N_325);
nand U7256 (N_7256,N_3302,N_2359);
nand U7257 (N_7257,N_2888,N_1476);
nor U7258 (N_7258,N_4935,N_1803);
or U7259 (N_7259,N_565,N_608);
nor U7260 (N_7260,N_2593,N_4922);
nand U7261 (N_7261,N_3334,N_88);
xor U7262 (N_7262,N_2382,N_601);
nand U7263 (N_7263,N_1534,N_2012);
and U7264 (N_7264,N_3189,N_2956);
nor U7265 (N_7265,N_2924,N_4955);
or U7266 (N_7266,N_1386,N_2671);
nor U7267 (N_7267,N_1059,N_2989);
and U7268 (N_7268,N_190,N_3494);
nor U7269 (N_7269,N_1668,N_1116);
xnor U7270 (N_7270,N_1615,N_467);
or U7271 (N_7271,N_206,N_1275);
or U7272 (N_7272,N_4435,N_1687);
or U7273 (N_7273,N_2741,N_4444);
nand U7274 (N_7274,N_1147,N_3467);
and U7275 (N_7275,N_1407,N_1690);
and U7276 (N_7276,N_688,N_403);
and U7277 (N_7277,N_2420,N_1235);
and U7278 (N_7278,N_2674,N_3136);
or U7279 (N_7279,N_4994,N_2103);
xor U7280 (N_7280,N_1000,N_446);
or U7281 (N_7281,N_103,N_1154);
nor U7282 (N_7282,N_2966,N_1481);
or U7283 (N_7283,N_630,N_213);
or U7284 (N_7284,N_4566,N_1525);
nand U7285 (N_7285,N_4607,N_2470);
nor U7286 (N_7286,N_4889,N_167);
nor U7287 (N_7287,N_3443,N_40);
or U7288 (N_7288,N_3361,N_4254);
nor U7289 (N_7289,N_338,N_1603);
and U7290 (N_7290,N_894,N_3784);
xor U7291 (N_7291,N_2865,N_700);
and U7292 (N_7292,N_3061,N_998);
or U7293 (N_7293,N_759,N_113);
and U7294 (N_7294,N_3150,N_1365);
or U7295 (N_7295,N_4116,N_4944);
nor U7296 (N_7296,N_2176,N_4665);
nor U7297 (N_7297,N_1320,N_739);
and U7298 (N_7298,N_3016,N_2334);
and U7299 (N_7299,N_3758,N_2096);
or U7300 (N_7300,N_815,N_4156);
nor U7301 (N_7301,N_3684,N_1931);
nor U7302 (N_7302,N_1882,N_3444);
nand U7303 (N_7303,N_369,N_4885);
and U7304 (N_7304,N_2637,N_1886);
and U7305 (N_7305,N_2840,N_3033);
nand U7306 (N_7306,N_1411,N_347);
nand U7307 (N_7307,N_934,N_588);
nor U7308 (N_7308,N_3882,N_1122);
xnor U7309 (N_7309,N_3459,N_3916);
and U7310 (N_7310,N_4279,N_4022);
nand U7311 (N_7311,N_3238,N_2780);
nor U7312 (N_7312,N_4223,N_610);
and U7313 (N_7313,N_3388,N_4053);
xnor U7314 (N_7314,N_2893,N_4705);
nor U7315 (N_7315,N_4723,N_3656);
nand U7316 (N_7316,N_2725,N_2532);
and U7317 (N_7317,N_4448,N_4103);
nand U7318 (N_7318,N_1195,N_4489);
nor U7319 (N_7319,N_2358,N_4109);
nand U7320 (N_7320,N_2680,N_817);
nand U7321 (N_7321,N_3947,N_905);
nor U7322 (N_7322,N_2705,N_22);
nand U7323 (N_7323,N_1780,N_3910);
nor U7324 (N_7324,N_4000,N_4881);
xor U7325 (N_7325,N_13,N_571);
xnor U7326 (N_7326,N_3610,N_3869);
nand U7327 (N_7327,N_3424,N_1343);
and U7328 (N_7328,N_862,N_1013);
nor U7329 (N_7329,N_1155,N_2443);
and U7330 (N_7330,N_2688,N_3955);
and U7331 (N_7331,N_2465,N_3425);
xor U7332 (N_7332,N_2494,N_1710);
nand U7333 (N_7333,N_810,N_4784);
nor U7334 (N_7334,N_4978,N_1363);
xor U7335 (N_7335,N_3026,N_4442);
and U7336 (N_7336,N_3549,N_2094);
and U7337 (N_7337,N_4260,N_626);
nor U7338 (N_7338,N_3269,N_2395);
or U7339 (N_7339,N_2811,N_3089);
or U7340 (N_7340,N_1692,N_2804);
and U7341 (N_7341,N_4826,N_3582);
nand U7342 (N_7342,N_4794,N_406);
nand U7343 (N_7343,N_4154,N_1032);
or U7344 (N_7344,N_3765,N_2792);
nand U7345 (N_7345,N_931,N_4913);
xnor U7346 (N_7346,N_3038,N_1894);
nor U7347 (N_7347,N_2184,N_126);
nand U7348 (N_7348,N_395,N_1619);
nor U7349 (N_7349,N_1260,N_159);
and U7350 (N_7350,N_1679,N_4041);
nand U7351 (N_7351,N_1232,N_3054);
and U7352 (N_7352,N_1902,N_2079);
xor U7353 (N_7353,N_4486,N_2080);
nand U7354 (N_7354,N_4535,N_2136);
or U7355 (N_7355,N_2170,N_3543);
xnor U7356 (N_7356,N_4932,N_814);
nand U7357 (N_7357,N_2119,N_4847);
and U7358 (N_7358,N_1975,N_625);
xnor U7359 (N_7359,N_1752,N_4062);
or U7360 (N_7360,N_4182,N_4832);
nand U7361 (N_7361,N_1970,N_1561);
nand U7362 (N_7362,N_2651,N_4118);
or U7363 (N_7363,N_595,N_92);
nor U7364 (N_7364,N_1321,N_2591);
or U7365 (N_7365,N_226,N_1797);
and U7366 (N_7366,N_480,N_566);
or U7367 (N_7367,N_1089,N_838);
nand U7368 (N_7368,N_2278,N_770);
and U7369 (N_7369,N_326,N_3998);
nand U7370 (N_7370,N_1250,N_2285);
or U7371 (N_7371,N_4858,N_1180);
nor U7372 (N_7372,N_2816,N_4141);
or U7373 (N_7373,N_742,N_879);
or U7374 (N_7374,N_643,N_2148);
and U7375 (N_7375,N_1093,N_2946);
nand U7376 (N_7376,N_2243,N_3727);
nand U7377 (N_7377,N_754,N_2551);
nor U7378 (N_7378,N_1377,N_1864);
and U7379 (N_7379,N_582,N_1048);
nand U7380 (N_7380,N_1079,N_3191);
nand U7381 (N_7381,N_2142,N_3004);
and U7382 (N_7382,N_2548,N_1508);
nor U7383 (N_7383,N_2323,N_950);
xor U7384 (N_7384,N_394,N_240);
nor U7385 (N_7385,N_3092,N_1912);
nor U7386 (N_7386,N_94,N_3457);
nor U7387 (N_7387,N_1362,N_3013);
nand U7388 (N_7388,N_2955,N_4884);
nor U7389 (N_7389,N_4441,N_605);
and U7390 (N_7390,N_4446,N_342);
or U7391 (N_7391,N_2684,N_1259);
and U7392 (N_7392,N_995,N_3229);
nor U7393 (N_7393,N_3399,N_2829);
nand U7394 (N_7394,N_44,N_1140);
nand U7395 (N_7395,N_976,N_2052);
nor U7396 (N_7396,N_735,N_3843);
nand U7397 (N_7397,N_2592,N_160);
nor U7398 (N_7398,N_855,N_4653);
nand U7399 (N_7399,N_577,N_2258);
nor U7400 (N_7400,N_3304,N_1157);
nand U7401 (N_7401,N_1782,N_2886);
xor U7402 (N_7402,N_4453,N_3615);
and U7403 (N_7403,N_2703,N_1505);
or U7404 (N_7404,N_896,N_2361);
or U7405 (N_7405,N_822,N_4517);
nor U7406 (N_7406,N_3228,N_4528);
nor U7407 (N_7407,N_4763,N_2858);
nand U7408 (N_7408,N_859,N_3260);
nor U7409 (N_7409,N_354,N_3528);
nand U7410 (N_7410,N_2539,N_1440);
nor U7411 (N_7411,N_3936,N_1049);
xor U7412 (N_7412,N_3917,N_2484);
nand U7413 (N_7413,N_3036,N_3144);
nand U7414 (N_7414,N_286,N_154);
nor U7415 (N_7415,N_2580,N_2279);
and U7416 (N_7416,N_3475,N_2862);
and U7417 (N_7417,N_941,N_4274);
nand U7418 (N_7418,N_3460,N_319);
xor U7419 (N_7419,N_4467,N_3042);
nor U7420 (N_7420,N_1011,N_3138);
and U7421 (N_7421,N_2708,N_3527);
nand U7422 (N_7422,N_4682,N_2376);
and U7423 (N_7423,N_2907,N_1889);
nand U7424 (N_7424,N_2690,N_1167);
and U7425 (N_7425,N_2315,N_4132);
nand U7426 (N_7426,N_1130,N_2527);
nand U7427 (N_7427,N_1312,N_3696);
and U7428 (N_7428,N_4926,N_1051);
nand U7429 (N_7429,N_3874,N_4821);
nor U7430 (N_7430,N_4098,N_4793);
nand U7431 (N_7431,N_2288,N_4280);
nand U7432 (N_7432,N_788,N_1683);
nand U7433 (N_7433,N_2806,N_4749);
and U7434 (N_7434,N_2238,N_2921);
and U7435 (N_7435,N_4769,N_4786);
nand U7436 (N_7436,N_2339,N_4026);
and U7437 (N_7437,N_3342,N_4685);
nor U7438 (N_7438,N_2874,N_55);
or U7439 (N_7439,N_1105,N_1225);
nor U7440 (N_7440,N_4002,N_4016);
xor U7441 (N_7441,N_3182,N_1839);
nand U7442 (N_7442,N_34,N_4552);
xor U7443 (N_7443,N_3559,N_2950);
xor U7444 (N_7444,N_2178,N_2468);
nand U7445 (N_7445,N_966,N_1352);
or U7446 (N_7446,N_3816,N_410);
nand U7447 (N_7447,N_874,N_2210);
nand U7448 (N_7448,N_4649,N_3497);
and U7449 (N_7449,N_2984,N_1345);
xor U7450 (N_7450,N_3134,N_691);
or U7451 (N_7451,N_3611,N_244);
nand U7452 (N_7452,N_3209,N_4755);
nor U7453 (N_7453,N_4521,N_2081);
or U7454 (N_7454,N_3500,N_3669);
or U7455 (N_7455,N_1885,N_3071);
or U7456 (N_7456,N_4012,N_96);
nand U7457 (N_7457,N_3196,N_1869);
nand U7458 (N_7458,N_4559,N_3504);
or U7459 (N_7459,N_4342,N_3650);
or U7460 (N_7460,N_3300,N_1562);
xor U7461 (N_7461,N_1814,N_3167);
or U7462 (N_7462,N_1728,N_3385);
nor U7463 (N_7463,N_4406,N_561);
nor U7464 (N_7464,N_4285,N_3455);
nand U7465 (N_7465,N_4151,N_2071);
or U7466 (N_7466,N_370,N_3711);
and U7467 (N_7467,N_3965,N_4365);
or U7468 (N_7468,N_2569,N_205);
nor U7469 (N_7469,N_2246,N_3236);
nand U7470 (N_7470,N_1551,N_2002);
and U7471 (N_7471,N_3899,N_1291);
or U7472 (N_7472,N_779,N_2824);
nor U7473 (N_7473,N_3332,N_4706);
nor U7474 (N_7474,N_4457,N_2357);
nor U7475 (N_7475,N_125,N_1575);
and U7476 (N_7476,N_3353,N_2586);
or U7477 (N_7477,N_1621,N_4327);
nand U7478 (N_7478,N_3551,N_4115);
or U7479 (N_7479,N_782,N_1205);
xnor U7480 (N_7480,N_1459,N_3404);
and U7481 (N_7481,N_1319,N_596);
nor U7482 (N_7482,N_487,N_3616);
and U7483 (N_7483,N_3833,N_4263);
and U7484 (N_7484,N_580,N_3720);
nor U7485 (N_7485,N_717,N_694);
xnor U7486 (N_7486,N_1053,N_3788);
xnor U7487 (N_7487,N_293,N_4759);
and U7488 (N_7488,N_2281,N_2133);
and U7489 (N_7489,N_4654,N_2844);
nand U7490 (N_7490,N_344,N_908);
nor U7491 (N_7491,N_2379,N_1311);
or U7492 (N_7492,N_4998,N_3950);
and U7493 (N_7493,N_155,N_4503);
and U7494 (N_7494,N_3511,N_4952);
nand U7495 (N_7495,N_1008,N_2986);
or U7496 (N_7496,N_3258,N_2932);
nand U7497 (N_7497,N_4958,N_435);
or U7498 (N_7498,N_3283,N_1572);
nor U7499 (N_7499,N_415,N_1189);
xnor U7500 (N_7500,N_2650,N_1524);
nand U7501 (N_7501,N_585,N_99);
or U7502 (N_7502,N_1364,N_4654);
nand U7503 (N_7503,N_4446,N_3941);
and U7504 (N_7504,N_859,N_3439);
xnor U7505 (N_7505,N_822,N_2681);
or U7506 (N_7506,N_24,N_1156);
xor U7507 (N_7507,N_203,N_4742);
or U7508 (N_7508,N_4788,N_4296);
or U7509 (N_7509,N_3497,N_1892);
nand U7510 (N_7510,N_3066,N_4920);
and U7511 (N_7511,N_4279,N_2683);
or U7512 (N_7512,N_3751,N_667);
and U7513 (N_7513,N_3598,N_237);
nand U7514 (N_7514,N_4607,N_2851);
or U7515 (N_7515,N_2163,N_490);
xor U7516 (N_7516,N_4463,N_3825);
nor U7517 (N_7517,N_1085,N_1210);
xnor U7518 (N_7518,N_401,N_4349);
nand U7519 (N_7519,N_3978,N_2883);
or U7520 (N_7520,N_3843,N_3413);
xnor U7521 (N_7521,N_3226,N_4251);
and U7522 (N_7522,N_4740,N_1871);
nand U7523 (N_7523,N_4411,N_521);
or U7524 (N_7524,N_2881,N_1270);
nor U7525 (N_7525,N_2968,N_3899);
nand U7526 (N_7526,N_1835,N_4516);
nand U7527 (N_7527,N_1497,N_1500);
or U7528 (N_7528,N_1875,N_3547);
nor U7529 (N_7529,N_1885,N_3277);
xor U7530 (N_7530,N_1961,N_3167);
nor U7531 (N_7531,N_4250,N_4952);
or U7532 (N_7532,N_253,N_2751);
nor U7533 (N_7533,N_3587,N_1274);
nand U7534 (N_7534,N_758,N_2037);
nor U7535 (N_7535,N_2057,N_3909);
and U7536 (N_7536,N_3257,N_1306);
nor U7537 (N_7537,N_2265,N_2917);
nor U7538 (N_7538,N_1956,N_1279);
nor U7539 (N_7539,N_1978,N_4796);
nand U7540 (N_7540,N_3606,N_1587);
nor U7541 (N_7541,N_1489,N_462);
and U7542 (N_7542,N_4412,N_3610);
nand U7543 (N_7543,N_4063,N_2530);
nor U7544 (N_7544,N_581,N_3422);
nand U7545 (N_7545,N_3981,N_3143);
nand U7546 (N_7546,N_382,N_592);
or U7547 (N_7547,N_2599,N_4997);
and U7548 (N_7548,N_1059,N_3393);
nand U7549 (N_7549,N_4050,N_4024);
nand U7550 (N_7550,N_4947,N_1688);
nand U7551 (N_7551,N_3917,N_4549);
and U7552 (N_7552,N_2659,N_2771);
or U7553 (N_7553,N_245,N_3646);
nor U7554 (N_7554,N_702,N_225);
and U7555 (N_7555,N_2713,N_2205);
nand U7556 (N_7556,N_3343,N_4019);
and U7557 (N_7557,N_46,N_2569);
or U7558 (N_7558,N_988,N_577);
nand U7559 (N_7559,N_4783,N_1619);
or U7560 (N_7560,N_2967,N_1808);
and U7561 (N_7561,N_4547,N_1852);
nand U7562 (N_7562,N_4232,N_1928);
nand U7563 (N_7563,N_3093,N_4222);
and U7564 (N_7564,N_3598,N_4570);
and U7565 (N_7565,N_3846,N_4622);
nor U7566 (N_7566,N_448,N_1026);
nor U7567 (N_7567,N_600,N_4617);
nor U7568 (N_7568,N_3177,N_4546);
and U7569 (N_7569,N_3173,N_1515);
nor U7570 (N_7570,N_4472,N_1151);
and U7571 (N_7571,N_2440,N_65);
or U7572 (N_7572,N_2026,N_4684);
and U7573 (N_7573,N_904,N_4660);
and U7574 (N_7574,N_644,N_3551);
and U7575 (N_7575,N_3444,N_3356);
or U7576 (N_7576,N_1502,N_2315);
and U7577 (N_7577,N_903,N_1299);
nor U7578 (N_7578,N_2181,N_1306);
nand U7579 (N_7579,N_2901,N_1388);
or U7580 (N_7580,N_547,N_2585);
nand U7581 (N_7581,N_688,N_4111);
nor U7582 (N_7582,N_3485,N_4030);
or U7583 (N_7583,N_4501,N_2538);
nor U7584 (N_7584,N_2578,N_1063);
and U7585 (N_7585,N_4967,N_4386);
nand U7586 (N_7586,N_1229,N_4833);
nand U7587 (N_7587,N_4742,N_2507);
nor U7588 (N_7588,N_4357,N_4773);
and U7589 (N_7589,N_3679,N_2477);
nand U7590 (N_7590,N_576,N_3298);
and U7591 (N_7591,N_4821,N_150);
nor U7592 (N_7592,N_2126,N_658);
nor U7593 (N_7593,N_555,N_1013);
nand U7594 (N_7594,N_517,N_1244);
and U7595 (N_7595,N_2833,N_2875);
or U7596 (N_7596,N_3631,N_1913);
nor U7597 (N_7597,N_1264,N_781);
xnor U7598 (N_7598,N_4141,N_3794);
or U7599 (N_7599,N_4041,N_2943);
nand U7600 (N_7600,N_4198,N_4589);
nand U7601 (N_7601,N_3129,N_488);
and U7602 (N_7602,N_2193,N_2185);
or U7603 (N_7603,N_3664,N_850);
and U7604 (N_7604,N_4068,N_2770);
nor U7605 (N_7605,N_3626,N_3642);
and U7606 (N_7606,N_44,N_619);
or U7607 (N_7607,N_4728,N_4727);
or U7608 (N_7608,N_3586,N_1378);
or U7609 (N_7609,N_975,N_4802);
nor U7610 (N_7610,N_1521,N_2594);
nand U7611 (N_7611,N_2350,N_1960);
nor U7612 (N_7612,N_1489,N_3621);
nand U7613 (N_7613,N_3177,N_1953);
or U7614 (N_7614,N_56,N_86);
nor U7615 (N_7615,N_4978,N_451);
nor U7616 (N_7616,N_2126,N_2675);
and U7617 (N_7617,N_761,N_4791);
and U7618 (N_7618,N_2537,N_1516);
or U7619 (N_7619,N_2039,N_951);
nand U7620 (N_7620,N_4552,N_1358);
xnor U7621 (N_7621,N_2006,N_4774);
nor U7622 (N_7622,N_2752,N_3511);
nor U7623 (N_7623,N_410,N_3386);
nand U7624 (N_7624,N_330,N_3375);
and U7625 (N_7625,N_1942,N_1974);
nand U7626 (N_7626,N_1647,N_3661);
and U7627 (N_7627,N_1329,N_3213);
nor U7628 (N_7628,N_2743,N_1012);
nand U7629 (N_7629,N_1498,N_4611);
and U7630 (N_7630,N_2951,N_945);
and U7631 (N_7631,N_3775,N_2432);
or U7632 (N_7632,N_1205,N_297);
or U7633 (N_7633,N_1474,N_1638);
nor U7634 (N_7634,N_1991,N_3787);
nand U7635 (N_7635,N_749,N_2329);
nand U7636 (N_7636,N_4840,N_1379);
nor U7637 (N_7637,N_2108,N_907);
nand U7638 (N_7638,N_3141,N_3719);
or U7639 (N_7639,N_705,N_1659);
or U7640 (N_7640,N_4210,N_2474);
nor U7641 (N_7641,N_1540,N_811);
and U7642 (N_7642,N_4122,N_4125);
and U7643 (N_7643,N_819,N_4567);
or U7644 (N_7644,N_4932,N_4961);
or U7645 (N_7645,N_677,N_731);
nor U7646 (N_7646,N_2603,N_4088);
and U7647 (N_7647,N_1561,N_3971);
nand U7648 (N_7648,N_1261,N_4189);
and U7649 (N_7649,N_3232,N_2312);
nor U7650 (N_7650,N_1376,N_1400);
nor U7651 (N_7651,N_690,N_1019);
or U7652 (N_7652,N_4823,N_1678);
and U7653 (N_7653,N_1751,N_1719);
nor U7654 (N_7654,N_3391,N_2746);
and U7655 (N_7655,N_1831,N_3031);
nor U7656 (N_7656,N_529,N_3012);
or U7657 (N_7657,N_3872,N_4941);
nand U7658 (N_7658,N_4725,N_3986);
nor U7659 (N_7659,N_4801,N_419);
and U7660 (N_7660,N_4041,N_487);
nand U7661 (N_7661,N_3834,N_3116);
nor U7662 (N_7662,N_2904,N_348);
nand U7663 (N_7663,N_1254,N_1140);
nand U7664 (N_7664,N_1812,N_529);
or U7665 (N_7665,N_2513,N_867);
and U7666 (N_7666,N_4596,N_2236);
and U7667 (N_7667,N_4911,N_522);
and U7668 (N_7668,N_2727,N_3995);
and U7669 (N_7669,N_2574,N_1415);
nor U7670 (N_7670,N_725,N_456);
or U7671 (N_7671,N_2872,N_4995);
and U7672 (N_7672,N_2156,N_2178);
and U7673 (N_7673,N_4823,N_159);
and U7674 (N_7674,N_2166,N_2956);
nand U7675 (N_7675,N_3074,N_521);
or U7676 (N_7676,N_4510,N_177);
or U7677 (N_7677,N_1785,N_3500);
and U7678 (N_7678,N_473,N_2428);
or U7679 (N_7679,N_3898,N_2846);
nand U7680 (N_7680,N_1151,N_1389);
nor U7681 (N_7681,N_2652,N_3324);
nor U7682 (N_7682,N_4090,N_4830);
xnor U7683 (N_7683,N_4438,N_284);
nor U7684 (N_7684,N_2073,N_1992);
nor U7685 (N_7685,N_2581,N_3218);
nor U7686 (N_7686,N_1604,N_2244);
xor U7687 (N_7687,N_2852,N_2788);
and U7688 (N_7688,N_2975,N_4675);
or U7689 (N_7689,N_138,N_1676);
or U7690 (N_7690,N_2019,N_3217);
and U7691 (N_7691,N_1416,N_2111);
or U7692 (N_7692,N_4326,N_3653);
or U7693 (N_7693,N_2398,N_56);
nand U7694 (N_7694,N_2790,N_3621);
nor U7695 (N_7695,N_2938,N_4534);
and U7696 (N_7696,N_466,N_4999);
nand U7697 (N_7697,N_189,N_1376);
or U7698 (N_7698,N_2803,N_2273);
and U7699 (N_7699,N_4468,N_4630);
or U7700 (N_7700,N_1172,N_1960);
nor U7701 (N_7701,N_1396,N_4257);
and U7702 (N_7702,N_3141,N_4925);
nand U7703 (N_7703,N_3698,N_638);
and U7704 (N_7704,N_2008,N_1911);
and U7705 (N_7705,N_1280,N_2619);
nand U7706 (N_7706,N_138,N_3878);
nor U7707 (N_7707,N_1847,N_1801);
or U7708 (N_7708,N_3506,N_285);
nand U7709 (N_7709,N_1704,N_4125);
xnor U7710 (N_7710,N_4676,N_3415);
or U7711 (N_7711,N_2130,N_1907);
nor U7712 (N_7712,N_1282,N_712);
nand U7713 (N_7713,N_2817,N_1334);
xnor U7714 (N_7714,N_3524,N_1761);
or U7715 (N_7715,N_2868,N_1089);
xor U7716 (N_7716,N_2867,N_3824);
nor U7717 (N_7717,N_2595,N_115);
xnor U7718 (N_7718,N_2639,N_418);
nor U7719 (N_7719,N_1884,N_2658);
nand U7720 (N_7720,N_3999,N_4456);
xor U7721 (N_7721,N_3912,N_3777);
or U7722 (N_7722,N_3860,N_3599);
nand U7723 (N_7723,N_3087,N_1085);
nor U7724 (N_7724,N_1470,N_2122);
xor U7725 (N_7725,N_2912,N_1247);
or U7726 (N_7726,N_2590,N_294);
or U7727 (N_7727,N_498,N_1775);
nor U7728 (N_7728,N_2785,N_627);
nor U7729 (N_7729,N_2986,N_4675);
and U7730 (N_7730,N_3443,N_2531);
nand U7731 (N_7731,N_122,N_735);
nand U7732 (N_7732,N_127,N_92);
and U7733 (N_7733,N_4310,N_2539);
or U7734 (N_7734,N_1200,N_1401);
xnor U7735 (N_7735,N_2539,N_2225);
nor U7736 (N_7736,N_2692,N_4566);
or U7737 (N_7737,N_2224,N_330);
or U7738 (N_7738,N_1332,N_539);
nor U7739 (N_7739,N_1967,N_2175);
nand U7740 (N_7740,N_2797,N_4092);
xnor U7741 (N_7741,N_3351,N_2397);
and U7742 (N_7742,N_246,N_2648);
or U7743 (N_7743,N_4427,N_402);
nor U7744 (N_7744,N_886,N_1025);
or U7745 (N_7745,N_4514,N_512);
nor U7746 (N_7746,N_3560,N_2397);
xnor U7747 (N_7747,N_169,N_1706);
nand U7748 (N_7748,N_2075,N_1750);
and U7749 (N_7749,N_4506,N_4785);
and U7750 (N_7750,N_279,N_1956);
or U7751 (N_7751,N_2835,N_4329);
or U7752 (N_7752,N_1302,N_2906);
and U7753 (N_7753,N_4557,N_640);
or U7754 (N_7754,N_1485,N_3462);
nand U7755 (N_7755,N_159,N_1122);
or U7756 (N_7756,N_741,N_1349);
nand U7757 (N_7757,N_379,N_1257);
or U7758 (N_7758,N_607,N_68);
or U7759 (N_7759,N_4160,N_1488);
or U7760 (N_7760,N_4235,N_2150);
nor U7761 (N_7761,N_4663,N_2650);
or U7762 (N_7762,N_2043,N_3582);
and U7763 (N_7763,N_3216,N_3545);
nor U7764 (N_7764,N_577,N_1571);
nand U7765 (N_7765,N_1850,N_3793);
and U7766 (N_7766,N_3471,N_1263);
nand U7767 (N_7767,N_3149,N_4468);
or U7768 (N_7768,N_864,N_543);
nand U7769 (N_7769,N_3333,N_3519);
and U7770 (N_7770,N_4284,N_4565);
or U7771 (N_7771,N_3991,N_4461);
xnor U7772 (N_7772,N_3726,N_862);
or U7773 (N_7773,N_235,N_2528);
nand U7774 (N_7774,N_2048,N_18);
and U7775 (N_7775,N_4965,N_1949);
nor U7776 (N_7776,N_4542,N_2787);
or U7777 (N_7777,N_2596,N_2613);
nand U7778 (N_7778,N_4972,N_3304);
nor U7779 (N_7779,N_3465,N_1993);
nand U7780 (N_7780,N_2076,N_25);
and U7781 (N_7781,N_4956,N_4877);
nand U7782 (N_7782,N_3126,N_907);
or U7783 (N_7783,N_2286,N_165);
nand U7784 (N_7784,N_613,N_4165);
and U7785 (N_7785,N_4032,N_1124);
nor U7786 (N_7786,N_3449,N_3944);
or U7787 (N_7787,N_594,N_978);
xnor U7788 (N_7788,N_2183,N_932);
and U7789 (N_7789,N_4880,N_4687);
nor U7790 (N_7790,N_3033,N_1322);
xor U7791 (N_7791,N_3097,N_2920);
nor U7792 (N_7792,N_234,N_3629);
and U7793 (N_7793,N_3887,N_1435);
nand U7794 (N_7794,N_2108,N_3209);
nor U7795 (N_7795,N_1052,N_50);
nand U7796 (N_7796,N_1812,N_1243);
or U7797 (N_7797,N_446,N_3389);
nand U7798 (N_7798,N_153,N_2551);
nor U7799 (N_7799,N_1814,N_2283);
nand U7800 (N_7800,N_2663,N_4754);
nor U7801 (N_7801,N_1992,N_436);
or U7802 (N_7802,N_4990,N_632);
and U7803 (N_7803,N_198,N_3589);
xnor U7804 (N_7804,N_4240,N_4274);
nand U7805 (N_7805,N_4044,N_3317);
xnor U7806 (N_7806,N_4366,N_1847);
or U7807 (N_7807,N_3485,N_1407);
nor U7808 (N_7808,N_284,N_1303);
and U7809 (N_7809,N_2589,N_4755);
nor U7810 (N_7810,N_2093,N_4471);
or U7811 (N_7811,N_4679,N_4231);
xnor U7812 (N_7812,N_1060,N_2617);
xnor U7813 (N_7813,N_1981,N_3488);
nand U7814 (N_7814,N_2564,N_3058);
nand U7815 (N_7815,N_808,N_2392);
and U7816 (N_7816,N_4239,N_4584);
nor U7817 (N_7817,N_3807,N_4570);
nand U7818 (N_7818,N_1128,N_4187);
nor U7819 (N_7819,N_3008,N_345);
and U7820 (N_7820,N_4108,N_1087);
xor U7821 (N_7821,N_1476,N_953);
nor U7822 (N_7822,N_3615,N_69);
nand U7823 (N_7823,N_2938,N_4358);
or U7824 (N_7824,N_1992,N_1783);
xnor U7825 (N_7825,N_1963,N_1805);
and U7826 (N_7826,N_1879,N_2600);
or U7827 (N_7827,N_2811,N_2389);
nor U7828 (N_7828,N_1412,N_2952);
nor U7829 (N_7829,N_2441,N_3454);
xnor U7830 (N_7830,N_1738,N_0);
or U7831 (N_7831,N_379,N_4269);
xor U7832 (N_7832,N_805,N_769);
nor U7833 (N_7833,N_4141,N_2426);
nand U7834 (N_7834,N_540,N_3526);
nand U7835 (N_7835,N_1472,N_4121);
and U7836 (N_7836,N_1500,N_933);
nand U7837 (N_7837,N_1263,N_4776);
nor U7838 (N_7838,N_373,N_3388);
nor U7839 (N_7839,N_221,N_2869);
or U7840 (N_7840,N_334,N_4124);
or U7841 (N_7841,N_701,N_1623);
xnor U7842 (N_7842,N_3370,N_1899);
nand U7843 (N_7843,N_907,N_4779);
and U7844 (N_7844,N_1189,N_517);
nor U7845 (N_7845,N_3027,N_4459);
or U7846 (N_7846,N_3646,N_724);
nand U7847 (N_7847,N_1340,N_4597);
or U7848 (N_7848,N_4114,N_4511);
nor U7849 (N_7849,N_672,N_102);
xnor U7850 (N_7850,N_1407,N_2981);
and U7851 (N_7851,N_2570,N_2352);
and U7852 (N_7852,N_2797,N_4281);
or U7853 (N_7853,N_3622,N_3873);
or U7854 (N_7854,N_4907,N_2091);
nor U7855 (N_7855,N_3337,N_4200);
nor U7856 (N_7856,N_3268,N_4385);
nor U7857 (N_7857,N_4897,N_4166);
nand U7858 (N_7858,N_1117,N_3232);
and U7859 (N_7859,N_4825,N_3211);
nor U7860 (N_7860,N_4843,N_3549);
or U7861 (N_7861,N_4016,N_3545);
or U7862 (N_7862,N_633,N_446);
nand U7863 (N_7863,N_4270,N_3966);
or U7864 (N_7864,N_839,N_671);
xnor U7865 (N_7865,N_4931,N_1443);
nand U7866 (N_7866,N_956,N_1440);
nand U7867 (N_7867,N_1314,N_2162);
and U7868 (N_7868,N_1052,N_2048);
or U7869 (N_7869,N_4916,N_3609);
nand U7870 (N_7870,N_1590,N_4715);
or U7871 (N_7871,N_17,N_2828);
nand U7872 (N_7872,N_3285,N_1766);
and U7873 (N_7873,N_4684,N_1521);
or U7874 (N_7874,N_4598,N_591);
or U7875 (N_7875,N_4670,N_4053);
and U7876 (N_7876,N_203,N_3267);
nor U7877 (N_7877,N_2969,N_498);
nor U7878 (N_7878,N_2263,N_1843);
nand U7879 (N_7879,N_2649,N_3949);
or U7880 (N_7880,N_4180,N_2019);
nor U7881 (N_7881,N_3879,N_3397);
nand U7882 (N_7882,N_1405,N_2885);
or U7883 (N_7883,N_2836,N_402);
nor U7884 (N_7884,N_4081,N_3149);
nor U7885 (N_7885,N_239,N_2048);
or U7886 (N_7886,N_4146,N_1989);
nor U7887 (N_7887,N_904,N_3085);
nor U7888 (N_7888,N_4773,N_1259);
and U7889 (N_7889,N_2834,N_68);
and U7890 (N_7890,N_4044,N_4713);
nand U7891 (N_7891,N_3964,N_1967);
or U7892 (N_7892,N_3633,N_4782);
nand U7893 (N_7893,N_2461,N_3459);
nor U7894 (N_7894,N_338,N_1577);
and U7895 (N_7895,N_2851,N_1197);
and U7896 (N_7896,N_4806,N_4023);
or U7897 (N_7897,N_3160,N_1850);
xnor U7898 (N_7898,N_2131,N_4648);
nor U7899 (N_7899,N_4479,N_4140);
and U7900 (N_7900,N_1181,N_1001);
and U7901 (N_7901,N_3724,N_145);
nor U7902 (N_7902,N_3503,N_2876);
nor U7903 (N_7903,N_4332,N_1687);
and U7904 (N_7904,N_2248,N_885);
or U7905 (N_7905,N_2841,N_2264);
nor U7906 (N_7906,N_43,N_2398);
and U7907 (N_7907,N_2159,N_616);
and U7908 (N_7908,N_2276,N_2534);
xnor U7909 (N_7909,N_3703,N_1083);
nand U7910 (N_7910,N_1923,N_307);
or U7911 (N_7911,N_2745,N_1444);
nor U7912 (N_7912,N_2412,N_322);
xnor U7913 (N_7913,N_2641,N_742);
or U7914 (N_7914,N_2928,N_1782);
or U7915 (N_7915,N_4664,N_2538);
and U7916 (N_7916,N_4767,N_127);
nand U7917 (N_7917,N_594,N_3915);
and U7918 (N_7918,N_4586,N_1429);
nand U7919 (N_7919,N_4520,N_3457);
or U7920 (N_7920,N_527,N_487);
nand U7921 (N_7921,N_3026,N_305);
nand U7922 (N_7922,N_2938,N_880);
nand U7923 (N_7923,N_3322,N_2684);
or U7924 (N_7924,N_3008,N_281);
and U7925 (N_7925,N_3899,N_4075);
and U7926 (N_7926,N_4357,N_4947);
and U7927 (N_7927,N_908,N_4865);
or U7928 (N_7928,N_1277,N_4617);
xor U7929 (N_7929,N_331,N_1207);
nor U7930 (N_7930,N_4119,N_2547);
nand U7931 (N_7931,N_759,N_885);
nand U7932 (N_7932,N_2883,N_2674);
nor U7933 (N_7933,N_2216,N_1664);
and U7934 (N_7934,N_289,N_2675);
nor U7935 (N_7935,N_1540,N_1446);
nor U7936 (N_7936,N_2965,N_3904);
and U7937 (N_7937,N_2084,N_1090);
nor U7938 (N_7938,N_1265,N_580);
or U7939 (N_7939,N_3838,N_183);
nor U7940 (N_7940,N_4759,N_1529);
or U7941 (N_7941,N_588,N_83);
or U7942 (N_7942,N_3576,N_1706);
xor U7943 (N_7943,N_3470,N_4473);
nand U7944 (N_7944,N_2411,N_511);
and U7945 (N_7945,N_3816,N_767);
and U7946 (N_7946,N_4129,N_3618);
and U7947 (N_7947,N_4883,N_3971);
and U7948 (N_7948,N_1713,N_2124);
or U7949 (N_7949,N_1373,N_3200);
xor U7950 (N_7950,N_4571,N_2542);
nor U7951 (N_7951,N_1058,N_3734);
or U7952 (N_7952,N_4067,N_473);
nand U7953 (N_7953,N_4205,N_577);
and U7954 (N_7954,N_1350,N_3258);
nand U7955 (N_7955,N_3356,N_836);
or U7956 (N_7956,N_480,N_1739);
nand U7957 (N_7957,N_2790,N_3293);
nor U7958 (N_7958,N_1731,N_2239);
nor U7959 (N_7959,N_1644,N_4892);
nor U7960 (N_7960,N_4103,N_329);
and U7961 (N_7961,N_4914,N_4432);
and U7962 (N_7962,N_3924,N_3088);
and U7963 (N_7963,N_2547,N_697);
nor U7964 (N_7964,N_3951,N_4415);
or U7965 (N_7965,N_2055,N_218);
nand U7966 (N_7966,N_357,N_1636);
nand U7967 (N_7967,N_4924,N_4733);
and U7968 (N_7968,N_3429,N_2219);
and U7969 (N_7969,N_833,N_4424);
or U7970 (N_7970,N_2529,N_3970);
nand U7971 (N_7971,N_2100,N_3971);
and U7972 (N_7972,N_2350,N_3484);
nand U7973 (N_7973,N_1278,N_3153);
nor U7974 (N_7974,N_2317,N_4530);
or U7975 (N_7975,N_3609,N_1889);
or U7976 (N_7976,N_494,N_3578);
and U7977 (N_7977,N_1325,N_2587);
nor U7978 (N_7978,N_1933,N_1087);
and U7979 (N_7979,N_316,N_1440);
or U7980 (N_7980,N_4399,N_709);
nand U7981 (N_7981,N_1658,N_138);
or U7982 (N_7982,N_3874,N_1795);
xor U7983 (N_7983,N_2031,N_4943);
nand U7984 (N_7984,N_4580,N_1269);
nor U7985 (N_7985,N_1822,N_1245);
or U7986 (N_7986,N_2072,N_63);
or U7987 (N_7987,N_1474,N_2184);
nand U7988 (N_7988,N_1280,N_3587);
xnor U7989 (N_7989,N_4637,N_726);
nor U7990 (N_7990,N_1612,N_4120);
and U7991 (N_7991,N_1036,N_55);
nor U7992 (N_7992,N_2815,N_998);
or U7993 (N_7993,N_2441,N_2172);
and U7994 (N_7994,N_1489,N_3101);
or U7995 (N_7995,N_3482,N_350);
nor U7996 (N_7996,N_786,N_3930);
and U7997 (N_7997,N_4979,N_4642);
nand U7998 (N_7998,N_4319,N_1000);
nor U7999 (N_7999,N_4109,N_3785);
nand U8000 (N_8000,N_2580,N_751);
or U8001 (N_8001,N_4057,N_1613);
or U8002 (N_8002,N_1725,N_2687);
or U8003 (N_8003,N_1800,N_4054);
nor U8004 (N_8004,N_1457,N_239);
nand U8005 (N_8005,N_2300,N_4183);
and U8006 (N_8006,N_3587,N_631);
and U8007 (N_8007,N_376,N_4690);
and U8008 (N_8008,N_1044,N_1606);
and U8009 (N_8009,N_240,N_2451);
and U8010 (N_8010,N_4406,N_580);
and U8011 (N_8011,N_3527,N_625);
nand U8012 (N_8012,N_1690,N_1177);
or U8013 (N_8013,N_1797,N_1284);
nand U8014 (N_8014,N_3072,N_3566);
nor U8015 (N_8015,N_2522,N_1603);
and U8016 (N_8016,N_833,N_2736);
xnor U8017 (N_8017,N_3835,N_1711);
or U8018 (N_8018,N_2088,N_741);
xor U8019 (N_8019,N_1521,N_1458);
xnor U8020 (N_8020,N_2433,N_803);
nor U8021 (N_8021,N_96,N_3807);
nand U8022 (N_8022,N_3355,N_3157);
nor U8023 (N_8023,N_4686,N_2374);
and U8024 (N_8024,N_340,N_3456);
or U8025 (N_8025,N_2470,N_130);
nor U8026 (N_8026,N_3902,N_3174);
or U8027 (N_8027,N_2123,N_2009);
nand U8028 (N_8028,N_4893,N_401);
and U8029 (N_8029,N_2656,N_4625);
nand U8030 (N_8030,N_1180,N_4570);
and U8031 (N_8031,N_1458,N_2364);
nand U8032 (N_8032,N_285,N_1274);
and U8033 (N_8033,N_1591,N_3976);
xor U8034 (N_8034,N_2178,N_1537);
nand U8035 (N_8035,N_494,N_1998);
nand U8036 (N_8036,N_2308,N_4369);
xor U8037 (N_8037,N_1969,N_933);
nand U8038 (N_8038,N_4290,N_3661);
nand U8039 (N_8039,N_2593,N_4950);
and U8040 (N_8040,N_18,N_1171);
and U8041 (N_8041,N_2471,N_793);
nand U8042 (N_8042,N_748,N_2274);
or U8043 (N_8043,N_4409,N_3855);
nand U8044 (N_8044,N_2079,N_4210);
nand U8045 (N_8045,N_812,N_3827);
xnor U8046 (N_8046,N_2470,N_3507);
nand U8047 (N_8047,N_1070,N_4977);
and U8048 (N_8048,N_1804,N_329);
nand U8049 (N_8049,N_240,N_1753);
or U8050 (N_8050,N_64,N_2713);
and U8051 (N_8051,N_518,N_169);
nand U8052 (N_8052,N_4475,N_3563);
nand U8053 (N_8053,N_4414,N_1590);
and U8054 (N_8054,N_3300,N_4618);
nand U8055 (N_8055,N_490,N_752);
nor U8056 (N_8056,N_1318,N_771);
nor U8057 (N_8057,N_3002,N_3798);
or U8058 (N_8058,N_4808,N_1006);
xnor U8059 (N_8059,N_4536,N_3832);
nor U8060 (N_8060,N_2112,N_389);
nor U8061 (N_8061,N_1770,N_1216);
nand U8062 (N_8062,N_2450,N_4014);
and U8063 (N_8063,N_4781,N_776);
xnor U8064 (N_8064,N_3563,N_3465);
nor U8065 (N_8065,N_1118,N_3696);
and U8066 (N_8066,N_540,N_2727);
or U8067 (N_8067,N_1322,N_1739);
and U8068 (N_8068,N_1722,N_4264);
or U8069 (N_8069,N_1239,N_154);
and U8070 (N_8070,N_2995,N_3454);
nand U8071 (N_8071,N_1911,N_2245);
xor U8072 (N_8072,N_1276,N_1781);
and U8073 (N_8073,N_3098,N_383);
or U8074 (N_8074,N_4637,N_3677);
and U8075 (N_8075,N_4903,N_858);
or U8076 (N_8076,N_2950,N_532);
nor U8077 (N_8077,N_4014,N_699);
and U8078 (N_8078,N_4354,N_2751);
nand U8079 (N_8079,N_2283,N_2311);
or U8080 (N_8080,N_1854,N_2719);
nand U8081 (N_8081,N_78,N_2773);
and U8082 (N_8082,N_2388,N_2734);
xnor U8083 (N_8083,N_377,N_1947);
and U8084 (N_8084,N_3850,N_1868);
and U8085 (N_8085,N_2987,N_2066);
nor U8086 (N_8086,N_790,N_1514);
and U8087 (N_8087,N_2795,N_2083);
nor U8088 (N_8088,N_4383,N_2629);
xnor U8089 (N_8089,N_3939,N_4662);
nor U8090 (N_8090,N_1633,N_2155);
xor U8091 (N_8091,N_1725,N_1301);
and U8092 (N_8092,N_1325,N_1547);
or U8093 (N_8093,N_4899,N_4718);
nor U8094 (N_8094,N_2944,N_2680);
nand U8095 (N_8095,N_4781,N_3059);
nor U8096 (N_8096,N_2296,N_4233);
or U8097 (N_8097,N_2955,N_2179);
nand U8098 (N_8098,N_2001,N_4574);
nand U8099 (N_8099,N_2418,N_1669);
and U8100 (N_8100,N_544,N_4068);
and U8101 (N_8101,N_847,N_3642);
and U8102 (N_8102,N_4847,N_3218);
and U8103 (N_8103,N_3604,N_264);
nor U8104 (N_8104,N_2092,N_2683);
nor U8105 (N_8105,N_544,N_2284);
nor U8106 (N_8106,N_3842,N_2300);
nand U8107 (N_8107,N_3088,N_2972);
nor U8108 (N_8108,N_4822,N_3491);
nor U8109 (N_8109,N_1608,N_2072);
and U8110 (N_8110,N_2843,N_347);
nor U8111 (N_8111,N_3286,N_151);
nor U8112 (N_8112,N_4230,N_2299);
and U8113 (N_8113,N_504,N_1010);
or U8114 (N_8114,N_3058,N_1823);
and U8115 (N_8115,N_4732,N_282);
nor U8116 (N_8116,N_83,N_273);
and U8117 (N_8117,N_3165,N_349);
nor U8118 (N_8118,N_2846,N_3120);
nor U8119 (N_8119,N_4073,N_427);
and U8120 (N_8120,N_1128,N_4858);
nand U8121 (N_8121,N_1305,N_1225);
xnor U8122 (N_8122,N_4595,N_429);
or U8123 (N_8123,N_3754,N_1468);
nand U8124 (N_8124,N_4759,N_792);
xnor U8125 (N_8125,N_673,N_3555);
xnor U8126 (N_8126,N_1204,N_211);
nor U8127 (N_8127,N_511,N_2063);
or U8128 (N_8128,N_1089,N_3164);
and U8129 (N_8129,N_3760,N_1641);
nand U8130 (N_8130,N_189,N_238);
nor U8131 (N_8131,N_2065,N_2004);
nand U8132 (N_8132,N_4897,N_4272);
and U8133 (N_8133,N_1555,N_404);
and U8134 (N_8134,N_3272,N_4917);
and U8135 (N_8135,N_2720,N_1695);
nor U8136 (N_8136,N_3905,N_1297);
nand U8137 (N_8137,N_4307,N_4546);
nand U8138 (N_8138,N_1595,N_4640);
or U8139 (N_8139,N_4007,N_4850);
nand U8140 (N_8140,N_4354,N_499);
or U8141 (N_8141,N_3012,N_862);
and U8142 (N_8142,N_2438,N_3166);
and U8143 (N_8143,N_2636,N_3342);
nor U8144 (N_8144,N_3684,N_1257);
xor U8145 (N_8145,N_547,N_3935);
or U8146 (N_8146,N_4009,N_1992);
nor U8147 (N_8147,N_446,N_864);
nand U8148 (N_8148,N_4451,N_4419);
nor U8149 (N_8149,N_3390,N_2943);
nand U8150 (N_8150,N_2592,N_2168);
and U8151 (N_8151,N_2870,N_3499);
nand U8152 (N_8152,N_2697,N_3588);
xnor U8153 (N_8153,N_3162,N_4758);
nor U8154 (N_8154,N_931,N_3831);
and U8155 (N_8155,N_2472,N_2824);
xor U8156 (N_8156,N_1564,N_3260);
and U8157 (N_8157,N_2506,N_3367);
nand U8158 (N_8158,N_1938,N_160);
or U8159 (N_8159,N_1983,N_2038);
nand U8160 (N_8160,N_877,N_682);
nand U8161 (N_8161,N_4153,N_3398);
and U8162 (N_8162,N_3017,N_3355);
and U8163 (N_8163,N_500,N_1212);
or U8164 (N_8164,N_1960,N_2027);
or U8165 (N_8165,N_2691,N_976);
xor U8166 (N_8166,N_3566,N_4355);
nor U8167 (N_8167,N_889,N_2524);
xor U8168 (N_8168,N_210,N_2710);
or U8169 (N_8169,N_3138,N_53);
xnor U8170 (N_8170,N_3632,N_3139);
nor U8171 (N_8171,N_1866,N_509);
nor U8172 (N_8172,N_749,N_4172);
nand U8173 (N_8173,N_3344,N_1212);
and U8174 (N_8174,N_4417,N_126);
and U8175 (N_8175,N_2800,N_1731);
nor U8176 (N_8176,N_554,N_3822);
xor U8177 (N_8177,N_615,N_1186);
nand U8178 (N_8178,N_2310,N_1654);
or U8179 (N_8179,N_1734,N_3587);
xnor U8180 (N_8180,N_4793,N_233);
xnor U8181 (N_8181,N_4129,N_2046);
nor U8182 (N_8182,N_114,N_3127);
nand U8183 (N_8183,N_529,N_1980);
and U8184 (N_8184,N_3553,N_2630);
or U8185 (N_8185,N_1876,N_2864);
nand U8186 (N_8186,N_2615,N_804);
nand U8187 (N_8187,N_2806,N_4129);
nor U8188 (N_8188,N_2147,N_2883);
nor U8189 (N_8189,N_50,N_380);
and U8190 (N_8190,N_4107,N_161);
and U8191 (N_8191,N_2198,N_1855);
and U8192 (N_8192,N_1200,N_2647);
or U8193 (N_8193,N_3603,N_3395);
nor U8194 (N_8194,N_2832,N_929);
nand U8195 (N_8195,N_2984,N_2264);
nor U8196 (N_8196,N_1140,N_4299);
nor U8197 (N_8197,N_2467,N_1427);
nor U8198 (N_8198,N_2920,N_2206);
xor U8199 (N_8199,N_1657,N_2235);
and U8200 (N_8200,N_3860,N_170);
and U8201 (N_8201,N_4763,N_693);
nor U8202 (N_8202,N_3450,N_4067);
or U8203 (N_8203,N_4358,N_1406);
nor U8204 (N_8204,N_2732,N_688);
and U8205 (N_8205,N_463,N_649);
and U8206 (N_8206,N_1100,N_4233);
nand U8207 (N_8207,N_3863,N_2004);
nor U8208 (N_8208,N_4236,N_1015);
nand U8209 (N_8209,N_1810,N_3183);
nor U8210 (N_8210,N_4239,N_3297);
or U8211 (N_8211,N_363,N_4704);
nor U8212 (N_8212,N_775,N_961);
and U8213 (N_8213,N_4263,N_1284);
or U8214 (N_8214,N_3791,N_4336);
or U8215 (N_8215,N_2223,N_2747);
and U8216 (N_8216,N_460,N_1312);
nor U8217 (N_8217,N_4736,N_2690);
nor U8218 (N_8218,N_4672,N_889);
and U8219 (N_8219,N_411,N_1815);
or U8220 (N_8220,N_4131,N_1322);
and U8221 (N_8221,N_570,N_2034);
nand U8222 (N_8222,N_981,N_1194);
or U8223 (N_8223,N_4147,N_3944);
and U8224 (N_8224,N_20,N_406);
xor U8225 (N_8225,N_2489,N_2595);
and U8226 (N_8226,N_3481,N_4932);
and U8227 (N_8227,N_1784,N_106);
nor U8228 (N_8228,N_1112,N_1705);
nor U8229 (N_8229,N_4108,N_643);
xnor U8230 (N_8230,N_3949,N_2706);
or U8231 (N_8231,N_1450,N_2237);
or U8232 (N_8232,N_3505,N_1656);
nand U8233 (N_8233,N_136,N_908);
nor U8234 (N_8234,N_2630,N_559);
nand U8235 (N_8235,N_1350,N_4658);
and U8236 (N_8236,N_3130,N_70);
or U8237 (N_8237,N_2514,N_4710);
nand U8238 (N_8238,N_587,N_4470);
xor U8239 (N_8239,N_1019,N_2562);
and U8240 (N_8240,N_2749,N_310);
nor U8241 (N_8241,N_4315,N_4943);
nor U8242 (N_8242,N_1188,N_4258);
and U8243 (N_8243,N_2877,N_4409);
nand U8244 (N_8244,N_3171,N_4154);
nor U8245 (N_8245,N_2007,N_4329);
and U8246 (N_8246,N_2754,N_380);
and U8247 (N_8247,N_1718,N_4820);
nand U8248 (N_8248,N_4832,N_4402);
xor U8249 (N_8249,N_4292,N_748);
and U8250 (N_8250,N_1322,N_3709);
and U8251 (N_8251,N_3505,N_118);
and U8252 (N_8252,N_1091,N_4876);
nor U8253 (N_8253,N_3276,N_4607);
and U8254 (N_8254,N_3889,N_2713);
and U8255 (N_8255,N_3152,N_4261);
nor U8256 (N_8256,N_1238,N_3798);
or U8257 (N_8257,N_2711,N_3783);
nand U8258 (N_8258,N_2935,N_4891);
nor U8259 (N_8259,N_5,N_1777);
nor U8260 (N_8260,N_2853,N_3826);
or U8261 (N_8261,N_4825,N_4085);
nor U8262 (N_8262,N_920,N_731);
xnor U8263 (N_8263,N_4276,N_3468);
xnor U8264 (N_8264,N_1405,N_4289);
or U8265 (N_8265,N_4196,N_3589);
or U8266 (N_8266,N_4541,N_2648);
nand U8267 (N_8267,N_3125,N_4375);
nand U8268 (N_8268,N_3562,N_278);
nor U8269 (N_8269,N_559,N_4675);
nor U8270 (N_8270,N_348,N_763);
nor U8271 (N_8271,N_2205,N_1977);
or U8272 (N_8272,N_4684,N_4675);
or U8273 (N_8273,N_350,N_3925);
nand U8274 (N_8274,N_1455,N_2591);
nand U8275 (N_8275,N_1198,N_694);
and U8276 (N_8276,N_1755,N_2228);
nor U8277 (N_8277,N_2878,N_769);
or U8278 (N_8278,N_4324,N_2093);
and U8279 (N_8279,N_4540,N_72);
nand U8280 (N_8280,N_4002,N_4222);
nand U8281 (N_8281,N_2728,N_1509);
and U8282 (N_8282,N_244,N_2149);
nor U8283 (N_8283,N_993,N_3987);
and U8284 (N_8284,N_3426,N_4344);
or U8285 (N_8285,N_2822,N_1567);
and U8286 (N_8286,N_1477,N_133);
and U8287 (N_8287,N_2296,N_936);
or U8288 (N_8288,N_2428,N_2463);
and U8289 (N_8289,N_4474,N_4041);
and U8290 (N_8290,N_628,N_2424);
nor U8291 (N_8291,N_479,N_2363);
xnor U8292 (N_8292,N_3033,N_4807);
and U8293 (N_8293,N_398,N_2884);
or U8294 (N_8294,N_567,N_4878);
or U8295 (N_8295,N_1084,N_1895);
nand U8296 (N_8296,N_4357,N_4592);
nor U8297 (N_8297,N_1964,N_20);
and U8298 (N_8298,N_4666,N_4088);
nor U8299 (N_8299,N_3323,N_3894);
or U8300 (N_8300,N_1190,N_4796);
and U8301 (N_8301,N_694,N_4027);
nand U8302 (N_8302,N_1172,N_1921);
and U8303 (N_8303,N_1047,N_4928);
and U8304 (N_8304,N_3949,N_4029);
and U8305 (N_8305,N_664,N_2352);
nor U8306 (N_8306,N_1151,N_510);
xor U8307 (N_8307,N_3690,N_4912);
nand U8308 (N_8308,N_2714,N_2420);
or U8309 (N_8309,N_1717,N_4584);
nor U8310 (N_8310,N_1794,N_4477);
nand U8311 (N_8311,N_3102,N_3191);
nand U8312 (N_8312,N_2915,N_923);
nand U8313 (N_8313,N_4053,N_1048);
and U8314 (N_8314,N_1605,N_4307);
nand U8315 (N_8315,N_1465,N_1623);
nor U8316 (N_8316,N_282,N_3447);
and U8317 (N_8317,N_1816,N_2915);
nor U8318 (N_8318,N_4657,N_2485);
and U8319 (N_8319,N_4609,N_3558);
or U8320 (N_8320,N_2765,N_1695);
and U8321 (N_8321,N_3245,N_4097);
and U8322 (N_8322,N_1677,N_4570);
nor U8323 (N_8323,N_3329,N_4431);
nand U8324 (N_8324,N_1952,N_3641);
and U8325 (N_8325,N_1572,N_3098);
or U8326 (N_8326,N_3004,N_36);
nor U8327 (N_8327,N_4493,N_1184);
nor U8328 (N_8328,N_453,N_2831);
nand U8329 (N_8329,N_355,N_1105);
nand U8330 (N_8330,N_231,N_2712);
nand U8331 (N_8331,N_2096,N_2242);
xnor U8332 (N_8332,N_336,N_4814);
nand U8333 (N_8333,N_4614,N_1271);
or U8334 (N_8334,N_3780,N_2752);
nand U8335 (N_8335,N_1222,N_3474);
nand U8336 (N_8336,N_4652,N_3142);
or U8337 (N_8337,N_4947,N_1707);
nand U8338 (N_8338,N_3827,N_2311);
nand U8339 (N_8339,N_4360,N_3095);
and U8340 (N_8340,N_3778,N_2841);
nand U8341 (N_8341,N_311,N_4196);
nor U8342 (N_8342,N_3291,N_1122);
xnor U8343 (N_8343,N_643,N_1728);
xnor U8344 (N_8344,N_904,N_4129);
nand U8345 (N_8345,N_724,N_3668);
or U8346 (N_8346,N_1303,N_2553);
nand U8347 (N_8347,N_859,N_1260);
and U8348 (N_8348,N_666,N_370);
or U8349 (N_8349,N_4793,N_2234);
or U8350 (N_8350,N_318,N_2812);
or U8351 (N_8351,N_156,N_2264);
nand U8352 (N_8352,N_4123,N_3710);
nor U8353 (N_8353,N_4293,N_1113);
nor U8354 (N_8354,N_4431,N_1303);
xnor U8355 (N_8355,N_3867,N_2378);
or U8356 (N_8356,N_3333,N_3712);
and U8357 (N_8357,N_2709,N_852);
or U8358 (N_8358,N_3683,N_1007);
nand U8359 (N_8359,N_2962,N_4515);
nor U8360 (N_8360,N_4048,N_2439);
nand U8361 (N_8361,N_84,N_3045);
or U8362 (N_8362,N_4679,N_229);
nor U8363 (N_8363,N_2636,N_3078);
or U8364 (N_8364,N_4754,N_1978);
xnor U8365 (N_8365,N_2857,N_3883);
nand U8366 (N_8366,N_2045,N_194);
nor U8367 (N_8367,N_4670,N_744);
nand U8368 (N_8368,N_332,N_2905);
nand U8369 (N_8369,N_4772,N_2636);
and U8370 (N_8370,N_3814,N_4853);
or U8371 (N_8371,N_426,N_2987);
or U8372 (N_8372,N_657,N_614);
or U8373 (N_8373,N_1678,N_3189);
xnor U8374 (N_8374,N_4055,N_3231);
nand U8375 (N_8375,N_4754,N_2931);
nor U8376 (N_8376,N_3772,N_288);
or U8377 (N_8377,N_2675,N_3095);
nor U8378 (N_8378,N_103,N_1986);
nor U8379 (N_8379,N_4254,N_3009);
nand U8380 (N_8380,N_1369,N_577);
or U8381 (N_8381,N_3299,N_4622);
nand U8382 (N_8382,N_4527,N_2322);
nor U8383 (N_8383,N_4862,N_4772);
nor U8384 (N_8384,N_1964,N_391);
nand U8385 (N_8385,N_2608,N_1952);
nand U8386 (N_8386,N_3334,N_2310);
and U8387 (N_8387,N_2358,N_175);
or U8388 (N_8388,N_4962,N_3811);
xor U8389 (N_8389,N_4813,N_2249);
nor U8390 (N_8390,N_1043,N_4840);
and U8391 (N_8391,N_1540,N_1230);
nand U8392 (N_8392,N_4456,N_509);
nand U8393 (N_8393,N_1509,N_2577);
nand U8394 (N_8394,N_4987,N_4984);
or U8395 (N_8395,N_2952,N_3024);
nand U8396 (N_8396,N_4014,N_2246);
nor U8397 (N_8397,N_3033,N_870);
xnor U8398 (N_8398,N_3430,N_930);
nand U8399 (N_8399,N_2778,N_953);
and U8400 (N_8400,N_227,N_997);
and U8401 (N_8401,N_2464,N_1558);
xnor U8402 (N_8402,N_3206,N_3649);
nand U8403 (N_8403,N_451,N_4746);
nor U8404 (N_8404,N_579,N_2654);
and U8405 (N_8405,N_1014,N_4345);
nor U8406 (N_8406,N_302,N_4856);
and U8407 (N_8407,N_4489,N_3686);
and U8408 (N_8408,N_958,N_4655);
or U8409 (N_8409,N_4462,N_2717);
nand U8410 (N_8410,N_510,N_2532);
nand U8411 (N_8411,N_1118,N_3760);
nor U8412 (N_8412,N_4450,N_3801);
nand U8413 (N_8413,N_18,N_847);
and U8414 (N_8414,N_187,N_1011);
or U8415 (N_8415,N_907,N_3897);
and U8416 (N_8416,N_1103,N_969);
xor U8417 (N_8417,N_1901,N_3496);
xor U8418 (N_8418,N_1666,N_4938);
or U8419 (N_8419,N_1114,N_3379);
nor U8420 (N_8420,N_1674,N_524);
nand U8421 (N_8421,N_2182,N_357);
nand U8422 (N_8422,N_1850,N_4840);
xor U8423 (N_8423,N_4709,N_926);
or U8424 (N_8424,N_959,N_4255);
and U8425 (N_8425,N_3982,N_2350);
nand U8426 (N_8426,N_2044,N_3334);
nor U8427 (N_8427,N_3670,N_3031);
or U8428 (N_8428,N_613,N_359);
nand U8429 (N_8429,N_2985,N_4423);
or U8430 (N_8430,N_1640,N_1511);
or U8431 (N_8431,N_2387,N_2983);
nand U8432 (N_8432,N_2795,N_1697);
nor U8433 (N_8433,N_3427,N_988);
or U8434 (N_8434,N_2950,N_3087);
or U8435 (N_8435,N_3833,N_3463);
nor U8436 (N_8436,N_1633,N_2039);
or U8437 (N_8437,N_3217,N_2177);
xor U8438 (N_8438,N_1311,N_3270);
and U8439 (N_8439,N_2074,N_1683);
and U8440 (N_8440,N_1219,N_2176);
or U8441 (N_8441,N_3616,N_2424);
xor U8442 (N_8442,N_4743,N_1559);
nand U8443 (N_8443,N_50,N_835);
nand U8444 (N_8444,N_492,N_2652);
or U8445 (N_8445,N_4821,N_2457);
or U8446 (N_8446,N_2519,N_1235);
nor U8447 (N_8447,N_2986,N_4105);
nor U8448 (N_8448,N_4245,N_379);
xor U8449 (N_8449,N_673,N_3493);
and U8450 (N_8450,N_2099,N_4619);
xnor U8451 (N_8451,N_3636,N_2090);
and U8452 (N_8452,N_3273,N_2493);
and U8453 (N_8453,N_608,N_4027);
nor U8454 (N_8454,N_4500,N_1329);
and U8455 (N_8455,N_1999,N_4826);
or U8456 (N_8456,N_1028,N_2920);
or U8457 (N_8457,N_1377,N_3437);
or U8458 (N_8458,N_887,N_4336);
or U8459 (N_8459,N_1431,N_4441);
or U8460 (N_8460,N_1333,N_4365);
and U8461 (N_8461,N_1520,N_3993);
xnor U8462 (N_8462,N_3755,N_3564);
and U8463 (N_8463,N_3458,N_1274);
nor U8464 (N_8464,N_3997,N_3290);
or U8465 (N_8465,N_2271,N_339);
xor U8466 (N_8466,N_2812,N_4173);
nor U8467 (N_8467,N_2835,N_1314);
or U8468 (N_8468,N_2411,N_2435);
and U8469 (N_8469,N_1038,N_4662);
nor U8470 (N_8470,N_1375,N_4777);
or U8471 (N_8471,N_2859,N_1467);
nor U8472 (N_8472,N_2898,N_2800);
nand U8473 (N_8473,N_2984,N_2547);
and U8474 (N_8474,N_1680,N_3102);
nand U8475 (N_8475,N_3930,N_278);
nor U8476 (N_8476,N_2115,N_1927);
or U8477 (N_8477,N_2771,N_2850);
and U8478 (N_8478,N_4035,N_3163);
or U8479 (N_8479,N_894,N_2733);
xor U8480 (N_8480,N_686,N_1182);
nor U8481 (N_8481,N_2001,N_4828);
nand U8482 (N_8482,N_2245,N_2011);
xor U8483 (N_8483,N_1978,N_4767);
nor U8484 (N_8484,N_3374,N_2482);
nand U8485 (N_8485,N_801,N_2496);
nand U8486 (N_8486,N_4195,N_4294);
nor U8487 (N_8487,N_1337,N_3065);
or U8488 (N_8488,N_2554,N_1202);
nand U8489 (N_8489,N_3651,N_1509);
and U8490 (N_8490,N_1811,N_3591);
or U8491 (N_8491,N_2731,N_1844);
and U8492 (N_8492,N_1409,N_625);
nor U8493 (N_8493,N_2439,N_2238);
and U8494 (N_8494,N_3889,N_2910);
nand U8495 (N_8495,N_3531,N_3629);
nor U8496 (N_8496,N_4128,N_753);
and U8497 (N_8497,N_2781,N_6);
nor U8498 (N_8498,N_210,N_651);
or U8499 (N_8499,N_4448,N_1726);
xor U8500 (N_8500,N_3715,N_3430);
or U8501 (N_8501,N_346,N_3024);
nand U8502 (N_8502,N_2770,N_1433);
nand U8503 (N_8503,N_3656,N_4674);
and U8504 (N_8504,N_4137,N_567);
or U8505 (N_8505,N_4380,N_2161);
and U8506 (N_8506,N_1203,N_441);
xnor U8507 (N_8507,N_4199,N_2373);
or U8508 (N_8508,N_1972,N_1322);
or U8509 (N_8509,N_2779,N_1435);
nand U8510 (N_8510,N_3211,N_4204);
nand U8511 (N_8511,N_316,N_2679);
or U8512 (N_8512,N_2064,N_3292);
or U8513 (N_8513,N_3115,N_4063);
and U8514 (N_8514,N_2506,N_3303);
and U8515 (N_8515,N_3555,N_4390);
nor U8516 (N_8516,N_4424,N_2819);
and U8517 (N_8517,N_799,N_3464);
or U8518 (N_8518,N_4802,N_472);
nor U8519 (N_8519,N_2956,N_2147);
and U8520 (N_8520,N_3978,N_4189);
or U8521 (N_8521,N_2091,N_786);
nand U8522 (N_8522,N_1586,N_2866);
nand U8523 (N_8523,N_4920,N_1084);
nand U8524 (N_8524,N_1676,N_1346);
nand U8525 (N_8525,N_172,N_755);
nand U8526 (N_8526,N_1838,N_505);
nand U8527 (N_8527,N_4076,N_605);
nor U8528 (N_8528,N_91,N_4344);
nand U8529 (N_8529,N_4338,N_3955);
nand U8530 (N_8530,N_620,N_2457);
nor U8531 (N_8531,N_4392,N_2310);
nor U8532 (N_8532,N_4361,N_3782);
nor U8533 (N_8533,N_4425,N_4703);
nor U8534 (N_8534,N_3785,N_59);
nor U8535 (N_8535,N_4780,N_889);
nand U8536 (N_8536,N_450,N_3453);
nor U8537 (N_8537,N_487,N_170);
or U8538 (N_8538,N_754,N_2708);
xor U8539 (N_8539,N_2499,N_395);
or U8540 (N_8540,N_3419,N_2581);
nor U8541 (N_8541,N_48,N_2509);
and U8542 (N_8542,N_4650,N_1488);
nor U8543 (N_8543,N_4,N_2281);
and U8544 (N_8544,N_268,N_3479);
and U8545 (N_8545,N_3562,N_410);
and U8546 (N_8546,N_3969,N_2485);
and U8547 (N_8547,N_1100,N_1923);
or U8548 (N_8548,N_3582,N_4731);
nor U8549 (N_8549,N_1958,N_2780);
and U8550 (N_8550,N_1490,N_3697);
or U8551 (N_8551,N_4313,N_3082);
nor U8552 (N_8552,N_3591,N_3985);
nand U8553 (N_8553,N_3204,N_1858);
xor U8554 (N_8554,N_4990,N_2089);
nor U8555 (N_8555,N_4422,N_3285);
or U8556 (N_8556,N_4364,N_2910);
and U8557 (N_8557,N_4430,N_4145);
or U8558 (N_8558,N_4378,N_1487);
nand U8559 (N_8559,N_4699,N_460);
or U8560 (N_8560,N_3907,N_3933);
and U8561 (N_8561,N_1893,N_1837);
nand U8562 (N_8562,N_3725,N_4911);
and U8563 (N_8563,N_4247,N_2359);
and U8564 (N_8564,N_4857,N_1574);
and U8565 (N_8565,N_977,N_2857);
and U8566 (N_8566,N_3161,N_3688);
or U8567 (N_8567,N_3770,N_3192);
xor U8568 (N_8568,N_186,N_1813);
and U8569 (N_8569,N_1635,N_2099);
or U8570 (N_8570,N_1672,N_455);
nand U8571 (N_8571,N_4299,N_2675);
or U8572 (N_8572,N_1539,N_551);
or U8573 (N_8573,N_3198,N_1093);
and U8574 (N_8574,N_984,N_524);
nand U8575 (N_8575,N_3259,N_4042);
nand U8576 (N_8576,N_3845,N_3911);
and U8577 (N_8577,N_1884,N_3540);
and U8578 (N_8578,N_902,N_4405);
nor U8579 (N_8579,N_3418,N_4442);
and U8580 (N_8580,N_97,N_1580);
or U8581 (N_8581,N_1419,N_403);
and U8582 (N_8582,N_1829,N_4595);
nand U8583 (N_8583,N_1211,N_3547);
and U8584 (N_8584,N_2199,N_1225);
and U8585 (N_8585,N_3835,N_981);
nand U8586 (N_8586,N_763,N_966);
nand U8587 (N_8587,N_233,N_2364);
nor U8588 (N_8588,N_2666,N_95);
or U8589 (N_8589,N_999,N_1680);
xnor U8590 (N_8590,N_174,N_1459);
nand U8591 (N_8591,N_3185,N_3285);
nor U8592 (N_8592,N_4174,N_1430);
or U8593 (N_8593,N_475,N_1451);
or U8594 (N_8594,N_4841,N_1907);
or U8595 (N_8595,N_3116,N_2280);
or U8596 (N_8596,N_1564,N_2425);
nor U8597 (N_8597,N_2914,N_4036);
or U8598 (N_8598,N_4877,N_2487);
nor U8599 (N_8599,N_4059,N_2153);
nand U8600 (N_8600,N_1381,N_4934);
nand U8601 (N_8601,N_4552,N_2404);
nor U8602 (N_8602,N_1495,N_2441);
nand U8603 (N_8603,N_318,N_2717);
nand U8604 (N_8604,N_2666,N_4841);
or U8605 (N_8605,N_3218,N_4546);
or U8606 (N_8606,N_3318,N_4672);
or U8607 (N_8607,N_3899,N_3260);
or U8608 (N_8608,N_4993,N_3649);
or U8609 (N_8609,N_829,N_1241);
and U8610 (N_8610,N_3781,N_1390);
nor U8611 (N_8611,N_3795,N_312);
nand U8612 (N_8612,N_969,N_3707);
nor U8613 (N_8613,N_2043,N_3986);
xnor U8614 (N_8614,N_430,N_2820);
xnor U8615 (N_8615,N_3423,N_2770);
and U8616 (N_8616,N_4820,N_4575);
nor U8617 (N_8617,N_433,N_2317);
nand U8618 (N_8618,N_815,N_1637);
and U8619 (N_8619,N_2280,N_2950);
xor U8620 (N_8620,N_1864,N_4008);
nor U8621 (N_8621,N_1089,N_4256);
or U8622 (N_8622,N_2893,N_2781);
and U8623 (N_8623,N_883,N_821);
nor U8624 (N_8624,N_374,N_1704);
xnor U8625 (N_8625,N_966,N_3386);
nand U8626 (N_8626,N_2731,N_2679);
or U8627 (N_8627,N_2802,N_4696);
and U8628 (N_8628,N_1239,N_2825);
xnor U8629 (N_8629,N_4325,N_2865);
nor U8630 (N_8630,N_4702,N_3867);
or U8631 (N_8631,N_1519,N_3809);
nand U8632 (N_8632,N_2778,N_4611);
nand U8633 (N_8633,N_130,N_674);
or U8634 (N_8634,N_1150,N_1086);
nor U8635 (N_8635,N_2482,N_2728);
nor U8636 (N_8636,N_4166,N_3429);
nand U8637 (N_8637,N_3925,N_3956);
nand U8638 (N_8638,N_166,N_2459);
nand U8639 (N_8639,N_2032,N_437);
or U8640 (N_8640,N_253,N_1693);
or U8641 (N_8641,N_496,N_1794);
or U8642 (N_8642,N_941,N_2645);
nand U8643 (N_8643,N_3009,N_1029);
or U8644 (N_8644,N_2898,N_4215);
nor U8645 (N_8645,N_2794,N_3782);
nand U8646 (N_8646,N_2329,N_4046);
and U8647 (N_8647,N_4994,N_4419);
and U8648 (N_8648,N_40,N_205);
xor U8649 (N_8649,N_1022,N_2424);
or U8650 (N_8650,N_238,N_2130);
or U8651 (N_8651,N_3045,N_1516);
nand U8652 (N_8652,N_2163,N_4510);
nor U8653 (N_8653,N_4635,N_409);
or U8654 (N_8654,N_605,N_1990);
xor U8655 (N_8655,N_3916,N_4820);
or U8656 (N_8656,N_1408,N_417);
or U8657 (N_8657,N_737,N_643);
nand U8658 (N_8658,N_4414,N_423);
and U8659 (N_8659,N_1880,N_2153);
or U8660 (N_8660,N_112,N_1408);
xor U8661 (N_8661,N_3383,N_3897);
xor U8662 (N_8662,N_3409,N_2322);
xor U8663 (N_8663,N_4876,N_3523);
or U8664 (N_8664,N_1015,N_4763);
or U8665 (N_8665,N_695,N_3861);
nand U8666 (N_8666,N_2012,N_506);
nand U8667 (N_8667,N_84,N_3379);
nand U8668 (N_8668,N_4603,N_814);
or U8669 (N_8669,N_3210,N_866);
nand U8670 (N_8670,N_491,N_3719);
and U8671 (N_8671,N_3077,N_1592);
and U8672 (N_8672,N_3339,N_2230);
nand U8673 (N_8673,N_879,N_2857);
and U8674 (N_8674,N_1507,N_2395);
and U8675 (N_8675,N_4122,N_371);
xnor U8676 (N_8676,N_2030,N_1948);
nor U8677 (N_8677,N_3929,N_989);
nor U8678 (N_8678,N_1692,N_424);
nand U8679 (N_8679,N_4438,N_2289);
and U8680 (N_8680,N_4272,N_293);
xnor U8681 (N_8681,N_1816,N_4412);
nor U8682 (N_8682,N_2054,N_437);
and U8683 (N_8683,N_4232,N_49);
or U8684 (N_8684,N_1716,N_1489);
and U8685 (N_8685,N_1198,N_4159);
and U8686 (N_8686,N_1506,N_4740);
nand U8687 (N_8687,N_1736,N_3262);
and U8688 (N_8688,N_638,N_1426);
xnor U8689 (N_8689,N_4172,N_4529);
nand U8690 (N_8690,N_27,N_2240);
and U8691 (N_8691,N_1961,N_3927);
nand U8692 (N_8692,N_3406,N_1382);
and U8693 (N_8693,N_2549,N_2687);
nor U8694 (N_8694,N_3699,N_2917);
nor U8695 (N_8695,N_1688,N_4182);
or U8696 (N_8696,N_978,N_3327);
nor U8697 (N_8697,N_2618,N_3510);
or U8698 (N_8698,N_276,N_1825);
and U8699 (N_8699,N_4083,N_2796);
or U8700 (N_8700,N_1078,N_756);
nand U8701 (N_8701,N_3965,N_2684);
and U8702 (N_8702,N_3884,N_1502);
nand U8703 (N_8703,N_1324,N_4682);
or U8704 (N_8704,N_3627,N_1921);
or U8705 (N_8705,N_2857,N_2672);
nand U8706 (N_8706,N_1018,N_1408);
nand U8707 (N_8707,N_955,N_2784);
or U8708 (N_8708,N_4619,N_2538);
xnor U8709 (N_8709,N_3215,N_2248);
nand U8710 (N_8710,N_2806,N_3047);
or U8711 (N_8711,N_44,N_1275);
nand U8712 (N_8712,N_944,N_2608);
xor U8713 (N_8713,N_321,N_747);
nand U8714 (N_8714,N_1508,N_1539);
nor U8715 (N_8715,N_2414,N_2687);
nand U8716 (N_8716,N_1299,N_1359);
or U8717 (N_8717,N_4558,N_4561);
and U8718 (N_8718,N_4753,N_3507);
and U8719 (N_8719,N_2740,N_1105);
or U8720 (N_8720,N_3856,N_3344);
and U8721 (N_8721,N_1496,N_1289);
nand U8722 (N_8722,N_1973,N_557);
or U8723 (N_8723,N_1096,N_4868);
nor U8724 (N_8724,N_1134,N_577);
xnor U8725 (N_8725,N_4135,N_4908);
nand U8726 (N_8726,N_1724,N_2436);
and U8727 (N_8727,N_2598,N_2093);
nor U8728 (N_8728,N_2014,N_2923);
nand U8729 (N_8729,N_150,N_3640);
xnor U8730 (N_8730,N_4185,N_4623);
nand U8731 (N_8731,N_4115,N_79);
nor U8732 (N_8732,N_3898,N_2519);
xor U8733 (N_8733,N_4418,N_4123);
or U8734 (N_8734,N_79,N_469);
and U8735 (N_8735,N_4358,N_2491);
nor U8736 (N_8736,N_995,N_1351);
and U8737 (N_8737,N_2395,N_2382);
nand U8738 (N_8738,N_2018,N_231);
and U8739 (N_8739,N_2182,N_2840);
or U8740 (N_8740,N_2503,N_204);
and U8741 (N_8741,N_3673,N_1845);
or U8742 (N_8742,N_2064,N_2333);
xnor U8743 (N_8743,N_2776,N_1589);
nor U8744 (N_8744,N_4703,N_4705);
or U8745 (N_8745,N_2573,N_4225);
and U8746 (N_8746,N_1478,N_2802);
or U8747 (N_8747,N_4861,N_4111);
and U8748 (N_8748,N_4221,N_3967);
or U8749 (N_8749,N_685,N_2877);
and U8750 (N_8750,N_1623,N_3042);
and U8751 (N_8751,N_3960,N_4512);
nand U8752 (N_8752,N_2804,N_329);
nand U8753 (N_8753,N_4231,N_2430);
xor U8754 (N_8754,N_1428,N_4590);
or U8755 (N_8755,N_1099,N_3416);
nor U8756 (N_8756,N_4921,N_488);
or U8757 (N_8757,N_4441,N_1899);
and U8758 (N_8758,N_2512,N_1953);
and U8759 (N_8759,N_3087,N_240);
and U8760 (N_8760,N_2117,N_1005);
and U8761 (N_8761,N_4455,N_4674);
or U8762 (N_8762,N_2150,N_2115);
nor U8763 (N_8763,N_1329,N_3563);
or U8764 (N_8764,N_4856,N_558);
nand U8765 (N_8765,N_1403,N_1750);
nor U8766 (N_8766,N_179,N_2905);
or U8767 (N_8767,N_1046,N_1633);
and U8768 (N_8768,N_2418,N_1504);
nor U8769 (N_8769,N_3239,N_3359);
and U8770 (N_8770,N_3918,N_1769);
nor U8771 (N_8771,N_4126,N_1089);
nand U8772 (N_8772,N_4102,N_4228);
or U8773 (N_8773,N_2570,N_730);
nand U8774 (N_8774,N_4907,N_3558);
nand U8775 (N_8775,N_4990,N_3262);
and U8776 (N_8776,N_2529,N_3864);
xnor U8777 (N_8777,N_2423,N_2383);
and U8778 (N_8778,N_3381,N_3900);
nor U8779 (N_8779,N_1913,N_128);
or U8780 (N_8780,N_2570,N_3);
xnor U8781 (N_8781,N_970,N_2203);
xnor U8782 (N_8782,N_4780,N_2688);
nand U8783 (N_8783,N_1632,N_784);
xor U8784 (N_8784,N_1400,N_399);
or U8785 (N_8785,N_3031,N_2035);
or U8786 (N_8786,N_636,N_1004);
and U8787 (N_8787,N_4611,N_2093);
or U8788 (N_8788,N_2791,N_2855);
nor U8789 (N_8789,N_47,N_2916);
nand U8790 (N_8790,N_3386,N_3861);
nor U8791 (N_8791,N_1508,N_2173);
and U8792 (N_8792,N_3940,N_3869);
and U8793 (N_8793,N_2940,N_3347);
and U8794 (N_8794,N_883,N_2733);
nor U8795 (N_8795,N_3711,N_204);
and U8796 (N_8796,N_726,N_4644);
or U8797 (N_8797,N_3561,N_3784);
xnor U8798 (N_8798,N_1532,N_1499);
nor U8799 (N_8799,N_1615,N_4444);
xor U8800 (N_8800,N_1072,N_1732);
nand U8801 (N_8801,N_3983,N_4121);
and U8802 (N_8802,N_3285,N_199);
xnor U8803 (N_8803,N_3528,N_1507);
xnor U8804 (N_8804,N_1215,N_2933);
nand U8805 (N_8805,N_4948,N_1068);
xnor U8806 (N_8806,N_3582,N_4678);
or U8807 (N_8807,N_3500,N_2752);
nand U8808 (N_8808,N_3112,N_3101);
nand U8809 (N_8809,N_1296,N_4044);
and U8810 (N_8810,N_3736,N_331);
nor U8811 (N_8811,N_636,N_3330);
xor U8812 (N_8812,N_1271,N_1193);
nor U8813 (N_8813,N_4570,N_1524);
and U8814 (N_8814,N_3781,N_1029);
or U8815 (N_8815,N_1883,N_4265);
and U8816 (N_8816,N_1498,N_4090);
and U8817 (N_8817,N_243,N_1799);
nor U8818 (N_8818,N_4161,N_4744);
or U8819 (N_8819,N_571,N_3984);
nand U8820 (N_8820,N_112,N_2470);
nand U8821 (N_8821,N_1269,N_9);
nand U8822 (N_8822,N_957,N_3955);
xor U8823 (N_8823,N_2641,N_758);
and U8824 (N_8824,N_2212,N_2069);
or U8825 (N_8825,N_56,N_3854);
or U8826 (N_8826,N_2566,N_2157);
nand U8827 (N_8827,N_946,N_741);
nand U8828 (N_8828,N_1855,N_3816);
or U8829 (N_8829,N_581,N_4161);
and U8830 (N_8830,N_4486,N_2156);
or U8831 (N_8831,N_4135,N_3347);
nand U8832 (N_8832,N_1797,N_729);
nand U8833 (N_8833,N_4583,N_4471);
or U8834 (N_8834,N_123,N_1327);
nand U8835 (N_8835,N_1003,N_919);
and U8836 (N_8836,N_1448,N_944);
xnor U8837 (N_8837,N_2655,N_2903);
nor U8838 (N_8838,N_3917,N_4846);
nor U8839 (N_8839,N_2322,N_2795);
nand U8840 (N_8840,N_3067,N_3021);
nor U8841 (N_8841,N_1787,N_2354);
nand U8842 (N_8842,N_1932,N_2039);
and U8843 (N_8843,N_31,N_2559);
or U8844 (N_8844,N_976,N_2385);
xnor U8845 (N_8845,N_863,N_2628);
nand U8846 (N_8846,N_1276,N_3545);
or U8847 (N_8847,N_3224,N_644);
nor U8848 (N_8848,N_4667,N_1009);
nor U8849 (N_8849,N_1773,N_764);
nand U8850 (N_8850,N_4097,N_4885);
nor U8851 (N_8851,N_2977,N_3068);
nand U8852 (N_8852,N_730,N_4794);
nor U8853 (N_8853,N_3098,N_376);
nand U8854 (N_8854,N_1164,N_1815);
xor U8855 (N_8855,N_4915,N_612);
nor U8856 (N_8856,N_1069,N_1992);
and U8857 (N_8857,N_4903,N_4165);
and U8858 (N_8858,N_3556,N_1506);
xnor U8859 (N_8859,N_1888,N_77);
nor U8860 (N_8860,N_1121,N_3937);
nor U8861 (N_8861,N_869,N_4378);
nor U8862 (N_8862,N_3082,N_653);
or U8863 (N_8863,N_4062,N_2309);
nand U8864 (N_8864,N_4806,N_793);
nor U8865 (N_8865,N_644,N_4941);
and U8866 (N_8866,N_1709,N_2997);
and U8867 (N_8867,N_4710,N_1606);
nor U8868 (N_8868,N_1305,N_4721);
and U8869 (N_8869,N_4512,N_819);
nor U8870 (N_8870,N_2904,N_4691);
and U8871 (N_8871,N_919,N_2087);
nor U8872 (N_8872,N_4068,N_3746);
nor U8873 (N_8873,N_1139,N_1916);
nor U8874 (N_8874,N_344,N_1303);
or U8875 (N_8875,N_1326,N_2621);
and U8876 (N_8876,N_4502,N_4956);
nand U8877 (N_8877,N_460,N_3818);
and U8878 (N_8878,N_468,N_3732);
nor U8879 (N_8879,N_3931,N_1439);
or U8880 (N_8880,N_2326,N_1110);
nor U8881 (N_8881,N_744,N_871);
or U8882 (N_8882,N_1865,N_3796);
xor U8883 (N_8883,N_4653,N_4601);
or U8884 (N_8884,N_2327,N_1823);
or U8885 (N_8885,N_2470,N_968);
and U8886 (N_8886,N_2423,N_2447);
nand U8887 (N_8887,N_637,N_1859);
and U8888 (N_8888,N_2857,N_1640);
nor U8889 (N_8889,N_2991,N_3279);
or U8890 (N_8890,N_4576,N_2764);
and U8891 (N_8891,N_4553,N_585);
or U8892 (N_8892,N_4150,N_1647);
and U8893 (N_8893,N_3059,N_1118);
nor U8894 (N_8894,N_233,N_2376);
and U8895 (N_8895,N_3282,N_3112);
and U8896 (N_8896,N_1973,N_2474);
nand U8897 (N_8897,N_3690,N_2590);
nor U8898 (N_8898,N_4667,N_3807);
nor U8899 (N_8899,N_4331,N_3020);
xnor U8900 (N_8900,N_3626,N_1967);
nand U8901 (N_8901,N_4424,N_1255);
nor U8902 (N_8902,N_1578,N_4066);
and U8903 (N_8903,N_1530,N_698);
and U8904 (N_8904,N_1926,N_1837);
and U8905 (N_8905,N_4518,N_271);
nand U8906 (N_8906,N_4235,N_4261);
xnor U8907 (N_8907,N_2927,N_4211);
nand U8908 (N_8908,N_4506,N_1633);
nand U8909 (N_8909,N_4114,N_2346);
or U8910 (N_8910,N_1147,N_2353);
or U8911 (N_8911,N_2845,N_20);
or U8912 (N_8912,N_1343,N_2467);
xor U8913 (N_8913,N_3295,N_3458);
and U8914 (N_8914,N_2813,N_4594);
nor U8915 (N_8915,N_4045,N_2101);
nand U8916 (N_8916,N_4639,N_4304);
nor U8917 (N_8917,N_4854,N_673);
nand U8918 (N_8918,N_662,N_960);
nand U8919 (N_8919,N_3031,N_1945);
or U8920 (N_8920,N_785,N_1653);
nor U8921 (N_8921,N_1592,N_3310);
nand U8922 (N_8922,N_2713,N_4875);
or U8923 (N_8923,N_446,N_504);
nor U8924 (N_8924,N_4527,N_1227);
or U8925 (N_8925,N_4228,N_207);
and U8926 (N_8926,N_516,N_798);
xnor U8927 (N_8927,N_2848,N_3918);
or U8928 (N_8928,N_3766,N_3276);
and U8929 (N_8929,N_2162,N_159);
nand U8930 (N_8930,N_1066,N_2878);
nor U8931 (N_8931,N_4730,N_4993);
or U8932 (N_8932,N_4855,N_4451);
nand U8933 (N_8933,N_1972,N_2221);
or U8934 (N_8934,N_3249,N_4885);
and U8935 (N_8935,N_641,N_3813);
and U8936 (N_8936,N_2720,N_4541);
and U8937 (N_8937,N_2729,N_3422);
nor U8938 (N_8938,N_4003,N_2188);
xor U8939 (N_8939,N_483,N_2834);
and U8940 (N_8940,N_1787,N_4483);
or U8941 (N_8941,N_4944,N_4951);
or U8942 (N_8942,N_686,N_2018);
nand U8943 (N_8943,N_3353,N_2395);
nand U8944 (N_8944,N_1033,N_39);
or U8945 (N_8945,N_2320,N_748);
nand U8946 (N_8946,N_524,N_3932);
and U8947 (N_8947,N_680,N_1141);
nor U8948 (N_8948,N_3,N_1692);
xor U8949 (N_8949,N_212,N_486);
xor U8950 (N_8950,N_3472,N_4667);
or U8951 (N_8951,N_1554,N_4577);
nor U8952 (N_8952,N_4799,N_3574);
nor U8953 (N_8953,N_1025,N_3397);
or U8954 (N_8954,N_1721,N_4515);
nand U8955 (N_8955,N_684,N_3321);
nand U8956 (N_8956,N_3198,N_3728);
nor U8957 (N_8957,N_1777,N_453);
nor U8958 (N_8958,N_3098,N_4708);
nand U8959 (N_8959,N_154,N_3266);
nand U8960 (N_8960,N_996,N_1117);
or U8961 (N_8961,N_4921,N_3659);
nand U8962 (N_8962,N_3344,N_4011);
nor U8963 (N_8963,N_4318,N_1329);
or U8964 (N_8964,N_4811,N_4018);
nand U8965 (N_8965,N_2804,N_1259);
nor U8966 (N_8966,N_4421,N_3361);
nor U8967 (N_8967,N_4750,N_1658);
and U8968 (N_8968,N_160,N_4724);
and U8969 (N_8969,N_4764,N_4196);
and U8970 (N_8970,N_3840,N_3768);
or U8971 (N_8971,N_4224,N_557);
nand U8972 (N_8972,N_4136,N_333);
or U8973 (N_8973,N_1428,N_350);
or U8974 (N_8974,N_2281,N_1301);
or U8975 (N_8975,N_983,N_3254);
nor U8976 (N_8976,N_1497,N_1238);
nand U8977 (N_8977,N_980,N_4855);
nor U8978 (N_8978,N_1745,N_430);
or U8979 (N_8979,N_4177,N_2061);
or U8980 (N_8980,N_980,N_2422);
nor U8981 (N_8981,N_3044,N_3421);
nor U8982 (N_8982,N_2901,N_2442);
xor U8983 (N_8983,N_1807,N_2040);
xnor U8984 (N_8984,N_2644,N_4522);
nand U8985 (N_8985,N_2355,N_3443);
nor U8986 (N_8986,N_1080,N_4919);
or U8987 (N_8987,N_425,N_3711);
nand U8988 (N_8988,N_4741,N_4985);
nor U8989 (N_8989,N_2651,N_2952);
nor U8990 (N_8990,N_4912,N_1129);
and U8991 (N_8991,N_1133,N_554);
nand U8992 (N_8992,N_4201,N_3101);
and U8993 (N_8993,N_2560,N_1542);
nor U8994 (N_8994,N_3865,N_1717);
or U8995 (N_8995,N_4800,N_1201);
nor U8996 (N_8996,N_4385,N_585);
nand U8997 (N_8997,N_1014,N_4829);
or U8998 (N_8998,N_342,N_1533);
nor U8999 (N_8999,N_4216,N_1172);
xnor U9000 (N_9000,N_1144,N_347);
and U9001 (N_9001,N_3210,N_281);
nor U9002 (N_9002,N_3344,N_517);
and U9003 (N_9003,N_1862,N_439);
nand U9004 (N_9004,N_2374,N_3749);
and U9005 (N_9005,N_4822,N_2229);
nor U9006 (N_9006,N_3195,N_566);
nand U9007 (N_9007,N_3158,N_3190);
or U9008 (N_9008,N_245,N_1836);
and U9009 (N_9009,N_4302,N_730);
and U9010 (N_9010,N_4546,N_3542);
nand U9011 (N_9011,N_4223,N_3682);
nand U9012 (N_9012,N_2257,N_4762);
nand U9013 (N_9013,N_1591,N_341);
and U9014 (N_9014,N_3185,N_1055);
nor U9015 (N_9015,N_2968,N_2113);
nor U9016 (N_9016,N_2147,N_972);
and U9017 (N_9017,N_1332,N_2832);
or U9018 (N_9018,N_1791,N_393);
nor U9019 (N_9019,N_310,N_168);
and U9020 (N_9020,N_1279,N_608);
and U9021 (N_9021,N_1753,N_978);
nor U9022 (N_9022,N_831,N_2308);
nand U9023 (N_9023,N_2207,N_362);
and U9024 (N_9024,N_2475,N_4321);
and U9025 (N_9025,N_3271,N_2061);
nand U9026 (N_9026,N_4131,N_1807);
and U9027 (N_9027,N_2617,N_620);
or U9028 (N_9028,N_3506,N_3495);
xnor U9029 (N_9029,N_3633,N_4426);
nor U9030 (N_9030,N_561,N_3842);
nand U9031 (N_9031,N_4778,N_4547);
nand U9032 (N_9032,N_1617,N_3262);
or U9033 (N_9033,N_3253,N_1699);
and U9034 (N_9034,N_3166,N_3330);
and U9035 (N_9035,N_3565,N_3289);
or U9036 (N_9036,N_1968,N_1971);
nor U9037 (N_9037,N_1403,N_1742);
nand U9038 (N_9038,N_3473,N_1255);
nor U9039 (N_9039,N_2959,N_4651);
or U9040 (N_9040,N_2493,N_3005);
and U9041 (N_9041,N_141,N_2601);
nor U9042 (N_9042,N_3750,N_1435);
or U9043 (N_9043,N_4863,N_398);
or U9044 (N_9044,N_200,N_2913);
xor U9045 (N_9045,N_3458,N_4283);
or U9046 (N_9046,N_2505,N_2133);
and U9047 (N_9047,N_2631,N_2911);
and U9048 (N_9048,N_1812,N_3489);
nor U9049 (N_9049,N_2015,N_1253);
or U9050 (N_9050,N_3817,N_3806);
nor U9051 (N_9051,N_2460,N_4963);
and U9052 (N_9052,N_3019,N_1684);
nor U9053 (N_9053,N_1361,N_4680);
and U9054 (N_9054,N_4416,N_3956);
nor U9055 (N_9055,N_4522,N_3965);
nor U9056 (N_9056,N_2598,N_46);
and U9057 (N_9057,N_3415,N_4197);
and U9058 (N_9058,N_4633,N_184);
or U9059 (N_9059,N_2881,N_1825);
nor U9060 (N_9060,N_666,N_3533);
and U9061 (N_9061,N_3340,N_3904);
nor U9062 (N_9062,N_2094,N_1707);
nand U9063 (N_9063,N_4124,N_1951);
nand U9064 (N_9064,N_120,N_3834);
and U9065 (N_9065,N_3302,N_3471);
and U9066 (N_9066,N_2211,N_647);
nor U9067 (N_9067,N_304,N_3594);
nand U9068 (N_9068,N_3492,N_3849);
nand U9069 (N_9069,N_483,N_7);
and U9070 (N_9070,N_54,N_2630);
and U9071 (N_9071,N_3903,N_1678);
nor U9072 (N_9072,N_3249,N_702);
nor U9073 (N_9073,N_4562,N_2557);
nor U9074 (N_9074,N_3922,N_2091);
xor U9075 (N_9075,N_2518,N_1896);
xnor U9076 (N_9076,N_1868,N_4111);
or U9077 (N_9077,N_4293,N_2766);
nand U9078 (N_9078,N_4696,N_1092);
or U9079 (N_9079,N_3904,N_3155);
nor U9080 (N_9080,N_3132,N_74);
nor U9081 (N_9081,N_2173,N_233);
nor U9082 (N_9082,N_1236,N_4149);
and U9083 (N_9083,N_1346,N_2704);
and U9084 (N_9084,N_4859,N_666);
nand U9085 (N_9085,N_4473,N_2706);
nor U9086 (N_9086,N_4523,N_982);
nand U9087 (N_9087,N_791,N_3630);
nor U9088 (N_9088,N_3395,N_3501);
nor U9089 (N_9089,N_4015,N_3032);
or U9090 (N_9090,N_571,N_520);
and U9091 (N_9091,N_1559,N_3668);
nand U9092 (N_9092,N_1645,N_1797);
nor U9093 (N_9093,N_1028,N_3462);
nand U9094 (N_9094,N_2885,N_1200);
or U9095 (N_9095,N_3649,N_52);
nand U9096 (N_9096,N_1290,N_3584);
nor U9097 (N_9097,N_2506,N_1588);
and U9098 (N_9098,N_2517,N_2476);
and U9099 (N_9099,N_4120,N_3895);
nand U9100 (N_9100,N_61,N_3541);
nor U9101 (N_9101,N_1553,N_4125);
nor U9102 (N_9102,N_3844,N_466);
and U9103 (N_9103,N_1863,N_3453);
and U9104 (N_9104,N_98,N_3349);
and U9105 (N_9105,N_4664,N_1609);
nand U9106 (N_9106,N_2912,N_4006);
nand U9107 (N_9107,N_306,N_1708);
and U9108 (N_9108,N_4926,N_733);
and U9109 (N_9109,N_77,N_3939);
and U9110 (N_9110,N_4509,N_3995);
and U9111 (N_9111,N_2880,N_717);
or U9112 (N_9112,N_1888,N_1019);
nor U9113 (N_9113,N_958,N_1794);
nor U9114 (N_9114,N_459,N_2568);
and U9115 (N_9115,N_2151,N_738);
nand U9116 (N_9116,N_3063,N_225);
nand U9117 (N_9117,N_1766,N_3735);
nor U9118 (N_9118,N_781,N_2779);
and U9119 (N_9119,N_1215,N_1295);
nor U9120 (N_9120,N_1644,N_4905);
nor U9121 (N_9121,N_1856,N_2661);
nand U9122 (N_9122,N_4302,N_2052);
nand U9123 (N_9123,N_2659,N_4135);
or U9124 (N_9124,N_780,N_286);
or U9125 (N_9125,N_434,N_3776);
nor U9126 (N_9126,N_984,N_3277);
xnor U9127 (N_9127,N_4004,N_308);
nand U9128 (N_9128,N_2157,N_3718);
nand U9129 (N_9129,N_1695,N_3352);
nor U9130 (N_9130,N_697,N_335);
nand U9131 (N_9131,N_10,N_76);
nor U9132 (N_9132,N_1101,N_387);
and U9133 (N_9133,N_4445,N_4186);
nand U9134 (N_9134,N_3177,N_1596);
nor U9135 (N_9135,N_4104,N_4622);
and U9136 (N_9136,N_16,N_1712);
and U9137 (N_9137,N_24,N_183);
or U9138 (N_9138,N_1914,N_57);
nand U9139 (N_9139,N_4285,N_3338);
and U9140 (N_9140,N_758,N_4557);
and U9141 (N_9141,N_2794,N_3808);
nor U9142 (N_9142,N_1498,N_1419);
and U9143 (N_9143,N_953,N_2188);
or U9144 (N_9144,N_118,N_4782);
nor U9145 (N_9145,N_444,N_1340);
nor U9146 (N_9146,N_2558,N_3740);
nor U9147 (N_9147,N_934,N_439);
xnor U9148 (N_9148,N_4570,N_4300);
nor U9149 (N_9149,N_4022,N_4080);
and U9150 (N_9150,N_4836,N_4314);
nor U9151 (N_9151,N_637,N_1538);
or U9152 (N_9152,N_790,N_3986);
and U9153 (N_9153,N_4684,N_3424);
or U9154 (N_9154,N_2711,N_944);
nand U9155 (N_9155,N_4546,N_3326);
or U9156 (N_9156,N_2141,N_3267);
or U9157 (N_9157,N_3194,N_1970);
or U9158 (N_9158,N_155,N_3605);
and U9159 (N_9159,N_4527,N_2904);
and U9160 (N_9160,N_2174,N_623);
nand U9161 (N_9161,N_434,N_4532);
and U9162 (N_9162,N_3236,N_406);
nor U9163 (N_9163,N_4264,N_3209);
or U9164 (N_9164,N_1487,N_4315);
nor U9165 (N_9165,N_1923,N_715);
and U9166 (N_9166,N_3204,N_4715);
nor U9167 (N_9167,N_3529,N_1763);
and U9168 (N_9168,N_1948,N_3467);
and U9169 (N_9169,N_4991,N_2533);
and U9170 (N_9170,N_1996,N_957);
nor U9171 (N_9171,N_2612,N_2053);
and U9172 (N_9172,N_3296,N_2314);
or U9173 (N_9173,N_3027,N_1687);
xor U9174 (N_9174,N_1928,N_3819);
nand U9175 (N_9175,N_4832,N_2473);
nand U9176 (N_9176,N_3022,N_4949);
xnor U9177 (N_9177,N_3495,N_688);
xnor U9178 (N_9178,N_3031,N_4580);
and U9179 (N_9179,N_3490,N_228);
and U9180 (N_9180,N_4212,N_2221);
xor U9181 (N_9181,N_3783,N_3631);
nor U9182 (N_9182,N_51,N_608);
and U9183 (N_9183,N_4547,N_4780);
xor U9184 (N_9184,N_16,N_172);
or U9185 (N_9185,N_2108,N_3531);
or U9186 (N_9186,N_4926,N_3104);
and U9187 (N_9187,N_2943,N_3857);
and U9188 (N_9188,N_4028,N_2817);
nor U9189 (N_9189,N_2771,N_883);
nor U9190 (N_9190,N_3537,N_3485);
and U9191 (N_9191,N_484,N_3426);
or U9192 (N_9192,N_4527,N_2009);
or U9193 (N_9193,N_522,N_2539);
xor U9194 (N_9194,N_1709,N_3205);
and U9195 (N_9195,N_2208,N_2885);
nor U9196 (N_9196,N_2751,N_174);
nand U9197 (N_9197,N_3158,N_4313);
nor U9198 (N_9198,N_3868,N_2319);
and U9199 (N_9199,N_4400,N_2921);
and U9200 (N_9200,N_2438,N_3586);
and U9201 (N_9201,N_2911,N_661);
and U9202 (N_9202,N_4269,N_1930);
nand U9203 (N_9203,N_3684,N_2902);
nand U9204 (N_9204,N_1243,N_3869);
or U9205 (N_9205,N_328,N_4800);
xnor U9206 (N_9206,N_1071,N_801);
or U9207 (N_9207,N_440,N_1781);
and U9208 (N_9208,N_4691,N_455);
nand U9209 (N_9209,N_3565,N_722);
and U9210 (N_9210,N_123,N_2611);
nand U9211 (N_9211,N_1744,N_876);
xor U9212 (N_9212,N_4742,N_3627);
and U9213 (N_9213,N_3848,N_3585);
nor U9214 (N_9214,N_632,N_1793);
or U9215 (N_9215,N_19,N_4994);
or U9216 (N_9216,N_2301,N_49);
and U9217 (N_9217,N_1174,N_467);
and U9218 (N_9218,N_3785,N_2431);
or U9219 (N_9219,N_362,N_4466);
nand U9220 (N_9220,N_2332,N_1308);
nor U9221 (N_9221,N_1666,N_1470);
and U9222 (N_9222,N_848,N_2955);
and U9223 (N_9223,N_4609,N_1508);
nand U9224 (N_9224,N_4879,N_1564);
and U9225 (N_9225,N_2169,N_2803);
nor U9226 (N_9226,N_4710,N_2933);
nor U9227 (N_9227,N_4610,N_2145);
and U9228 (N_9228,N_2231,N_4913);
nand U9229 (N_9229,N_3949,N_4190);
or U9230 (N_9230,N_343,N_4958);
or U9231 (N_9231,N_4191,N_1798);
or U9232 (N_9232,N_4987,N_1540);
nand U9233 (N_9233,N_3892,N_3166);
nor U9234 (N_9234,N_2814,N_3637);
and U9235 (N_9235,N_2834,N_45);
and U9236 (N_9236,N_2395,N_4268);
nand U9237 (N_9237,N_2622,N_1612);
and U9238 (N_9238,N_202,N_3837);
nor U9239 (N_9239,N_28,N_3570);
and U9240 (N_9240,N_695,N_3729);
nand U9241 (N_9241,N_1696,N_1708);
and U9242 (N_9242,N_2577,N_2105);
and U9243 (N_9243,N_393,N_4513);
nor U9244 (N_9244,N_3807,N_154);
nor U9245 (N_9245,N_2930,N_95);
or U9246 (N_9246,N_158,N_3239);
nand U9247 (N_9247,N_3527,N_4151);
nor U9248 (N_9248,N_4922,N_1615);
and U9249 (N_9249,N_1821,N_97);
nand U9250 (N_9250,N_94,N_3605);
and U9251 (N_9251,N_3246,N_3567);
or U9252 (N_9252,N_3287,N_3924);
nand U9253 (N_9253,N_1460,N_3769);
nand U9254 (N_9254,N_1444,N_4405);
nand U9255 (N_9255,N_2120,N_647);
nand U9256 (N_9256,N_4041,N_1215);
nor U9257 (N_9257,N_1368,N_967);
or U9258 (N_9258,N_4951,N_917);
nand U9259 (N_9259,N_2736,N_2804);
and U9260 (N_9260,N_3105,N_2461);
and U9261 (N_9261,N_360,N_455);
nand U9262 (N_9262,N_2611,N_2701);
or U9263 (N_9263,N_4640,N_1302);
nor U9264 (N_9264,N_3542,N_4003);
and U9265 (N_9265,N_3219,N_676);
nor U9266 (N_9266,N_3168,N_1479);
nand U9267 (N_9267,N_4923,N_4787);
nor U9268 (N_9268,N_4770,N_2938);
nand U9269 (N_9269,N_4174,N_251);
or U9270 (N_9270,N_4264,N_194);
and U9271 (N_9271,N_3541,N_2712);
or U9272 (N_9272,N_578,N_1039);
nand U9273 (N_9273,N_2451,N_4759);
and U9274 (N_9274,N_542,N_4839);
and U9275 (N_9275,N_3198,N_2758);
or U9276 (N_9276,N_2433,N_1253);
nand U9277 (N_9277,N_2717,N_3306);
or U9278 (N_9278,N_2304,N_1075);
or U9279 (N_9279,N_3881,N_1916);
xor U9280 (N_9280,N_1925,N_3841);
and U9281 (N_9281,N_1447,N_4300);
or U9282 (N_9282,N_92,N_2056);
or U9283 (N_9283,N_170,N_3282);
nand U9284 (N_9284,N_997,N_3242);
nand U9285 (N_9285,N_4897,N_1756);
xor U9286 (N_9286,N_2014,N_119);
or U9287 (N_9287,N_4347,N_220);
and U9288 (N_9288,N_3996,N_343);
nand U9289 (N_9289,N_284,N_153);
nor U9290 (N_9290,N_3266,N_230);
xnor U9291 (N_9291,N_1986,N_3563);
or U9292 (N_9292,N_4047,N_2316);
nand U9293 (N_9293,N_1623,N_3498);
or U9294 (N_9294,N_2246,N_4739);
nand U9295 (N_9295,N_86,N_1425);
or U9296 (N_9296,N_1618,N_2275);
or U9297 (N_9297,N_629,N_3167);
or U9298 (N_9298,N_1047,N_4340);
and U9299 (N_9299,N_964,N_2316);
nand U9300 (N_9300,N_1963,N_3041);
and U9301 (N_9301,N_1297,N_3265);
nor U9302 (N_9302,N_4240,N_579);
nand U9303 (N_9303,N_1170,N_911);
xor U9304 (N_9304,N_4078,N_2043);
or U9305 (N_9305,N_4271,N_2550);
nor U9306 (N_9306,N_1599,N_2277);
nor U9307 (N_9307,N_3208,N_3270);
and U9308 (N_9308,N_1250,N_1591);
and U9309 (N_9309,N_4968,N_1245);
nor U9310 (N_9310,N_3849,N_1682);
or U9311 (N_9311,N_2631,N_787);
or U9312 (N_9312,N_314,N_4064);
xor U9313 (N_9313,N_97,N_1547);
nand U9314 (N_9314,N_1155,N_1669);
or U9315 (N_9315,N_2795,N_799);
nor U9316 (N_9316,N_2499,N_2864);
and U9317 (N_9317,N_1037,N_585);
nor U9318 (N_9318,N_4939,N_2307);
or U9319 (N_9319,N_3752,N_2869);
and U9320 (N_9320,N_4048,N_4177);
nor U9321 (N_9321,N_4436,N_4224);
nand U9322 (N_9322,N_1664,N_1421);
nor U9323 (N_9323,N_2368,N_3701);
xnor U9324 (N_9324,N_4322,N_82);
and U9325 (N_9325,N_4467,N_494);
nor U9326 (N_9326,N_2245,N_4765);
and U9327 (N_9327,N_1518,N_2694);
nor U9328 (N_9328,N_3453,N_2588);
nor U9329 (N_9329,N_2225,N_176);
nor U9330 (N_9330,N_4931,N_446);
nand U9331 (N_9331,N_4504,N_2901);
nand U9332 (N_9332,N_4093,N_933);
nand U9333 (N_9333,N_2502,N_4278);
nand U9334 (N_9334,N_3807,N_4983);
xor U9335 (N_9335,N_2554,N_2858);
or U9336 (N_9336,N_4105,N_4100);
nand U9337 (N_9337,N_856,N_2443);
and U9338 (N_9338,N_4565,N_2001);
and U9339 (N_9339,N_107,N_2894);
xnor U9340 (N_9340,N_122,N_1110);
nand U9341 (N_9341,N_1437,N_2564);
nor U9342 (N_9342,N_2017,N_4667);
nand U9343 (N_9343,N_1996,N_2674);
and U9344 (N_9344,N_1860,N_306);
or U9345 (N_9345,N_1211,N_3943);
or U9346 (N_9346,N_4362,N_1978);
nor U9347 (N_9347,N_3603,N_2553);
or U9348 (N_9348,N_1898,N_4367);
nor U9349 (N_9349,N_4918,N_4636);
or U9350 (N_9350,N_1370,N_414);
nand U9351 (N_9351,N_1126,N_4030);
or U9352 (N_9352,N_3162,N_1254);
or U9353 (N_9353,N_1302,N_3922);
and U9354 (N_9354,N_4365,N_1681);
nand U9355 (N_9355,N_4511,N_3933);
or U9356 (N_9356,N_1361,N_2799);
nor U9357 (N_9357,N_1837,N_968);
nand U9358 (N_9358,N_3238,N_4974);
nor U9359 (N_9359,N_4878,N_4999);
xnor U9360 (N_9360,N_2018,N_292);
or U9361 (N_9361,N_1362,N_3676);
nand U9362 (N_9362,N_987,N_549);
or U9363 (N_9363,N_2684,N_3353);
nor U9364 (N_9364,N_3514,N_947);
nor U9365 (N_9365,N_2842,N_2966);
or U9366 (N_9366,N_3654,N_4248);
nand U9367 (N_9367,N_2499,N_2900);
and U9368 (N_9368,N_2965,N_3610);
and U9369 (N_9369,N_383,N_581);
or U9370 (N_9370,N_118,N_1178);
nand U9371 (N_9371,N_3391,N_2829);
nand U9372 (N_9372,N_4921,N_2607);
or U9373 (N_9373,N_1687,N_3777);
nand U9374 (N_9374,N_195,N_1219);
or U9375 (N_9375,N_3479,N_3765);
nor U9376 (N_9376,N_3744,N_1350);
or U9377 (N_9377,N_4943,N_3710);
or U9378 (N_9378,N_303,N_776);
nand U9379 (N_9379,N_4651,N_14);
nand U9380 (N_9380,N_3254,N_4802);
or U9381 (N_9381,N_1478,N_2469);
xor U9382 (N_9382,N_3606,N_1742);
and U9383 (N_9383,N_4074,N_815);
nor U9384 (N_9384,N_4827,N_2708);
nand U9385 (N_9385,N_3964,N_3371);
xor U9386 (N_9386,N_3028,N_4411);
and U9387 (N_9387,N_3889,N_4198);
or U9388 (N_9388,N_289,N_3001);
xnor U9389 (N_9389,N_1163,N_3591);
and U9390 (N_9390,N_4393,N_1404);
and U9391 (N_9391,N_4310,N_3877);
nand U9392 (N_9392,N_906,N_2484);
and U9393 (N_9393,N_4710,N_1967);
xnor U9394 (N_9394,N_3963,N_1426);
and U9395 (N_9395,N_3945,N_2369);
nor U9396 (N_9396,N_3957,N_2596);
or U9397 (N_9397,N_77,N_1166);
or U9398 (N_9398,N_1002,N_165);
or U9399 (N_9399,N_3864,N_421);
nor U9400 (N_9400,N_542,N_3696);
nor U9401 (N_9401,N_962,N_2069);
nor U9402 (N_9402,N_677,N_1029);
and U9403 (N_9403,N_4779,N_3877);
or U9404 (N_9404,N_2377,N_471);
nand U9405 (N_9405,N_945,N_1724);
nor U9406 (N_9406,N_526,N_3790);
nor U9407 (N_9407,N_2645,N_3562);
and U9408 (N_9408,N_2975,N_1999);
xnor U9409 (N_9409,N_387,N_4666);
and U9410 (N_9410,N_2849,N_143);
nor U9411 (N_9411,N_2286,N_2650);
and U9412 (N_9412,N_1770,N_525);
and U9413 (N_9413,N_4071,N_1641);
or U9414 (N_9414,N_1441,N_2475);
nand U9415 (N_9415,N_423,N_2440);
and U9416 (N_9416,N_1318,N_1754);
or U9417 (N_9417,N_1421,N_309);
or U9418 (N_9418,N_615,N_4388);
or U9419 (N_9419,N_3196,N_2729);
nor U9420 (N_9420,N_3792,N_1903);
or U9421 (N_9421,N_2237,N_1161);
nand U9422 (N_9422,N_2549,N_3619);
or U9423 (N_9423,N_819,N_4766);
nand U9424 (N_9424,N_1511,N_2640);
and U9425 (N_9425,N_1682,N_437);
or U9426 (N_9426,N_4621,N_705);
nor U9427 (N_9427,N_2999,N_3352);
nor U9428 (N_9428,N_1968,N_1738);
or U9429 (N_9429,N_4250,N_4728);
and U9430 (N_9430,N_2162,N_609);
and U9431 (N_9431,N_384,N_2944);
xnor U9432 (N_9432,N_2275,N_4350);
xor U9433 (N_9433,N_1113,N_3924);
and U9434 (N_9434,N_4209,N_4774);
or U9435 (N_9435,N_1935,N_3684);
nand U9436 (N_9436,N_2671,N_3628);
nand U9437 (N_9437,N_3826,N_623);
nor U9438 (N_9438,N_628,N_982);
and U9439 (N_9439,N_1635,N_2085);
xor U9440 (N_9440,N_1684,N_4066);
nor U9441 (N_9441,N_4732,N_4527);
and U9442 (N_9442,N_1508,N_3428);
or U9443 (N_9443,N_2906,N_2669);
nor U9444 (N_9444,N_2688,N_1912);
nand U9445 (N_9445,N_4748,N_3955);
nor U9446 (N_9446,N_4555,N_3559);
nor U9447 (N_9447,N_4978,N_264);
nor U9448 (N_9448,N_355,N_4829);
or U9449 (N_9449,N_1632,N_4231);
or U9450 (N_9450,N_2792,N_4292);
or U9451 (N_9451,N_3718,N_4285);
or U9452 (N_9452,N_244,N_1095);
nor U9453 (N_9453,N_1196,N_4672);
or U9454 (N_9454,N_2655,N_605);
and U9455 (N_9455,N_917,N_624);
and U9456 (N_9456,N_47,N_4604);
nand U9457 (N_9457,N_4501,N_3266);
and U9458 (N_9458,N_2857,N_1839);
nor U9459 (N_9459,N_4025,N_1498);
xnor U9460 (N_9460,N_1233,N_2435);
or U9461 (N_9461,N_2991,N_4482);
xnor U9462 (N_9462,N_4738,N_1769);
nand U9463 (N_9463,N_4620,N_3280);
nand U9464 (N_9464,N_4205,N_1116);
and U9465 (N_9465,N_4591,N_2180);
nor U9466 (N_9466,N_2731,N_2572);
and U9467 (N_9467,N_4649,N_2505);
or U9468 (N_9468,N_3523,N_1775);
or U9469 (N_9469,N_1364,N_3131);
nand U9470 (N_9470,N_4170,N_1634);
nor U9471 (N_9471,N_2948,N_4569);
nor U9472 (N_9472,N_3577,N_255);
or U9473 (N_9473,N_2224,N_455);
nor U9474 (N_9474,N_273,N_526);
or U9475 (N_9475,N_667,N_1187);
and U9476 (N_9476,N_4703,N_4330);
nor U9477 (N_9477,N_3966,N_1335);
and U9478 (N_9478,N_4703,N_1572);
or U9479 (N_9479,N_2000,N_3441);
and U9480 (N_9480,N_833,N_2732);
nor U9481 (N_9481,N_439,N_1780);
or U9482 (N_9482,N_1024,N_2208);
and U9483 (N_9483,N_3816,N_1008);
nand U9484 (N_9484,N_4559,N_1869);
nor U9485 (N_9485,N_3227,N_60);
or U9486 (N_9486,N_4466,N_4303);
nor U9487 (N_9487,N_1511,N_810);
nor U9488 (N_9488,N_4495,N_4749);
or U9489 (N_9489,N_2058,N_1937);
nor U9490 (N_9490,N_2669,N_3917);
nand U9491 (N_9491,N_1185,N_2533);
or U9492 (N_9492,N_3092,N_1364);
nor U9493 (N_9493,N_4585,N_1207);
or U9494 (N_9494,N_321,N_2442);
nand U9495 (N_9495,N_316,N_1175);
nand U9496 (N_9496,N_525,N_2685);
and U9497 (N_9497,N_4880,N_3751);
nor U9498 (N_9498,N_4416,N_126);
nand U9499 (N_9499,N_3183,N_2008);
or U9500 (N_9500,N_1313,N_4095);
xor U9501 (N_9501,N_1941,N_3910);
nor U9502 (N_9502,N_2701,N_336);
and U9503 (N_9503,N_3146,N_2272);
and U9504 (N_9504,N_4738,N_3572);
xnor U9505 (N_9505,N_3267,N_1354);
nor U9506 (N_9506,N_1376,N_2969);
or U9507 (N_9507,N_1083,N_1380);
nand U9508 (N_9508,N_3232,N_3543);
or U9509 (N_9509,N_1033,N_4119);
or U9510 (N_9510,N_4321,N_4232);
and U9511 (N_9511,N_3785,N_3016);
and U9512 (N_9512,N_1401,N_4182);
and U9513 (N_9513,N_1648,N_3740);
or U9514 (N_9514,N_4109,N_473);
or U9515 (N_9515,N_3269,N_3501);
nor U9516 (N_9516,N_1085,N_113);
and U9517 (N_9517,N_4942,N_2226);
nor U9518 (N_9518,N_4000,N_1340);
and U9519 (N_9519,N_2426,N_28);
nor U9520 (N_9520,N_1258,N_808);
nand U9521 (N_9521,N_4892,N_3568);
or U9522 (N_9522,N_4022,N_4609);
nand U9523 (N_9523,N_4216,N_4719);
and U9524 (N_9524,N_2743,N_1594);
xnor U9525 (N_9525,N_4692,N_3374);
and U9526 (N_9526,N_1642,N_4434);
nor U9527 (N_9527,N_3261,N_1210);
nor U9528 (N_9528,N_1628,N_4929);
nor U9529 (N_9529,N_3380,N_959);
or U9530 (N_9530,N_2816,N_3340);
and U9531 (N_9531,N_3157,N_1781);
nand U9532 (N_9532,N_3818,N_1372);
or U9533 (N_9533,N_2233,N_3241);
nor U9534 (N_9534,N_513,N_2119);
or U9535 (N_9535,N_1124,N_4222);
nor U9536 (N_9536,N_1655,N_2169);
and U9537 (N_9537,N_476,N_4433);
nand U9538 (N_9538,N_283,N_1366);
nand U9539 (N_9539,N_371,N_1279);
nand U9540 (N_9540,N_908,N_1995);
and U9541 (N_9541,N_765,N_1115);
and U9542 (N_9542,N_3175,N_1145);
xnor U9543 (N_9543,N_733,N_903);
nor U9544 (N_9544,N_196,N_2116);
and U9545 (N_9545,N_4814,N_426);
and U9546 (N_9546,N_3701,N_4838);
nor U9547 (N_9547,N_537,N_930);
or U9548 (N_9548,N_781,N_3689);
or U9549 (N_9549,N_4907,N_3024);
and U9550 (N_9550,N_3164,N_2950);
nor U9551 (N_9551,N_2528,N_2897);
or U9552 (N_9552,N_4627,N_304);
and U9553 (N_9553,N_1341,N_1176);
xnor U9554 (N_9554,N_2977,N_1761);
nand U9555 (N_9555,N_3984,N_4073);
nand U9556 (N_9556,N_2328,N_978);
nor U9557 (N_9557,N_855,N_4305);
nand U9558 (N_9558,N_692,N_2282);
or U9559 (N_9559,N_3483,N_4587);
nor U9560 (N_9560,N_382,N_1925);
or U9561 (N_9561,N_3919,N_187);
nor U9562 (N_9562,N_4776,N_1953);
or U9563 (N_9563,N_4198,N_4626);
nor U9564 (N_9564,N_636,N_3027);
nand U9565 (N_9565,N_412,N_1360);
nor U9566 (N_9566,N_2019,N_1428);
or U9567 (N_9567,N_1189,N_3474);
xnor U9568 (N_9568,N_3613,N_2516);
nand U9569 (N_9569,N_3354,N_1935);
nand U9570 (N_9570,N_1145,N_1297);
nor U9571 (N_9571,N_3197,N_964);
and U9572 (N_9572,N_1532,N_4877);
nor U9573 (N_9573,N_2471,N_3575);
or U9574 (N_9574,N_3905,N_331);
nand U9575 (N_9575,N_433,N_20);
or U9576 (N_9576,N_2517,N_1281);
or U9577 (N_9577,N_2466,N_382);
xnor U9578 (N_9578,N_767,N_3305);
nand U9579 (N_9579,N_2051,N_3347);
nor U9580 (N_9580,N_129,N_2000);
or U9581 (N_9581,N_2208,N_3306);
or U9582 (N_9582,N_4222,N_120);
nor U9583 (N_9583,N_3442,N_4872);
and U9584 (N_9584,N_3938,N_3618);
nand U9585 (N_9585,N_3192,N_1259);
nand U9586 (N_9586,N_3268,N_3833);
and U9587 (N_9587,N_3647,N_2680);
nor U9588 (N_9588,N_3026,N_3464);
nor U9589 (N_9589,N_2666,N_790);
nand U9590 (N_9590,N_574,N_4478);
and U9591 (N_9591,N_307,N_838);
and U9592 (N_9592,N_2446,N_272);
or U9593 (N_9593,N_2515,N_4587);
nor U9594 (N_9594,N_1857,N_865);
or U9595 (N_9595,N_2646,N_239);
nand U9596 (N_9596,N_115,N_902);
and U9597 (N_9597,N_4475,N_2052);
or U9598 (N_9598,N_2439,N_2295);
nor U9599 (N_9599,N_1493,N_3541);
nor U9600 (N_9600,N_960,N_978);
and U9601 (N_9601,N_4371,N_553);
nand U9602 (N_9602,N_1229,N_4117);
or U9603 (N_9603,N_429,N_3057);
nor U9604 (N_9604,N_1430,N_3898);
or U9605 (N_9605,N_2205,N_763);
xnor U9606 (N_9606,N_1250,N_2565);
xor U9607 (N_9607,N_1385,N_1596);
nor U9608 (N_9608,N_2676,N_1372);
nor U9609 (N_9609,N_4908,N_1788);
and U9610 (N_9610,N_1856,N_1047);
nand U9611 (N_9611,N_4231,N_34);
nand U9612 (N_9612,N_1440,N_2497);
or U9613 (N_9613,N_3800,N_3231);
and U9614 (N_9614,N_3047,N_3886);
nor U9615 (N_9615,N_1598,N_4559);
or U9616 (N_9616,N_881,N_2137);
nor U9617 (N_9617,N_4170,N_1357);
nor U9618 (N_9618,N_3641,N_1833);
nand U9619 (N_9619,N_2654,N_2726);
and U9620 (N_9620,N_356,N_2716);
nand U9621 (N_9621,N_3833,N_1535);
and U9622 (N_9622,N_375,N_3361);
and U9623 (N_9623,N_2477,N_1302);
or U9624 (N_9624,N_2841,N_3254);
nand U9625 (N_9625,N_407,N_594);
nor U9626 (N_9626,N_1784,N_4053);
and U9627 (N_9627,N_4723,N_4578);
xnor U9628 (N_9628,N_4291,N_1679);
nor U9629 (N_9629,N_2014,N_1893);
and U9630 (N_9630,N_3458,N_580);
and U9631 (N_9631,N_4938,N_2003);
nand U9632 (N_9632,N_3852,N_2905);
and U9633 (N_9633,N_1649,N_2992);
xnor U9634 (N_9634,N_3665,N_1958);
or U9635 (N_9635,N_3689,N_1989);
nand U9636 (N_9636,N_3909,N_4580);
or U9637 (N_9637,N_194,N_1491);
and U9638 (N_9638,N_2907,N_3574);
nor U9639 (N_9639,N_4780,N_2644);
or U9640 (N_9640,N_2214,N_236);
or U9641 (N_9641,N_1417,N_1790);
nor U9642 (N_9642,N_918,N_4227);
or U9643 (N_9643,N_4119,N_3420);
nor U9644 (N_9644,N_2965,N_398);
and U9645 (N_9645,N_3531,N_3238);
nor U9646 (N_9646,N_3448,N_1271);
nor U9647 (N_9647,N_2659,N_3301);
and U9648 (N_9648,N_3247,N_4644);
or U9649 (N_9649,N_4997,N_4998);
nor U9650 (N_9650,N_189,N_3534);
nand U9651 (N_9651,N_1643,N_316);
nand U9652 (N_9652,N_685,N_4009);
nor U9653 (N_9653,N_4457,N_3486);
and U9654 (N_9654,N_3666,N_4512);
and U9655 (N_9655,N_146,N_2266);
nor U9656 (N_9656,N_848,N_79);
and U9657 (N_9657,N_1954,N_4880);
and U9658 (N_9658,N_3713,N_3621);
xor U9659 (N_9659,N_1851,N_937);
xnor U9660 (N_9660,N_3218,N_2706);
xnor U9661 (N_9661,N_2712,N_2925);
xor U9662 (N_9662,N_2904,N_3393);
nor U9663 (N_9663,N_1197,N_4810);
and U9664 (N_9664,N_3858,N_3094);
or U9665 (N_9665,N_633,N_4705);
or U9666 (N_9666,N_4235,N_4911);
or U9667 (N_9667,N_255,N_2097);
or U9668 (N_9668,N_1558,N_3899);
nor U9669 (N_9669,N_4123,N_4243);
nor U9670 (N_9670,N_3804,N_3138);
nor U9671 (N_9671,N_3175,N_4863);
or U9672 (N_9672,N_3279,N_3085);
nand U9673 (N_9673,N_1236,N_1701);
or U9674 (N_9674,N_194,N_4874);
or U9675 (N_9675,N_4799,N_3803);
nand U9676 (N_9676,N_4536,N_1208);
and U9677 (N_9677,N_51,N_4560);
or U9678 (N_9678,N_1434,N_804);
nand U9679 (N_9679,N_3921,N_391);
nand U9680 (N_9680,N_3764,N_498);
and U9681 (N_9681,N_1342,N_2362);
or U9682 (N_9682,N_4174,N_3876);
and U9683 (N_9683,N_3806,N_1071);
nor U9684 (N_9684,N_4868,N_3854);
or U9685 (N_9685,N_945,N_4956);
nand U9686 (N_9686,N_2633,N_1894);
nand U9687 (N_9687,N_3605,N_1572);
and U9688 (N_9688,N_1834,N_3436);
or U9689 (N_9689,N_4343,N_1724);
nand U9690 (N_9690,N_4307,N_4962);
and U9691 (N_9691,N_3993,N_2052);
xor U9692 (N_9692,N_1243,N_633);
nor U9693 (N_9693,N_685,N_2795);
nor U9694 (N_9694,N_298,N_1618);
nor U9695 (N_9695,N_2423,N_956);
nor U9696 (N_9696,N_3766,N_1468);
and U9697 (N_9697,N_4178,N_3985);
xor U9698 (N_9698,N_997,N_1846);
nor U9699 (N_9699,N_2592,N_3509);
xor U9700 (N_9700,N_1395,N_4689);
nand U9701 (N_9701,N_2423,N_2352);
and U9702 (N_9702,N_4452,N_1457);
or U9703 (N_9703,N_4873,N_1684);
or U9704 (N_9704,N_4246,N_949);
and U9705 (N_9705,N_1056,N_4155);
and U9706 (N_9706,N_2724,N_1242);
and U9707 (N_9707,N_110,N_785);
or U9708 (N_9708,N_1462,N_124);
or U9709 (N_9709,N_55,N_728);
xor U9710 (N_9710,N_1600,N_103);
xor U9711 (N_9711,N_4026,N_4404);
xnor U9712 (N_9712,N_1004,N_786);
or U9713 (N_9713,N_733,N_1270);
nand U9714 (N_9714,N_414,N_1130);
and U9715 (N_9715,N_2463,N_4258);
or U9716 (N_9716,N_4980,N_2851);
nand U9717 (N_9717,N_3352,N_3256);
nor U9718 (N_9718,N_2393,N_1527);
xor U9719 (N_9719,N_681,N_1837);
xnor U9720 (N_9720,N_915,N_4079);
nor U9721 (N_9721,N_4852,N_4753);
nand U9722 (N_9722,N_2365,N_3400);
or U9723 (N_9723,N_3668,N_87);
nand U9724 (N_9724,N_3078,N_3827);
or U9725 (N_9725,N_4244,N_2504);
xor U9726 (N_9726,N_465,N_3338);
nor U9727 (N_9727,N_1000,N_1264);
or U9728 (N_9728,N_2441,N_1780);
or U9729 (N_9729,N_1958,N_294);
nand U9730 (N_9730,N_3708,N_2893);
nor U9731 (N_9731,N_435,N_2893);
nand U9732 (N_9732,N_2497,N_395);
nand U9733 (N_9733,N_584,N_4680);
or U9734 (N_9734,N_3637,N_616);
nand U9735 (N_9735,N_3007,N_422);
and U9736 (N_9736,N_3807,N_2137);
or U9737 (N_9737,N_4955,N_4253);
nor U9738 (N_9738,N_2393,N_2345);
xor U9739 (N_9739,N_512,N_4319);
xnor U9740 (N_9740,N_1086,N_3545);
and U9741 (N_9741,N_3647,N_590);
nor U9742 (N_9742,N_1391,N_861);
nor U9743 (N_9743,N_4467,N_4484);
nor U9744 (N_9744,N_1670,N_3437);
nor U9745 (N_9745,N_1459,N_3933);
nor U9746 (N_9746,N_933,N_3005);
or U9747 (N_9747,N_2168,N_4021);
and U9748 (N_9748,N_3472,N_4124);
xor U9749 (N_9749,N_3934,N_161);
or U9750 (N_9750,N_4345,N_924);
nor U9751 (N_9751,N_4699,N_1500);
nor U9752 (N_9752,N_702,N_3852);
and U9753 (N_9753,N_3021,N_3956);
or U9754 (N_9754,N_3723,N_433);
and U9755 (N_9755,N_1643,N_2431);
nand U9756 (N_9756,N_4984,N_4974);
xor U9757 (N_9757,N_2416,N_4818);
nand U9758 (N_9758,N_25,N_1826);
or U9759 (N_9759,N_3559,N_2294);
nand U9760 (N_9760,N_3560,N_3064);
and U9761 (N_9761,N_3604,N_1615);
nand U9762 (N_9762,N_849,N_1319);
nor U9763 (N_9763,N_4821,N_276);
xor U9764 (N_9764,N_2999,N_3458);
or U9765 (N_9765,N_4211,N_2123);
and U9766 (N_9766,N_4135,N_1983);
or U9767 (N_9767,N_3812,N_2082);
or U9768 (N_9768,N_2827,N_4094);
nand U9769 (N_9769,N_2603,N_791);
nor U9770 (N_9770,N_4857,N_1482);
xor U9771 (N_9771,N_4095,N_4045);
or U9772 (N_9772,N_1641,N_2521);
or U9773 (N_9773,N_2430,N_268);
and U9774 (N_9774,N_4654,N_4842);
and U9775 (N_9775,N_1550,N_3659);
or U9776 (N_9776,N_3903,N_836);
and U9777 (N_9777,N_3331,N_3219);
or U9778 (N_9778,N_11,N_1771);
or U9779 (N_9779,N_2416,N_4994);
or U9780 (N_9780,N_1047,N_2632);
nand U9781 (N_9781,N_2862,N_1739);
or U9782 (N_9782,N_3103,N_2599);
and U9783 (N_9783,N_1668,N_4152);
nor U9784 (N_9784,N_3199,N_3627);
or U9785 (N_9785,N_222,N_633);
and U9786 (N_9786,N_570,N_1728);
or U9787 (N_9787,N_1179,N_325);
and U9788 (N_9788,N_4557,N_1035);
and U9789 (N_9789,N_2625,N_4163);
and U9790 (N_9790,N_1027,N_2542);
xor U9791 (N_9791,N_342,N_814);
nand U9792 (N_9792,N_3289,N_1151);
and U9793 (N_9793,N_4673,N_338);
and U9794 (N_9794,N_4746,N_1828);
nand U9795 (N_9795,N_2265,N_937);
or U9796 (N_9796,N_2981,N_2537);
and U9797 (N_9797,N_3354,N_3402);
xnor U9798 (N_9798,N_2867,N_4280);
or U9799 (N_9799,N_211,N_1374);
nand U9800 (N_9800,N_1893,N_2079);
nor U9801 (N_9801,N_44,N_1322);
nand U9802 (N_9802,N_4576,N_2059);
nand U9803 (N_9803,N_3187,N_4310);
and U9804 (N_9804,N_1298,N_149);
nor U9805 (N_9805,N_319,N_2425);
nor U9806 (N_9806,N_889,N_3636);
nand U9807 (N_9807,N_989,N_4080);
xnor U9808 (N_9808,N_3570,N_4699);
or U9809 (N_9809,N_2454,N_597);
or U9810 (N_9810,N_1302,N_2655);
nand U9811 (N_9811,N_4514,N_3094);
and U9812 (N_9812,N_2739,N_1386);
nand U9813 (N_9813,N_2804,N_1310);
or U9814 (N_9814,N_370,N_4043);
nor U9815 (N_9815,N_3238,N_1904);
or U9816 (N_9816,N_3743,N_696);
and U9817 (N_9817,N_3142,N_1506);
nor U9818 (N_9818,N_4908,N_1655);
nor U9819 (N_9819,N_4583,N_1254);
nand U9820 (N_9820,N_1760,N_2127);
nor U9821 (N_9821,N_1312,N_2621);
nor U9822 (N_9822,N_2034,N_4886);
or U9823 (N_9823,N_2014,N_2916);
nor U9824 (N_9824,N_1246,N_928);
or U9825 (N_9825,N_4486,N_2178);
nand U9826 (N_9826,N_1501,N_1009);
xnor U9827 (N_9827,N_658,N_2994);
or U9828 (N_9828,N_3943,N_4705);
and U9829 (N_9829,N_3538,N_3913);
nor U9830 (N_9830,N_2572,N_4734);
or U9831 (N_9831,N_1776,N_2974);
and U9832 (N_9832,N_3077,N_4981);
nor U9833 (N_9833,N_3136,N_1450);
nor U9834 (N_9834,N_3269,N_1985);
or U9835 (N_9835,N_3733,N_2293);
and U9836 (N_9836,N_451,N_3907);
nor U9837 (N_9837,N_1774,N_3503);
nand U9838 (N_9838,N_3249,N_318);
or U9839 (N_9839,N_3744,N_1588);
and U9840 (N_9840,N_628,N_4834);
nor U9841 (N_9841,N_3012,N_1488);
and U9842 (N_9842,N_175,N_3377);
and U9843 (N_9843,N_3569,N_2992);
nand U9844 (N_9844,N_4702,N_3408);
or U9845 (N_9845,N_988,N_973);
or U9846 (N_9846,N_246,N_2610);
or U9847 (N_9847,N_520,N_2481);
and U9848 (N_9848,N_2383,N_2892);
and U9849 (N_9849,N_296,N_2414);
or U9850 (N_9850,N_3832,N_3513);
and U9851 (N_9851,N_4595,N_4815);
nor U9852 (N_9852,N_2340,N_2742);
nor U9853 (N_9853,N_902,N_562);
and U9854 (N_9854,N_2206,N_1697);
nand U9855 (N_9855,N_2882,N_2838);
nor U9856 (N_9856,N_1516,N_3959);
or U9857 (N_9857,N_2609,N_143);
nor U9858 (N_9858,N_4936,N_3211);
nor U9859 (N_9859,N_2765,N_779);
nor U9860 (N_9860,N_1582,N_3004);
and U9861 (N_9861,N_3103,N_1305);
nor U9862 (N_9862,N_4589,N_1205);
or U9863 (N_9863,N_714,N_1879);
nor U9864 (N_9864,N_4852,N_4173);
nor U9865 (N_9865,N_4772,N_4842);
nand U9866 (N_9866,N_4171,N_2821);
and U9867 (N_9867,N_3838,N_4717);
xor U9868 (N_9868,N_2328,N_2798);
xnor U9869 (N_9869,N_1198,N_1174);
nor U9870 (N_9870,N_1601,N_4132);
nor U9871 (N_9871,N_3165,N_3029);
nand U9872 (N_9872,N_800,N_3378);
nand U9873 (N_9873,N_1369,N_4742);
nand U9874 (N_9874,N_4731,N_4832);
and U9875 (N_9875,N_3974,N_221);
and U9876 (N_9876,N_2489,N_1010);
or U9877 (N_9877,N_3456,N_3360);
or U9878 (N_9878,N_4429,N_404);
and U9879 (N_9879,N_4360,N_3501);
or U9880 (N_9880,N_2435,N_894);
xor U9881 (N_9881,N_399,N_2126);
or U9882 (N_9882,N_4533,N_4166);
xor U9883 (N_9883,N_2740,N_1624);
or U9884 (N_9884,N_1112,N_3766);
nand U9885 (N_9885,N_2727,N_3198);
nor U9886 (N_9886,N_4615,N_2350);
nor U9887 (N_9887,N_4229,N_2440);
nor U9888 (N_9888,N_4129,N_952);
or U9889 (N_9889,N_3040,N_1131);
nor U9890 (N_9890,N_4948,N_291);
xor U9891 (N_9891,N_3237,N_648);
nand U9892 (N_9892,N_3074,N_69);
or U9893 (N_9893,N_2921,N_2826);
nor U9894 (N_9894,N_2606,N_2278);
nor U9895 (N_9895,N_2035,N_449);
nand U9896 (N_9896,N_964,N_1000);
nand U9897 (N_9897,N_3648,N_2029);
nand U9898 (N_9898,N_1020,N_2033);
and U9899 (N_9899,N_1794,N_3478);
nor U9900 (N_9900,N_4619,N_3718);
and U9901 (N_9901,N_2434,N_182);
nor U9902 (N_9902,N_1576,N_549);
nand U9903 (N_9903,N_4329,N_4991);
or U9904 (N_9904,N_3106,N_920);
nor U9905 (N_9905,N_3823,N_4518);
and U9906 (N_9906,N_2845,N_1767);
and U9907 (N_9907,N_2831,N_3346);
or U9908 (N_9908,N_4513,N_3716);
nand U9909 (N_9909,N_568,N_1331);
and U9910 (N_9910,N_3158,N_3575);
nor U9911 (N_9911,N_3638,N_3933);
or U9912 (N_9912,N_4144,N_4283);
or U9913 (N_9913,N_216,N_361);
xnor U9914 (N_9914,N_430,N_427);
or U9915 (N_9915,N_1888,N_1653);
xor U9916 (N_9916,N_586,N_900);
nand U9917 (N_9917,N_2872,N_953);
and U9918 (N_9918,N_2455,N_1418);
nand U9919 (N_9919,N_4710,N_3105);
or U9920 (N_9920,N_4895,N_4270);
or U9921 (N_9921,N_1542,N_4367);
nor U9922 (N_9922,N_3169,N_1004);
nand U9923 (N_9923,N_3028,N_2476);
xnor U9924 (N_9924,N_757,N_4522);
nand U9925 (N_9925,N_3591,N_621);
nand U9926 (N_9926,N_3078,N_4482);
or U9927 (N_9927,N_3152,N_1324);
nand U9928 (N_9928,N_1115,N_3810);
nor U9929 (N_9929,N_1057,N_4849);
xnor U9930 (N_9930,N_3095,N_272);
xnor U9931 (N_9931,N_3324,N_1310);
and U9932 (N_9932,N_1943,N_2304);
nand U9933 (N_9933,N_3578,N_2454);
nor U9934 (N_9934,N_4930,N_3237);
or U9935 (N_9935,N_161,N_2725);
or U9936 (N_9936,N_2375,N_2285);
nand U9937 (N_9937,N_467,N_1467);
nor U9938 (N_9938,N_2567,N_1481);
and U9939 (N_9939,N_632,N_2304);
and U9940 (N_9940,N_1094,N_957);
and U9941 (N_9941,N_2831,N_3983);
or U9942 (N_9942,N_2516,N_3546);
nor U9943 (N_9943,N_2605,N_1691);
nor U9944 (N_9944,N_1730,N_304);
and U9945 (N_9945,N_4101,N_3208);
nand U9946 (N_9946,N_4049,N_1852);
and U9947 (N_9947,N_1051,N_4523);
nand U9948 (N_9948,N_3658,N_2850);
and U9949 (N_9949,N_2709,N_4710);
nand U9950 (N_9950,N_2625,N_4728);
nand U9951 (N_9951,N_221,N_4229);
or U9952 (N_9952,N_1682,N_2881);
nor U9953 (N_9953,N_733,N_743);
or U9954 (N_9954,N_430,N_4132);
nand U9955 (N_9955,N_2763,N_3102);
nor U9956 (N_9956,N_4418,N_2767);
nand U9957 (N_9957,N_2063,N_2573);
and U9958 (N_9958,N_2370,N_4149);
xnor U9959 (N_9959,N_1011,N_959);
nand U9960 (N_9960,N_547,N_2825);
and U9961 (N_9961,N_3192,N_345);
xnor U9962 (N_9962,N_4045,N_3033);
nor U9963 (N_9963,N_4181,N_2236);
or U9964 (N_9964,N_4301,N_364);
and U9965 (N_9965,N_1477,N_1325);
and U9966 (N_9966,N_941,N_1527);
nand U9967 (N_9967,N_3622,N_4490);
nor U9968 (N_9968,N_4548,N_2975);
nor U9969 (N_9969,N_189,N_4635);
and U9970 (N_9970,N_2410,N_4948);
or U9971 (N_9971,N_3438,N_2649);
and U9972 (N_9972,N_704,N_1491);
nor U9973 (N_9973,N_4975,N_4070);
nor U9974 (N_9974,N_2829,N_1500);
xor U9975 (N_9975,N_3262,N_206);
nand U9976 (N_9976,N_4689,N_620);
or U9977 (N_9977,N_1109,N_4318);
nand U9978 (N_9978,N_1189,N_2503);
and U9979 (N_9979,N_2480,N_2115);
nor U9980 (N_9980,N_2559,N_162);
nand U9981 (N_9981,N_4829,N_3384);
or U9982 (N_9982,N_4510,N_3973);
or U9983 (N_9983,N_3533,N_2752);
and U9984 (N_9984,N_4393,N_1107);
nand U9985 (N_9985,N_147,N_2910);
and U9986 (N_9986,N_418,N_1170);
nand U9987 (N_9987,N_3748,N_2343);
xor U9988 (N_9988,N_4305,N_4657);
or U9989 (N_9989,N_2335,N_4555);
nand U9990 (N_9990,N_2464,N_2245);
nand U9991 (N_9991,N_1339,N_2470);
nand U9992 (N_9992,N_2997,N_1204);
or U9993 (N_9993,N_4213,N_4250);
nand U9994 (N_9994,N_616,N_2787);
xnor U9995 (N_9995,N_2498,N_3222);
nor U9996 (N_9996,N_4639,N_397);
nor U9997 (N_9997,N_2936,N_703);
nand U9998 (N_9998,N_4577,N_197);
nor U9999 (N_9999,N_4869,N_2192);
or U10000 (N_10000,N_6375,N_8707);
nand U10001 (N_10001,N_8361,N_5258);
or U10002 (N_10002,N_9159,N_8632);
nor U10003 (N_10003,N_8991,N_5180);
nor U10004 (N_10004,N_8536,N_6984);
nor U10005 (N_10005,N_9619,N_6223);
xnor U10006 (N_10006,N_6393,N_6362);
nand U10007 (N_10007,N_6724,N_9585);
or U10008 (N_10008,N_9995,N_7950);
nor U10009 (N_10009,N_7514,N_6266);
xor U10010 (N_10010,N_8326,N_6317);
and U10011 (N_10011,N_7595,N_8734);
xnor U10012 (N_10012,N_9312,N_8495);
nand U10013 (N_10013,N_5420,N_6775);
and U10014 (N_10014,N_9766,N_8784);
and U10015 (N_10015,N_8910,N_9216);
xor U10016 (N_10016,N_7622,N_6033);
or U10017 (N_10017,N_6229,N_8235);
and U10018 (N_10018,N_5221,N_7850);
or U10019 (N_10019,N_8723,N_8846);
nand U10020 (N_10020,N_5036,N_6730);
or U10021 (N_10021,N_9526,N_5170);
nand U10022 (N_10022,N_6830,N_8420);
nor U10023 (N_10023,N_6626,N_9869);
and U10024 (N_10024,N_8436,N_7503);
or U10025 (N_10025,N_5421,N_6779);
nor U10026 (N_10026,N_8544,N_9945);
and U10027 (N_10027,N_5386,N_9790);
and U10028 (N_10028,N_9334,N_9286);
and U10029 (N_10029,N_7464,N_5827);
nor U10030 (N_10030,N_6566,N_7977);
nand U10031 (N_10031,N_7927,N_9803);
nor U10032 (N_10032,N_8921,N_7285);
xor U10033 (N_10033,N_8912,N_8643);
nand U10034 (N_10034,N_9400,N_7088);
and U10035 (N_10035,N_7478,N_6662);
or U10036 (N_10036,N_5492,N_8011);
and U10037 (N_10037,N_7846,N_5133);
nand U10038 (N_10038,N_7426,N_9249);
and U10039 (N_10039,N_5068,N_8700);
nor U10040 (N_10040,N_6803,N_5515);
nand U10041 (N_10041,N_9788,N_8785);
nor U10042 (N_10042,N_5164,N_6133);
and U10043 (N_10043,N_8229,N_5882);
nand U10044 (N_10044,N_8849,N_6621);
nor U10045 (N_10045,N_6006,N_8301);
nand U10046 (N_10046,N_6915,N_9771);
or U10047 (N_10047,N_7283,N_7300);
or U10048 (N_10048,N_9465,N_8965);
nand U10049 (N_10049,N_5497,N_8597);
nor U10050 (N_10050,N_5601,N_8382);
and U10051 (N_10051,N_5796,N_6822);
nand U10052 (N_10052,N_8101,N_6208);
nand U10053 (N_10053,N_9376,N_8903);
and U10054 (N_10054,N_7101,N_5625);
xnor U10055 (N_10055,N_8896,N_7284);
nand U10056 (N_10056,N_5504,N_6173);
nand U10057 (N_10057,N_6806,N_8687);
and U10058 (N_10058,N_8561,N_6354);
or U10059 (N_10059,N_7576,N_6076);
and U10060 (N_10060,N_6828,N_6609);
and U10061 (N_10061,N_6794,N_7791);
nor U10062 (N_10062,N_7396,N_5220);
nor U10063 (N_10063,N_7868,N_6212);
nor U10064 (N_10064,N_7308,N_8188);
or U10065 (N_10065,N_6183,N_7705);
xnor U10066 (N_10066,N_6257,N_6811);
and U10067 (N_10067,N_5501,N_9475);
and U10068 (N_10068,N_8464,N_9503);
nand U10069 (N_10069,N_6572,N_9816);
or U10070 (N_10070,N_5849,N_9714);
and U10071 (N_10071,N_8907,N_7481);
nand U10072 (N_10072,N_6979,N_5554);
xor U10073 (N_10073,N_5673,N_8883);
or U10074 (N_10074,N_7356,N_5433);
xnor U10075 (N_10075,N_9494,N_8506);
nor U10076 (N_10076,N_5087,N_8322);
or U10077 (N_10077,N_8054,N_5716);
nor U10078 (N_10078,N_9117,N_7301);
and U10079 (N_10079,N_7193,N_5630);
nand U10080 (N_10080,N_6324,N_9954);
nor U10081 (N_10081,N_7804,N_6597);
nand U10082 (N_10082,N_8678,N_8198);
and U10083 (N_10083,N_9891,N_7382);
nand U10084 (N_10084,N_7392,N_5527);
and U10085 (N_10085,N_6792,N_7614);
nor U10086 (N_10086,N_5779,N_7240);
or U10087 (N_10087,N_8456,N_8060);
and U10088 (N_10088,N_7185,N_6941);
nand U10089 (N_10089,N_7035,N_7414);
or U10090 (N_10090,N_6922,N_5464);
nand U10091 (N_10091,N_5281,N_7482);
nand U10092 (N_10092,N_6969,N_6882);
nand U10093 (N_10093,N_6648,N_9586);
nand U10094 (N_10094,N_7402,N_5029);
or U10095 (N_10095,N_5418,N_8321);
or U10096 (N_10096,N_5413,N_6715);
nand U10097 (N_10097,N_9674,N_5776);
and U10098 (N_10098,N_5968,N_9584);
or U10099 (N_10099,N_6176,N_8016);
nand U10100 (N_10100,N_8547,N_9907);
nor U10101 (N_10101,N_7377,N_6505);
and U10102 (N_10102,N_7974,N_5586);
or U10103 (N_10103,N_8167,N_5282);
and U10104 (N_10104,N_5631,N_6047);
or U10105 (N_10105,N_5992,N_7855);
nand U10106 (N_10106,N_9225,N_5686);
nand U10107 (N_10107,N_7215,N_7948);
and U10108 (N_10108,N_8617,N_8049);
nand U10109 (N_10109,N_9377,N_7197);
or U10110 (N_10110,N_9611,N_5910);
and U10111 (N_10111,N_6744,N_8862);
nand U10112 (N_10112,N_6040,N_5090);
nor U10113 (N_10113,N_7555,N_5046);
nor U10114 (N_10114,N_6222,N_8172);
nor U10115 (N_10115,N_5193,N_5949);
nand U10116 (N_10116,N_7174,N_5300);
or U10117 (N_10117,N_7628,N_5664);
nor U10118 (N_10118,N_8150,N_6459);
and U10119 (N_10119,N_6330,N_6655);
nand U10120 (N_10120,N_7731,N_7632);
nand U10121 (N_10121,N_7202,N_9588);
and U10122 (N_10122,N_5127,N_5031);
and U10123 (N_10123,N_7933,N_6771);
nand U10124 (N_10124,N_9232,N_6042);
nor U10125 (N_10125,N_5764,N_6313);
nand U10126 (N_10126,N_6968,N_9612);
or U10127 (N_10127,N_7996,N_8341);
nand U10128 (N_10128,N_5793,N_6365);
nand U10129 (N_10129,N_9917,N_5409);
xnor U10130 (N_10130,N_7781,N_6109);
nand U10131 (N_10131,N_5357,N_5248);
or U10132 (N_10132,N_5195,N_7609);
and U10133 (N_10133,N_6370,N_9574);
or U10134 (N_10134,N_7867,N_6675);
and U10135 (N_10135,N_5295,N_8760);
nand U10136 (N_10136,N_7316,N_8942);
and U10137 (N_10137,N_8758,N_5502);
or U10138 (N_10138,N_7347,N_7582);
nand U10139 (N_10139,N_6963,N_9221);
and U10140 (N_10140,N_7673,N_8124);
nand U10141 (N_10141,N_6301,N_8268);
or U10142 (N_10142,N_5028,N_7373);
xor U10143 (N_10143,N_8541,N_9784);
nor U10144 (N_10144,N_5675,N_7122);
and U10145 (N_10145,N_5839,N_6419);
or U10146 (N_10146,N_8486,N_7750);
or U10147 (N_10147,N_9902,N_8433);
nor U10148 (N_10148,N_9825,N_9536);
nand U10149 (N_10149,N_6914,N_9212);
nand U10150 (N_10150,N_9818,N_5639);
and U10151 (N_10151,N_6574,N_7754);
nand U10152 (N_10152,N_5561,N_7799);
xor U10153 (N_10153,N_6933,N_7567);
nand U10154 (N_10154,N_7932,N_5469);
and U10155 (N_10155,N_5247,N_8162);
and U10156 (N_10156,N_5438,N_7383);
nor U10157 (N_10157,N_8540,N_6015);
nor U10158 (N_10158,N_5157,N_5013);
nand U10159 (N_10159,N_7938,N_5712);
or U10160 (N_10160,N_5027,N_5547);
nor U10161 (N_10161,N_5808,N_7633);
nand U10162 (N_10162,N_5002,N_7753);
or U10163 (N_10163,N_6778,N_7689);
and U10164 (N_10164,N_9920,N_7230);
xor U10165 (N_10165,N_9914,N_8961);
or U10166 (N_10166,N_6220,N_6050);
nand U10167 (N_10167,N_9994,N_8572);
nand U10168 (N_10168,N_7447,N_8193);
xnor U10169 (N_10169,N_7898,N_8745);
and U10170 (N_10170,N_6619,N_8287);
and U10171 (N_10171,N_7142,N_9557);
and U10172 (N_10172,N_8851,N_7231);
nand U10173 (N_10173,N_7683,N_8738);
or U10174 (N_10174,N_7528,N_8444);
or U10175 (N_10175,N_5478,N_7442);
and U10176 (N_10176,N_9164,N_8946);
or U10177 (N_10177,N_9723,N_5312);
xnor U10178 (N_10178,N_7430,N_6820);
and U10179 (N_10179,N_7236,N_5941);
or U10180 (N_10180,N_8880,N_8206);
nand U10181 (N_10181,N_9116,N_9455);
nor U10182 (N_10182,N_8189,N_8674);
nor U10183 (N_10183,N_9260,N_8209);
and U10184 (N_10184,N_9856,N_9928);
nor U10185 (N_10185,N_8007,N_7335);
or U10186 (N_10186,N_8087,N_6353);
nand U10187 (N_10187,N_7972,N_9686);
and U10188 (N_10188,N_9796,N_9009);
nor U10189 (N_10189,N_8574,N_5495);
or U10190 (N_10190,N_7304,N_7278);
nor U10191 (N_10191,N_7601,N_8146);
nand U10192 (N_10192,N_7794,N_9390);
nor U10193 (N_10193,N_7295,N_8283);
and U10194 (N_10194,N_7217,N_8783);
and U10195 (N_10195,N_7186,N_5050);
xnor U10196 (N_10196,N_5823,N_8499);
nand U10197 (N_10197,N_5939,N_9942);
and U10198 (N_10198,N_7890,N_6136);
and U10199 (N_10199,N_5475,N_5679);
nor U10200 (N_10200,N_6360,N_8663);
nand U10201 (N_10201,N_5177,N_8267);
nor U10202 (N_10202,N_5626,N_7533);
or U10203 (N_10203,N_5961,N_8040);
nor U10204 (N_10204,N_5965,N_7145);
nand U10205 (N_10205,N_6578,N_6287);
nor U10206 (N_10206,N_7672,N_9798);
or U10207 (N_10207,N_5655,N_5113);
and U10208 (N_10208,N_7554,N_5393);
nand U10209 (N_10209,N_8048,N_7138);
and U10210 (N_10210,N_7027,N_8667);
nand U10211 (N_10211,N_8050,N_5471);
and U10212 (N_10212,N_7674,N_5889);
or U10213 (N_10213,N_8699,N_6777);
or U10214 (N_10214,N_9348,N_8688);
or U10215 (N_10215,N_6760,N_9805);
or U10216 (N_10216,N_6474,N_5905);
and U10217 (N_10217,N_5765,N_7748);
or U10218 (N_10218,N_6009,N_9428);
and U10219 (N_10219,N_7262,N_7963);
nor U10220 (N_10220,N_8219,N_7235);
nor U10221 (N_10221,N_5301,N_6003);
nand U10222 (N_10222,N_7654,N_7289);
or U10223 (N_10223,N_8164,N_6396);
and U10224 (N_10224,N_8794,N_6711);
and U10225 (N_10225,N_9861,N_6315);
nand U10226 (N_10226,N_7515,N_5804);
or U10227 (N_10227,N_8523,N_6157);
and U10228 (N_10228,N_6286,N_9191);
nand U10229 (N_10229,N_9495,N_7976);
or U10230 (N_10230,N_8207,N_5314);
nand U10231 (N_10231,N_8014,N_8036);
and U10232 (N_10232,N_7579,N_7086);
or U10233 (N_10233,N_6096,N_7448);
or U10234 (N_10234,N_8295,N_9090);
nand U10235 (N_10235,N_9183,N_7495);
xnor U10236 (N_10236,N_6861,N_6320);
or U10237 (N_10237,N_8119,N_7054);
and U10238 (N_10238,N_7733,N_6978);
or U10239 (N_10239,N_7372,N_9243);
and U10240 (N_10240,N_5855,N_9336);
nand U10241 (N_10241,N_8842,N_5480);
nand U10242 (N_10242,N_6603,N_8416);
or U10243 (N_10243,N_7046,N_9020);
and U10244 (N_10244,N_5709,N_8709);
and U10245 (N_10245,N_6568,N_8804);
nor U10246 (N_10246,N_8461,N_5840);
or U10247 (N_10247,N_9975,N_9765);
and U10248 (N_10248,N_6823,N_7181);
nand U10249 (N_10249,N_9036,N_7825);
or U10250 (N_10250,N_7268,N_8122);
nand U10251 (N_10251,N_9114,N_9882);
and U10252 (N_10252,N_5197,N_8155);
nor U10253 (N_10253,N_6007,N_8931);
nand U10254 (N_10254,N_8276,N_6649);
nor U10255 (N_10255,N_9808,N_5881);
nor U10256 (N_10256,N_8479,N_5754);
or U10257 (N_10257,N_8197,N_5848);
nor U10258 (N_10258,N_8117,N_8303);
nor U10259 (N_10259,N_5482,N_7715);
or U10260 (N_10260,N_9072,N_9357);
nand U10261 (N_10261,N_7605,N_6293);
or U10262 (N_10262,N_9346,N_9100);
and U10263 (N_10263,N_7324,N_8533);
nand U10264 (N_10264,N_5878,N_8520);
and U10265 (N_10265,N_9950,N_6254);
and U10266 (N_10266,N_5629,N_7840);
or U10267 (N_10267,N_7995,N_6769);
or U10268 (N_10268,N_5638,N_7374);
or U10269 (N_10269,N_6247,N_9614);
and U10270 (N_10270,N_7886,N_7258);
nand U10271 (N_10271,N_6659,N_9595);
nor U10272 (N_10272,N_7379,N_7204);
nor U10273 (N_10273,N_7108,N_9649);
and U10274 (N_10274,N_8236,N_6366);
xor U10275 (N_10275,N_6196,N_5940);
or U10276 (N_10276,N_8998,N_5244);
nor U10277 (N_10277,N_5147,N_8775);
nor U10278 (N_10278,N_6858,N_9038);
or U10279 (N_10279,N_5742,N_5703);
nand U10280 (N_10280,N_7588,N_7550);
nand U10281 (N_10281,N_5700,N_8681);
or U10282 (N_10282,N_8010,N_8598);
and U10283 (N_10283,N_6110,N_7617);
and U10284 (N_10284,N_7330,N_5137);
nor U10285 (N_10285,N_8988,N_6904);
nand U10286 (N_10286,N_9507,N_9043);
and U10287 (N_10287,N_5242,N_9845);
nand U10288 (N_10288,N_8993,N_8161);
nand U10289 (N_10289,N_7786,N_5611);
nor U10290 (N_10290,N_9449,N_9145);
xor U10291 (N_10291,N_9452,N_7012);
nor U10292 (N_10292,N_9393,N_7969);
and U10293 (N_10293,N_9366,N_5929);
nand U10294 (N_10294,N_7249,N_7759);
xnor U10295 (N_10295,N_6054,N_5101);
xor U10296 (N_10296,N_6795,N_7676);
and U10297 (N_10297,N_9931,N_8884);
and U10298 (N_10298,N_8447,N_7028);
nand U10299 (N_10299,N_9015,N_6939);
and U10300 (N_10300,N_5057,N_7057);
and U10301 (N_10301,N_8743,N_9958);
and U10302 (N_10302,N_6340,N_7650);
nand U10303 (N_10303,N_7862,N_6906);
and U10304 (N_10304,N_6886,N_5191);
xor U10305 (N_10305,N_8127,N_5782);
nand U10306 (N_10306,N_7707,N_8195);
xor U10307 (N_10307,N_8366,N_7656);
or U10308 (N_10308,N_9591,N_7162);
or U10309 (N_10309,N_9335,N_9441);
and U10310 (N_10310,N_5368,N_7973);
and U10311 (N_10311,N_5389,N_9172);
nand U10312 (N_10312,N_8485,N_7111);
nand U10313 (N_10313,N_5020,N_6121);
nand U10314 (N_10314,N_7302,N_7728);
nand U10315 (N_10315,N_8690,N_6781);
nand U10316 (N_10316,N_7878,N_6759);
nor U10317 (N_10317,N_9606,N_9035);
nor U10318 (N_10318,N_7698,N_8868);
xor U10319 (N_10319,N_9760,N_9434);
or U10320 (N_10320,N_7851,N_9941);
or U10321 (N_10321,N_5531,N_6788);
or U10322 (N_10322,N_5023,N_7755);
nor U10323 (N_10323,N_9559,N_8962);
nand U10324 (N_10324,N_8364,N_9740);
nor U10325 (N_10325,N_7487,N_8424);
nor U10326 (N_10326,N_8185,N_9399);
nor U10327 (N_10327,N_8771,N_7100);
xor U10328 (N_10328,N_5642,N_9696);
nand U10329 (N_10329,N_6761,N_5158);
nor U10330 (N_10330,N_7102,N_5388);
nand U10331 (N_10331,N_9860,N_9565);
and U10332 (N_10332,N_8062,N_5483);
and U10333 (N_10333,N_9309,N_6390);
nor U10334 (N_10334,N_7847,N_9040);
nand U10335 (N_10335,N_7079,N_8953);
nor U10336 (N_10336,N_6462,N_9398);
nor U10337 (N_10337,N_9240,N_8889);
nand U10338 (N_10338,N_9669,N_5770);
and U10339 (N_10339,N_6402,N_8857);
nor U10340 (N_10340,N_8067,N_7954);
xnor U10341 (N_10341,N_7675,N_9829);
nand U10342 (N_10342,N_8419,N_5865);
and U10343 (N_10343,N_7504,N_6277);
xnor U10344 (N_10344,N_6782,N_5188);
or U10345 (N_10345,N_5085,N_5916);
nand U10346 (N_10346,N_9733,N_5277);
and U10347 (N_10347,N_8736,N_6727);
and U10348 (N_10348,N_9343,N_7522);
nor U10349 (N_10349,N_5318,N_7099);
nand U10350 (N_10350,N_7915,N_6668);
or U10351 (N_10351,N_6556,N_8782);
nor U10352 (N_10352,N_8952,N_7148);
or U10353 (N_10353,N_9098,N_7920);
or U10354 (N_10354,N_6833,N_9888);
nand U10355 (N_10355,N_5359,N_5648);
and U10356 (N_10356,N_9572,N_9124);
xor U10357 (N_10357,N_5181,N_8627);
xnor U10358 (N_10358,N_6610,N_5959);
nor U10359 (N_10359,N_6106,N_8901);
and U10360 (N_10360,N_9424,N_9084);
nand U10361 (N_10361,N_7690,N_8645);
nand U10362 (N_10362,N_5066,N_5333);
and U10363 (N_10363,N_9724,N_9178);
nand U10364 (N_10364,N_8171,N_6584);
and U10365 (N_10365,N_8201,N_7121);
or U10366 (N_10366,N_8414,N_8452);
nor U10367 (N_10367,N_6916,N_6528);
nand U10368 (N_10368,N_5985,N_5896);
and U10369 (N_10369,N_7808,N_8400);
or U10370 (N_10370,N_8780,N_6569);
nand U10371 (N_10371,N_7282,N_6664);
xor U10372 (N_10372,N_5903,N_6087);
or U10373 (N_10373,N_9016,N_8555);
and U10374 (N_10374,N_9039,N_6726);
xnor U10375 (N_10375,N_9474,N_8345);
and U10376 (N_10376,N_7376,N_5832);
or U10377 (N_10377,N_9073,N_8939);
xor U10378 (N_10378,N_7171,N_6465);
and U10379 (N_10379,N_7062,N_5913);
or U10380 (N_10380,N_9139,N_8802);
and U10381 (N_10381,N_8554,N_7050);
nand U10382 (N_10382,N_5211,N_7516);
nand U10383 (N_10383,N_5500,N_9986);
nand U10384 (N_10384,N_6912,N_6897);
and U10385 (N_10385,N_9290,N_9151);
nor U10386 (N_10386,N_6486,N_6723);
and U10387 (N_10387,N_8739,N_7055);
and U10388 (N_10388,N_7361,N_5542);
nor U10389 (N_10389,N_6321,N_7022);
and U10390 (N_10390,N_5689,N_6546);
nand U10391 (N_10391,N_5407,N_8240);
and U10392 (N_10392,N_6080,N_7228);
xnor U10393 (N_10393,N_7668,N_6355);
nor U10394 (N_10394,N_5185,N_9857);
nand U10395 (N_10395,N_7745,N_9838);
and U10396 (N_10396,N_8956,N_8537);
nand U10397 (N_10397,N_6034,N_9456);
nor U10398 (N_10398,N_8886,N_8353);
and U10399 (N_10399,N_5831,N_6826);
nor U10400 (N_10400,N_6159,N_5073);
or U10401 (N_10401,N_5982,N_6774);
or U10402 (N_10402,N_6174,N_6517);
or U10403 (N_10403,N_5996,N_9013);
and U10404 (N_10404,N_8347,N_8019);
nor U10405 (N_10405,N_7941,N_6398);
nand U10406 (N_10406,N_9905,N_9079);
nor U10407 (N_10407,N_8034,N_9822);
and U10408 (N_10408,N_5463,N_8811);
nor U10409 (N_10409,N_7732,N_6078);
or U10410 (N_10410,N_8113,N_7990);
and U10411 (N_10411,N_6068,N_7742);
nand U10412 (N_10412,N_7010,N_6364);
nand U10413 (N_10413,N_6520,N_7470);
nand U10414 (N_10414,N_5476,N_7313);
xnor U10415 (N_10415,N_9638,N_7272);
nand U10416 (N_10416,N_5795,N_9830);
nand U10417 (N_10417,N_7993,N_5098);
or U10418 (N_10418,N_9149,N_8312);
or U10419 (N_10419,N_5752,N_6890);
or U10420 (N_10420,N_5222,N_7222);
and U10421 (N_10421,N_7777,N_6108);
or U10422 (N_10422,N_6154,N_7000);
nor U10423 (N_10423,N_5826,N_9528);
xor U10424 (N_10424,N_9851,N_6498);
or U10425 (N_10425,N_5788,N_6225);
nor U10426 (N_10426,N_5890,N_5160);
or U10427 (N_10427,N_9508,N_5498);
and U10428 (N_10428,N_6385,N_6156);
or U10429 (N_10429,N_7998,N_7439);
nand U10430 (N_10430,N_9438,N_7457);
nor U10431 (N_10431,N_9444,N_7934);
xor U10432 (N_10432,N_8876,N_5640);
or U10433 (N_10433,N_9094,N_7255);
and U10434 (N_10434,N_6435,N_9450);
and U10435 (N_10435,N_5313,N_8875);
or U10436 (N_10436,N_5837,N_9021);
or U10437 (N_10437,N_6669,N_7018);
nand U10438 (N_10438,N_7252,N_8418);
or U10439 (N_10439,N_9432,N_8649);
nor U10440 (N_10440,N_8483,N_6606);
nor U10441 (N_10441,N_7548,N_8354);
or U10442 (N_10442,N_8257,N_8503);
or U10443 (N_10443,N_7139,N_6294);
or U10444 (N_10444,N_6495,N_7149);
nand U10445 (N_10445,N_8916,N_6526);
or U10446 (N_10446,N_9575,N_5490);
nor U10447 (N_10447,N_7835,N_9533);
nand U10448 (N_10448,N_6338,N_9248);
nor U10449 (N_10449,N_8539,N_6622);
xor U10450 (N_10450,N_5614,N_5459);
xnor U10451 (N_10451,N_6678,N_6024);
and U10452 (N_10452,N_5392,N_5694);
or U10453 (N_10453,N_7485,N_5385);
and U10454 (N_10454,N_9246,N_5159);
and U10455 (N_10455,N_9319,N_9935);
and U10456 (N_10456,N_9513,N_6937);
nand U10457 (N_10457,N_9439,N_7917);
nor U10458 (N_10458,N_7093,N_7491);
xnor U10459 (N_10459,N_5736,N_8484);
nand U10460 (N_10460,N_9717,N_5390);
or U10461 (N_10461,N_5403,N_6309);
and U10462 (N_10462,N_9997,N_5844);
and U10463 (N_10463,N_9102,N_7869);
and U10464 (N_10464,N_8032,N_6644);
and U10465 (N_10465,N_9453,N_7856);
nor U10466 (N_10466,N_8378,N_6306);
or U10467 (N_10467,N_6586,N_9978);
nor U10468 (N_10468,N_8824,N_6525);
nor U10469 (N_10469,N_6071,N_5914);
or U10470 (N_10470,N_6815,N_9321);
nand U10471 (N_10471,N_9814,N_9362);
and U10472 (N_10472,N_5944,N_5962);
and U10473 (N_10473,N_9197,N_6227);
and U10474 (N_10474,N_9989,N_7233);
and U10475 (N_10475,N_7418,N_6756);
and U10476 (N_10476,N_7410,N_9835);
or U10477 (N_10477,N_5095,N_8894);
xor U10478 (N_10478,N_5327,N_9943);
nand U10479 (N_10479,N_5039,N_7544);
nand U10480 (N_10480,N_8560,N_5064);
nand U10481 (N_10481,N_7957,N_8075);
or U10482 (N_10482,N_8575,N_8204);
xor U10483 (N_10483,N_7106,N_5874);
nand U10484 (N_10484,N_9929,N_7445);
nor U10485 (N_10485,N_6607,N_6630);
or U10486 (N_10486,N_8764,N_9990);
or U10487 (N_10487,N_6262,N_5074);
and U10488 (N_10488,N_9150,N_6384);
nor U10489 (N_10489,N_7572,N_5083);
nor U10490 (N_10490,N_5030,N_9486);
or U10491 (N_10491,N_5316,N_9537);
nor U10492 (N_10492,N_9984,N_8566);
and U10493 (N_10493,N_8149,N_8489);
nor U10494 (N_10494,N_8830,N_5275);
nor U10495 (N_10495,N_7349,N_9932);
nor U10496 (N_10496,N_8589,N_9464);
nor U10497 (N_10497,N_7147,N_6902);
nand U10498 (N_10498,N_6747,N_7961);
or U10499 (N_10499,N_9473,N_9480);
nand U10500 (N_10500,N_8021,N_8975);
and U10501 (N_10501,N_6395,N_6274);
or U10502 (N_10502,N_9632,N_7765);
nand U10503 (N_10503,N_6799,N_6834);
or U10504 (N_10504,N_8337,N_5529);
xnor U10505 (N_10505,N_6460,N_5192);
and U10506 (N_10506,N_5223,N_5194);
nor U10507 (N_10507,N_7205,N_7717);
nor U10508 (N_10508,N_9687,N_7944);
or U10509 (N_10509,N_7436,N_7505);
and U10510 (N_10510,N_8922,N_6976);
nor U10511 (N_10511,N_9824,N_8066);
xnor U10512 (N_10512,N_7011,N_6860);
and U10513 (N_10513,N_8105,N_5011);
nand U10514 (N_10514,N_9001,N_9018);
nor U10515 (N_10515,N_8937,N_7734);
or U10516 (N_10516,N_6408,N_6591);
nand U10517 (N_10517,N_6178,N_5202);
nor U10518 (N_10518,N_5341,N_7469);
nand U10519 (N_10519,N_7743,N_9185);
nand U10520 (N_10520,N_9846,N_7506);
or U10521 (N_10521,N_7471,N_9388);
nor U10522 (N_10522,N_6344,N_9715);
nor U10523 (N_10523,N_5723,N_6786);
nand U10524 (N_10524,N_6887,N_9599);
nor U10525 (N_10525,N_8613,N_7083);
and U10526 (N_10526,N_7247,N_6986);
nand U10527 (N_10527,N_9898,N_9590);
or U10528 (N_10528,N_6256,N_8675);
nand U10529 (N_10529,N_7701,N_6944);
xnor U10530 (N_10530,N_5190,N_9878);
or U10531 (N_10531,N_9792,N_5128);
and U10532 (N_10532,N_8064,N_5102);
or U10533 (N_10533,N_7433,N_7746);
nand U10534 (N_10534,N_8137,N_8821);
or U10535 (N_10535,N_7201,N_6182);
or U10536 (N_10536,N_7161,N_9443);
nor U10537 (N_10537,N_9304,N_9957);
or U10538 (N_10538,N_5382,N_7921);
nor U10539 (N_10539,N_6989,N_7807);
nor U10540 (N_10540,N_9332,N_7239);
and U10541 (N_10541,N_5659,N_7651);
nor U10542 (N_10542,N_6144,N_7169);
nor U10543 (N_10543,N_7594,N_7760);
or U10544 (N_10544,N_6379,N_9204);
or U10545 (N_10545,N_8328,N_6634);
nor U10546 (N_10546,N_6328,N_6875);
nor U10547 (N_10547,N_8976,N_7530);
nor U10548 (N_10548,N_9126,N_8384);
nor U10549 (N_10549,N_5344,N_5336);
xor U10550 (N_10550,N_7687,N_8581);
nand U10551 (N_10551,N_8228,N_9604);
or U10552 (N_10552,N_7646,N_6950);
and U10553 (N_10553,N_5843,N_9363);
nand U10554 (N_10554,N_5454,N_6595);
nand U10555 (N_10555,N_8805,N_8728);
nor U10556 (N_10556,N_5111,N_9296);
and U10557 (N_10557,N_6478,N_7558);
or U10558 (N_10558,N_7493,N_6911);
and U10559 (N_10559,N_5287,N_6554);
xor U10560 (N_10560,N_8427,N_8092);
or U10561 (N_10561,N_6907,N_8877);
or U10562 (N_10562,N_7340,N_7679);
and U10563 (N_10563,N_8273,N_5431);
nor U10564 (N_10564,N_8951,N_5605);
xnor U10565 (N_10565,N_7838,N_6899);
xnor U10566 (N_10566,N_5835,N_6020);
nor U10567 (N_10567,N_9677,N_7883);
and U10568 (N_10568,N_6111,N_7118);
or U10569 (N_10569,N_8263,N_6800);
or U10570 (N_10570,N_5789,N_6236);
nor U10571 (N_10571,N_5885,N_8259);
and U10572 (N_10572,N_6139,N_8072);
and U10573 (N_10573,N_9168,N_8925);
nor U10574 (N_10574,N_6038,N_8985);
nand U10575 (N_10575,N_6248,N_7114);
xnor U10576 (N_10576,N_7253,N_7077);
or U10577 (N_10577,N_6158,N_6129);
xor U10578 (N_10578,N_8936,N_6436);
nand U10579 (N_10579,N_6743,N_9412);
xnor U10580 (N_10580,N_7386,N_6311);
and U10581 (N_10581,N_9341,N_9779);
or U10582 (N_10582,N_7811,N_5850);
or U10583 (N_10583,N_8213,N_5854);
and U10584 (N_10584,N_5582,N_9370);
or U10585 (N_10585,N_8677,N_9551);
and U10586 (N_10586,N_8254,N_8654);
nand U10587 (N_10587,N_7492,N_7428);
and U10588 (N_10588,N_9051,N_7385);
nor U10589 (N_10589,N_7094,N_8439);
nor U10590 (N_10590,N_5836,N_8143);
and U10591 (N_10591,N_7703,N_6927);
nor U10592 (N_10592,N_9916,N_9196);
or U10593 (N_10593,N_8053,N_9809);
and U10594 (N_10594,N_5481,N_6695);
and U10595 (N_10595,N_5141,N_6135);
and U10596 (N_10596,N_7798,N_9981);
or U10597 (N_10597,N_5725,N_7306);
nand U10598 (N_10598,N_5720,N_8116);
and U10599 (N_10599,N_5489,N_9692);
and U10600 (N_10600,N_6682,N_5760);
or U10601 (N_10601,N_8660,N_8035);
nor U10602 (N_10602,N_8766,N_5484);
nand U10603 (N_10603,N_7132,N_5510);
nand U10604 (N_10604,N_6893,N_6443);
and U10605 (N_10605,N_7696,N_8157);
nand U10606 (N_10606,N_7784,N_8314);
and U10607 (N_10607,N_9275,N_8817);
nand U10608 (N_10608,N_6600,N_6991);
or U10609 (N_10609,N_5240,N_7165);
or U10610 (N_10610,N_5171,N_6650);
and U10611 (N_10611,N_7153,N_5315);
nand U10612 (N_10612,N_8665,N_7190);
and U10613 (N_10613,N_6671,N_5270);
nor U10614 (N_10614,N_9328,N_5451);
xnor U10615 (N_10615,N_9181,N_8417);
nor U10616 (N_10616,N_8604,N_8199);
nand U10617 (N_10617,N_8924,N_9429);
nor U10618 (N_10618,N_8855,N_5165);
nor U10619 (N_10619,N_6325,N_6753);
or U10620 (N_10620,N_7865,N_8080);
and U10621 (N_10621,N_8803,N_8338);
and U10622 (N_10622,N_8897,N_7509);
nor U10623 (N_10623,N_9976,N_6055);
and U10624 (N_10624,N_9128,N_9287);
and U10625 (N_10625,N_7423,N_6210);
nor U10626 (N_10626,N_6895,N_8871);
or U10627 (N_10627,N_9741,N_5766);
and U10628 (N_10628,N_5246,N_8602);
and U10629 (N_10629,N_6909,N_6039);
nand U10630 (N_10630,N_5862,N_6417);
nand U10631 (N_10631,N_5280,N_7317);
nand U10632 (N_10632,N_7133,N_7359);
nand U10633 (N_10633,N_8630,N_9777);
nand U10634 (N_10634,N_5565,N_5410);
nor U10635 (N_10635,N_9266,N_7643);
nand U10636 (N_10636,N_5260,N_7790);
xor U10637 (N_10637,N_8658,N_7805);
or U10638 (N_10638,N_8650,N_7060);
nor U10639 (N_10639,N_6694,N_5587);
nand U10640 (N_10640,N_9889,N_5268);
nand U10641 (N_10641,N_7183,N_9756);
xnor U10642 (N_10642,N_9245,N_8573);
or U10643 (N_10643,N_8239,N_7297);
nor U10644 (N_10644,N_9676,N_7841);
nand U10645 (N_10645,N_6160,N_8446);
nor U10646 (N_10646,N_9104,N_5551);
and U10647 (N_10647,N_8527,N_8234);
and U10648 (N_10648,N_5600,N_8248);
or U10649 (N_10649,N_9647,N_5001);
or U10650 (N_10650,N_7722,N_6657);
nor U10651 (N_10651,N_7971,N_9826);
and U10652 (N_10652,N_6975,N_8243);
nand U10653 (N_10653,N_6807,N_9730);
xor U10654 (N_10654,N_8631,N_7246);
and U10655 (N_10655,N_8642,N_9538);
and U10656 (N_10656,N_8829,N_5530);
and U10657 (N_10657,N_8297,N_5866);
and U10658 (N_10658,N_6114,N_9720);
or U10659 (N_10659,N_5494,N_8398);
or U10660 (N_10660,N_6290,N_7511);
and U10661 (N_10661,N_5156,N_9743);
nor U10662 (N_10662,N_9939,N_9229);
nor U10663 (N_10663,N_9293,N_8730);
nor U10664 (N_10664,N_8571,N_8579);
or U10665 (N_10665,N_6312,N_5952);
nand U10666 (N_10666,N_9310,N_7871);
nand U10667 (N_10667,N_5458,N_6030);
or U10668 (N_10668,N_8950,N_8448);
nor U10669 (N_10669,N_8106,N_6837);
or U10670 (N_10670,N_5512,N_7144);
nor U10671 (N_10671,N_9547,N_5201);
nor U10672 (N_10672,N_8357,N_5124);
and U10673 (N_10673,N_6484,N_9877);
nand U10674 (N_10674,N_6148,N_5460);
xnor U10675 (N_10675,N_7466,N_5537);
nor U10676 (N_10676,N_7508,N_8721);
nand U10677 (N_10677,N_6430,N_7842);
nor U10678 (N_10678,N_7970,N_5983);
xnor U10679 (N_10679,N_5805,N_5618);
xnor U10680 (N_10680,N_6138,N_8000);
or U10681 (N_10681,N_6702,N_8142);
and U10682 (N_10682,N_9774,N_9919);
or U10683 (N_10683,N_6322,N_9823);
nand U10684 (N_10684,N_8989,N_7958);
nand U10685 (N_10685,N_5065,N_6037);
xnor U10686 (N_10686,N_6031,N_9037);
or U10687 (N_10687,N_6614,N_7036);
nor U10688 (N_10688,N_8963,N_7488);
or U10689 (N_10689,N_6757,N_6994);
and U10690 (N_10690,N_9996,N_8763);
and U10691 (N_10691,N_9280,N_6061);
or U10692 (N_10692,N_7574,N_7724);
nand U10693 (N_10693,N_7237,N_9786);
or U10694 (N_10694,N_8233,N_7105);
nor U10695 (N_10695,N_6251,N_5886);
nor U10696 (N_10696,N_9522,N_7926);
nand U10697 (N_10697,N_9207,N_8208);
nand U10698 (N_10698,N_8980,N_6284);
nor U10699 (N_10699,N_8947,N_9731);
nor U10700 (N_10700,N_7350,N_8094);
or U10701 (N_10701,N_6056,N_9921);
and U10702 (N_10702,N_9719,N_9500);
nor U10703 (N_10703,N_5594,N_8787);
or U10704 (N_10704,N_5767,N_5990);
and U10705 (N_10705,N_6797,N_6596);
nor U10706 (N_10706,N_9333,N_8902);
or U10707 (N_10707,N_5577,N_9447);
nor U10708 (N_10708,N_7894,N_9030);
or U10709 (N_10709,N_6487,N_7366);
or U10710 (N_10710,N_5126,N_8968);
nor U10711 (N_10711,N_9772,N_9867);
nand U10712 (N_10712,N_5635,N_7983);
or U10713 (N_10713,N_5091,N_6928);
or U10714 (N_10714,N_8609,N_6374);
and U10715 (N_10715,N_5330,N_7056);
nand U10716 (N_10716,N_7814,N_8455);
or U10717 (N_10717,N_6116,N_8893);
nand U10718 (N_10718,N_7642,N_7325);
or U10719 (N_10719,N_5414,N_6368);
and U10720 (N_10720,N_8744,N_8168);
and U10721 (N_10721,N_7949,N_5021);
nor U10722 (N_10722,N_5811,N_9392);
or U10723 (N_10723,N_6429,N_6864);
nor U10724 (N_10724,N_8496,N_6224);
xor U10725 (N_10725,N_6549,N_7180);
nor U10726 (N_10726,N_7502,N_7198);
or U10727 (N_10727,N_9257,N_6400);
and U10728 (N_10728,N_5685,N_6200);
or U10729 (N_10729,N_6589,N_5262);
and U10730 (N_10730,N_9340,N_8471);
nand U10731 (N_10731,N_7685,N_6252);
nor U10732 (N_10732,N_9074,N_6618);
nor U10733 (N_10733,N_5933,N_7820);
or U10734 (N_10734,N_6000,N_7882);
nor U10735 (N_10735,N_5364,N_5334);
and U10736 (N_10736,N_6188,N_8285);
nor U10737 (N_10737,N_5973,N_8881);
nor U10738 (N_10738,N_6641,N_8576);
or U10739 (N_10739,N_9645,N_9406);
xnor U10740 (N_10740,N_7085,N_9353);
nor U10741 (N_10741,N_5930,N_7053);
xor U10742 (N_10742,N_5544,N_9670);
or U10743 (N_10743,N_6696,N_8336);
or U10744 (N_10744,N_6921,N_6545);
nand U10745 (N_10745,N_6326,N_8065);
nor U10746 (N_10746,N_8655,N_8765);
and U10747 (N_10747,N_9430,N_7725);
and U10748 (N_10748,N_6688,N_7070);
and U10749 (N_10749,N_9345,N_7048);
and U10750 (N_10750,N_9270,N_9662);
and U10751 (N_10751,N_7251,N_8684);
and U10752 (N_10752,N_7591,N_6804);
nor U10753 (N_10753,N_5535,N_5233);
nand U10754 (N_10754,N_8279,N_9054);
nand U10755 (N_10755,N_5589,N_8004);
nor U10756 (N_10756,N_6722,N_8487);
xor U10757 (N_10757,N_7901,N_7160);
xnor U10758 (N_10758,N_7420,N_8469);
xor U10759 (N_10759,N_6701,N_5871);
or U10760 (N_10760,N_6725,N_5319);
and U10761 (N_10761,N_6932,N_5439);
and U10762 (N_10762,N_7892,N_7072);
or U10763 (N_10763,N_7793,N_5014);
or U10764 (N_10764,N_9855,N_5486);
nor U10765 (N_10765,N_7040,N_7776);
nor U10766 (N_10766,N_6084,N_8362);
nand U10767 (N_10767,N_5666,N_8624);
nand U10768 (N_10768,N_5566,N_9325);
or U10769 (N_10769,N_7126,N_6440);
xor U10770 (N_10770,N_8731,N_9580);
nand U10771 (N_10771,N_6085,N_7163);
and U10772 (N_10772,N_5213,N_9617);
or U10773 (N_10773,N_9361,N_6289);
or U10774 (N_10774,N_6557,N_8086);
and U10775 (N_10775,N_9521,N_9089);
or U10776 (N_10776,N_9874,N_9849);
nor U10777 (N_10777,N_5289,N_5806);
and U10778 (N_10778,N_8304,N_7797);
and U10779 (N_10779,N_6062,N_9195);
and U10780 (N_10780,N_8735,N_7788);
xor U10781 (N_10781,N_8160,N_5667);
or U10782 (N_10782,N_7716,N_6101);
xnor U10783 (N_10783,N_6707,N_8841);
or U10784 (N_10784,N_8669,N_7059);
nand U10785 (N_10785,N_6534,N_6966);
or U10786 (N_10786,N_6530,N_8465);
and U10787 (N_10787,N_9481,N_5511);
xnor U10788 (N_10788,N_8190,N_8371);
or U10789 (N_10789,N_7017,N_5994);
nor U10790 (N_10790,N_6872,N_9254);
or U10791 (N_10791,N_8791,N_7991);
and U10792 (N_10792,N_5422,N_8724);
and U10793 (N_10793,N_7422,N_7919);
xor U10794 (N_10794,N_6693,N_6892);
or U10795 (N_10795,N_8929,N_8015);
and U10796 (N_10796,N_6608,N_6177);
nor U10797 (N_10797,N_7307,N_6480);
xnor U10798 (N_10798,N_5224,N_9305);
and U10799 (N_10799,N_7719,N_8271);
nand U10800 (N_10800,N_6098,N_7738);
and U10801 (N_10801,N_6013,N_9800);
or U10802 (N_10802,N_5801,N_9592);
or U10803 (N_10803,N_6145,N_8826);
or U10804 (N_10804,N_7864,N_5532);
nor U10805 (N_10805,N_5468,N_5907);
and U10806 (N_10806,N_7521,N_9214);
nand U10807 (N_10807,N_6332,N_6216);
and U10808 (N_10808,N_9554,N_8847);
nand U10809 (N_10809,N_9175,N_9799);
or U10810 (N_10810,N_8568,N_8538);
nand U10811 (N_10811,N_5817,N_6851);
nor U10812 (N_10812,N_9652,N_7935);
xor U10813 (N_10813,N_9658,N_9689);
nand U10814 (N_10814,N_9187,N_8196);
and U10815 (N_10815,N_5123,N_5225);
and U10816 (N_10816,N_9839,N_8934);
or U10817 (N_10817,N_6741,N_9966);
or U10818 (N_10818,N_8009,N_7303);
or U10819 (N_10819,N_8899,N_7021);
nor U10820 (N_10820,N_9987,N_7296);
xor U10821 (N_10821,N_7904,N_9265);
nor U10822 (N_10822,N_7095,N_6333);
nor U10823 (N_10823,N_5938,N_7600);
nand U10824 (N_10824,N_8940,N_8612);
nand U10825 (N_10825,N_5691,N_6414);
and U10826 (N_10826,N_6300,N_8680);
and U10827 (N_10827,N_6751,N_5129);
nand U10828 (N_10828,N_9189,N_7120);
and U10829 (N_10829,N_5833,N_9458);
and U10830 (N_10830,N_5773,N_9776);
nand U10831 (N_10831,N_9306,N_8443);
xor U10832 (N_10832,N_6022,N_9525);
nand U10833 (N_10833,N_9262,N_5496);
nor U10834 (N_10834,N_9478,N_6754);
or U10835 (N_10835,N_5324,N_9022);
and U10836 (N_10836,N_7667,N_5620);
nand U10837 (N_10837,N_7836,N_5713);
nand U10838 (N_10838,N_8076,N_7568);
or U10839 (N_10839,N_5974,N_5075);
and U10840 (N_10840,N_7119,N_9206);
and U10841 (N_10841,N_9057,N_6065);
nor U10842 (N_10842,N_6102,N_7839);
nand U10843 (N_10843,N_8701,N_6249);
nor U10844 (N_10844,N_6790,N_6259);
nand U10845 (N_10845,N_8406,N_6439);
nand U10846 (N_10846,N_6345,N_7620);
nor U10847 (N_10847,N_5397,N_5234);
nor U10848 (N_10848,N_6559,N_9906);
nor U10849 (N_10849,N_6658,N_7782);
and U10850 (N_10850,N_5149,N_7876);
or U10851 (N_10851,N_7329,N_6611);
nand U10852 (N_10852,N_7024,N_5989);
nor U10853 (N_10853,N_6553,N_6667);
nor U10854 (N_10854,N_9871,N_8392);
or U10855 (N_10855,N_6232,N_7006);
nand U10856 (N_10856,N_6471,N_8282);
nand U10857 (N_10857,N_5743,N_7880);
nand U10858 (N_10858,N_9140,N_5633);
or U10859 (N_10859,N_9161,N_8324);
nand U10860 (N_10860,N_7520,N_6548);
nor U10861 (N_10861,N_5596,N_9233);
nand U10862 (N_10862,N_6381,N_8553);
and U10863 (N_10863,N_6555,N_8063);
nand U10864 (N_10864,N_9840,N_6394);
nand U10865 (N_10865,N_6599,N_5876);
xnor U10866 (N_10866,N_6812,N_8360);
and U10867 (N_10867,N_7353,N_7443);
nor U10868 (N_10868,N_6560,N_7735);
nor U10869 (N_10869,N_7497,N_6550);
or U10870 (N_10870,N_8955,N_8375);
and U10871 (N_10871,N_8020,N_7291);
nand U10872 (N_10872,N_9383,N_6714);
nor U10873 (N_10873,N_5231,N_9622);
or U10874 (N_10874,N_7564,N_8129);
and U10875 (N_10875,N_8746,N_6043);
and U10876 (N_10876,N_7004,N_6235);
nor U10877 (N_10877,N_5019,N_9339);
nand U10878 (N_10878,N_7913,N_6406);
nor U10879 (N_10879,N_5726,N_7887);
nand U10880 (N_10880,N_5453,N_9913);
or U10881 (N_10881,N_5851,N_7456);
nand U10882 (N_10882,N_9813,N_5053);
nand U10883 (N_10883,N_8451,N_5506);
nand U10884 (N_10884,N_9451,N_5183);
xor U10885 (N_10885,N_6153,N_9529);
xor U10886 (N_10886,N_6493,N_8742);
nor U10887 (N_10887,N_9077,N_7796);
nand U10888 (N_10888,N_6112,N_9228);
nand U10889 (N_10889,N_9801,N_6780);
nand U10890 (N_10890,N_7714,N_6411);
and U10891 (N_10891,N_5493,N_6297);
nand U10892 (N_10892,N_6242,N_6011);
nor U10893 (N_10893,N_9725,N_9524);
nand U10894 (N_10894,N_6423,N_8879);
and U10895 (N_10895,N_8247,N_9184);
nor U10896 (N_10896,N_7319,N_5829);
or U10897 (N_10897,N_6458,N_9496);
and U10898 (N_10898,N_6226,N_7404);
nand U10899 (N_10899,N_5533,N_5015);
nand U10900 (N_10900,N_8999,N_7729);
nor U10901 (N_10901,N_6704,N_9010);
or U10902 (N_10902,N_6996,N_8813);
and U10903 (N_10903,N_7486,N_5017);
and U10904 (N_10904,N_6187,N_9003);
nor U10905 (N_10905,N_6501,N_5114);
or U10906 (N_10906,N_6877,N_9252);
nor U10907 (N_10907,N_8974,N_7792);
or U10908 (N_10908,N_5634,N_6845);
nand U10909 (N_10909,N_7460,N_9352);
or U10910 (N_10910,N_7030,N_8722);
and U10911 (N_10911,N_8662,N_8379);
nand U10912 (N_10912,N_5963,N_8028);
or U10913 (N_10913,N_7137,N_8530);
and U10914 (N_10914,N_9303,N_8697);
nor U10915 (N_10915,N_7924,N_5557);
nand U10916 (N_10916,N_9408,N_7803);
nor U10917 (N_10917,N_7463,N_6281);
or U10918 (N_10918,N_7517,N_8863);
nand U10919 (N_10919,N_8610,N_6954);
nor U10920 (N_10920,N_7837,N_5442);
nand U10921 (N_10921,N_6169,N_7467);
and U10922 (N_10922,N_5088,N_7593);
nand U10923 (N_10923,N_5103,N_8558);
nor U10924 (N_10924,N_5900,N_6124);
xnor U10925 (N_10925,N_5794,N_8964);
or U10926 (N_10926,N_7425,N_5861);
nand U10927 (N_10927,N_6204,N_6841);
and U10928 (N_10928,N_9244,N_7214);
or U10929 (N_10929,N_8833,N_9631);
nor U10930 (N_10930,N_5927,N_5731);
xor U10931 (N_10931,N_5366,N_6942);
or U10932 (N_10932,N_8434,N_5578);
nand U10933 (N_10933,N_5581,N_5774);
nand U10934 (N_10934,N_5536,N_7647);
nand U10935 (N_10935,N_8269,N_7536);
nand U10936 (N_10936,N_6512,N_7206);
nand U10937 (N_10937,N_8981,N_5762);
and U10938 (N_10938,N_5718,N_6057);
nand U10939 (N_10939,N_7390,N_6378);
nor U10940 (N_10940,N_8629,N_6871);
and U10941 (N_10941,N_5249,N_5893);
xnor U10942 (N_10942,N_5323,N_5682);
and U10943 (N_10943,N_8532,N_6097);
xor U10944 (N_10944,N_7634,N_5687);
nand U10945 (N_10945,N_5172,N_6784);
nor U10946 (N_10946,N_9082,N_5541);
nand U10947 (N_10947,N_6929,N_9267);
nor U10948 (N_10948,N_8867,N_7479);
or U10949 (N_10949,N_9142,N_7636);
xnor U10950 (N_10950,N_9160,N_7821);
nand U10951 (N_10951,N_8715,N_6770);
nor U10952 (N_10952,N_6041,N_5901);
or U10953 (N_10953,N_8156,N_8906);
and U10954 (N_10954,N_8056,N_5367);
or U10955 (N_10955,N_9258,N_6477);
or U10956 (N_10956,N_8203,N_7985);
nand U10957 (N_10957,N_9176,N_7911);
nand U10958 (N_10958,N_6516,N_7465);
xnor U10959 (N_10959,N_9501,N_9682);
nand U10960 (N_10960,N_6651,N_7721);
nand U10961 (N_10961,N_8165,N_7682);
nand U10962 (N_10962,N_6791,N_7220);
nor U10963 (N_10963,N_7980,N_7401);
and U10964 (N_10964,N_6866,N_9250);
and U10965 (N_10965,N_6064,N_5155);
or U10966 (N_10966,N_9103,N_9271);
and U10967 (N_10967,N_9431,N_5584);
xnor U10968 (N_10968,N_7020,N_7136);
and U10969 (N_10969,N_8673,N_6661);
nand U10970 (N_10970,N_8422,N_8714);
or U10971 (N_10971,N_5107,N_9912);
xor U10972 (N_10972,N_6706,N_9831);
or U10973 (N_10973,N_5859,N_8848);
nor U10974 (N_10974,N_8686,N_8342);
or U10975 (N_10975,N_5271,N_5024);
xor U10976 (N_10976,N_5748,N_9885);
and U10977 (N_10977,N_8348,N_8402);
and U10978 (N_10978,N_8408,N_5148);
or U10979 (N_10979,N_7875,N_6537);
nor U10980 (N_10980,N_8797,N_7769);
and U10981 (N_10981,N_9884,N_6142);
or U10982 (N_10982,N_7182,N_8470);
xnor U10983 (N_10983,N_8104,N_6255);
nor U10984 (N_10984,N_5802,N_8885);
nor U10985 (N_10985,N_8997,N_6146);
nor U10986 (N_10986,N_9460,N_5727);
or U10987 (N_10987,N_8623,N_7860);
nand U10988 (N_10988,N_5756,N_6699);
and U10989 (N_10989,N_5984,N_8003);
xor U10990 (N_10990,N_8103,N_7128);
nand U10991 (N_10991,N_5254,N_6341);
or U10992 (N_10992,N_9418,N_7270);
nand U10993 (N_10993,N_5182,N_9998);
xor U10994 (N_10994,N_5474,N_9282);
or U10995 (N_10995,N_9227,N_6888);
nor U10996 (N_10996,N_5853,N_6134);
nor U10997 (N_10997,N_5467,N_6570);
nor U10998 (N_10998,N_8175,N_5947);
and U10999 (N_10999,N_7348,N_5971);
nand U11000 (N_11000,N_9198,N_8151);
or U11001 (N_11001,N_5524,N_9354);
nand U11002 (N_11002,N_6479,N_6310);
and U11003 (N_11003,N_5216,N_6758);
or U11004 (N_11004,N_6518,N_9793);
and U11005 (N_11005,N_7244,N_7653);
or U11006 (N_11006,N_5100,N_5003);
nand U11007 (N_11007,N_6917,N_8853);
nand U11008 (N_11008,N_7637,N_8027);
nand U11009 (N_11009,N_9739,N_5340);
nor U11010 (N_11010,N_8918,N_9778);
nor U11011 (N_11011,N_5175,N_5787);
nor U11012 (N_11012,N_9794,N_5346);
and U11013 (N_11013,N_9042,N_8274);
or U11014 (N_11014,N_9628,N_6231);
nor U11015 (N_11015,N_9834,N_7704);
nand U11016 (N_11016,N_8217,N_9025);
nand U11017 (N_11017,N_6444,N_7708);
nor U11018 (N_11018,N_7438,N_9864);
xor U11019 (N_11019,N_6785,N_6593);
nor U11020 (N_11020,N_7552,N_6513);
xor U11021 (N_11021,N_5306,N_9041);
or U11022 (N_11022,N_7853,N_5479);
xor U11023 (N_11023,N_9681,N_6551);
nor U11024 (N_11024,N_7819,N_9616);
nor U11025 (N_11025,N_8557,N_5352);
nand U11026 (N_11026,N_5521,N_6507);
nor U11027 (N_11027,N_5653,N_9085);
and U11028 (N_11028,N_5915,N_7449);
or U11029 (N_11029,N_5035,N_5549);
or U11030 (N_11030,N_9893,N_6025);
and U11031 (N_11031,N_5781,N_6983);
nor U11032 (N_11032,N_8778,N_8110);
and U11033 (N_11033,N_9510,N_5022);
or U11034 (N_11034,N_5239,N_9484);
xnor U11035 (N_11035,N_5538,N_7014);
xor U11036 (N_11036,N_9283,N_7752);
and U11037 (N_11037,N_8814,N_6103);
and U11038 (N_11038,N_6437,N_9955);
xor U11039 (N_11039,N_8178,N_5934);
nor U11040 (N_11040,N_9697,N_9568);
nand U11041 (N_11041,N_8777,N_5563);
and U11042 (N_11042,N_6234,N_6233);
xnor U11043 (N_11043,N_9937,N_7939);
nand U11044 (N_11044,N_6175,N_7810);
and U11045 (N_11045,N_7741,N_5153);
nand U11046 (N_11046,N_6673,N_8832);
nand U11047 (N_11047,N_6180,N_5956);
or U11048 (N_11048,N_7686,N_9520);
or U11049 (N_11049,N_6982,N_6637);
nand U11050 (N_11050,N_9561,N_6476);
nor U11051 (N_11051,N_9061,N_8079);
nand U11052 (N_11052,N_5858,N_7542);
or U11053 (N_11053,N_9519,N_5797);
nand U11054 (N_11054,N_5173,N_7065);
or U11055 (N_11055,N_9736,N_5513);
or U11056 (N_11056,N_6970,N_9048);
nand U11057 (N_11057,N_5351,N_9747);
nor U11058 (N_11058,N_5369,N_6817);
and U11059 (N_11059,N_7293,N_9137);
and U11060 (N_11060,N_9515,N_9887);
nand U11061 (N_11061,N_9815,N_7388);
nand U11062 (N_11062,N_6666,N_6612);
nand U11063 (N_11063,N_5728,N_5906);
and U11064 (N_11064,N_5860,N_7966);
nor U11065 (N_11065,N_9382,N_5006);
nor U11066 (N_11066,N_8453,N_9947);
nand U11067 (N_11067,N_8403,N_7931);
nand U11068 (N_11068,N_5981,N_9728);
nor U11069 (N_11069,N_9024,N_9177);
nor U11070 (N_11070,N_8411,N_5228);
or U11071 (N_11071,N_8755,N_7712);
nand U11072 (N_11072,N_6624,N_7242);
nor U11073 (N_11073,N_9454,N_6742);
nor U11074 (N_11074,N_6319,N_8838);
xor U11075 (N_11075,N_7416,N_5332);
nand U11076 (N_11076,N_9337,N_8801);
xnor U11077 (N_11077,N_5693,N_9380);
nand U11078 (N_11078,N_9426,N_8531);
xor U11079 (N_11079,N_8377,N_6640);
or U11080 (N_11080,N_7280,N_5991);
nor U11081 (N_11081,N_5217,N_5263);
nand U11082 (N_11082,N_9737,N_6582);
and U11083 (N_11083,N_6461,N_9131);
or U11084 (N_11084,N_7559,N_6852);
and U11085 (N_11085,N_8512,N_7843);
or U11086 (N_11086,N_9795,N_9386);
and U11087 (N_11087,N_8442,N_7394);
nand U11088 (N_11088,N_7824,N_6371);
or U11089 (N_11089,N_9964,N_7720);
nand U11090 (N_11090,N_6850,N_8308);
and U11091 (N_11091,N_7967,N_5267);
nand U11092 (N_11092,N_9579,N_7757);
nor U11093 (N_11093,N_5353,N_6636);
nand U11094 (N_11094,N_6283,N_7736);
nand U11095 (N_11095,N_5146,N_5624);
nor U11096 (N_11096,N_5964,N_6719);
nand U11097 (N_11097,N_8488,N_9404);
nor U11098 (N_11098,N_8661,N_6990);
or U11099 (N_11099,N_9461,N_9751);
or U11100 (N_11100,N_5702,N_7489);
and U11101 (N_11101,N_9014,N_5665);
nor U11102 (N_11102,N_9364,N_9713);
nor U11103 (N_11103,N_9302,N_9203);
and U11104 (N_11104,N_7154,N_9504);
and U11105 (N_11105,N_9491,N_6067);
nand U11106 (N_11106,N_6027,N_5238);
and U11107 (N_11107,N_5924,N_5658);
xor U11108 (N_11108,N_7713,N_6848);
nor U11109 (N_11109,N_7968,N_8621);
or U11110 (N_11110,N_5488,N_7512);
nand U11111 (N_11111,N_9865,N_6985);
and U11112 (N_11112,N_9107,N_5707);
nor U11113 (N_11113,N_5747,N_9956);
nor U11114 (N_11114,N_9180,N_8251);
nand U11115 (N_11115,N_7639,N_6412);
or U11116 (N_11116,N_5771,N_6620);
nand U11117 (N_11117,N_5714,N_8519);
nand U11118 (N_11118,N_7727,N_7071);
or U11119 (N_11119,N_8253,N_6239);
and U11120 (N_11120,N_5923,N_8018);
xor U11121 (N_11121,N_8221,N_8310);
nand U11122 (N_11122,N_9264,N_7212);
and U11123 (N_11123,N_9753,N_9127);
nand U11124 (N_11124,N_5034,N_6245);
or U11125 (N_11125,N_9567,N_5662);
nor U11126 (N_11126,N_7749,N_9044);
nand U11127 (N_11127,N_8069,N_8138);
and U11128 (N_11128,N_8659,N_9927);
nor U11129 (N_11129,N_7323,N_6403);
nand U11130 (N_11130,N_5376,N_6335);
and U11131 (N_11131,N_6564,N_5526);
xor U11132 (N_11132,N_7577,N_7321);
nand U11133 (N_11133,N_8905,N_6772);
or U11134 (N_11134,N_5178,N_6026);
and U11135 (N_11135,N_5360,N_8748);
and U11136 (N_11136,N_5293,N_7274);
or U11137 (N_11137,N_7570,N_8584);
or U11138 (N_11138,N_9768,N_5711);
or U11139 (N_11139,N_9959,N_8107);
and U11140 (N_11140,N_5617,N_8635);
or U11141 (N_11141,N_6765,N_9169);
or U11142 (N_11142,N_8820,N_8895);
or U11143 (N_11143,N_7922,N_8052);
nand U11144 (N_11144,N_5619,N_7702);
or U11145 (N_11145,N_7399,N_6705);
nor U11146 (N_11146,N_6426,N_6839);
and U11147 (N_11147,N_6604,N_5018);
nor U11148 (N_11148,N_8012,N_7200);
and U11149 (N_11149,N_9096,N_6143);
or U11150 (N_11150,N_6825,N_7473);
nor U11151 (N_11151,N_8325,N_7135);
or U11152 (N_11152,N_7806,N_7822);
nand U11153 (N_11153,N_9583,N_6147);
and U11154 (N_11154,N_5986,N_7315);
nor U11155 (N_11155,N_8601,N_8024);
nor U11156 (N_11156,N_6836,N_7510);
nor U11157 (N_11157,N_5710,N_8509);
or U11158 (N_11158,N_7612,N_5864);
nand U11159 (N_11159,N_9075,N_7229);
and U11160 (N_11160,N_9482,N_9006);
nand U11161 (N_11161,N_6470,N_8085);
or U11162 (N_11162,N_6167,N_7346);
nor U11163 (N_11163,N_6483,N_5729);
or U11164 (N_11164,N_8982,N_7351);
and U11165 (N_11165,N_9179,N_6238);
and U11166 (N_11166,N_5071,N_8737);
nor U11167 (N_11167,N_6431,N_5701);
nor U11168 (N_11168,N_5455,N_5960);
nor U11169 (N_11169,N_9718,N_7134);
and U11170 (N_11170,N_7266,N_8074);
and U11171 (N_11171,N_7946,N_5089);
and U11172 (N_11172,N_8047,N_6581);
or U11173 (N_11173,N_5375,N_9235);
or U11174 (N_11174,N_9872,N_9726);
xor U11175 (N_11175,N_5445,N_8013);
and U11176 (N_11176,N_7960,N_8501);
nand U11177 (N_11177,N_5348,N_9563);
and U11178 (N_11178,N_5695,N_7309);
nand U11179 (N_11179,N_6454,N_6576);
or U11180 (N_11180,N_9278,N_7625);
nand U11181 (N_11181,N_9759,N_6988);
and U11182 (N_11182,N_6258,N_9071);
nand U11183 (N_11183,N_7365,N_9477);
nand U11184 (N_11184,N_6292,N_5813);
nor U11185 (N_11185,N_9892,N_8505);
and U11186 (N_11186,N_8732,N_6166);
and U11187 (N_11187,N_8477,N_7937);
or U11188 (N_11188,N_5899,N_9710);
and U11189 (N_11189,N_8494,N_7453);
nor U11190 (N_11190,N_9313,N_9605);
and U11191 (N_11191,N_5235,N_5604);
nor U11192 (N_11192,N_6529,N_5199);
nand U11193 (N_11193,N_9194,N_7081);
nand U11194 (N_11194,N_5443,N_8693);
or U11195 (N_11195,N_7870,N_9058);
and U11196 (N_11196,N_7408,N_5783);
nor U11197 (N_11197,N_9165,N_9597);
xor U11198 (N_11198,N_8158,N_8413);
and U11199 (N_11199,N_7832,N_6561);
nor U11200 (N_11200,N_5739,N_5540);
or U11201 (N_11201,N_9385,N_6199);
nand U11202 (N_11202,N_5895,N_6773);
nor U11203 (N_11203,N_5080,N_5622);
nor U11204 (N_11204,N_6997,N_5063);
nor U11205 (N_11205,N_7936,N_6473);
nor U11206 (N_11206,N_6481,N_8033);
nor U11207 (N_11207,N_5138,N_9780);
nor U11208 (N_11208,N_7833,N_6712);
nand U11209 (N_11209,N_5256,N_9147);
xor U11210 (N_11210,N_6126,N_8595);
xor U11211 (N_11211,N_8389,N_6107);
xor U11212 (N_11212,N_8995,N_7167);
nand U11213 (N_11213,N_6827,N_7336);
and U11214 (N_11214,N_8386,N_6434);
nand U11215 (N_11215,N_6958,N_9236);
nand U11216 (N_11216,N_5200,N_6798);
nand U11217 (N_11217,N_7730,N_6358);
nand U11218 (N_11218,N_9980,N_5884);
and U11219 (N_11219,N_9802,N_8475);
nand U11220 (N_11220,N_6857,N_7592);
nand U11221 (N_11221,N_8339,N_9379);
and U11222 (N_11222,N_6407,N_7872);
nand U11223 (N_11223,N_9413,N_6733);
or U11224 (N_11224,N_7483,N_9656);
nor U11225 (N_11225,N_9047,N_5426);
nor U11226 (N_11226,N_9653,N_5250);
nor U11227 (N_11227,N_5715,N_8580);
or U11228 (N_11228,N_8711,N_9263);
or U11229 (N_11229,N_7038,N_8154);
xnor U11230 (N_11230,N_7412,N_6413);
and U11231 (N_11231,N_6951,N_9069);
xnor U11232 (N_11232,N_6464,N_8712);
and U11233 (N_11233,N_5967,N_7454);
and U11234 (N_11234,N_8806,N_5038);
xnor U11235 (N_11235,N_8205,N_5051);
nor U11236 (N_11236,N_8524,N_7587);
or U11237 (N_11237,N_8121,N_9422);
nor U11238 (N_11238,N_6137,N_8493);
nand U11239 (N_11239,N_9032,N_5550);
or U11240 (N_11240,N_8300,N_6977);
nand U11241 (N_11241,N_8194,N_5408);
and U11242 (N_11242,N_5215,N_5746);
or U11243 (N_11243,N_5775,N_5892);
xnor U11244 (N_11244,N_8577,N_9381);
nor U11245 (N_11245,N_8139,N_8095);
nor U11246 (N_11246,N_8747,N_7874);
and U11247 (N_11247,N_6282,N_8834);
or U11248 (N_11248,N_8037,N_5184);
nand U11249 (N_11249,N_7213,N_9534);
nand U11250 (N_11250,N_7795,N_7866);
nor U11251 (N_11251,N_9369,N_9752);
nand U11252 (N_11252,N_5569,N_5966);
nand U11253 (N_11253,N_8570,N_6069);
nand U11254 (N_11254,N_6731,N_9569);
nand U11255 (N_11255,N_7532,N_7358);
or U11256 (N_11256,N_8333,N_5435);
nor U11257 (N_11257,N_9371,N_9427);
or U11258 (N_11258,N_8807,N_9700);
or U11259 (N_11259,N_8096,N_8226);
nand U11260 (N_11260,N_6750,N_5612);
xnor U11261 (N_11261,N_6616,N_5863);
nand U11262 (N_11262,N_5086,N_9092);
or U11263 (N_11263,N_8676,N_8526);
or U11264 (N_11264,N_7829,N_6422);
nand U11265 (N_11265,N_9291,N_9279);
xnor U11266 (N_11266,N_9163,N_5880);
nor U11267 (N_11267,N_7238,N_8944);
or U11268 (N_11268,N_6214,N_9876);
and U11269 (N_11269,N_7844,N_5406);
nor U11270 (N_11270,N_6438,N_9553);
nand U11271 (N_11271,N_8767,N_9208);
nor U11272 (N_11272,N_7415,N_9153);
and U11273 (N_11273,N_9115,N_7885);
nor U11274 (N_11274,N_5269,N_9008);
nor U11275 (N_11275,N_9977,N_8421);
xor U11276 (N_11276,N_8808,N_8926);
xnor U11277 (N_11277,N_8128,N_5054);
and U11278 (N_11278,N_7575,N_5778);
and U11279 (N_11279,N_8083,N_7421);
and U11280 (N_11280,N_7534,N_5033);
nand U11281 (N_11281,N_9836,N_5918);
nand U11282 (N_11282,N_6535,N_9272);
nand U11283 (N_11283,N_6372,N_6424);
nor U11284 (N_11284,N_7409,N_5345);
nand U11285 (N_11285,N_7563,N_8202);
nor U11286 (N_11286,N_9403,N_9442);
nor U11287 (N_11287,N_5379,N_7981);
or U11288 (N_11288,N_6253,N_5321);
nand U11289 (N_11289,N_5957,N_6993);
or U11290 (N_11290,N_7115,N_8039);
xnor U11291 (N_11291,N_9953,N_7774);
or U11292 (N_11292,N_8145,N_5621);
nand U11293 (N_11293,N_5401,N_8230);
nand U11294 (N_11294,N_6677,N_8923);
and U11295 (N_11295,N_7172,N_5363);
nand U11296 (N_11296,N_7928,N_9543);
and U11297 (N_11297,N_7815,N_9610);
or U11298 (N_11298,N_6856,N_9440);
or U11299 (N_11299,N_8585,N_6801);
or U11300 (N_11300,N_8586,N_5257);
nand U11301 (N_11301,N_7450,N_9329);
or U11302 (N_11302,N_6709,N_8166);
and U11303 (N_11303,N_8258,N_8425);
or U11304 (N_11304,N_9842,N_8517);
nand U11305 (N_11305,N_6615,N_7273);
nor U11306 (N_11306,N_8187,N_8332);
and U11307 (N_11307,N_9555,N_5909);
and U11308 (N_11308,N_8682,N_6280);
xnor U11309 (N_11309,N_9678,N_6059);
nor U11310 (N_11310,N_7858,N_8242);
and U11311 (N_11311,N_8261,N_5656);
or U11312 (N_11312,N_7659,N_9256);
nand U11313 (N_11313,N_7173,N_5134);
or U11314 (N_11314,N_5226,N_6348);
nor U11315 (N_11315,N_6074,N_7834);
or U11316 (N_11316,N_9903,N_8270);
nand U11317 (N_11317,N_6499,N_7260);
nand U11318 (N_11318,N_8522,N_5299);
nand U11319 (N_11319,N_6367,N_7631);
nor U11320 (N_11320,N_6489,N_8789);
xnor U11321 (N_11321,N_5668,N_6323);
nor U11322 (N_11322,N_7879,N_7498);
xor U11323 (N_11323,N_7943,N_5179);
or U11324 (N_11324,N_8432,N_6995);
and U11325 (N_11325,N_6879,N_8340);
and U11326 (N_11326,N_5883,N_9900);
or U11327 (N_11327,N_8294,N_7337);
nor U11328 (N_11328,N_8511,N_8720);
nor U11329 (N_11329,N_9342,N_8795);
and U11330 (N_11330,N_9623,N_7177);
or U11331 (N_11331,N_8182,N_7232);
or U11332 (N_11332,N_9215,N_7545);
and U11333 (N_11333,N_9699,N_6151);
nand U11334 (N_11334,N_5005,N_5814);
nor U11335 (N_11335,N_9640,N_6452);
xnor U11336 (N_11336,N_5606,N_5097);
nor U11337 (N_11337,N_8774,N_6352);
and U11338 (N_11338,N_8466,N_5646);
or U11339 (N_11339,N_9210,N_8043);
nand U11340 (N_11340,N_7210,N_5058);
and U11341 (N_11341,N_9238,N_5356);
xor U11342 (N_11342,N_6884,N_5436);
nor U11343 (N_11343,N_8534,N_8596);
and U11344 (N_11344,N_5214,N_6472);
and U11345 (N_11345,N_8860,N_7661);
or U11346 (N_11346,N_7603,N_5810);
or U11347 (N_11347,N_5590,N_8055);
and U11348 (N_11348,N_9446,N_9492);
nor U11349 (N_11349,N_9911,N_6492);
nor U11350 (N_11350,N_7546,N_8727);
xnor U11351 (N_11351,N_7903,N_6511);
or U11352 (N_11352,N_8383,N_7031);
and U11353 (N_11353,N_9292,N_8224);
nand U11354 (N_11354,N_8245,N_6613);
or U11355 (N_11355,N_5135,N_9190);
and U11356 (N_11356,N_8656,N_5487);
and U11357 (N_11357,N_9946,N_6032);
nor U11358 (N_11358,N_5007,N_7802);
or U11359 (N_11359,N_5921,N_5187);
and U11360 (N_11360,N_6089,N_5325);
nand U11361 (N_11361,N_6494,N_7758);
nand U11362 (N_11362,N_5758,N_6100);
nand U11363 (N_11363,N_8170,N_5902);
or U11364 (N_11364,N_6508,N_6448);
or U11365 (N_11365,N_6558,N_8705);
xnor U11366 (N_11366,N_5784,N_6949);
and U11367 (N_11367,N_5750,N_7540);
or U11368 (N_11368,N_5161,N_8358);
or U11369 (N_11369,N_9577,N_6118);
nand U11370 (N_11370,N_6710,N_7779);
or U11371 (N_11371,N_7744,N_8996);
nand U11372 (N_11372,N_5288,N_8979);
and U11373 (N_11373,N_7245,N_9123);
nor U11374 (N_11374,N_9011,N_8637);
xor U11375 (N_11375,N_8391,N_9890);
and U11376 (N_11376,N_6201,N_5868);
or U11377 (N_11377,N_6017,N_8927);
nor U11378 (N_11378,N_6674,N_8220);
nand U11379 (N_11379,N_6973,N_6509);
nor U11380 (N_11380,N_8754,N_9708);
or U11381 (N_11381,N_8237,N_7191);
xnor U11382 (N_11382,N_7398,N_5647);
nor U11383 (N_11383,N_7395,N_9241);
and U11384 (N_11384,N_9436,N_7884);
or U11385 (N_11385,N_5800,N_6605);
or U11386 (N_11386,N_7863,N_5291);
and U11387 (N_11387,N_8435,N_5466);
or U11388 (N_11388,N_9471,N_6959);
xnor U11389 (N_11389,N_9416,N_9070);
and U11390 (N_11390,N_5585,N_6215);
and U11391 (N_11391,N_8550,N_5253);
nand U11392 (N_11392,N_7526,N_5574);
and U11393 (N_11393,N_9742,N_8696);
and U11394 (N_11394,N_9166,N_8082);
nor U11395 (N_11395,N_8943,N_9307);
nand U11396 (N_11396,N_8445,N_7726);
and U11397 (N_11397,N_9738,N_7789);
and U11398 (N_11398,N_8994,N_6670);
xnor U11399 (N_11399,N_7569,N_5602);
nor U11400 (N_11400,N_5473,N_7218);
nor U11401 (N_11401,N_8211,N_8845);
and U11402 (N_11402,N_7751,N_8394);
and U11403 (N_11403,N_8525,N_6218);
nor U11404 (N_11404,N_8307,N_9219);
nand U11405 (N_11405,N_5232,N_7519);
and U11406 (N_11406,N_9129,N_8822);
nand U11407 (N_11407,N_8551,N_9972);
or U11408 (N_11408,N_7695,N_5518);
xnor U11409 (N_11409,N_8288,N_8972);
nor U11410 (N_11410,N_9318,N_5786);
nand U11411 (N_11411,N_5632,N_8218);
nor U11412 (N_11412,N_8395,N_6563);
nand U11413 (N_11413,N_6583,N_6910);
xor U11414 (N_11414,N_6192,N_6938);
nand U11415 (N_11415,N_6350,N_7170);
and U11416 (N_11416,N_8462,N_8365);
or U11417 (N_11417,N_6805,N_9690);
xor U11418 (N_11418,N_9630,N_9560);
nand U11419 (N_11419,N_9607,N_5499);
nor U11420 (N_11420,N_8284,N_7982);
or U11421 (N_11421,N_6653,N_8672);
nand U11422 (N_11422,N_8441,N_9666);
or U11423 (N_11423,N_9420,N_5998);
and U11424 (N_11424,N_8836,N_6447);
nand U11425 (N_11425,N_6739,N_6562);
and U11426 (N_11426,N_5790,N_5447);
nor U11427 (N_11427,N_8319,N_8958);
nand U11428 (N_11428,N_5444,N_6515);
xor U11429 (N_11429,N_6161,N_5641);
or U11430 (N_11430,N_8265,N_9106);
or U11431 (N_11431,N_7912,N_5660);
and U11432 (N_11432,N_9111,N_5763);
or U11433 (N_11433,N_9925,N_7068);
nand U11434 (N_11434,N_6863,N_6818);
nand U11435 (N_11435,N_5398,N_5461);
nand U11436 (N_11436,N_5198,N_7257);
nand U11437 (N_11437,N_8986,N_7092);
and U11438 (N_11438,N_6628,N_7942);
or U11439 (N_11439,N_5652,N_9055);
nor U11440 (N_11440,N_7818,N_6896);
nor U11441 (N_11441,N_7826,N_5042);
and U11442 (N_11442,N_9497,N_7008);
or U11443 (N_11443,N_8798,N_7459);
and U11444 (N_11444,N_6632,N_7893);
nand U11445 (N_11445,N_8022,N_7369);
nand U11446 (N_11446,N_6342,N_8619);
and U11447 (N_11447,N_7900,N_8038);
and U11448 (N_11448,N_5151,N_9338);
nand U11449 (N_11449,N_5434,N_6847);
nand U11450 (N_11450,N_9635,N_9789);
nor U11451 (N_11451,N_8668,N_7076);
nand U11452 (N_11452,N_5105,N_7986);
or U11453 (N_11453,N_5294,N_7455);
and U11454 (N_11454,N_7663,N_7352);
nor U11455 (N_11455,N_9050,N_9218);
nand U11456 (N_11456,N_6194,N_6115);
nor U11457 (N_11457,N_6072,N_9750);
or U11458 (N_11458,N_5593,N_9045);
nor U11459 (N_11459,N_8865,N_5040);
nand U11460 (N_11460,N_6002,N_6221);
nor U11461 (N_11461,N_5559,N_6005);
or U11462 (N_11462,N_6401,N_5266);
or U11463 (N_11463,N_9157,N_6263);
xor U11464 (N_11464,N_6679,N_5092);
nor U11465 (N_11465,N_9746,N_9411);
nor U11466 (N_11466,N_9251,N_7087);
and U11467 (N_11467,N_6343,N_6244);
nand U11468 (N_11468,N_5699,N_5450);
or U11469 (N_11469,N_6405,N_8153);
nand U11470 (N_11470,N_8238,N_6749);
xor U11471 (N_11471,N_7152,N_9171);
and U11472 (N_11472,N_6934,N_9895);
nand U11473 (N_11473,N_9298,N_9213);
nand U11474 (N_11474,N_5070,N_6125);
and U11475 (N_11475,N_8401,N_5570);
nand U11476 (N_11476,N_9897,N_6987);
nand U11477 (N_11477,N_9086,N_9915);
nand U11478 (N_11478,N_8904,N_7196);
and U11479 (N_11479,N_6729,N_9936);
and U11480 (N_11480,N_5846,N_6278);
or U11481 (N_11481,N_6418,N_6646);
and U11482 (N_11482,N_8289,N_6919);
xor U11483 (N_11483,N_8636,N_5326);
or U11484 (N_11484,N_9850,N_7561);
nand U11485 (N_11485,N_8497,N_8147);
nand U11486 (N_11486,N_8607,N_9034);
and U11487 (N_11487,N_6463,N_5809);
nor U11488 (N_11488,N_6336,N_6814);
or U11489 (N_11489,N_5688,N_7043);
or U11490 (N_11490,N_6140,N_6967);
nor U11491 (N_11491,N_7551,N_9922);
or U11492 (N_11492,N_5822,N_6363);
and U11493 (N_11493,N_9783,N_6734);
nor U11494 (N_11494,N_5920,N_7669);
xor U11495 (N_11495,N_7189,N_9712);
nand U11496 (N_11496,N_7342,N_6881);
or U11497 (N_11497,N_7905,N_8583);
and U11498 (N_11498,N_6122,N_9255);
and U11499 (N_11499,N_9023,N_9099);
nand U11500 (N_11500,N_5615,N_7657);
or U11501 (N_11501,N_8467,N_9087);
nand U11502 (N_11502,N_9556,N_7155);
xor U11503 (N_11503,N_9804,N_8134);
or U11504 (N_11504,N_7243,N_7616);
and U11505 (N_11505,N_9971,N_9360);
nor U11506 (N_11506,N_7709,N_6930);
xor U11507 (N_11507,N_5207,N_6346);
nor U11508 (N_11508,N_6482,N_6058);
and U11509 (N_11509,N_9625,N_8374);
or U11510 (N_11510,N_8320,N_9004);
nor U11511 (N_11511,N_7925,N_5010);
nor U11512 (N_11512,N_7334,N_8478);
or U11513 (N_11513,N_8818,N_8222);
and U11514 (N_11514,N_8873,N_7357);
xnor U11515 (N_11515,N_5251,N_6380);
nor U11516 (N_11516,N_8250,N_9675);
or U11517 (N_11517,N_9633,N_9909);
nor U11518 (N_11518,N_7747,N_7940);
nor U11519 (N_11519,N_8231,N_8892);
or U11520 (N_11520,N_8703,N_6243);
and U11521 (N_11521,N_7809,N_5564);
nor U11522 (N_11522,N_6357,N_6585);
nand U11523 (N_11523,N_5358,N_9231);
xor U11524 (N_11524,N_8454,N_6295);
and U11525 (N_11525,N_5012,N_7648);
or U11526 (N_11526,N_9642,N_5274);
nor U11527 (N_11527,N_7387,N_9433);
nor U11528 (N_11528,N_6573,N_7638);
nand U11529 (N_11529,N_8125,N_8148);
nor U11530 (N_11530,N_9512,N_5608);
nor U11531 (N_11531,N_7207,N_5307);
nand U11532 (N_11532,N_9566,N_6952);
or U11533 (N_11533,N_5387,N_9923);
and U11534 (N_11534,N_6580,N_5061);
and U11535 (N_11535,N_5099,N_9940);
nand U11536 (N_11536,N_7067,N_5505);
and U11537 (N_11537,N_5792,N_8407);
and U11538 (N_11538,N_9539,N_8223);
nand U11539 (N_11539,N_6762,N_5932);
nor U11540 (N_11540,N_6865,N_5821);
nor U11541 (N_11541,N_6318,N_9289);
nor U11542 (N_11542,N_6427,N_8216);
xnor U11543 (N_11543,N_6894,N_7281);
and U11544 (N_11544,N_8173,N_8468);
and U11545 (N_11545,N_5597,N_8887);
nor U11546 (N_11546,N_9810,N_5255);
and U11547 (N_11547,N_7524,N_6940);
nand U11548 (N_11548,N_8317,N_8515);
nand U11549 (N_11549,N_7655,N_8772);
or U11550 (N_11550,N_5218,N_6392);
nor U11551 (N_11551,N_6207,N_5678);
and U11552 (N_11552,N_9314,N_7693);
nand U11553 (N_11553,N_9933,N_7063);
nand U11554 (N_11554,N_9650,N_9581);
or U11555 (N_11555,N_7507,N_7199);
or U11556 (N_11556,N_8334,N_6305);
and U11557 (N_11557,N_5144,N_7254);
nor U11558 (N_11558,N_7764,N_8569);
nor U11559 (N_11559,N_9705,N_6094);
or U11560 (N_11560,N_5152,N_6008);
nor U11561 (N_11561,N_8987,N_5872);
and U11562 (N_11562,N_8935,N_8232);
xor U11563 (N_11563,N_6918,N_9226);
and U11564 (N_11564,N_5636,N_9119);
or U11565 (N_11565,N_5096,N_7264);
xor U11566 (N_11566,N_7697,N_8098);
and U11567 (N_11567,N_9654,N_5265);
nor U11568 (N_11568,N_9068,N_7906);
and U11569 (N_11569,N_6874,N_5931);
nand U11570 (N_11570,N_7194,N_6981);
nand U11571 (N_11571,N_6036,N_5698);
nor U11572 (N_11572,N_7626,N_6191);
and U11573 (N_11573,N_8152,N_7299);
xor U11574 (N_11574,N_8556,N_9540);
nand U11575 (N_11575,N_9134,N_7541);
or U11576 (N_11576,N_6404,N_8840);
nand U11577 (N_11577,N_8068,N_6361);
xor U11578 (N_11578,N_6813,N_8118);
or U11579 (N_11579,N_5657,N_7069);
nor U11580 (N_11580,N_7756,N_7854);
nor U11581 (N_11581,N_9791,N_6913);
nand U11582 (N_11582,N_9019,N_9472);
or U11583 (N_11583,N_6291,N_6264);
xor U11584 (N_11584,N_9394,N_9745);
or U11585 (N_11585,N_8293,N_6170);
or U11586 (N_11586,N_9854,N_7310);
and U11587 (N_11587,N_5595,N_7458);
nand U11588 (N_11588,N_9769,N_6211);
nor U11589 (N_11589,N_5661,N_6633);
or U11590 (N_11590,N_6764,N_5371);
nor U11591 (N_11591,N_5654,N_7857);
nor U11592 (N_11592,N_7891,N_9896);
nor U11593 (N_11593,N_6905,N_7930);
and U11594 (N_11594,N_8126,N_6832);
and U11595 (N_11595,N_8633,N_6965);
nor U11596 (N_11596,N_5567,N_5339);
nor U11597 (N_11597,N_7518,N_7623);
xor U11598 (N_11598,N_6010,N_8839);
nand U11599 (N_11599,N_7130,N_9405);
and U11600 (N_11600,N_7608,N_6992);
nand U11601 (N_11601,N_5169,N_7098);
nand U11602 (N_11602,N_7535,N_6539);
and U11603 (N_11603,N_6260,N_8698);
nand U11604 (N_11604,N_5697,N_9667);
nand U11605 (N_11605,N_7446,N_9109);
and U11606 (N_11606,N_6268,N_8123);
or U11607 (N_11607,N_7539,N_7256);
nand U11608 (N_11608,N_5081,N_9688);
nor U11609 (N_11609,N_6601,N_5365);
xnor U11610 (N_11610,N_9960,N_6998);
or U11611 (N_11611,N_6691,N_6531);
and U11612 (N_11612,N_7881,N_8685);
nand U11613 (N_11613,N_7131,N_9060);
and U11614 (N_11614,N_9274,N_7305);
nand U11615 (N_11615,N_6388,N_8611);
xnor U11616 (N_11616,N_5937,N_7271);
and U11617 (N_11617,N_7129,N_8041);
nand U11618 (N_11618,N_8057,N_9620);
nor U11619 (N_11619,N_9239,N_8949);
or U11620 (N_11620,N_5082,N_7338);
xnor U11621 (N_11621,N_6947,N_9881);
nand U11622 (N_11622,N_5645,N_8603);
and U11623 (N_11623,N_6763,N_9209);
nor U11624 (N_11624,N_5432,N_5452);
and U11625 (N_11625,N_8244,N_6598);
and U11626 (N_11626,N_8135,N_9999);
or U11627 (N_11627,N_7413,N_8112);
nand U11628 (N_11628,N_7525,N_9858);
and U11629 (N_11629,N_7580,N_7740);
and U11630 (N_11630,N_7345,N_6117);
and U11631 (N_11631,N_8159,N_9193);
nor U11632 (N_11632,N_9173,N_7908);
or U11633 (N_11633,N_7763,N_5059);
or U11634 (N_11634,N_9143,N_9659);
nor U11635 (N_11635,N_6016,N_6163);
or U11636 (N_11636,N_8666,N_5503);
xnor U11637 (N_11637,N_6543,N_8460);
nand U11638 (N_11638,N_9199,N_7684);
nor U11639 (N_11639,N_9644,N_9901);
or U11640 (N_11640,N_7029,N_6186);
and U11641 (N_11641,N_7945,N_7461);
or U11642 (N_11642,N_5926,N_9148);
nand U11643 (N_11643,N_6532,N_5663);
xor U11644 (N_11644,N_7341,N_6303);
or U11645 (N_11645,N_7355,N_7275);
xor U11646 (N_11646,N_6420,N_7662);
or U11647 (N_11647,N_9754,N_9974);
nor U11648 (N_11648,N_9395,N_8492);
or U11649 (N_11649,N_7216,N_5416);
nor U11650 (N_11650,N_5942,N_5708);
or U11651 (N_11651,N_6018,N_9067);
nor U11652 (N_11652,N_7610,N_8131);
nand U11653 (N_11653,N_5026,N_8917);
nor U11654 (N_11654,N_5507,N_7384);
nand U11655 (N_11655,N_5610,N_8428);
and U11656 (N_11656,N_6205,N_7298);
nor U11657 (N_11657,N_9767,N_5419);
or U11658 (N_11658,N_7678,N_5616);
nand U11659 (N_11659,N_9220,N_9410);
nand U11660 (N_11660,N_6485,N_5139);
and U11661 (N_11661,N_6308,N_8329);
and U11662 (N_11662,N_5067,N_6840);
nor U11663 (N_11663,N_7371,N_5298);
nand U11664 (N_11664,N_7598,N_6120);
nand U11665 (N_11665,N_6421,N_7694);
or U11666 (N_11666,N_5684,N_6903);
nand U11667 (N_11667,N_9844,N_8481);
and U11668 (N_11668,N_6665,N_9948);
or U11669 (N_11669,N_7125,N_5650);
and U11670 (N_11670,N_8552,N_5670);
nand U11671 (N_11671,N_5888,N_9324);
nor U11672 (N_11672,N_7381,N_9033);
or U11673 (N_11673,N_6416,N_6279);
nand U11674 (N_11674,N_6870,N_9883);
nand U11675 (N_11675,N_9673,N_8367);
nor U11676 (N_11676,N_6838,N_7823);
nand U11677 (N_11677,N_9634,N_5044);
xor U11678 (N_11678,N_7328,N_8316);
nor U11679 (N_11679,N_9374,N_9934);
or U11680 (N_11680,N_8592,N_7585);
nand U11681 (N_11681,N_5928,N_6776);
nand U11682 (N_11682,N_7852,N_6051);
or U11683 (N_11683,N_6299,N_8480);
or U11684 (N_11684,N_8073,N_9655);
xor U11685 (N_11685,N_6623,N_7468);
and U11686 (N_11686,N_5045,N_7660);
xnor U11687 (N_11687,N_9468,N_9237);
or U11688 (N_11688,N_8866,N_6088);
nand U11689 (N_11689,N_8174,N_6964);
nand U11690 (N_11690,N_7061,N_7902);
nand U11691 (N_11691,N_6150,N_6737);
nand U11692 (N_11692,N_9083,N_5391);
or U11693 (N_11693,N_9118,N_9660);
xnor U11694 (N_11694,N_7710,N_6105);
nand U11695 (N_11695,N_7159,N_6241);
and U11696 (N_11696,N_7537,N_6519);
or U11697 (N_11697,N_9511,N_7670);
xor U11698 (N_11698,N_5206,N_5598);
nor U11699 (N_11699,N_6091,N_9317);
xnor U11700 (N_11700,N_8405,N_6802);
or U11701 (N_11701,N_5825,N_8620);
nand U11702 (N_11702,N_5674,N_5477);
and U11703 (N_11703,N_7583,N_8719);
xnor U11704 (N_11704,N_9926,N_9499);
or U11705 (N_11705,N_6063,N_8393);
nor U11706 (N_11706,N_5037,N_5643);
nor U11707 (N_11707,N_7952,N_9646);
nor U11708 (N_11708,N_9217,N_7259);
or U11709 (N_11709,N_5284,N_6768);
nand U11710 (N_11710,N_5241,N_5970);
nand U11711 (N_11711,N_6643,N_7192);
nand U11712 (N_11712,N_8692,N_7117);
or U11713 (N_11713,N_9387,N_6491);
nand U11714 (N_11714,N_5690,N_9136);
nor U11715 (N_11715,N_8647,N_9820);
and U11716 (N_11716,N_5599,N_5799);
nor U11717 (N_11717,N_6542,N_8914);
or U11718 (N_11718,N_7613,N_5252);
and U11719 (N_11719,N_6961,N_5680);
and U11720 (N_11720,N_5008,N_9615);
nor U11721 (N_11721,N_5523,N_6972);
or U11722 (N_11722,N_9425,N_7311);
nand U11723 (N_11723,N_8740,N_8409);
nor U11724 (N_11724,N_7360,N_5545);
nand U11725 (N_11725,N_9397,N_7451);
nor U11726 (N_11726,N_8516,N_8970);
nand U11727 (N_11727,N_6962,N_5121);
nand U11728 (N_11728,N_8176,N_9027);
nand U11729 (N_11729,N_6755,N_8582);
or U11730 (N_11730,N_9558,N_6092);
or U11731 (N_11731,N_8938,N_8634);
or U11732 (N_11732,N_5361,N_6099);
xor U11733 (N_11733,N_5162,N_5163);
nand U11734 (N_11734,N_6410,N_9596);
or U11735 (N_11735,N_9550,N_5591);
nand U11736 (N_11736,N_6387,N_7034);
or U11737 (N_11737,N_8005,N_7538);
or U11738 (N_11738,N_9437,N_7618);
nor U11739 (N_11739,N_9727,N_5887);
or U11740 (N_11740,N_8476,N_5988);
or U11741 (N_11741,N_8978,N_8490);
xnor U11742 (N_11742,N_9613,N_9156);
and U11743 (N_11743,N_7166,N_5972);
nand U11744 (N_11744,N_6171,N_5791);
nand U11745 (N_11745,N_9344,N_8945);
nand U11746 (N_11746,N_8948,N_8136);
or U11747 (N_11747,N_8600,N_9026);
or U11748 (N_11748,N_9828,N_8133);
xnor U11749 (N_11749,N_5925,N_7005);
nand U11750 (N_11750,N_6104,N_8837);
nand U11751 (N_11751,N_8792,N_9875);
nand U11752 (N_11752,N_7500,N_8591);
nand U11753 (N_11753,N_9423,N_7560);
and U11754 (N_11754,N_6066,N_5429);
nor U11755 (N_11755,N_8502,N_8615);
xor U11756 (N_11756,N_5768,N_7596);
or U11757 (N_11757,N_9288,N_7225);
or U11758 (N_11758,N_8508,N_8277);
nor U11759 (N_11759,N_6457,N_9706);
nor U11760 (N_11760,N_7339,N_8827);
or U11761 (N_11761,N_5543,N_5798);
nor U11762 (N_11762,N_5897,N_6810);
and U11763 (N_11763,N_6544,N_7767);
or U11764 (N_11764,N_7224,N_5954);
and U11765 (N_11765,N_9562,N_6377);
nor U11766 (N_11766,N_6506,N_7047);
nor U11767 (N_11767,N_7150,N_9415);
and U11768 (N_11768,N_6081,N_5613);
or U11769 (N_11769,N_6001,N_5052);
or U11770 (N_11770,N_8059,N_8928);
nor U11771 (N_11771,N_9125,N_8144);
nor U11772 (N_11772,N_8959,N_5076);
or U11773 (N_11773,N_7800,N_5912);
nand U11774 (N_11774,N_5310,N_7772);
or U11775 (N_11775,N_8616,N_6697);
nand U11776 (N_11776,N_6004,N_5681);
or U11777 (N_11777,N_8264,N_5125);
and U11778 (N_11778,N_5732,N_8331);
or U11779 (N_11779,N_8920,N_8864);
and U11780 (N_11780,N_5016,N_8180);
or U11781 (N_11781,N_5856,N_5209);
or U11782 (N_11782,N_9421,N_9132);
nand U11783 (N_11783,N_5945,N_8567);
and U11784 (N_11784,N_8093,N_9300);
and U11785 (N_11785,N_7557,N_6351);
and U11786 (N_11786,N_5210,N_6428);
nand U11787 (N_11787,N_8070,N_9355);
nor U11788 (N_11788,N_9097,N_9535);
nor U11789 (N_11789,N_9847,N_5936);
and U11790 (N_11790,N_8770,N_7023);
nand U11791 (N_11791,N_9505,N_5308);
xnor U11792 (N_11792,N_9062,N_6672);
or U11793 (N_11793,N_5120,N_8967);
and U11794 (N_11794,N_6536,N_7080);
xnor U11795 (N_11795,N_5894,N_7074);
nor U11796 (N_11796,N_9782,N_8109);
or U11797 (N_11797,N_8751,N_6829);
and U11798 (N_11798,N_7393,N_8545);
nor U11799 (N_11799,N_5987,N_9259);
nand U11800 (N_11800,N_9152,N_7078);
xor U11801 (N_11801,N_6783,N_5812);
or U11802 (N_11802,N_7110,N_7042);
xnor U11803 (N_11803,N_7073,N_5749);
and U11804 (N_11804,N_7143,N_7861);
and U11805 (N_11805,N_8823,N_6878);
nand U11806 (N_11806,N_5078,N_8535);
and U11807 (N_11807,N_8343,N_5077);
nand U11808 (N_11808,N_8305,N_6687);
nor U11809 (N_11809,N_6873,N_9459);
or U11810 (N_11810,N_8614,N_8828);
nand U11811 (N_11811,N_5449,N_5411);
nand U11812 (N_11812,N_9080,N_7203);
nor U11813 (N_11813,N_5651,N_9827);
and U11814 (N_11814,N_8891,N_7269);
nand U11815 (N_11815,N_7097,N_6579);
nor U11816 (N_11816,N_6713,N_5174);
or U11817 (N_11817,N_7209,N_6021);
and U11818 (N_11818,N_6450,N_8542);
nand U11819 (N_11819,N_5722,N_9028);
and U11820 (N_11820,N_5204,N_9409);
or U11821 (N_11821,N_5302,N_8210);
nand U11822 (N_11822,N_8909,N_9005);
and U11823 (N_11823,N_7082,N_7084);
nor U11824 (N_11824,N_9417,N_9918);
and U11825 (N_11825,N_8759,N_8491);
nand U11826 (N_11826,N_7671,N_5917);
nor U11827 (N_11827,N_8768,N_6217);
and U11828 (N_11828,N_8812,N_6456);
nand U11829 (N_11829,N_5999,N_7658);
nand U11830 (N_11830,N_5122,N_8249);
xnor U11831 (N_11831,N_6475,N_8757);
nand U11832 (N_11832,N_9702,N_6172);
nand U11833 (N_11833,N_8120,N_5383);
nor U11834 (N_11834,N_9859,N_5237);
and U11835 (N_11835,N_5769,N_5404);
nor U11836 (N_11836,N_9285,N_7292);
or U11837 (N_11837,N_5803,N_5227);
and U11838 (N_11838,N_9356,N_7127);
and U11839 (N_11839,N_7025,N_6809);
nor U11840 (N_11840,N_5867,N_9787);
nor U11841 (N_11841,N_8646,N_6980);
nor U11842 (N_11842,N_8323,N_9174);
and U11843 (N_11843,N_5000,N_5953);
and U11844 (N_11844,N_8410,N_5847);
nor U11845 (N_11845,N_6077,N_8313);
nand U11846 (N_11846,N_5525,N_6824);
nor U11847 (N_11847,N_9930,N_7737);
nor U11848 (N_11848,N_5628,N_6272);
and U11849 (N_11849,N_8933,N_8017);
nand U11850 (N_11850,N_8177,N_7211);
xor U11851 (N_11851,N_7331,N_5683);
nor U11852 (N_11852,N_7400,N_9108);
or U11853 (N_11853,N_5457,N_7141);
or U11854 (N_11854,N_6155,N_5108);
and U11855 (N_11855,N_5116,N_7664);
nor U11856 (N_11856,N_9323,N_9326);
or U11857 (N_11857,N_6502,N_8671);
or U11858 (N_11858,N_9732,N_8786);
and U11859 (N_11859,N_7477,N_6467);
or U11860 (N_11860,N_5109,N_9600);
nand U11861 (N_11861,N_5056,N_8280);
nand U11862 (N_11862,N_5753,N_9277);
or U11863 (N_11863,N_5845,N_7918);
and U11864 (N_11864,N_6716,N_9407);
nand U11865 (N_11865,N_5283,N_9093);
and U11866 (N_11866,N_9944,N_8498);
or U11867 (N_11867,N_5219,N_8081);
nor U11868 (N_11868,N_9463,N_6522);
or U11869 (N_11869,N_6752,N_7112);
xor U11870 (N_11870,N_7549,N_6028);
or U11871 (N_11871,N_7831,N_6090);
nor U11872 (N_11872,N_8513,N_6948);
xor U11873 (N_11873,N_6900,N_5118);
and U11874 (N_11874,N_5993,N_9701);
nor U11875 (N_11875,N_6082,N_6504);
or U11876 (N_11876,N_8256,N_8335);
or U11877 (N_11877,N_8977,N_5230);
nand U11878 (N_11878,N_6128,N_9053);
nor U11879 (N_11879,N_9518,N_7378);
and U11880 (N_11880,N_5004,N_7562);
or U11881 (N_11881,N_5384,N_9299);
and U11882 (N_11882,N_8108,N_5824);
and U11883 (N_11883,N_8652,N_8548);
nand U11884 (N_11884,N_5607,N_5395);
nor U11885 (N_11885,N_6700,N_5264);
or U11886 (N_11886,N_9052,N_5508);
and U11887 (N_11887,N_6132,N_7250);
xor U11888 (N_11888,N_5719,N_5355);
and U11889 (N_11889,N_7314,N_9138);
nor U11890 (N_11890,N_5285,N_5279);
and U11891 (N_11891,N_9135,N_8691);
or U11892 (N_11892,N_9273,N_6269);
nor U11893 (N_11893,N_8044,N_6466);
nor U11894 (N_11894,N_8761,N_6660);
or U11895 (N_11895,N_7547,N_7226);
and U11896 (N_11896,N_8664,N_5229);
and U11897 (N_11897,N_8045,N_8831);
or U11898 (N_11898,N_8559,N_7287);
nor U11899 (N_11899,N_8099,N_7241);
and U11900 (N_11900,N_8599,N_8725);
nor U11901 (N_11901,N_5588,N_6488);
and U11902 (N_11902,N_7499,N_6060);
nor U11903 (N_11903,N_9749,N_5402);
and U11904 (N_11904,N_7089,N_8169);
nor U11905 (N_11905,N_5131,N_7375);
nor U11906 (N_11906,N_5055,N_7999);
and U11907 (N_11907,N_8298,N_5877);
and U11908 (N_11908,N_7333,N_6206);
nor U11909 (N_11909,N_9076,N_6267);
or U11910 (N_11910,N_7184,N_7649);
or U11911 (N_11911,N_5948,N_6787);
and U11912 (N_11912,N_9017,N_7771);
nor U11913 (N_11913,N_8514,N_9351);
nor U11914 (N_11914,N_6859,N_8749);
or U11915 (N_11915,N_5834,N_5955);
or U11916 (N_11916,N_7929,N_5733);
and U11917 (N_11917,N_9602,N_6349);
or U11918 (N_11918,N_5446,N_9488);
and U11919 (N_11919,N_6023,N_9548);
nor U11920 (N_11920,N_8140,N_9224);
and U11921 (N_11921,N_6846,N_6433);
or U11922 (N_11922,N_9748,N_6168);
nor U11923 (N_11923,N_7003,N_6123);
nand U11924 (N_11924,N_5140,N_9029);
nor U11925 (N_11925,N_5815,N_9991);
and U11926 (N_11926,N_9564,N_7607);
nand U11927 (N_11927,N_7380,N_7584);
nor U11928 (N_11928,N_9672,N_8186);
or U11929 (N_11929,N_5322,N_9367);
nand U11930 (N_11930,N_9462,N_8042);
or U11931 (N_11931,N_8521,N_9049);
nor U11932 (N_11932,N_6184,N_7391);
nand U11933 (N_11933,N_9532,N_7007);
nor U11934 (N_11934,N_9899,N_8641);
or U11935 (N_11935,N_9671,N_8309);
or U11936 (N_11936,N_9549,N_5734);
nor U11937 (N_11937,N_9598,N_9880);
nor U11938 (N_11938,N_6796,N_9868);
xnor U11939 (N_11939,N_6240,N_8006);
and U11940 (N_11940,N_8843,N_5196);
or U11941 (N_11941,N_7475,N_9186);
and U11942 (N_11942,N_8077,N_9316);
or U11943 (N_11943,N_5047,N_9498);
nor U11944 (N_11944,N_6029,N_9832);
or U11945 (N_11945,N_7816,N_9812);
nand U11946 (N_11946,N_5167,N_7109);
xnor U11947 (N_11947,N_5869,N_7956);
or U11948 (N_11948,N_6676,N_9573);
nor U11949 (N_11949,N_5150,N_7813);
xor U11950 (N_11950,N_6296,N_5671);
nand U11951 (N_11951,N_7571,N_6708);
nand U11952 (N_11952,N_6195,N_8861);
nor U11953 (N_11953,N_8973,N_5772);
or U11954 (N_11954,N_7045,N_7151);
and U11955 (N_11955,N_9848,N_6179);
xor U11956 (N_11956,N_6908,N_8385);
nand U11957 (N_11957,N_9002,N_5627);
or U11958 (N_11958,N_8741,N_9201);
nand U11959 (N_11959,N_7531,N_9531);
or U11960 (N_11960,N_9744,N_5997);
nand U11961 (N_11961,N_6152,N_8071);
or U11962 (N_11962,N_6891,N_7318);
xor U11963 (N_11963,N_9797,N_8061);
and U11964 (N_11964,N_8657,N_9527);
nor U11965 (N_11965,N_8510,N_8528);
nand U11966 (N_11966,N_5761,N_7523);
and U11967 (N_11967,N_8718,N_7015);
nor U11968 (N_11968,N_5400,N_6510);
and U11969 (N_11969,N_5534,N_8192);
and U11970 (N_11970,N_6446,N_7096);
or U11971 (N_11971,N_8626,N_7362);
nand U11972 (N_11972,N_5119,N_8844);
or U11973 (N_11973,N_5320,N_6250);
or U11974 (N_11974,N_6130,N_8769);
xnor U11975 (N_11975,N_9414,N_9483);
nor U11976 (N_11976,N_5841,N_5870);
nand U11977 (N_11977,N_8184,N_6808);
and U11978 (N_11978,N_5558,N_6073);
and U11979 (N_11979,N_9626,N_8437);
and U11980 (N_11980,N_9284,N_5879);
and U11981 (N_11981,N_8796,N_9685);
and U11982 (N_11982,N_7091,N_6230);
and U11983 (N_11983,N_5338,N_5644);
nand U11984 (N_11984,N_7640,N_6285);
nor U11985 (N_11985,N_6432,N_6736);
nor U11986 (N_11986,N_9347,N_8290);
nor U11987 (N_11987,N_8426,N_7962);
xor U11988 (N_11988,N_5568,N_8605);
nand U11989 (N_11989,N_7234,N_9695);
or U11990 (N_11990,N_7965,N_5104);
nand U11991 (N_11991,N_8474,N_7039);
and U11992 (N_11992,N_9657,N_5842);
nor U11993 (N_11993,N_5456,N_6552);
nand U11994 (N_11994,N_7009,N_7370);
nand U11995 (N_11995,N_9470,N_9031);
nand U11996 (N_11996,N_9624,N_8799);
xnor U11997 (N_11997,N_7770,N_9331);
xnor U11998 (N_11998,N_8717,N_6298);
and U11999 (N_11999,N_9046,N_8344);
xor U12000 (N_12000,N_9063,N_7286);
and U12001 (N_12001,N_9938,N_7019);
and U12002 (N_12002,N_5539,N_6514);
or U12003 (N_12003,N_8299,N_6923);
nor U12004 (N_12004,N_5465,N_8588);
and U12005 (N_12005,N_8815,N_8726);
or U12006 (N_12006,N_9843,N_9349);
nand U12007 (N_12007,N_7848,N_6523);
and U12008 (N_12008,N_7989,N_8046);
nor U12009 (N_12009,N_6304,N_5189);
and U12010 (N_12010,N_9594,N_8957);
or U12011 (N_12011,N_9709,N_8315);
and U12012 (N_12012,N_6049,N_8565);
and U12013 (N_12013,N_6397,N_9485);
and U12014 (N_12014,N_8252,N_8352);
nor U12015 (N_12015,N_8302,N_8262);
nand U12016 (N_12016,N_7828,N_6920);
or U12017 (N_12017,N_9211,N_5911);
nand U12018 (N_12018,N_7146,N_6732);
or U12019 (N_12019,N_8363,N_9679);
nand U12020 (N_12020,N_7987,N_5415);
xnor U12021 (N_12021,N_7762,N_8111);
xor U12022 (N_12022,N_8356,N_5696);
or U12023 (N_12023,N_5236,N_7873);
and U12024 (N_12024,N_6953,N_6451);
nand U12025 (N_12025,N_8415,N_5979);
and U12026 (N_12026,N_5730,N_6835);
or U12027 (N_12027,N_6625,N_9969);
xnor U12028 (N_12028,N_9967,N_9373);
nand U12029 (N_12029,N_8756,N_6577);
nand U12030 (N_12030,N_5329,N_9056);
nor U12031 (N_12031,N_5943,N_5744);
and U12032 (N_12032,N_9301,N_6496);
nor U12033 (N_12033,N_7066,N_9276);
nand U12034 (N_12034,N_8438,N_5562);
nor U12035 (N_12035,N_9636,N_5819);
nand U12036 (N_12036,N_8115,N_7787);
xnor U12037 (N_12037,N_9988,N_6720);
or U12038 (N_12038,N_9545,N_6113);
nor U12039 (N_12039,N_8404,N_7437);
nand U12040 (N_12040,N_5552,N_8606);
nor U12041 (N_12041,N_8628,N_6565);
nor U12042 (N_12042,N_7652,N_5373);
xor U12043 (N_12043,N_9297,N_7179);
and U12044 (N_12044,N_8272,N_6567);
nor U12045 (N_12045,N_8708,N_5603);
or U12046 (N_12046,N_8430,N_5009);
or U12047 (N_12047,N_5820,N_7267);
or U12048 (N_12048,N_7123,N_8919);
nand U12049 (N_12049,N_5573,N_5669);
and U12050 (N_12050,N_5516,N_5935);
or U12051 (N_12051,N_9593,N_6960);
or U12052 (N_12052,N_7691,N_9120);
and U12053 (N_12053,N_5412,N_6594);
xor U12054 (N_12054,N_5424,N_8639);
nand U12055 (N_12055,N_6974,N_7979);
nand U12056 (N_12056,N_5130,N_8200);
nand U12057 (N_12057,N_7706,N_7288);
and U12058 (N_12058,N_7290,N_8992);
and U12059 (N_12059,N_6745,N_9952);
and U12060 (N_12060,N_6575,N_7959);
and U12061 (N_12061,N_6209,N_6999);
nor U12062 (N_12062,N_9122,N_6717);
nand U12063 (N_12063,N_8373,N_7997);
or U12064 (N_12064,N_8651,N_5350);
nor U12065 (N_12065,N_7766,N_6276);
nor U12066 (N_12066,N_5908,N_5546);
and U12067 (N_12067,N_7064,N_5423);
nor U12068 (N_12068,N_9467,N_7484);
and U12069 (N_12069,N_9680,N_6876);
or U12070 (N_12070,N_5168,N_8869);
xnor U12071 (N_12071,N_6497,N_6012);
or U12072 (N_12072,N_9294,N_5724);
or U12073 (N_12073,N_6048,N_5592);
xor U12074 (N_12074,N_5555,N_9968);
nand U12075 (N_12075,N_7389,N_8563);
or U12076 (N_12076,N_9330,N_9770);
nor U12077 (N_12077,N_5919,N_9703);
and U12078 (N_12078,N_6880,N_8132);
nor U12079 (N_12079,N_6819,N_7641);
or U12080 (N_12080,N_8390,N_6149);
nand U12081 (N_12081,N_9963,N_7026);
and U12082 (N_12082,N_6468,N_8084);
and U12083 (N_12083,N_9506,N_6957);
nor U12084 (N_12084,N_5304,N_8969);
nand U12085 (N_12085,N_8710,N_7951);
and U12086 (N_12086,N_5623,N_7116);
xnor U12087 (N_12087,N_8372,N_9603);
and U12088 (N_12088,N_8114,N_5575);
nor U12089 (N_12089,N_9490,N_6391);
nand U12090 (N_12090,N_6540,N_6645);
and U12091 (N_12091,N_5305,N_9476);
or U12092 (N_12092,N_7775,N_7964);
nand U12093 (N_12093,N_9663,N_5377);
nor U12094 (N_12094,N_5738,N_8291);
and U12095 (N_12095,N_6127,N_8564);
or U12096 (N_12096,N_9866,N_7427);
nor U12097 (N_12097,N_6527,N_9716);
or U12098 (N_12098,N_7599,N_8457);
or U12099 (N_12099,N_9234,N_5261);
and U12100 (N_12100,N_6441,N_8689);
nor U12101 (N_12101,N_5110,N_7294);
nor U12102 (N_12102,N_8275,N_5462);
or U12103 (N_12103,N_5354,N_7441);
nor U12104 (N_12104,N_5517,N_5041);
nor U12105 (N_12105,N_7909,N_8179);
and U12106 (N_12106,N_7090,N_8590);
xnor U12107 (N_12107,N_6382,N_6602);
nand U12108 (N_12108,N_6083,N_5785);
nor U12109 (N_12109,N_5084,N_7768);
nor U12110 (N_12110,N_7896,N_8001);
nor U12111 (N_12111,N_6246,N_8670);
and U12112 (N_12112,N_5203,N_7494);
nor U12113 (N_12113,N_8212,N_8733);
xnor U12114 (N_12114,N_7444,N_8713);
nor U12115 (N_12115,N_6638,N_9269);
or U12116 (N_12116,N_6376,N_5115);
and U12117 (N_12117,N_6685,N_8941);
nand U12118 (N_12118,N_9230,N_9973);
nor U12119 (N_12119,N_9639,N_7344);
xor U12120 (N_12120,N_7490,N_6383);
xnor U12121 (N_12121,N_8368,N_9146);
or U12122 (N_12122,N_9985,N_9870);
and U12123 (N_12123,N_7403,N_8463);
and U12124 (N_12124,N_6237,N_6198);
and U12125 (N_12125,N_5245,N_8026);
xor U12126 (N_12126,N_9764,N_5259);
nor U12127 (N_12127,N_5717,N_7261);
and U12128 (N_12128,N_6821,N_7419);
nor U12129 (N_12129,N_5106,N_7263);
nand U12130 (N_12130,N_7431,N_8900);
and U12131 (N_12131,N_7907,N_9651);
nor U12132 (N_12132,N_7075,N_5043);
nor U12133 (N_12133,N_7897,N_8679);
nor U12134 (N_12134,N_5303,N_6689);
or U12135 (N_12135,N_9541,N_8878);
xor U12136 (N_12136,N_8622,N_5309);
nand U12137 (N_12137,N_5980,N_9457);
and U12138 (N_12138,N_6469,N_5335);
nor U12139 (N_12139,N_8702,N_9375);
nor U12140 (N_12140,N_6271,N_5751);
nor U12141 (N_12141,N_5818,N_8625);
and U12142 (N_12142,N_7953,N_6663);
and U12143 (N_12143,N_9530,N_5208);
and U12144 (N_12144,N_5425,N_9095);
nand U12145 (N_12145,N_8781,N_5405);
nand U12146 (N_12146,N_6642,N_6767);
or U12147 (N_12147,N_7978,N_7354);
nand U12148 (N_12148,N_7265,N_5757);
nor U12149 (N_12149,N_9311,N_8809);
and U12150 (N_12150,N_9908,N_6314);
nor U12151 (N_12151,N_7429,N_9365);
or U12152 (N_12152,N_5136,N_9253);
nand U12153 (N_12153,N_9781,N_6869);
or U12154 (N_12154,N_5740,N_5132);
and U12155 (N_12155,N_6680,N_8858);
or U12156 (N_12156,N_8473,N_5069);
nor U12157 (N_12157,N_7602,N_7168);
or U12158 (N_12158,N_5838,N_7049);
nor U12159 (N_12159,N_9121,N_7630);
and U12160 (N_12160,N_7013,N_8638);
or U12161 (N_12161,N_7320,N_6337);
nor U12162 (N_12162,N_6070,N_6925);
xnor U12163 (N_12163,N_8089,N_5976);
and U12164 (N_12164,N_7877,N_8752);
xor U12165 (N_12165,N_8500,N_6356);
and U12166 (N_12166,N_7785,N_9359);
xnor U12167 (N_12167,N_7107,N_6095);
nand U12168 (N_12168,N_9711,N_6698);
nand U12169 (N_12169,N_5427,N_9648);
xor U12170 (N_12170,N_8908,N_6164);
or U12171 (N_12171,N_7188,N_7223);
or U12172 (N_12172,N_7597,N_9691);
or U12173 (N_12173,N_9162,N_8504);
or U12174 (N_12174,N_9065,N_8396);
nor U12175 (N_12175,N_9863,N_9965);
nor U12176 (N_12176,N_9110,N_8002);
nor U12177 (N_12177,N_6844,N_6141);
nor U12178 (N_12178,N_7699,N_8311);
and U12179 (N_12179,N_8793,N_8954);
and U12180 (N_12180,N_5759,N_8025);
or U12181 (N_12181,N_6853,N_9601);
or U12182 (N_12182,N_7556,N_6588);
or U12183 (N_12183,N_9158,N_8729);
and U12184 (N_12184,N_8549,N_6652);
or U12185 (N_12185,N_6924,N_6789);
or U12186 (N_12186,N_5852,N_9962);
nor U12187 (N_12187,N_6842,N_9064);
nor U12188 (N_12188,N_9113,N_5951);
nor U12189 (N_12189,N_7859,N_7680);
or U12190 (N_12190,N_9668,N_6415);
xnor U12191 (N_12191,N_9081,N_7761);
or U12192 (N_12192,N_8355,N_7364);
or U12193 (N_12193,N_8330,N_5556);
nand U12194 (N_12194,N_6086,N_8191);
and U12195 (N_12195,N_9188,N_9372);
nand U12196 (N_12196,N_5672,N_9105);
nor U12197 (N_12197,N_8370,N_5317);
nand U12198 (N_12198,N_8776,N_9391);
and U12199 (N_12199,N_7975,N_8859);
nor U12200 (N_12200,N_7627,N_6587);
and U12201 (N_12201,N_6316,N_9979);
nand U12202 (N_12202,N_7619,N_8359);
nand U12203 (N_12203,N_7723,N_7124);
nor U12204 (N_12204,N_9205,N_7326);
or U12205 (N_12205,N_8412,N_9735);
or U12206 (N_12206,N_8327,N_9130);
nand U12207 (N_12207,N_5311,N_9641);
nand U12208 (N_12208,N_6862,N_7604);
or U12209 (N_12209,N_8215,N_5328);
or U12210 (N_12210,N_6766,N_7947);
nand U12211 (N_12211,N_6093,N_5969);
nand U12212 (N_12212,N_6334,N_5176);
and U12213 (N_12213,N_9684,N_7589);
and U12214 (N_12214,N_8790,N_9833);
nor U12215 (N_12215,N_5060,N_8773);
xor U12216 (N_12216,N_7406,N_7397);
nor U12217 (N_12217,N_6442,N_9000);
or U12218 (N_12218,N_5721,N_6684);
nor U12219 (N_12219,N_5958,N_6181);
or U12220 (N_12220,N_5609,N_6738);
or U12221 (N_12221,N_6867,N_7277);
and U12222 (N_12222,N_5243,N_9698);
or U12223 (N_12223,N_6331,N_7279);
xnor U12224 (N_12224,N_8648,N_6503);
nor U12225 (N_12225,N_8854,N_6868);
nor U12226 (N_12226,N_5380,N_7845);
nand U12227 (N_12227,N_9144,N_5579);
nor U12228 (N_12228,N_8429,N_6631);
or U12229 (N_12229,N_9773,N_9514);
nand U12230 (N_12230,N_7276,N_5509);
and U12231 (N_12231,N_9059,N_8351);
nor U12232 (N_12232,N_6854,N_7164);
nand U12233 (N_12233,N_6079,N_6926);
nand U12234 (N_12234,N_7586,N_5830);
nand U12235 (N_12235,N_9192,N_9133);
nand U12236 (N_12236,N_5485,N_8608);
or U12237 (N_12237,N_8529,N_8181);
and U12238 (N_12238,N_7681,N_8350);
and U12239 (N_12239,N_8023,N_5472);
and U12240 (N_12240,N_9643,N_5637);
nor U12241 (N_12241,N_9078,N_9721);
or U12242 (N_12242,N_9261,N_5816);
xnor U12243 (N_12243,N_9637,N_9509);
nor U12244 (N_12244,N_9012,N_5296);
nand U12245 (N_12245,N_6019,N_6347);
xnor U12246 (N_12246,N_6202,N_7432);
nand U12247 (N_12247,N_8380,N_9517);
xnor U12248 (N_12248,N_6721,N_9322);
or U12249 (N_12249,N_9401,N_5374);
nor U12250 (N_12250,N_5528,N_7611);
nor U12251 (N_12251,N_7343,N_5522);
and U12252 (N_12252,N_6193,N_5904);
nor U12253 (N_12253,N_7994,N_8594);
nor U12254 (N_12254,N_5898,N_8762);
or U12255 (N_12255,N_9862,N_8102);
nand U12256 (N_12256,N_7955,N_9775);
or U12257 (N_12257,N_9570,N_5922);
and U12258 (N_12258,N_8640,N_5580);
nand U12259 (N_12259,N_8874,N_9837);
or U12260 (N_12260,N_9493,N_8225);
nor U12261 (N_12261,N_5145,N_9665);
and U12262 (N_12262,N_7984,N_5278);
or U12263 (N_12263,N_8882,N_8546);
nor U12264 (N_12264,N_9970,N_5735);
and U12265 (N_12265,N_5186,N_7899);
and U12266 (N_12266,N_9378,N_6883);
nand U12267 (N_12267,N_9112,N_6683);
xor U12268 (N_12268,N_6885,N_6399);
xnor U12269 (N_12269,N_7368,N_6816);
or U12270 (N_12270,N_5342,N_6275);
nand U12271 (N_12271,N_9664,N_9308);
nand U12272 (N_12272,N_5343,N_7434);
xnor U12273 (N_12273,N_5048,N_9088);
xnor U12274 (N_12274,N_9807,N_9516);
xor U12275 (N_12275,N_9993,N_5519);
and U12276 (N_12276,N_7363,N_5677);
nand U12277 (N_12277,N_6490,N_9785);
nor U12278 (N_12278,N_6075,N_7566);
nand U12279 (N_12279,N_9396,N_9544);
nor U12280 (N_12280,N_9983,N_8091);
nor U12281 (N_12281,N_8318,N_8644);
nand U12282 (N_12282,N_8090,N_7113);
and U12283 (N_12283,N_9761,N_9101);
xnor U12284 (N_12284,N_6197,N_8788);
and U12285 (N_12285,N_5437,N_9327);
nor U12286 (N_12286,N_8753,N_6617);
nor U12287 (N_12287,N_6955,N_8888);
or U12288 (N_12288,N_5276,N_6359);
nor U12289 (N_12289,N_5273,N_8423);
nor U12290 (N_12290,N_6654,N_8683);
and U12291 (N_12291,N_9707,N_9466);
or U12292 (N_12292,N_7817,N_6288);
nand U12293 (N_12293,N_6746,N_7812);
or U12294 (N_12294,N_6386,N_7665);
and U12295 (N_12295,N_6946,N_9608);
nand U12296 (N_12296,N_6889,N_8440);
nor U12297 (N_12297,N_7910,N_5995);
or U12298 (N_12298,N_8388,N_5520);
nor U12299 (N_12299,N_9223,N_5649);
nor U12300 (N_12300,N_5946,N_9247);
and U12301 (N_12301,N_5399,N_5025);
nand U12302 (N_12302,N_5470,N_6445);
nor U12303 (N_12303,N_5875,N_6935);
and U12304 (N_12304,N_9066,N_8255);
nor U12305 (N_12305,N_7992,N_6793);
xnor U12306 (N_12306,N_5441,N_8983);
nor U12307 (N_12307,N_6943,N_7158);
or U12308 (N_12308,N_6369,N_9242);
nor U12309 (N_12309,N_9694,N_5396);
and U12310 (N_12310,N_7849,N_7227);
nand U12311 (N_12311,N_8399,N_7103);
xor U12312 (N_12312,N_5286,N_9350);
xor U12313 (N_12313,N_6740,N_7140);
or U12314 (N_12314,N_5514,N_6265);
and U12315 (N_12315,N_9582,N_8482);
nand U12316 (N_12316,N_7778,N_5704);
or U12317 (N_12317,N_8051,N_9435);
nor U12318 (N_12318,N_8819,N_9758);
nor U12319 (N_12319,N_9627,N_5571);
nor U12320 (N_12320,N_5292,N_8587);
xor U12321 (N_12321,N_5576,N_8286);
nor U12322 (N_12322,N_8346,N_8852);
nand U12323 (N_12323,N_8825,N_9886);
nand U12324 (N_12324,N_5370,N_8930);
and U12325 (N_12325,N_8960,N_6373);
and U12326 (N_12326,N_8030,N_7914);
and U12327 (N_12327,N_5828,N_5079);
xor U12328 (N_12328,N_5755,N_7480);
nand U12329 (N_12329,N_7700,N_8971);
or U12330 (N_12330,N_8990,N_7645);
or U12331 (N_12331,N_8543,N_5154);
nor U12332 (N_12332,N_7176,N_8241);
and U12333 (N_12333,N_5381,N_5745);
nor U12334 (N_12334,N_7677,N_6592);
and U12335 (N_12335,N_7032,N_5777);
xor U12336 (N_12336,N_8163,N_8381);
or U12337 (N_12337,N_9924,N_7780);
and U12338 (N_12338,N_6035,N_5337);
nor U12339 (N_12339,N_8227,N_5977);
nor U12340 (N_12340,N_5891,N_5448);
or U12341 (N_12341,N_6686,N_6339);
nand U12342 (N_12342,N_9222,N_6936);
and U12343 (N_12343,N_6307,N_9154);
nand U12344 (N_12344,N_5491,N_5741);
and U12345 (N_12345,N_6898,N_8518);
nand U12346 (N_12346,N_6931,N_6692);
nor U12347 (N_12347,N_8507,N_9806);
or U12348 (N_12348,N_6189,N_8872);
xnor U12349 (N_12349,N_8984,N_6647);
and U12350 (N_12350,N_5676,N_6855);
or U12351 (N_12351,N_6219,N_6849);
or U12352 (N_12352,N_9982,N_9894);
nand U12353 (N_12353,N_8397,N_9629);
nor U12354 (N_12354,N_9502,N_6728);
or U12355 (N_12355,N_8097,N_8706);
or U12356 (N_12356,N_9167,N_5362);
xor U12357 (N_12357,N_7044,N_8562);
and U12358 (N_12358,N_9571,N_5706);
xor U12359 (N_12359,N_5062,N_5331);
nor U12360 (N_12360,N_6541,N_6270);
or U12361 (N_12361,N_8653,N_8695);
and U12362 (N_12362,N_7624,N_9523);
and U12363 (N_12363,N_7037,N_6203);
nor U12364 (N_12364,N_8141,N_5705);
nor U12365 (N_12365,N_7248,N_6690);
nor U12366 (N_12366,N_6547,N_9621);
xnor U12367 (N_12367,N_7219,N_6500);
nor U12368 (N_12368,N_7496,N_8449);
or U12369 (N_12369,N_9576,N_8296);
or U12370 (N_12370,N_6703,N_7332);
or U12371 (N_12371,N_5430,N_9155);
or U12372 (N_12372,N_7606,N_7590);
nand U12373 (N_12373,N_7051,N_9419);
nor U12374 (N_12374,N_8450,N_9358);
nand U12375 (N_12375,N_8281,N_7462);
nor U12376 (N_12376,N_8266,N_6329);
and U12377 (N_12377,N_6656,N_9295);
or U12378 (N_12378,N_5347,N_9762);
xor U12379 (N_12379,N_7058,N_5032);
xnor U12380 (N_12380,N_7889,N_8750);
nor U12381 (N_12381,N_7178,N_9448);
and U12382 (N_12382,N_8915,N_9542);
or U12383 (N_12383,N_5378,N_9951);
or U12384 (N_12384,N_8870,N_7801);
xor U12385 (N_12385,N_6046,N_9182);
and U12386 (N_12386,N_7002,N_9841);
or U12387 (N_12387,N_5417,N_8008);
or U12388 (N_12388,N_6635,N_9469);
or U12389 (N_12389,N_6045,N_7367);
xor U12390 (N_12390,N_7688,N_6044);
nor U12391 (N_12391,N_7827,N_7692);
nand U12392 (N_12392,N_7452,N_6571);
or U12393 (N_12393,N_8088,N_7476);
and U12394 (N_12394,N_8593,N_8913);
and U12395 (N_12395,N_7157,N_9763);
and U12396 (N_12396,N_6119,N_8816);
or U12397 (N_12397,N_7195,N_5094);
and U12398 (N_12398,N_8932,N_7033);
nand U12399 (N_12399,N_8835,N_9202);
nor U12400 (N_12400,N_9693,N_8618);
nand U12401 (N_12401,N_8966,N_8800);
xnor U12402 (N_12402,N_5780,N_6162);
or U12403 (N_12403,N_9910,N_8694);
and U12404 (N_12404,N_9853,N_8349);
nor U12405 (N_12405,N_7573,N_7553);
nor U12406 (N_12406,N_5072,N_5290);
xnor U12407 (N_12407,N_7565,N_7322);
or U12408 (N_12408,N_6524,N_8890);
or U12409 (N_12409,N_9729,N_9268);
or U12410 (N_12410,N_9873,N_8810);
and U12411 (N_12411,N_9007,N_7175);
or U12412 (N_12412,N_6971,N_7529);
and U12413 (N_12413,N_6273,N_9281);
or U12414 (N_12414,N_5583,N_5117);
xor U12415 (N_12415,N_5166,N_5143);
nand U12416 (N_12416,N_7988,N_7635);
and U12417 (N_12417,N_9852,N_9589);
or U12418 (N_12418,N_7527,N_7104);
nor U12419 (N_12419,N_8214,N_8130);
or U12420 (N_12420,N_6538,N_7405);
nand U12421 (N_12421,N_6165,N_7830);
nand U12422 (N_12422,N_6627,N_6052);
and U12423 (N_12423,N_9170,N_9200);
nand U12424 (N_12424,N_6453,N_9817);
and U12425 (N_12425,N_8779,N_8078);
and U12426 (N_12426,N_7578,N_8716);
nand U12427 (N_12427,N_8856,N_7052);
or U12428 (N_12428,N_9587,N_5548);
or U12429 (N_12429,N_6901,N_9811);
nand U12430 (N_12430,N_9879,N_7208);
or U12431 (N_12431,N_7327,N_5440);
nand U12432 (N_12432,N_6185,N_9609);
xnor U12433 (N_12433,N_6409,N_7001);
or U12434 (N_12434,N_8578,N_6590);
and U12435 (N_12435,N_5212,N_5950);
and U12436 (N_12436,N_6228,N_6261);
or U12437 (N_12437,N_8100,N_5857);
nand U12438 (N_12438,N_7718,N_6748);
nor U12439 (N_12439,N_8911,N_6327);
nand U12440 (N_12440,N_9315,N_7629);
and U12441 (N_12441,N_9961,N_7474);
nor U12442 (N_12442,N_6455,N_5205);
nor U12443 (N_12443,N_7621,N_7711);
and U12444 (N_12444,N_8898,N_7644);
nand U12445 (N_12445,N_7312,N_8704);
nor U12446 (N_12446,N_7016,N_7513);
nor U12447 (N_12447,N_7581,N_8431);
or U12448 (N_12448,N_7923,N_6629);
or U12449 (N_12449,N_7041,N_9091);
and U12450 (N_12450,N_9445,N_9755);
or U12451 (N_12451,N_9722,N_7739);
or U12452 (N_12452,N_5978,N_9389);
nand U12453 (N_12453,N_8031,N_9734);
nor U12454 (N_12454,N_8459,N_8376);
and U12455 (N_12455,N_9821,N_7187);
and U12456 (N_12456,N_8472,N_8278);
and U12457 (N_12457,N_8306,N_9320);
nor U12458 (N_12458,N_7666,N_6639);
nand U12459 (N_12459,N_7501,N_9704);
xor U12460 (N_12460,N_6945,N_7221);
or U12461 (N_12461,N_8458,N_7435);
and U12462 (N_12462,N_9618,N_6521);
or U12463 (N_12463,N_7411,N_5372);
and U12464 (N_12464,N_9661,N_7543);
and U12465 (N_12465,N_7472,N_7615);
nand U12466 (N_12466,N_8850,N_6956);
nor U12467 (N_12467,N_5873,N_5737);
nand U12468 (N_12468,N_5975,N_7407);
nand U12469 (N_12469,N_5112,N_8058);
or U12470 (N_12470,N_9479,N_8183);
and U12471 (N_12471,N_5807,N_9757);
nor U12472 (N_12472,N_9368,N_5142);
nor U12473 (N_12473,N_7773,N_6302);
and U12474 (N_12474,N_5692,N_9552);
or U12475 (N_12475,N_5349,N_9578);
and U12476 (N_12476,N_9384,N_8369);
or U12477 (N_12477,N_6843,N_7156);
nand U12478 (N_12478,N_9819,N_9683);
or U12479 (N_12479,N_5049,N_9992);
or U12480 (N_12480,N_6831,N_6213);
or U12481 (N_12481,N_7783,N_5428);
nand U12482 (N_12482,N_7895,N_6425);
nand U12483 (N_12483,N_7424,N_9489);
and U12484 (N_12484,N_9904,N_8246);
and U12485 (N_12485,N_5093,N_5572);
or U12486 (N_12486,N_6190,N_6681);
nor U12487 (N_12487,N_7440,N_7888);
or U12488 (N_12488,N_6131,N_9949);
and U12489 (N_12489,N_5297,N_5560);
nand U12490 (N_12490,N_8387,N_6389);
nand U12491 (N_12491,N_6718,N_8260);
xor U12492 (N_12492,N_9402,N_6533);
or U12493 (N_12493,N_6053,N_6735);
and U12494 (N_12494,N_9546,N_7916);
or U12495 (N_12495,N_5553,N_6449);
nand U12496 (N_12496,N_7417,N_9141);
and U12497 (N_12497,N_9487,N_5272);
and U12498 (N_12498,N_6014,N_8029);
or U12499 (N_12499,N_5394,N_8292);
nand U12500 (N_12500,N_6746,N_5406);
nand U12501 (N_12501,N_6355,N_6752);
xor U12502 (N_12502,N_5848,N_6398);
and U12503 (N_12503,N_9327,N_8286);
nor U12504 (N_12504,N_7149,N_5831);
nor U12505 (N_12505,N_8853,N_5613);
xor U12506 (N_12506,N_8551,N_8844);
nand U12507 (N_12507,N_6029,N_6113);
or U12508 (N_12508,N_8383,N_5770);
nor U12509 (N_12509,N_9844,N_9851);
or U12510 (N_12510,N_7005,N_7821);
and U12511 (N_12511,N_5551,N_8599);
or U12512 (N_12512,N_7645,N_9187);
or U12513 (N_12513,N_6871,N_7483);
nand U12514 (N_12514,N_9048,N_9900);
nand U12515 (N_12515,N_6846,N_7443);
or U12516 (N_12516,N_8673,N_5935);
or U12517 (N_12517,N_6264,N_5124);
and U12518 (N_12518,N_8882,N_8896);
or U12519 (N_12519,N_9709,N_8882);
xnor U12520 (N_12520,N_9207,N_5574);
nand U12521 (N_12521,N_6924,N_6074);
and U12522 (N_12522,N_7468,N_5136);
or U12523 (N_12523,N_5376,N_5272);
or U12524 (N_12524,N_6702,N_9162);
xor U12525 (N_12525,N_7540,N_6664);
xnor U12526 (N_12526,N_7748,N_9603);
nor U12527 (N_12527,N_7259,N_5962);
or U12528 (N_12528,N_5844,N_5076);
or U12529 (N_12529,N_8247,N_7468);
or U12530 (N_12530,N_8099,N_5809);
nor U12531 (N_12531,N_5631,N_5500);
nor U12532 (N_12532,N_9451,N_9670);
nor U12533 (N_12533,N_5372,N_6185);
nor U12534 (N_12534,N_8605,N_6423);
and U12535 (N_12535,N_5177,N_9945);
or U12536 (N_12536,N_5894,N_7320);
nand U12537 (N_12537,N_5336,N_9185);
nand U12538 (N_12538,N_5182,N_5583);
or U12539 (N_12539,N_5738,N_8686);
xnor U12540 (N_12540,N_8506,N_8440);
and U12541 (N_12541,N_7522,N_7575);
nand U12542 (N_12542,N_6676,N_8096);
and U12543 (N_12543,N_6572,N_6217);
and U12544 (N_12544,N_8114,N_8669);
nand U12545 (N_12545,N_8120,N_7505);
or U12546 (N_12546,N_9597,N_7875);
and U12547 (N_12547,N_9339,N_8201);
or U12548 (N_12548,N_9587,N_7697);
nor U12549 (N_12549,N_6622,N_9483);
and U12550 (N_12550,N_7957,N_7968);
xnor U12551 (N_12551,N_7376,N_7414);
nand U12552 (N_12552,N_6557,N_7541);
nor U12553 (N_12553,N_6322,N_7005);
and U12554 (N_12554,N_5114,N_6377);
nand U12555 (N_12555,N_8515,N_8726);
nand U12556 (N_12556,N_7672,N_6994);
xnor U12557 (N_12557,N_7959,N_7231);
nand U12558 (N_12558,N_5381,N_7110);
or U12559 (N_12559,N_5883,N_6871);
or U12560 (N_12560,N_7362,N_5736);
and U12561 (N_12561,N_9864,N_7057);
xor U12562 (N_12562,N_8221,N_7342);
or U12563 (N_12563,N_8892,N_9132);
and U12564 (N_12564,N_7815,N_8321);
nor U12565 (N_12565,N_6907,N_5747);
nand U12566 (N_12566,N_9648,N_7989);
nor U12567 (N_12567,N_8958,N_5057);
nor U12568 (N_12568,N_6680,N_7841);
or U12569 (N_12569,N_8447,N_7166);
nor U12570 (N_12570,N_7659,N_7657);
and U12571 (N_12571,N_7783,N_5784);
xor U12572 (N_12572,N_7334,N_7157);
nor U12573 (N_12573,N_5957,N_5950);
nand U12574 (N_12574,N_9068,N_7082);
or U12575 (N_12575,N_8320,N_6235);
and U12576 (N_12576,N_6344,N_7641);
and U12577 (N_12577,N_8125,N_8540);
xnor U12578 (N_12578,N_7464,N_6768);
nand U12579 (N_12579,N_8944,N_8190);
or U12580 (N_12580,N_9058,N_5849);
nand U12581 (N_12581,N_8234,N_9519);
or U12582 (N_12582,N_6228,N_5970);
or U12583 (N_12583,N_9007,N_6278);
nand U12584 (N_12584,N_7409,N_7719);
and U12585 (N_12585,N_9119,N_6149);
and U12586 (N_12586,N_8832,N_6355);
nor U12587 (N_12587,N_5217,N_5510);
or U12588 (N_12588,N_9825,N_5579);
and U12589 (N_12589,N_8541,N_5770);
and U12590 (N_12590,N_8574,N_7247);
and U12591 (N_12591,N_6868,N_5886);
nor U12592 (N_12592,N_8386,N_7675);
nand U12593 (N_12593,N_5413,N_8432);
or U12594 (N_12594,N_8132,N_8540);
nor U12595 (N_12595,N_9528,N_6607);
nor U12596 (N_12596,N_8656,N_8581);
nor U12597 (N_12597,N_7027,N_7478);
nand U12598 (N_12598,N_9740,N_5523);
and U12599 (N_12599,N_9318,N_7094);
or U12600 (N_12600,N_5732,N_9739);
or U12601 (N_12601,N_8072,N_7208);
and U12602 (N_12602,N_8436,N_6818);
nor U12603 (N_12603,N_5630,N_9245);
xor U12604 (N_12604,N_6388,N_8025);
or U12605 (N_12605,N_5614,N_7937);
and U12606 (N_12606,N_9368,N_9854);
nor U12607 (N_12607,N_5450,N_7299);
nor U12608 (N_12608,N_5467,N_8037);
nand U12609 (N_12609,N_7456,N_9836);
nand U12610 (N_12610,N_5270,N_9994);
or U12611 (N_12611,N_6709,N_9626);
nor U12612 (N_12612,N_9204,N_7844);
nand U12613 (N_12613,N_8395,N_8895);
and U12614 (N_12614,N_5106,N_9192);
xor U12615 (N_12615,N_5162,N_8111);
nor U12616 (N_12616,N_6017,N_7421);
xor U12617 (N_12617,N_5595,N_7219);
and U12618 (N_12618,N_7178,N_9288);
nand U12619 (N_12619,N_6047,N_5205);
or U12620 (N_12620,N_7649,N_8816);
or U12621 (N_12621,N_9048,N_7392);
or U12622 (N_12622,N_6326,N_7986);
nand U12623 (N_12623,N_8699,N_7150);
nor U12624 (N_12624,N_7040,N_5580);
or U12625 (N_12625,N_7268,N_7592);
nand U12626 (N_12626,N_9318,N_9213);
nand U12627 (N_12627,N_6649,N_9341);
nor U12628 (N_12628,N_7484,N_6596);
and U12629 (N_12629,N_6677,N_6400);
nand U12630 (N_12630,N_9682,N_5617);
nor U12631 (N_12631,N_9101,N_8480);
nand U12632 (N_12632,N_8113,N_5236);
and U12633 (N_12633,N_9663,N_7076);
or U12634 (N_12634,N_6432,N_5074);
or U12635 (N_12635,N_7993,N_6466);
or U12636 (N_12636,N_7519,N_8279);
and U12637 (N_12637,N_5494,N_5121);
nand U12638 (N_12638,N_9757,N_8266);
nor U12639 (N_12639,N_8058,N_7635);
or U12640 (N_12640,N_9277,N_9518);
or U12641 (N_12641,N_8738,N_6163);
nand U12642 (N_12642,N_6395,N_6185);
nand U12643 (N_12643,N_9598,N_7195);
or U12644 (N_12644,N_9308,N_8241);
or U12645 (N_12645,N_9288,N_5473);
nand U12646 (N_12646,N_5964,N_9903);
or U12647 (N_12647,N_9656,N_9568);
nand U12648 (N_12648,N_6007,N_8646);
and U12649 (N_12649,N_8379,N_6416);
nand U12650 (N_12650,N_5770,N_9298);
nand U12651 (N_12651,N_6403,N_6839);
xnor U12652 (N_12652,N_7379,N_9886);
or U12653 (N_12653,N_5285,N_7112);
xor U12654 (N_12654,N_6060,N_7951);
nor U12655 (N_12655,N_8934,N_7956);
nor U12656 (N_12656,N_9119,N_6365);
xor U12657 (N_12657,N_8045,N_9645);
nand U12658 (N_12658,N_7199,N_8189);
nor U12659 (N_12659,N_5307,N_5790);
nor U12660 (N_12660,N_9341,N_7612);
or U12661 (N_12661,N_8349,N_6553);
nor U12662 (N_12662,N_7465,N_9367);
and U12663 (N_12663,N_9149,N_8850);
or U12664 (N_12664,N_5560,N_7011);
nand U12665 (N_12665,N_8191,N_5740);
nand U12666 (N_12666,N_5471,N_6293);
nor U12667 (N_12667,N_9187,N_9981);
nor U12668 (N_12668,N_9233,N_8753);
nor U12669 (N_12669,N_6255,N_7907);
xor U12670 (N_12670,N_9433,N_6996);
nand U12671 (N_12671,N_8017,N_7510);
or U12672 (N_12672,N_6796,N_8875);
nand U12673 (N_12673,N_8135,N_9646);
xor U12674 (N_12674,N_6156,N_7226);
or U12675 (N_12675,N_8870,N_9459);
nor U12676 (N_12676,N_7454,N_7293);
nor U12677 (N_12677,N_5349,N_7606);
or U12678 (N_12678,N_8573,N_7732);
nor U12679 (N_12679,N_8301,N_5042);
nand U12680 (N_12680,N_8573,N_6584);
nor U12681 (N_12681,N_7516,N_5730);
xor U12682 (N_12682,N_5966,N_7944);
xnor U12683 (N_12683,N_7238,N_8368);
or U12684 (N_12684,N_6985,N_8304);
nand U12685 (N_12685,N_9969,N_5515);
nor U12686 (N_12686,N_9178,N_9680);
nor U12687 (N_12687,N_8455,N_5125);
nor U12688 (N_12688,N_9705,N_5321);
and U12689 (N_12689,N_9316,N_6775);
or U12690 (N_12690,N_5121,N_5083);
and U12691 (N_12691,N_6191,N_8619);
nand U12692 (N_12692,N_8117,N_8359);
and U12693 (N_12693,N_5721,N_9318);
nand U12694 (N_12694,N_6216,N_5690);
nand U12695 (N_12695,N_8252,N_8694);
and U12696 (N_12696,N_7935,N_5149);
nand U12697 (N_12697,N_6105,N_7899);
nor U12698 (N_12698,N_6502,N_8471);
or U12699 (N_12699,N_5734,N_7438);
or U12700 (N_12700,N_6811,N_7192);
nand U12701 (N_12701,N_5109,N_6804);
and U12702 (N_12702,N_9560,N_9795);
or U12703 (N_12703,N_5429,N_5590);
nor U12704 (N_12704,N_9690,N_6516);
and U12705 (N_12705,N_8210,N_7198);
nor U12706 (N_12706,N_5826,N_5665);
or U12707 (N_12707,N_7863,N_9974);
or U12708 (N_12708,N_7982,N_9486);
or U12709 (N_12709,N_8425,N_8552);
and U12710 (N_12710,N_8201,N_8717);
or U12711 (N_12711,N_6609,N_9430);
or U12712 (N_12712,N_8515,N_8187);
and U12713 (N_12713,N_9620,N_6479);
nor U12714 (N_12714,N_9620,N_7774);
nand U12715 (N_12715,N_6378,N_6164);
nand U12716 (N_12716,N_9120,N_9437);
or U12717 (N_12717,N_9888,N_7692);
or U12718 (N_12718,N_9542,N_7908);
nor U12719 (N_12719,N_8685,N_8924);
or U12720 (N_12720,N_5156,N_9570);
nor U12721 (N_12721,N_9001,N_7756);
nand U12722 (N_12722,N_9005,N_7948);
and U12723 (N_12723,N_8763,N_6757);
or U12724 (N_12724,N_5633,N_7208);
or U12725 (N_12725,N_5678,N_8076);
and U12726 (N_12726,N_7223,N_6553);
nand U12727 (N_12727,N_8856,N_8925);
nand U12728 (N_12728,N_7939,N_9092);
or U12729 (N_12729,N_7307,N_8322);
nand U12730 (N_12730,N_9049,N_9384);
nand U12731 (N_12731,N_7814,N_7993);
nand U12732 (N_12732,N_6761,N_5427);
nand U12733 (N_12733,N_9483,N_5923);
nand U12734 (N_12734,N_9311,N_6343);
xnor U12735 (N_12735,N_7811,N_5971);
nor U12736 (N_12736,N_6644,N_8569);
and U12737 (N_12737,N_7688,N_8406);
and U12738 (N_12738,N_9407,N_7616);
and U12739 (N_12739,N_6767,N_9653);
and U12740 (N_12740,N_6032,N_9636);
and U12741 (N_12741,N_9238,N_5705);
nand U12742 (N_12742,N_9981,N_5827);
nand U12743 (N_12743,N_9439,N_9669);
and U12744 (N_12744,N_9906,N_7881);
and U12745 (N_12745,N_9921,N_9010);
nor U12746 (N_12746,N_6925,N_9979);
nand U12747 (N_12747,N_8786,N_9175);
or U12748 (N_12748,N_6496,N_8517);
and U12749 (N_12749,N_7619,N_5942);
nor U12750 (N_12750,N_5239,N_5003);
nand U12751 (N_12751,N_9296,N_5731);
or U12752 (N_12752,N_9943,N_8005);
and U12753 (N_12753,N_6654,N_9654);
or U12754 (N_12754,N_9506,N_7014);
and U12755 (N_12755,N_9636,N_9377);
or U12756 (N_12756,N_9766,N_5359);
and U12757 (N_12757,N_9120,N_5159);
and U12758 (N_12758,N_9509,N_9011);
nand U12759 (N_12759,N_9033,N_9306);
nand U12760 (N_12760,N_7724,N_8567);
or U12761 (N_12761,N_8728,N_7086);
and U12762 (N_12762,N_7240,N_7652);
or U12763 (N_12763,N_9614,N_5921);
and U12764 (N_12764,N_7237,N_6083);
nand U12765 (N_12765,N_6624,N_7273);
nand U12766 (N_12766,N_7331,N_8514);
nor U12767 (N_12767,N_5405,N_7142);
or U12768 (N_12768,N_9453,N_8995);
or U12769 (N_12769,N_6399,N_9232);
and U12770 (N_12770,N_6140,N_9809);
nand U12771 (N_12771,N_6522,N_7709);
nand U12772 (N_12772,N_9802,N_6140);
and U12773 (N_12773,N_8095,N_8613);
nand U12774 (N_12774,N_8698,N_7367);
xor U12775 (N_12775,N_6428,N_8558);
or U12776 (N_12776,N_7027,N_7527);
and U12777 (N_12777,N_9856,N_7778);
or U12778 (N_12778,N_7782,N_7680);
and U12779 (N_12779,N_8190,N_7614);
xnor U12780 (N_12780,N_5300,N_7456);
or U12781 (N_12781,N_9662,N_8290);
xnor U12782 (N_12782,N_6514,N_5164);
nand U12783 (N_12783,N_8042,N_6697);
and U12784 (N_12784,N_8511,N_7051);
nor U12785 (N_12785,N_8032,N_7893);
nand U12786 (N_12786,N_7583,N_5017);
nand U12787 (N_12787,N_7445,N_7683);
nor U12788 (N_12788,N_7602,N_6850);
or U12789 (N_12789,N_7254,N_9420);
and U12790 (N_12790,N_8524,N_6716);
nor U12791 (N_12791,N_5580,N_7970);
or U12792 (N_12792,N_5163,N_7614);
nand U12793 (N_12793,N_7300,N_6596);
nor U12794 (N_12794,N_6430,N_6785);
nor U12795 (N_12795,N_9338,N_7007);
nand U12796 (N_12796,N_8082,N_6580);
or U12797 (N_12797,N_7817,N_5075);
nor U12798 (N_12798,N_7843,N_8161);
xnor U12799 (N_12799,N_8932,N_6629);
nand U12800 (N_12800,N_6397,N_9737);
nand U12801 (N_12801,N_7017,N_9457);
nor U12802 (N_12802,N_5700,N_7159);
and U12803 (N_12803,N_8489,N_9305);
nand U12804 (N_12804,N_5726,N_6490);
and U12805 (N_12805,N_8498,N_5228);
nor U12806 (N_12806,N_5823,N_7769);
or U12807 (N_12807,N_5692,N_7582);
or U12808 (N_12808,N_9622,N_8834);
xor U12809 (N_12809,N_8314,N_5926);
nor U12810 (N_12810,N_5000,N_7912);
nor U12811 (N_12811,N_9702,N_5786);
nand U12812 (N_12812,N_7257,N_9258);
xor U12813 (N_12813,N_8037,N_9559);
nor U12814 (N_12814,N_6770,N_9563);
nor U12815 (N_12815,N_5783,N_7250);
and U12816 (N_12816,N_7659,N_7328);
and U12817 (N_12817,N_7285,N_9226);
or U12818 (N_12818,N_7376,N_9506);
nor U12819 (N_12819,N_7370,N_8041);
and U12820 (N_12820,N_6573,N_6614);
or U12821 (N_12821,N_8037,N_9859);
nand U12822 (N_12822,N_8406,N_7966);
or U12823 (N_12823,N_9730,N_7675);
and U12824 (N_12824,N_9759,N_8721);
or U12825 (N_12825,N_9470,N_5936);
and U12826 (N_12826,N_6197,N_5571);
and U12827 (N_12827,N_8178,N_8374);
nand U12828 (N_12828,N_5652,N_7685);
nor U12829 (N_12829,N_8519,N_6868);
nand U12830 (N_12830,N_5990,N_8772);
and U12831 (N_12831,N_5144,N_8344);
nand U12832 (N_12832,N_8390,N_9253);
nand U12833 (N_12833,N_6744,N_7837);
nand U12834 (N_12834,N_8118,N_6388);
nand U12835 (N_12835,N_5489,N_8528);
nor U12836 (N_12836,N_9646,N_7145);
nor U12837 (N_12837,N_6297,N_5865);
and U12838 (N_12838,N_6917,N_9720);
or U12839 (N_12839,N_5756,N_9473);
and U12840 (N_12840,N_5823,N_6711);
nand U12841 (N_12841,N_5763,N_8028);
and U12842 (N_12842,N_8109,N_8643);
or U12843 (N_12843,N_8991,N_9091);
or U12844 (N_12844,N_7415,N_8895);
and U12845 (N_12845,N_8518,N_6864);
nor U12846 (N_12846,N_5414,N_9493);
nand U12847 (N_12847,N_6976,N_6696);
and U12848 (N_12848,N_7080,N_9911);
or U12849 (N_12849,N_6962,N_8253);
nor U12850 (N_12850,N_9642,N_8137);
nor U12851 (N_12851,N_7896,N_6406);
or U12852 (N_12852,N_8823,N_8266);
and U12853 (N_12853,N_8624,N_8192);
nand U12854 (N_12854,N_9789,N_6894);
or U12855 (N_12855,N_8097,N_6990);
nor U12856 (N_12856,N_9558,N_6740);
nand U12857 (N_12857,N_8804,N_8083);
or U12858 (N_12858,N_9303,N_7299);
or U12859 (N_12859,N_6264,N_6232);
and U12860 (N_12860,N_5353,N_5666);
nor U12861 (N_12861,N_5445,N_5980);
or U12862 (N_12862,N_5477,N_9209);
and U12863 (N_12863,N_6499,N_7562);
nand U12864 (N_12864,N_8232,N_8670);
nand U12865 (N_12865,N_5059,N_7083);
and U12866 (N_12866,N_9362,N_9729);
nor U12867 (N_12867,N_9598,N_6029);
xor U12868 (N_12868,N_5463,N_6422);
xor U12869 (N_12869,N_6686,N_8875);
nor U12870 (N_12870,N_6823,N_6355);
nor U12871 (N_12871,N_8677,N_5985);
and U12872 (N_12872,N_7608,N_7979);
or U12873 (N_12873,N_5089,N_9459);
and U12874 (N_12874,N_9314,N_5350);
nor U12875 (N_12875,N_5223,N_9907);
nor U12876 (N_12876,N_9335,N_6869);
or U12877 (N_12877,N_7660,N_7804);
nand U12878 (N_12878,N_8316,N_5184);
nand U12879 (N_12879,N_9500,N_7700);
or U12880 (N_12880,N_9186,N_9479);
nand U12881 (N_12881,N_6882,N_8359);
nand U12882 (N_12882,N_5867,N_8240);
xnor U12883 (N_12883,N_9100,N_6457);
nor U12884 (N_12884,N_8495,N_5734);
nor U12885 (N_12885,N_5781,N_8046);
nor U12886 (N_12886,N_9216,N_8908);
nor U12887 (N_12887,N_5939,N_6545);
nor U12888 (N_12888,N_8743,N_9763);
nor U12889 (N_12889,N_8853,N_8040);
xor U12890 (N_12890,N_8637,N_8510);
xor U12891 (N_12891,N_6969,N_8196);
or U12892 (N_12892,N_9253,N_6063);
or U12893 (N_12893,N_7186,N_8416);
nor U12894 (N_12894,N_7807,N_6717);
and U12895 (N_12895,N_6003,N_7191);
and U12896 (N_12896,N_7841,N_8928);
nand U12897 (N_12897,N_8168,N_6916);
and U12898 (N_12898,N_9208,N_9476);
and U12899 (N_12899,N_5997,N_6858);
or U12900 (N_12900,N_7069,N_5716);
nor U12901 (N_12901,N_6922,N_8506);
or U12902 (N_12902,N_8335,N_5624);
nand U12903 (N_12903,N_5463,N_8948);
and U12904 (N_12904,N_8705,N_7263);
nor U12905 (N_12905,N_5350,N_9416);
nand U12906 (N_12906,N_6627,N_6283);
nor U12907 (N_12907,N_7395,N_5837);
nand U12908 (N_12908,N_9167,N_6335);
and U12909 (N_12909,N_9995,N_6149);
xor U12910 (N_12910,N_7706,N_7295);
nand U12911 (N_12911,N_7249,N_8973);
or U12912 (N_12912,N_7072,N_7618);
nand U12913 (N_12913,N_8413,N_8271);
and U12914 (N_12914,N_9179,N_6061);
xor U12915 (N_12915,N_8359,N_7329);
nor U12916 (N_12916,N_8328,N_6955);
nand U12917 (N_12917,N_8466,N_9913);
nand U12918 (N_12918,N_6959,N_5202);
nor U12919 (N_12919,N_9551,N_8050);
or U12920 (N_12920,N_6739,N_7192);
xnor U12921 (N_12921,N_5849,N_8648);
and U12922 (N_12922,N_7310,N_8502);
xor U12923 (N_12923,N_7975,N_9330);
nand U12924 (N_12924,N_9115,N_7458);
nand U12925 (N_12925,N_9032,N_8453);
and U12926 (N_12926,N_6359,N_5260);
xnor U12927 (N_12927,N_9853,N_8976);
and U12928 (N_12928,N_5767,N_9047);
nand U12929 (N_12929,N_9334,N_7280);
nor U12930 (N_12930,N_5820,N_8352);
nand U12931 (N_12931,N_8996,N_6870);
and U12932 (N_12932,N_6431,N_6576);
xnor U12933 (N_12933,N_8834,N_9343);
nand U12934 (N_12934,N_9884,N_5244);
nand U12935 (N_12935,N_8663,N_8172);
nor U12936 (N_12936,N_7286,N_7601);
and U12937 (N_12937,N_6779,N_9764);
nor U12938 (N_12938,N_9247,N_9039);
nor U12939 (N_12939,N_7694,N_9114);
nor U12940 (N_12940,N_5515,N_9345);
and U12941 (N_12941,N_7398,N_8372);
xor U12942 (N_12942,N_8824,N_9682);
or U12943 (N_12943,N_5269,N_7469);
and U12944 (N_12944,N_9702,N_8426);
and U12945 (N_12945,N_7134,N_6843);
or U12946 (N_12946,N_7564,N_6430);
xor U12947 (N_12947,N_7696,N_8655);
xnor U12948 (N_12948,N_6883,N_7196);
nor U12949 (N_12949,N_6682,N_7421);
or U12950 (N_12950,N_5633,N_8817);
and U12951 (N_12951,N_6098,N_6184);
nand U12952 (N_12952,N_8390,N_5852);
nor U12953 (N_12953,N_9922,N_5830);
nor U12954 (N_12954,N_5960,N_6944);
or U12955 (N_12955,N_8377,N_8519);
or U12956 (N_12956,N_5152,N_6280);
nor U12957 (N_12957,N_9663,N_6057);
or U12958 (N_12958,N_5149,N_9248);
or U12959 (N_12959,N_7990,N_6333);
or U12960 (N_12960,N_5193,N_9624);
or U12961 (N_12961,N_5727,N_8155);
nor U12962 (N_12962,N_6934,N_8284);
nand U12963 (N_12963,N_6133,N_8273);
and U12964 (N_12964,N_6109,N_8168);
nand U12965 (N_12965,N_7496,N_8694);
nor U12966 (N_12966,N_7081,N_8391);
or U12967 (N_12967,N_7380,N_6376);
nor U12968 (N_12968,N_9573,N_6933);
nand U12969 (N_12969,N_7983,N_9022);
or U12970 (N_12970,N_6718,N_6232);
xor U12971 (N_12971,N_7906,N_8580);
or U12972 (N_12972,N_7927,N_8412);
nor U12973 (N_12973,N_7528,N_8006);
nor U12974 (N_12974,N_6830,N_8785);
nor U12975 (N_12975,N_7995,N_9101);
nand U12976 (N_12976,N_7681,N_9225);
nor U12977 (N_12977,N_5666,N_9581);
xnor U12978 (N_12978,N_5514,N_9902);
or U12979 (N_12979,N_6642,N_7201);
nor U12980 (N_12980,N_7755,N_6704);
nand U12981 (N_12981,N_8903,N_9615);
nand U12982 (N_12982,N_6568,N_5843);
and U12983 (N_12983,N_9903,N_6293);
nand U12984 (N_12984,N_9845,N_9579);
nor U12985 (N_12985,N_6777,N_6550);
and U12986 (N_12986,N_5182,N_9597);
or U12987 (N_12987,N_8715,N_9359);
and U12988 (N_12988,N_8351,N_7972);
nor U12989 (N_12989,N_6073,N_7757);
or U12990 (N_12990,N_5527,N_5493);
nor U12991 (N_12991,N_5489,N_8591);
and U12992 (N_12992,N_7939,N_8850);
and U12993 (N_12993,N_7930,N_8535);
nor U12994 (N_12994,N_5159,N_9066);
nand U12995 (N_12995,N_9450,N_9128);
and U12996 (N_12996,N_9935,N_8487);
and U12997 (N_12997,N_7186,N_5433);
nor U12998 (N_12998,N_7123,N_7708);
xnor U12999 (N_12999,N_9500,N_6125);
or U13000 (N_13000,N_9185,N_7009);
nor U13001 (N_13001,N_9747,N_8082);
and U13002 (N_13002,N_5998,N_7117);
nand U13003 (N_13003,N_7176,N_8264);
nor U13004 (N_13004,N_9377,N_6427);
nand U13005 (N_13005,N_6919,N_6496);
xor U13006 (N_13006,N_8197,N_8745);
and U13007 (N_13007,N_6236,N_5945);
nand U13008 (N_13008,N_8531,N_9821);
nand U13009 (N_13009,N_6026,N_8566);
xor U13010 (N_13010,N_6197,N_5907);
or U13011 (N_13011,N_7651,N_7579);
and U13012 (N_13012,N_6469,N_7470);
or U13013 (N_13013,N_9455,N_5954);
and U13014 (N_13014,N_5880,N_8096);
and U13015 (N_13015,N_8897,N_6117);
and U13016 (N_13016,N_7298,N_9752);
or U13017 (N_13017,N_8107,N_9726);
and U13018 (N_13018,N_5239,N_6123);
and U13019 (N_13019,N_6231,N_8916);
and U13020 (N_13020,N_5174,N_9756);
nand U13021 (N_13021,N_5140,N_5867);
and U13022 (N_13022,N_7514,N_6184);
or U13023 (N_13023,N_9005,N_7692);
nor U13024 (N_13024,N_5881,N_6128);
and U13025 (N_13025,N_6600,N_6424);
xor U13026 (N_13026,N_8462,N_9671);
nor U13027 (N_13027,N_9037,N_8851);
xor U13028 (N_13028,N_5342,N_8913);
or U13029 (N_13029,N_8362,N_6599);
or U13030 (N_13030,N_7832,N_8784);
nor U13031 (N_13031,N_6855,N_7288);
nor U13032 (N_13032,N_6927,N_7301);
nand U13033 (N_13033,N_5409,N_8879);
and U13034 (N_13034,N_6609,N_8266);
nand U13035 (N_13035,N_5374,N_9216);
or U13036 (N_13036,N_7242,N_5257);
and U13037 (N_13037,N_7339,N_8287);
nor U13038 (N_13038,N_6979,N_7244);
nand U13039 (N_13039,N_5678,N_6311);
nand U13040 (N_13040,N_5071,N_6229);
and U13041 (N_13041,N_9985,N_9755);
nand U13042 (N_13042,N_8375,N_8506);
nor U13043 (N_13043,N_9980,N_7821);
nand U13044 (N_13044,N_5291,N_7359);
and U13045 (N_13045,N_5137,N_9051);
nand U13046 (N_13046,N_6160,N_7038);
or U13047 (N_13047,N_7884,N_7193);
nand U13048 (N_13048,N_9553,N_6077);
xnor U13049 (N_13049,N_6650,N_5970);
nand U13050 (N_13050,N_7014,N_7137);
xnor U13051 (N_13051,N_6922,N_8079);
nor U13052 (N_13052,N_5051,N_6760);
nor U13053 (N_13053,N_9586,N_8919);
nor U13054 (N_13054,N_7380,N_6973);
nor U13055 (N_13055,N_6041,N_5836);
nor U13056 (N_13056,N_7025,N_5605);
nor U13057 (N_13057,N_5416,N_6202);
xnor U13058 (N_13058,N_5284,N_7481);
or U13059 (N_13059,N_6675,N_7629);
and U13060 (N_13060,N_8632,N_7972);
or U13061 (N_13061,N_9395,N_5535);
nor U13062 (N_13062,N_8596,N_5841);
and U13063 (N_13063,N_5677,N_7212);
and U13064 (N_13064,N_7271,N_9366);
nand U13065 (N_13065,N_5116,N_7565);
and U13066 (N_13066,N_9490,N_7544);
nor U13067 (N_13067,N_6582,N_5580);
and U13068 (N_13068,N_8531,N_5879);
or U13069 (N_13069,N_6131,N_8490);
xnor U13070 (N_13070,N_8605,N_5301);
and U13071 (N_13071,N_9131,N_5809);
nor U13072 (N_13072,N_5939,N_7362);
nand U13073 (N_13073,N_9861,N_7811);
nor U13074 (N_13074,N_6492,N_9734);
or U13075 (N_13075,N_7385,N_5019);
or U13076 (N_13076,N_9524,N_7129);
xnor U13077 (N_13077,N_5224,N_5934);
nand U13078 (N_13078,N_6219,N_8501);
or U13079 (N_13079,N_6806,N_7806);
or U13080 (N_13080,N_9081,N_7990);
and U13081 (N_13081,N_6455,N_6559);
and U13082 (N_13082,N_9811,N_6763);
nor U13083 (N_13083,N_5444,N_9810);
and U13084 (N_13084,N_9511,N_9938);
nand U13085 (N_13085,N_7742,N_8049);
and U13086 (N_13086,N_7831,N_5041);
and U13087 (N_13087,N_8824,N_9275);
or U13088 (N_13088,N_7227,N_5584);
or U13089 (N_13089,N_8022,N_9513);
nor U13090 (N_13090,N_6030,N_6763);
nand U13091 (N_13091,N_5981,N_8383);
nand U13092 (N_13092,N_5530,N_7593);
and U13093 (N_13093,N_9023,N_6227);
or U13094 (N_13094,N_5095,N_5155);
nand U13095 (N_13095,N_5009,N_5455);
and U13096 (N_13096,N_7479,N_7242);
nand U13097 (N_13097,N_6388,N_8603);
nand U13098 (N_13098,N_8530,N_9406);
nor U13099 (N_13099,N_8884,N_7002);
or U13100 (N_13100,N_9838,N_7347);
nor U13101 (N_13101,N_7998,N_9572);
nor U13102 (N_13102,N_9085,N_8229);
nand U13103 (N_13103,N_7738,N_8673);
nor U13104 (N_13104,N_9351,N_8662);
nor U13105 (N_13105,N_9929,N_6372);
and U13106 (N_13106,N_8877,N_5856);
nand U13107 (N_13107,N_6927,N_5645);
and U13108 (N_13108,N_6594,N_6090);
or U13109 (N_13109,N_5531,N_9322);
and U13110 (N_13110,N_9892,N_5880);
nor U13111 (N_13111,N_7073,N_7891);
nand U13112 (N_13112,N_8962,N_5841);
nand U13113 (N_13113,N_6644,N_6465);
nand U13114 (N_13114,N_5013,N_8725);
and U13115 (N_13115,N_8532,N_5271);
and U13116 (N_13116,N_6182,N_8249);
xnor U13117 (N_13117,N_7897,N_6629);
nor U13118 (N_13118,N_8432,N_9895);
nor U13119 (N_13119,N_7437,N_7984);
nand U13120 (N_13120,N_7434,N_9073);
nand U13121 (N_13121,N_9966,N_7125);
xnor U13122 (N_13122,N_9336,N_5792);
nand U13123 (N_13123,N_9335,N_6637);
or U13124 (N_13124,N_9821,N_6947);
or U13125 (N_13125,N_7662,N_7411);
nand U13126 (N_13126,N_6027,N_6897);
or U13127 (N_13127,N_5490,N_9039);
or U13128 (N_13128,N_7991,N_5707);
nand U13129 (N_13129,N_9805,N_7584);
nand U13130 (N_13130,N_9823,N_9963);
nor U13131 (N_13131,N_8871,N_5578);
nor U13132 (N_13132,N_7683,N_7192);
or U13133 (N_13133,N_5630,N_6130);
or U13134 (N_13134,N_9340,N_7866);
nor U13135 (N_13135,N_6531,N_6512);
or U13136 (N_13136,N_9810,N_7870);
or U13137 (N_13137,N_7662,N_6685);
or U13138 (N_13138,N_8283,N_5433);
nand U13139 (N_13139,N_9899,N_7939);
xnor U13140 (N_13140,N_7580,N_6366);
nor U13141 (N_13141,N_7595,N_8137);
nor U13142 (N_13142,N_7032,N_7088);
or U13143 (N_13143,N_7875,N_7053);
nand U13144 (N_13144,N_9507,N_9249);
nor U13145 (N_13145,N_5988,N_9814);
and U13146 (N_13146,N_9413,N_6577);
nand U13147 (N_13147,N_9188,N_9460);
or U13148 (N_13148,N_5025,N_9096);
nor U13149 (N_13149,N_5771,N_7613);
nor U13150 (N_13150,N_9372,N_9106);
and U13151 (N_13151,N_8743,N_9686);
xnor U13152 (N_13152,N_5214,N_7457);
and U13153 (N_13153,N_6571,N_9232);
and U13154 (N_13154,N_7688,N_8831);
nor U13155 (N_13155,N_5110,N_7959);
nor U13156 (N_13156,N_7745,N_5283);
nand U13157 (N_13157,N_9012,N_5365);
and U13158 (N_13158,N_5847,N_6334);
nand U13159 (N_13159,N_6388,N_5172);
nand U13160 (N_13160,N_6043,N_7120);
nor U13161 (N_13161,N_7681,N_7480);
nor U13162 (N_13162,N_8146,N_6642);
and U13163 (N_13163,N_8408,N_8089);
and U13164 (N_13164,N_7447,N_6105);
xor U13165 (N_13165,N_5125,N_9705);
nand U13166 (N_13166,N_6870,N_5322);
nor U13167 (N_13167,N_8537,N_7935);
nor U13168 (N_13168,N_5783,N_7757);
and U13169 (N_13169,N_9133,N_5225);
nor U13170 (N_13170,N_8380,N_8597);
nor U13171 (N_13171,N_7453,N_7360);
and U13172 (N_13172,N_6257,N_6154);
nor U13173 (N_13173,N_8031,N_7223);
nor U13174 (N_13174,N_8705,N_8006);
or U13175 (N_13175,N_7523,N_8312);
or U13176 (N_13176,N_7139,N_9043);
xor U13177 (N_13177,N_9754,N_5087);
or U13178 (N_13178,N_8666,N_9268);
and U13179 (N_13179,N_5315,N_6100);
and U13180 (N_13180,N_5674,N_5972);
nand U13181 (N_13181,N_8843,N_7285);
and U13182 (N_13182,N_5237,N_6525);
nand U13183 (N_13183,N_7896,N_9454);
or U13184 (N_13184,N_9561,N_9832);
and U13185 (N_13185,N_9733,N_7137);
or U13186 (N_13186,N_8116,N_6066);
nor U13187 (N_13187,N_9772,N_9232);
xor U13188 (N_13188,N_8053,N_6741);
or U13189 (N_13189,N_6651,N_8327);
nand U13190 (N_13190,N_5373,N_7658);
and U13191 (N_13191,N_6501,N_6790);
and U13192 (N_13192,N_6091,N_8893);
nand U13193 (N_13193,N_8710,N_7394);
and U13194 (N_13194,N_5056,N_7771);
nand U13195 (N_13195,N_5206,N_7369);
or U13196 (N_13196,N_8813,N_5155);
or U13197 (N_13197,N_9672,N_7555);
nor U13198 (N_13198,N_8882,N_8285);
and U13199 (N_13199,N_5192,N_7622);
or U13200 (N_13200,N_6595,N_5202);
or U13201 (N_13201,N_7899,N_6060);
and U13202 (N_13202,N_8216,N_5960);
or U13203 (N_13203,N_6854,N_5933);
and U13204 (N_13204,N_8459,N_5331);
and U13205 (N_13205,N_6313,N_8559);
or U13206 (N_13206,N_7118,N_5002);
or U13207 (N_13207,N_8861,N_8088);
or U13208 (N_13208,N_8645,N_9191);
nor U13209 (N_13209,N_6083,N_9897);
and U13210 (N_13210,N_7139,N_6467);
nor U13211 (N_13211,N_6222,N_7100);
and U13212 (N_13212,N_7799,N_7806);
nor U13213 (N_13213,N_6922,N_6574);
and U13214 (N_13214,N_7955,N_6824);
nand U13215 (N_13215,N_5463,N_9806);
xnor U13216 (N_13216,N_9223,N_9090);
nor U13217 (N_13217,N_8548,N_5256);
nand U13218 (N_13218,N_6553,N_9498);
xnor U13219 (N_13219,N_6032,N_8851);
nor U13220 (N_13220,N_9042,N_7997);
or U13221 (N_13221,N_6144,N_5998);
xor U13222 (N_13222,N_9169,N_5169);
or U13223 (N_13223,N_5382,N_8760);
nor U13224 (N_13224,N_5175,N_6065);
nand U13225 (N_13225,N_8226,N_6991);
nand U13226 (N_13226,N_7252,N_6107);
nand U13227 (N_13227,N_9148,N_7046);
nor U13228 (N_13228,N_5952,N_7044);
and U13229 (N_13229,N_8302,N_8269);
or U13230 (N_13230,N_9600,N_6379);
or U13231 (N_13231,N_5685,N_7937);
nand U13232 (N_13232,N_5866,N_8468);
and U13233 (N_13233,N_9115,N_9276);
or U13234 (N_13234,N_6501,N_6569);
nor U13235 (N_13235,N_6919,N_7788);
and U13236 (N_13236,N_7525,N_5398);
and U13237 (N_13237,N_9230,N_7829);
and U13238 (N_13238,N_9671,N_6423);
xor U13239 (N_13239,N_6245,N_6267);
and U13240 (N_13240,N_6341,N_8887);
and U13241 (N_13241,N_6271,N_9035);
xnor U13242 (N_13242,N_9329,N_8088);
xor U13243 (N_13243,N_5660,N_6411);
and U13244 (N_13244,N_6086,N_9713);
xor U13245 (N_13245,N_7366,N_6392);
nand U13246 (N_13246,N_8330,N_9738);
and U13247 (N_13247,N_5110,N_6102);
nor U13248 (N_13248,N_6699,N_7756);
nor U13249 (N_13249,N_9458,N_7593);
and U13250 (N_13250,N_5773,N_6205);
nand U13251 (N_13251,N_6161,N_8943);
nor U13252 (N_13252,N_9841,N_9130);
nand U13253 (N_13253,N_6570,N_5631);
nand U13254 (N_13254,N_7392,N_7733);
or U13255 (N_13255,N_9017,N_5680);
and U13256 (N_13256,N_7804,N_5871);
and U13257 (N_13257,N_6792,N_5339);
or U13258 (N_13258,N_8390,N_6086);
and U13259 (N_13259,N_6606,N_8838);
and U13260 (N_13260,N_8744,N_5748);
xor U13261 (N_13261,N_5726,N_7492);
and U13262 (N_13262,N_8008,N_7492);
and U13263 (N_13263,N_6301,N_6160);
nand U13264 (N_13264,N_7844,N_5609);
xor U13265 (N_13265,N_6085,N_9741);
and U13266 (N_13266,N_5574,N_9562);
or U13267 (N_13267,N_5523,N_7333);
nand U13268 (N_13268,N_8951,N_5389);
or U13269 (N_13269,N_7051,N_9478);
xor U13270 (N_13270,N_5143,N_5242);
nand U13271 (N_13271,N_9443,N_9897);
nor U13272 (N_13272,N_9623,N_5002);
xor U13273 (N_13273,N_7437,N_9282);
or U13274 (N_13274,N_5660,N_7917);
or U13275 (N_13275,N_7662,N_9279);
nor U13276 (N_13276,N_7610,N_9127);
and U13277 (N_13277,N_9827,N_9574);
nor U13278 (N_13278,N_7577,N_6750);
and U13279 (N_13279,N_5733,N_9180);
or U13280 (N_13280,N_6530,N_9096);
or U13281 (N_13281,N_8518,N_8707);
nand U13282 (N_13282,N_5808,N_5533);
nand U13283 (N_13283,N_6481,N_8932);
nor U13284 (N_13284,N_8012,N_5851);
and U13285 (N_13285,N_9158,N_9618);
nand U13286 (N_13286,N_9033,N_5243);
or U13287 (N_13287,N_7351,N_8904);
nor U13288 (N_13288,N_8516,N_7516);
nor U13289 (N_13289,N_9505,N_5857);
nor U13290 (N_13290,N_7335,N_6302);
and U13291 (N_13291,N_9368,N_8758);
xor U13292 (N_13292,N_5561,N_5524);
or U13293 (N_13293,N_9343,N_7850);
nor U13294 (N_13294,N_9256,N_6334);
nor U13295 (N_13295,N_8102,N_7820);
and U13296 (N_13296,N_7021,N_6910);
or U13297 (N_13297,N_5625,N_5353);
nand U13298 (N_13298,N_8505,N_7780);
or U13299 (N_13299,N_5657,N_9249);
or U13300 (N_13300,N_8797,N_6257);
xnor U13301 (N_13301,N_9644,N_9160);
or U13302 (N_13302,N_9341,N_8042);
xor U13303 (N_13303,N_5287,N_6088);
or U13304 (N_13304,N_8510,N_8176);
nor U13305 (N_13305,N_8119,N_8273);
nor U13306 (N_13306,N_5913,N_5123);
nand U13307 (N_13307,N_6151,N_8945);
xor U13308 (N_13308,N_6840,N_6772);
nor U13309 (N_13309,N_8368,N_6318);
and U13310 (N_13310,N_9102,N_6220);
and U13311 (N_13311,N_9544,N_7499);
xnor U13312 (N_13312,N_8778,N_9244);
nand U13313 (N_13313,N_8119,N_8277);
or U13314 (N_13314,N_8443,N_5611);
nand U13315 (N_13315,N_8067,N_6854);
nor U13316 (N_13316,N_6705,N_6053);
or U13317 (N_13317,N_8019,N_9012);
and U13318 (N_13318,N_8014,N_6855);
and U13319 (N_13319,N_5571,N_8583);
nand U13320 (N_13320,N_8410,N_8376);
nor U13321 (N_13321,N_5089,N_8647);
nand U13322 (N_13322,N_5021,N_5592);
nand U13323 (N_13323,N_9542,N_6846);
nor U13324 (N_13324,N_8064,N_8796);
and U13325 (N_13325,N_5955,N_8594);
and U13326 (N_13326,N_6549,N_7469);
and U13327 (N_13327,N_5441,N_6740);
or U13328 (N_13328,N_7457,N_8380);
nor U13329 (N_13329,N_5177,N_6469);
or U13330 (N_13330,N_7353,N_6990);
or U13331 (N_13331,N_6094,N_8541);
nor U13332 (N_13332,N_5049,N_7609);
xor U13333 (N_13333,N_9961,N_5999);
nor U13334 (N_13334,N_8350,N_9082);
nand U13335 (N_13335,N_6409,N_7102);
or U13336 (N_13336,N_7237,N_6017);
nor U13337 (N_13337,N_8974,N_8635);
and U13338 (N_13338,N_5949,N_7124);
nand U13339 (N_13339,N_7836,N_5770);
nor U13340 (N_13340,N_7518,N_8728);
xnor U13341 (N_13341,N_9543,N_7147);
nand U13342 (N_13342,N_7827,N_6275);
nand U13343 (N_13343,N_8912,N_5548);
nor U13344 (N_13344,N_6064,N_8776);
nor U13345 (N_13345,N_9111,N_8176);
and U13346 (N_13346,N_8397,N_6824);
nor U13347 (N_13347,N_5177,N_7378);
nand U13348 (N_13348,N_6605,N_8654);
nand U13349 (N_13349,N_9850,N_9140);
nand U13350 (N_13350,N_6441,N_9626);
nor U13351 (N_13351,N_8734,N_9627);
or U13352 (N_13352,N_5438,N_6724);
or U13353 (N_13353,N_9139,N_8769);
nand U13354 (N_13354,N_8418,N_5412);
nand U13355 (N_13355,N_8993,N_6425);
and U13356 (N_13356,N_6495,N_9144);
nand U13357 (N_13357,N_9238,N_6874);
or U13358 (N_13358,N_5521,N_8289);
nor U13359 (N_13359,N_5855,N_5637);
nor U13360 (N_13360,N_6180,N_8187);
nor U13361 (N_13361,N_6451,N_8013);
and U13362 (N_13362,N_5071,N_7151);
or U13363 (N_13363,N_8659,N_8564);
nor U13364 (N_13364,N_5893,N_5729);
or U13365 (N_13365,N_7328,N_9910);
nor U13366 (N_13366,N_5580,N_6746);
or U13367 (N_13367,N_7782,N_6007);
nand U13368 (N_13368,N_9276,N_8235);
nor U13369 (N_13369,N_9488,N_6837);
and U13370 (N_13370,N_9784,N_9843);
and U13371 (N_13371,N_8307,N_5333);
and U13372 (N_13372,N_7653,N_8092);
and U13373 (N_13373,N_9225,N_6593);
nand U13374 (N_13374,N_6316,N_7535);
and U13375 (N_13375,N_7281,N_5811);
and U13376 (N_13376,N_8849,N_9734);
xor U13377 (N_13377,N_8539,N_6044);
xor U13378 (N_13378,N_9333,N_9105);
and U13379 (N_13379,N_5188,N_7820);
and U13380 (N_13380,N_5586,N_9227);
nor U13381 (N_13381,N_9378,N_9717);
or U13382 (N_13382,N_9830,N_8131);
nor U13383 (N_13383,N_8446,N_6869);
nand U13384 (N_13384,N_9969,N_5570);
or U13385 (N_13385,N_7412,N_6587);
and U13386 (N_13386,N_9403,N_8949);
nand U13387 (N_13387,N_8648,N_7806);
nor U13388 (N_13388,N_8281,N_7450);
nand U13389 (N_13389,N_6758,N_6569);
and U13390 (N_13390,N_9761,N_9682);
or U13391 (N_13391,N_5187,N_8340);
or U13392 (N_13392,N_6933,N_7329);
or U13393 (N_13393,N_8541,N_8890);
or U13394 (N_13394,N_5075,N_7756);
nand U13395 (N_13395,N_6393,N_6476);
nand U13396 (N_13396,N_6241,N_6464);
and U13397 (N_13397,N_8443,N_5107);
or U13398 (N_13398,N_7022,N_8420);
or U13399 (N_13399,N_9549,N_7109);
nor U13400 (N_13400,N_6867,N_6960);
or U13401 (N_13401,N_5193,N_8449);
nand U13402 (N_13402,N_5586,N_5996);
or U13403 (N_13403,N_9163,N_7367);
or U13404 (N_13404,N_6361,N_6745);
and U13405 (N_13405,N_6598,N_7731);
and U13406 (N_13406,N_9855,N_6693);
nand U13407 (N_13407,N_9357,N_7236);
or U13408 (N_13408,N_6733,N_6275);
nor U13409 (N_13409,N_8926,N_8647);
nand U13410 (N_13410,N_8339,N_6744);
nor U13411 (N_13411,N_8191,N_9446);
and U13412 (N_13412,N_9401,N_5592);
and U13413 (N_13413,N_9881,N_9530);
nand U13414 (N_13414,N_8219,N_5092);
xnor U13415 (N_13415,N_9735,N_9295);
and U13416 (N_13416,N_7490,N_6723);
nor U13417 (N_13417,N_9140,N_9888);
nand U13418 (N_13418,N_9267,N_5916);
nor U13419 (N_13419,N_7190,N_8781);
xor U13420 (N_13420,N_6392,N_7718);
nand U13421 (N_13421,N_6014,N_8110);
nor U13422 (N_13422,N_7703,N_8560);
and U13423 (N_13423,N_7410,N_5266);
xor U13424 (N_13424,N_5267,N_6208);
nand U13425 (N_13425,N_6449,N_8408);
xnor U13426 (N_13426,N_9348,N_5404);
nor U13427 (N_13427,N_8228,N_6051);
or U13428 (N_13428,N_8682,N_8556);
xnor U13429 (N_13429,N_9491,N_8793);
nand U13430 (N_13430,N_5095,N_8830);
nor U13431 (N_13431,N_8990,N_5135);
nand U13432 (N_13432,N_9347,N_9825);
xor U13433 (N_13433,N_8183,N_7002);
nand U13434 (N_13434,N_8151,N_5983);
or U13435 (N_13435,N_7975,N_6306);
or U13436 (N_13436,N_8984,N_9537);
or U13437 (N_13437,N_5541,N_6867);
and U13438 (N_13438,N_5945,N_6095);
nor U13439 (N_13439,N_6441,N_7928);
nor U13440 (N_13440,N_5112,N_9778);
nand U13441 (N_13441,N_9747,N_5968);
nand U13442 (N_13442,N_9124,N_8821);
nand U13443 (N_13443,N_8920,N_5372);
nor U13444 (N_13444,N_5385,N_7247);
or U13445 (N_13445,N_8325,N_8548);
xnor U13446 (N_13446,N_5186,N_7715);
xnor U13447 (N_13447,N_8797,N_5071);
nand U13448 (N_13448,N_6663,N_8807);
or U13449 (N_13449,N_8151,N_9728);
nand U13450 (N_13450,N_9760,N_7368);
nor U13451 (N_13451,N_8345,N_6048);
and U13452 (N_13452,N_5722,N_9469);
nor U13453 (N_13453,N_8065,N_6965);
or U13454 (N_13454,N_6842,N_9363);
and U13455 (N_13455,N_6472,N_7883);
and U13456 (N_13456,N_7600,N_6478);
or U13457 (N_13457,N_9595,N_5803);
xor U13458 (N_13458,N_9694,N_9473);
nand U13459 (N_13459,N_8957,N_8666);
or U13460 (N_13460,N_5889,N_5399);
nor U13461 (N_13461,N_7218,N_5577);
or U13462 (N_13462,N_9388,N_9865);
nor U13463 (N_13463,N_7880,N_6960);
or U13464 (N_13464,N_8293,N_9817);
nor U13465 (N_13465,N_8689,N_7884);
or U13466 (N_13466,N_8619,N_5743);
nand U13467 (N_13467,N_7328,N_7070);
nor U13468 (N_13468,N_8055,N_6876);
nand U13469 (N_13469,N_7325,N_6965);
and U13470 (N_13470,N_5210,N_7296);
nand U13471 (N_13471,N_5490,N_5712);
or U13472 (N_13472,N_6656,N_6979);
and U13473 (N_13473,N_7599,N_5836);
and U13474 (N_13474,N_5727,N_6143);
xor U13475 (N_13475,N_5570,N_8741);
nand U13476 (N_13476,N_9013,N_5743);
nand U13477 (N_13477,N_7188,N_8199);
nand U13478 (N_13478,N_6292,N_5673);
nor U13479 (N_13479,N_7356,N_5300);
or U13480 (N_13480,N_9210,N_8399);
nor U13481 (N_13481,N_8456,N_9813);
or U13482 (N_13482,N_8050,N_8234);
nand U13483 (N_13483,N_8558,N_9610);
nor U13484 (N_13484,N_5764,N_6287);
nand U13485 (N_13485,N_7024,N_6247);
nor U13486 (N_13486,N_6077,N_5917);
xor U13487 (N_13487,N_7249,N_9179);
nor U13488 (N_13488,N_7013,N_9638);
nand U13489 (N_13489,N_9738,N_5221);
and U13490 (N_13490,N_8341,N_5104);
and U13491 (N_13491,N_6997,N_7745);
nor U13492 (N_13492,N_6592,N_8781);
or U13493 (N_13493,N_6019,N_6555);
or U13494 (N_13494,N_6742,N_9860);
nor U13495 (N_13495,N_6529,N_8843);
or U13496 (N_13496,N_6062,N_9194);
or U13497 (N_13497,N_7082,N_9087);
nor U13498 (N_13498,N_7046,N_9950);
or U13499 (N_13499,N_9300,N_5965);
nand U13500 (N_13500,N_8159,N_8030);
nand U13501 (N_13501,N_8725,N_6502);
and U13502 (N_13502,N_6185,N_7070);
xnor U13503 (N_13503,N_8473,N_5954);
and U13504 (N_13504,N_7755,N_8378);
nor U13505 (N_13505,N_9999,N_8585);
nor U13506 (N_13506,N_7806,N_8750);
nand U13507 (N_13507,N_5475,N_7028);
xnor U13508 (N_13508,N_9145,N_6473);
nand U13509 (N_13509,N_5096,N_9900);
nand U13510 (N_13510,N_9654,N_8227);
or U13511 (N_13511,N_9054,N_7081);
nand U13512 (N_13512,N_8429,N_5694);
or U13513 (N_13513,N_9007,N_9900);
xnor U13514 (N_13514,N_7600,N_8775);
nor U13515 (N_13515,N_8886,N_8925);
nor U13516 (N_13516,N_7137,N_9805);
nand U13517 (N_13517,N_8580,N_7070);
nand U13518 (N_13518,N_5279,N_7917);
nor U13519 (N_13519,N_6717,N_5891);
or U13520 (N_13520,N_6913,N_9464);
nand U13521 (N_13521,N_9038,N_6163);
nand U13522 (N_13522,N_5182,N_8469);
and U13523 (N_13523,N_7656,N_5435);
and U13524 (N_13524,N_5459,N_7090);
nand U13525 (N_13525,N_6577,N_9673);
or U13526 (N_13526,N_6844,N_9039);
or U13527 (N_13527,N_7634,N_5610);
and U13528 (N_13528,N_9346,N_7224);
nor U13529 (N_13529,N_7960,N_6929);
nor U13530 (N_13530,N_5561,N_8747);
or U13531 (N_13531,N_9844,N_5910);
or U13532 (N_13532,N_7711,N_7311);
nand U13533 (N_13533,N_9836,N_5187);
nand U13534 (N_13534,N_6763,N_6467);
or U13535 (N_13535,N_9664,N_7787);
nand U13536 (N_13536,N_9382,N_6894);
nor U13537 (N_13537,N_6006,N_8460);
xnor U13538 (N_13538,N_6913,N_5512);
xnor U13539 (N_13539,N_7045,N_9340);
xnor U13540 (N_13540,N_8860,N_5605);
or U13541 (N_13541,N_7564,N_6023);
and U13542 (N_13542,N_8962,N_9170);
or U13543 (N_13543,N_7803,N_5491);
nand U13544 (N_13544,N_9214,N_5983);
nand U13545 (N_13545,N_6320,N_6269);
or U13546 (N_13546,N_6701,N_9221);
nor U13547 (N_13547,N_7947,N_6342);
nand U13548 (N_13548,N_8367,N_5444);
xor U13549 (N_13549,N_9383,N_7037);
or U13550 (N_13550,N_9062,N_5375);
or U13551 (N_13551,N_6141,N_6980);
or U13552 (N_13552,N_5764,N_6945);
nand U13553 (N_13553,N_7876,N_5642);
nor U13554 (N_13554,N_5691,N_9173);
nor U13555 (N_13555,N_9975,N_5778);
xor U13556 (N_13556,N_6034,N_6629);
nor U13557 (N_13557,N_6364,N_5490);
or U13558 (N_13558,N_8866,N_5422);
nor U13559 (N_13559,N_9079,N_9356);
and U13560 (N_13560,N_6794,N_6879);
xor U13561 (N_13561,N_8597,N_6586);
nand U13562 (N_13562,N_7585,N_5688);
nor U13563 (N_13563,N_9542,N_7065);
nor U13564 (N_13564,N_9612,N_6131);
or U13565 (N_13565,N_5982,N_5477);
and U13566 (N_13566,N_6460,N_9301);
and U13567 (N_13567,N_6099,N_6849);
and U13568 (N_13568,N_7706,N_6972);
or U13569 (N_13569,N_7774,N_8524);
nand U13570 (N_13570,N_9203,N_6608);
or U13571 (N_13571,N_5407,N_5108);
nor U13572 (N_13572,N_8171,N_6709);
or U13573 (N_13573,N_7495,N_9244);
or U13574 (N_13574,N_8304,N_8510);
or U13575 (N_13575,N_5005,N_7178);
nand U13576 (N_13576,N_9452,N_9524);
nand U13577 (N_13577,N_7164,N_9840);
and U13578 (N_13578,N_8583,N_6674);
nor U13579 (N_13579,N_5751,N_7817);
nor U13580 (N_13580,N_8123,N_9981);
or U13581 (N_13581,N_8486,N_5148);
nand U13582 (N_13582,N_5524,N_8798);
nor U13583 (N_13583,N_7099,N_9557);
or U13584 (N_13584,N_5869,N_7119);
or U13585 (N_13585,N_7914,N_9363);
or U13586 (N_13586,N_7912,N_8738);
nand U13587 (N_13587,N_8081,N_8349);
nor U13588 (N_13588,N_6257,N_8384);
and U13589 (N_13589,N_6982,N_7995);
xnor U13590 (N_13590,N_8922,N_5510);
or U13591 (N_13591,N_8758,N_7280);
or U13592 (N_13592,N_5053,N_8115);
nand U13593 (N_13593,N_6995,N_6713);
or U13594 (N_13594,N_9631,N_5229);
and U13595 (N_13595,N_7445,N_9551);
nand U13596 (N_13596,N_7130,N_7700);
xnor U13597 (N_13597,N_9301,N_9912);
or U13598 (N_13598,N_7939,N_6099);
or U13599 (N_13599,N_8945,N_5954);
and U13600 (N_13600,N_6594,N_5463);
nand U13601 (N_13601,N_5592,N_5945);
nor U13602 (N_13602,N_7431,N_5511);
or U13603 (N_13603,N_6870,N_9105);
or U13604 (N_13604,N_9546,N_8956);
nor U13605 (N_13605,N_5874,N_6179);
and U13606 (N_13606,N_6871,N_5349);
nor U13607 (N_13607,N_6206,N_5052);
nand U13608 (N_13608,N_6691,N_6369);
nor U13609 (N_13609,N_5947,N_8460);
and U13610 (N_13610,N_8116,N_8410);
or U13611 (N_13611,N_9243,N_5615);
xor U13612 (N_13612,N_8034,N_6194);
nor U13613 (N_13613,N_5229,N_7744);
or U13614 (N_13614,N_8822,N_9274);
nand U13615 (N_13615,N_8629,N_6458);
nor U13616 (N_13616,N_9695,N_7281);
and U13617 (N_13617,N_6994,N_5488);
or U13618 (N_13618,N_6906,N_9587);
nor U13619 (N_13619,N_9206,N_5442);
nand U13620 (N_13620,N_8349,N_6620);
or U13621 (N_13621,N_8902,N_7728);
or U13622 (N_13622,N_8402,N_6064);
nor U13623 (N_13623,N_6415,N_8524);
nand U13624 (N_13624,N_7457,N_8162);
nor U13625 (N_13625,N_5755,N_5956);
nand U13626 (N_13626,N_8102,N_8877);
nand U13627 (N_13627,N_8538,N_6699);
nand U13628 (N_13628,N_9686,N_7355);
xnor U13629 (N_13629,N_5568,N_9667);
nand U13630 (N_13630,N_5533,N_6438);
and U13631 (N_13631,N_7567,N_7627);
or U13632 (N_13632,N_8530,N_6668);
nor U13633 (N_13633,N_9257,N_9199);
or U13634 (N_13634,N_8521,N_8528);
nor U13635 (N_13635,N_7533,N_7324);
nand U13636 (N_13636,N_7127,N_5500);
or U13637 (N_13637,N_5268,N_8006);
and U13638 (N_13638,N_7094,N_5120);
nand U13639 (N_13639,N_7845,N_8136);
nand U13640 (N_13640,N_9028,N_8095);
and U13641 (N_13641,N_9893,N_9593);
or U13642 (N_13642,N_8059,N_7651);
xor U13643 (N_13643,N_5009,N_9456);
or U13644 (N_13644,N_5655,N_6658);
and U13645 (N_13645,N_6520,N_8610);
and U13646 (N_13646,N_5074,N_7630);
or U13647 (N_13647,N_9353,N_5267);
or U13648 (N_13648,N_5846,N_6231);
or U13649 (N_13649,N_8520,N_5075);
or U13650 (N_13650,N_5921,N_6265);
and U13651 (N_13651,N_9901,N_6421);
nor U13652 (N_13652,N_6495,N_8783);
or U13653 (N_13653,N_9726,N_8154);
and U13654 (N_13654,N_7321,N_5650);
nor U13655 (N_13655,N_9367,N_5938);
xnor U13656 (N_13656,N_5657,N_6240);
nand U13657 (N_13657,N_6446,N_9488);
xnor U13658 (N_13658,N_5600,N_8771);
or U13659 (N_13659,N_8079,N_5935);
nor U13660 (N_13660,N_5495,N_9186);
nor U13661 (N_13661,N_9017,N_9686);
xnor U13662 (N_13662,N_5808,N_9704);
or U13663 (N_13663,N_7798,N_5064);
nand U13664 (N_13664,N_5803,N_8785);
nand U13665 (N_13665,N_6551,N_7800);
xor U13666 (N_13666,N_9974,N_6205);
and U13667 (N_13667,N_8693,N_7217);
or U13668 (N_13668,N_8564,N_8231);
nor U13669 (N_13669,N_8754,N_7774);
nand U13670 (N_13670,N_5534,N_7682);
nor U13671 (N_13671,N_7098,N_9488);
nand U13672 (N_13672,N_8697,N_6128);
and U13673 (N_13673,N_8738,N_9363);
and U13674 (N_13674,N_6404,N_6707);
and U13675 (N_13675,N_7237,N_8027);
and U13676 (N_13676,N_5276,N_8279);
or U13677 (N_13677,N_8410,N_9651);
nor U13678 (N_13678,N_5857,N_8445);
xor U13679 (N_13679,N_8530,N_8069);
or U13680 (N_13680,N_8275,N_9223);
nor U13681 (N_13681,N_5167,N_7955);
and U13682 (N_13682,N_5743,N_6787);
nor U13683 (N_13683,N_6066,N_7402);
and U13684 (N_13684,N_8842,N_8701);
or U13685 (N_13685,N_5762,N_9530);
and U13686 (N_13686,N_7302,N_7079);
nand U13687 (N_13687,N_5785,N_5858);
and U13688 (N_13688,N_6363,N_9130);
or U13689 (N_13689,N_7412,N_7567);
or U13690 (N_13690,N_5032,N_8715);
and U13691 (N_13691,N_7611,N_5431);
or U13692 (N_13692,N_5966,N_6033);
nand U13693 (N_13693,N_7778,N_6899);
xnor U13694 (N_13694,N_6329,N_9110);
or U13695 (N_13695,N_5199,N_6613);
xnor U13696 (N_13696,N_5946,N_9330);
nor U13697 (N_13697,N_5897,N_7952);
nor U13698 (N_13698,N_9497,N_8929);
and U13699 (N_13699,N_5414,N_5157);
nor U13700 (N_13700,N_8341,N_5086);
nand U13701 (N_13701,N_5330,N_5226);
nand U13702 (N_13702,N_6065,N_5996);
nor U13703 (N_13703,N_8923,N_9366);
or U13704 (N_13704,N_9637,N_6620);
nand U13705 (N_13705,N_5336,N_8934);
and U13706 (N_13706,N_6508,N_5272);
nor U13707 (N_13707,N_8668,N_6266);
and U13708 (N_13708,N_5629,N_7627);
or U13709 (N_13709,N_6199,N_5616);
or U13710 (N_13710,N_7452,N_6123);
nand U13711 (N_13711,N_5516,N_9746);
nand U13712 (N_13712,N_8877,N_8272);
nand U13713 (N_13713,N_7473,N_6587);
or U13714 (N_13714,N_7127,N_8641);
or U13715 (N_13715,N_5794,N_6103);
xnor U13716 (N_13716,N_8256,N_8486);
nand U13717 (N_13717,N_8453,N_6212);
or U13718 (N_13718,N_5644,N_5590);
and U13719 (N_13719,N_6010,N_9203);
or U13720 (N_13720,N_7299,N_5201);
xnor U13721 (N_13721,N_6542,N_8806);
and U13722 (N_13722,N_6008,N_8112);
nor U13723 (N_13723,N_7460,N_5772);
and U13724 (N_13724,N_7849,N_8280);
nand U13725 (N_13725,N_6878,N_8544);
nor U13726 (N_13726,N_8156,N_8215);
nor U13727 (N_13727,N_8707,N_8117);
and U13728 (N_13728,N_8924,N_9293);
nor U13729 (N_13729,N_9487,N_7842);
or U13730 (N_13730,N_6263,N_5548);
and U13731 (N_13731,N_9545,N_7974);
xnor U13732 (N_13732,N_9706,N_5354);
nand U13733 (N_13733,N_9412,N_7115);
and U13734 (N_13734,N_9262,N_7736);
and U13735 (N_13735,N_9312,N_9420);
nand U13736 (N_13736,N_6164,N_9068);
nor U13737 (N_13737,N_5694,N_8389);
xor U13738 (N_13738,N_7111,N_9692);
and U13739 (N_13739,N_8257,N_8778);
and U13740 (N_13740,N_9654,N_7869);
and U13741 (N_13741,N_7928,N_6367);
or U13742 (N_13742,N_6808,N_6290);
nor U13743 (N_13743,N_5531,N_8320);
nor U13744 (N_13744,N_5957,N_7642);
nand U13745 (N_13745,N_5876,N_7194);
and U13746 (N_13746,N_6046,N_8172);
or U13747 (N_13747,N_9248,N_7509);
nand U13748 (N_13748,N_8640,N_6494);
or U13749 (N_13749,N_8021,N_8478);
xor U13750 (N_13750,N_5171,N_8985);
nor U13751 (N_13751,N_8718,N_6200);
and U13752 (N_13752,N_9907,N_6498);
xor U13753 (N_13753,N_5227,N_7380);
and U13754 (N_13754,N_5187,N_5780);
and U13755 (N_13755,N_9792,N_6761);
nand U13756 (N_13756,N_7461,N_7465);
nor U13757 (N_13757,N_8776,N_5024);
and U13758 (N_13758,N_5578,N_8114);
xor U13759 (N_13759,N_8693,N_8655);
or U13760 (N_13760,N_8798,N_8601);
and U13761 (N_13761,N_5075,N_6366);
or U13762 (N_13762,N_6338,N_7482);
or U13763 (N_13763,N_5211,N_7222);
and U13764 (N_13764,N_5828,N_7617);
xor U13765 (N_13765,N_9582,N_6421);
or U13766 (N_13766,N_5781,N_9321);
or U13767 (N_13767,N_7352,N_6541);
xnor U13768 (N_13768,N_7491,N_7365);
xnor U13769 (N_13769,N_8718,N_5981);
nor U13770 (N_13770,N_7021,N_7317);
or U13771 (N_13771,N_9714,N_7299);
nand U13772 (N_13772,N_9588,N_9124);
or U13773 (N_13773,N_9340,N_6131);
or U13774 (N_13774,N_8749,N_7296);
nand U13775 (N_13775,N_9008,N_9700);
nand U13776 (N_13776,N_9618,N_7312);
nor U13777 (N_13777,N_6493,N_6294);
or U13778 (N_13778,N_9007,N_5331);
xnor U13779 (N_13779,N_5819,N_6598);
nand U13780 (N_13780,N_9757,N_5946);
nand U13781 (N_13781,N_8604,N_8399);
nor U13782 (N_13782,N_5117,N_7335);
nor U13783 (N_13783,N_9259,N_8927);
and U13784 (N_13784,N_7238,N_7661);
and U13785 (N_13785,N_8703,N_6473);
xor U13786 (N_13786,N_6820,N_6238);
and U13787 (N_13787,N_9282,N_5932);
or U13788 (N_13788,N_6282,N_8239);
nor U13789 (N_13789,N_8372,N_8422);
and U13790 (N_13790,N_6009,N_6741);
and U13791 (N_13791,N_5156,N_8079);
or U13792 (N_13792,N_8573,N_8387);
or U13793 (N_13793,N_6662,N_6512);
and U13794 (N_13794,N_5298,N_9383);
and U13795 (N_13795,N_7733,N_6826);
and U13796 (N_13796,N_8289,N_7207);
and U13797 (N_13797,N_5883,N_7785);
and U13798 (N_13798,N_6028,N_9534);
xor U13799 (N_13799,N_6165,N_9592);
or U13800 (N_13800,N_7363,N_8062);
nor U13801 (N_13801,N_7750,N_8021);
nand U13802 (N_13802,N_7286,N_8074);
nand U13803 (N_13803,N_7422,N_9645);
xnor U13804 (N_13804,N_7232,N_8597);
nor U13805 (N_13805,N_7929,N_7974);
nand U13806 (N_13806,N_8677,N_9645);
nor U13807 (N_13807,N_6734,N_6043);
nor U13808 (N_13808,N_6512,N_9769);
nand U13809 (N_13809,N_7018,N_6877);
or U13810 (N_13810,N_6696,N_8569);
nand U13811 (N_13811,N_6977,N_8692);
nor U13812 (N_13812,N_6306,N_6041);
nor U13813 (N_13813,N_5711,N_5636);
nor U13814 (N_13814,N_7628,N_6770);
or U13815 (N_13815,N_7691,N_8690);
xnor U13816 (N_13816,N_9582,N_8135);
nand U13817 (N_13817,N_6323,N_7059);
nor U13818 (N_13818,N_7538,N_6421);
nor U13819 (N_13819,N_6115,N_6105);
nand U13820 (N_13820,N_8046,N_8634);
or U13821 (N_13821,N_8809,N_6575);
nor U13822 (N_13822,N_7875,N_6755);
nand U13823 (N_13823,N_8014,N_9331);
or U13824 (N_13824,N_7472,N_5227);
or U13825 (N_13825,N_9033,N_8840);
nor U13826 (N_13826,N_7912,N_8811);
and U13827 (N_13827,N_5846,N_7463);
nand U13828 (N_13828,N_6600,N_5979);
nor U13829 (N_13829,N_8318,N_8772);
nor U13830 (N_13830,N_6249,N_6532);
xor U13831 (N_13831,N_9234,N_8743);
nor U13832 (N_13832,N_9383,N_7338);
xor U13833 (N_13833,N_9722,N_9683);
and U13834 (N_13834,N_9611,N_9038);
or U13835 (N_13835,N_7065,N_8121);
and U13836 (N_13836,N_6926,N_9256);
or U13837 (N_13837,N_9616,N_5851);
or U13838 (N_13838,N_9779,N_8740);
nor U13839 (N_13839,N_6022,N_9110);
and U13840 (N_13840,N_5716,N_9943);
nor U13841 (N_13841,N_9898,N_8857);
or U13842 (N_13842,N_8859,N_9091);
or U13843 (N_13843,N_9539,N_6634);
nor U13844 (N_13844,N_6663,N_9696);
nor U13845 (N_13845,N_9460,N_9268);
nor U13846 (N_13846,N_7856,N_5353);
nand U13847 (N_13847,N_5221,N_9676);
and U13848 (N_13848,N_6991,N_5886);
nand U13849 (N_13849,N_9722,N_8795);
nor U13850 (N_13850,N_8222,N_7958);
xor U13851 (N_13851,N_6903,N_6345);
and U13852 (N_13852,N_8346,N_5558);
nand U13853 (N_13853,N_9407,N_9077);
nor U13854 (N_13854,N_8080,N_7059);
nor U13855 (N_13855,N_8116,N_7925);
nand U13856 (N_13856,N_9396,N_8125);
nand U13857 (N_13857,N_9121,N_6744);
xnor U13858 (N_13858,N_5473,N_9620);
and U13859 (N_13859,N_9570,N_9365);
nor U13860 (N_13860,N_5054,N_7472);
or U13861 (N_13861,N_9832,N_7664);
nor U13862 (N_13862,N_5753,N_6896);
nor U13863 (N_13863,N_9676,N_8516);
nor U13864 (N_13864,N_8358,N_7137);
nor U13865 (N_13865,N_5257,N_5371);
nor U13866 (N_13866,N_7127,N_5462);
xnor U13867 (N_13867,N_6943,N_5641);
and U13868 (N_13868,N_6003,N_9111);
nor U13869 (N_13869,N_9324,N_7573);
or U13870 (N_13870,N_5757,N_8096);
nor U13871 (N_13871,N_8479,N_5598);
nand U13872 (N_13872,N_6605,N_9314);
nor U13873 (N_13873,N_9893,N_8540);
nand U13874 (N_13874,N_9246,N_5545);
xnor U13875 (N_13875,N_5151,N_5685);
nand U13876 (N_13876,N_8224,N_7250);
or U13877 (N_13877,N_7215,N_6085);
and U13878 (N_13878,N_5802,N_7616);
nor U13879 (N_13879,N_7153,N_7526);
or U13880 (N_13880,N_6784,N_7214);
nand U13881 (N_13881,N_5904,N_7113);
and U13882 (N_13882,N_7574,N_9095);
nor U13883 (N_13883,N_8934,N_6657);
nand U13884 (N_13884,N_9490,N_6413);
xnor U13885 (N_13885,N_6607,N_6943);
and U13886 (N_13886,N_8214,N_7313);
nor U13887 (N_13887,N_5880,N_6362);
nand U13888 (N_13888,N_6650,N_7710);
nand U13889 (N_13889,N_5763,N_7931);
or U13890 (N_13890,N_9057,N_6896);
and U13891 (N_13891,N_7588,N_8303);
and U13892 (N_13892,N_9972,N_8931);
nor U13893 (N_13893,N_8502,N_8524);
or U13894 (N_13894,N_5085,N_6272);
xor U13895 (N_13895,N_5024,N_9946);
or U13896 (N_13896,N_7842,N_9461);
and U13897 (N_13897,N_9557,N_9617);
or U13898 (N_13898,N_7891,N_5072);
nor U13899 (N_13899,N_6685,N_5066);
and U13900 (N_13900,N_6032,N_7378);
and U13901 (N_13901,N_7554,N_5500);
nand U13902 (N_13902,N_5926,N_8479);
xor U13903 (N_13903,N_5062,N_5811);
and U13904 (N_13904,N_9982,N_8307);
and U13905 (N_13905,N_8919,N_9190);
nand U13906 (N_13906,N_6036,N_6258);
or U13907 (N_13907,N_9029,N_5684);
nand U13908 (N_13908,N_7252,N_7586);
nand U13909 (N_13909,N_5752,N_6640);
nor U13910 (N_13910,N_5181,N_7790);
or U13911 (N_13911,N_6132,N_5154);
nor U13912 (N_13912,N_6042,N_8103);
and U13913 (N_13913,N_9935,N_8282);
nand U13914 (N_13914,N_6228,N_7857);
nand U13915 (N_13915,N_5473,N_9042);
or U13916 (N_13916,N_8413,N_8959);
nand U13917 (N_13917,N_6066,N_8579);
and U13918 (N_13918,N_7097,N_6815);
or U13919 (N_13919,N_5468,N_5340);
nor U13920 (N_13920,N_6995,N_5909);
and U13921 (N_13921,N_5316,N_9910);
nand U13922 (N_13922,N_5388,N_5978);
nor U13923 (N_13923,N_9584,N_5588);
and U13924 (N_13924,N_7550,N_9459);
or U13925 (N_13925,N_8346,N_7959);
nor U13926 (N_13926,N_6496,N_8190);
nand U13927 (N_13927,N_8352,N_8217);
nor U13928 (N_13928,N_9495,N_9970);
xnor U13929 (N_13929,N_5730,N_6369);
and U13930 (N_13930,N_9765,N_9787);
or U13931 (N_13931,N_8073,N_6995);
nand U13932 (N_13932,N_5743,N_5367);
nand U13933 (N_13933,N_5880,N_8023);
or U13934 (N_13934,N_6848,N_9717);
nand U13935 (N_13935,N_8864,N_7997);
or U13936 (N_13936,N_6685,N_5156);
nor U13937 (N_13937,N_6350,N_5306);
nor U13938 (N_13938,N_7307,N_6547);
nand U13939 (N_13939,N_8424,N_7001);
nand U13940 (N_13940,N_7729,N_9548);
xnor U13941 (N_13941,N_6282,N_5402);
or U13942 (N_13942,N_5606,N_7875);
and U13943 (N_13943,N_5754,N_5390);
nor U13944 (N_13944,N_9256,N_9772);
xor U13945 (N_13945,N_7671,N_9925);
nor U13946 (N_13946,N_7815,N_5929);
nor U13947 (N_13947,N_7441,N_9546);
nor U13948 (N_13948,N_8445,N_7741);
and U13949 (N_13949,N_7167,N_7520);
nand U13950 (N_13950,N_9293,N_7282);
and U13951 (N_13951,N_6836,N_9125);
or U13952 (N_13952,N_9167,N_8857);
nor U13953 (N_13953,N_7375,N_9368);
xor U13954 (N_13954,N_9006,N_6325);
nor U13955 (N_13955,N_6739,N_9172);
or U13956 (N_13956,N_8158,N_6833);
xnor U13957 (N_13957,N_9840,N_6576);
and U13958 (N_13958,N_8532,N_6286);
xor U13959 (N_13959,N_5620,N_8509);
nor U13960 (N_13960,N_6589,N_6676);
nor U13961 (N_13961,N_9939,N_8904);
nor U13962 (N_13962,N_8377,N_5894);
and U13963 (N_13963,N_9699,N_7879);
nor U13964 (N_13964,N_8076,N_7110);
or U13965 (N_13965,N_9425,N_9363);
nor U13966 (N_13966,N_6826,N_5722);
xnor U13967 (N_13967,N_9151,N_5457);
nand U13968 (N_13968,N_5477,N_9097);
and U13969 (N_13969,N_9910,N_5382);
nand U13970 (N_13970,N_8267,N_8952);
and U13971 (N_13971,N_8571,N_9247);
or U13972 (N_13972,N_8761,N_6124);
and U13973 (N_13973,N_6530,N_9716);
or U13974 (N_13974,N_6925,N_7474);
nand U13975 (N_13975,N_5057,N_8305);
nand U13976 (N_13976,N_9127,N_5615);
nand U13977 (N_13977,N_7220,N_5740);
and U13978 (N_13978,N_5451,N_5318);
nor U13979 (N_13979,N_9846,N_7572);
nand U13980 (N_13980,N_5107,N_5088);
or U13981 (N_13981,N_8771,N_9651);
or U13982 (N_13982,N_6880,N_6495);
nor U13983 (N_13983,N_5686,N_8372);
and U13984 (N_13984,N_6264,N_5651);
and U13985 (N_13985,N_9329,N_5500);
nor U13986 (N_13986,N_5975,N_6262);
nor U13987 (N_13987,N_6178,N_9531);
nor U13988 (N_13988,N_8894,N_6209);
and U13989 (N_13989,N_5895,N_7517);
xnor U13990 (N_13990,N_7736,N_8938);
nand U13991 (N_13991,N_6135,N_9737);
and U13992 (N_13992,N_5147,N_8439);
or U13993 (N_13993,N_8106,N_5319);
nand U13994 (N_13994,N_5543,N_7294);
nand U13995 (N_13995,N_9823,N_9528);
or U13996 (N_13996,N_6052,N_8434);
nand U13997 (N_13997,N_6151,N_7686);
nor U13998 (N_13998,N_6006,N_7405);
or U13999 (N_13999,N_8650,N_6204);
nor U14000 (N_14000,N_5136,N_9757);
or U14001 (N_14001,N_6389,N_7861);
or U14002 (N_14002,N_8346,N_7119);
nor U14003 (N_14003,N_7737,N_6567);
or U14004 (N_14004,N_7329,N_7309);
and U14005 (N_14005,N_8338,N_8334);
nand U14006 (N_14006,N_7090,N_6576);
or U14007 (N_14007,N_5481,N_8876);
and U14008 (N_14008,N_6796,N_9085);
nor U14009 (N_14009,N_9222,N_5491);
and U14010 (N_14010,N_5484,N_8135);
xnor U14011 (N_14011,N_8263,N_6551);
nand U14012 (N_14012,N_7102,N_9926);
or U14013 (N_14013,N_7840,N_9142);
and U14014 (N_14014,N_8361,N_8448);
or U14015 (N_14015,N_7802,N_9853);
and U14016 (N_14016,N_6237,N_9877);
and U14017 (N_14017,N_6208,N_6951);
and U14018 (N_14018,N_9984,N_8021);
and U14019 (N_14019,N_8688,N_6524);
nor U14020 (N_14020,N_7577,N_9142);
and U14021 (N_14021,N_7254,N_5386);
and U14022 (N_14022,N_9317,N_5912);
xor U14023 (N_14023,N_8994,N_8134);
nand U14024 (N_14024,N_9412,N_9383);
nor U14025 (N_14025,N_7174,N_7475);
or U14026 (N_14026,N_7197,N_7400);
xor U14027 (N_14027,N_5894,N_6636);
nand U14028 (N_14028,N_8551,N_5112);
and U14029 (N_14029,N_6194,N_7074);
and U14030 (N_14030,N_8402,N_7842);
nor U14031 (N_14031,N_6658,N_6185);
or U14032 (N_14032,N_5851,N_9019);
or U14033 (N_14033,N_6306,N_7206);
nor U14034 (N_14034,N_5801,N_9482);
nand U14035 (N_14035,N_5660,N_5439);
and U14036 (N_14036,N_5909,N_5777);
nand U14037 (N_14037,N_9879,N_9490);
or U14038 (N_14038,N_5865,N_8268);
nand U14039 (N_14039,N_8962,N_7602);
or U14040 (N_14040,N_9620,N_9707);
and U14041 (N_14041,N_8723,N_5309);
xor U14042 (N_14042,N_5379,N_7595);
or U14043 (N_14043,N_7486,N_9436);
and U14044 (N_14044,N_7389,N_5704);
nand U14045 (N_14045,N_8697,N_6436);
nand U14046 (N_14046,N_7945,N_6583);
and U14047 (N_14047,N_7118,N_9286);
xnor U14048 (N_14048,N_5662,N_6714);
or U14049 (N_14049,N_9939,N_9544);
nor U14050 (N_14050,N_8447,N_7619);
and U14051 (N_14051,N_5647,N_9527);
nand U14052 (N_14052,N_5197,N_5495);
nor U14053 (N_14053,N_9929,N_9582);
and U14054 (N_14054,N_9260,N_6060);
nand U14055 (N_14055,N_5135,N_8844);
and U14056 (N_14056,N_7331,N_5956);
or U14057 (N_14057,N_6050,N_5834);
and U14058 (N_14058,N_5462,N_5763);
and U14059 (N_14059,N_9055,N_7168);
nor U14060 (N_14060,N_7625,N_6011);
and U14061 (N_14061,N_9493,N_6006);
or U14062 (N_14062,N_8245,N_7693);
nor U14063 (N_14063,N_9962,N_7051);
nand U14064 (N_14064,N_7060,N_9675);
and U14065 (N_14065,N_7029,N_8245);
nand U14066 (N_14066,N_7444,N_8456);
nand U14067 (N_14067,N_7778,N_9381);
nand U14068 (N_14068,N_8228,N_6295);
nor U14069 (N_14069,N_6144,N_5618);
and U14070 (N_14070,N_6618,N_7200);
nor U14071 (N_14071,N_6255,N_9821);
or U14072 (N_14072,N_6347,N_5488);
nand U14073 (N_14073,N_5906,N_6401);
nor U14074 (N_14074,N_9085,N_8827);
and U14075 (N_14075,N_9476,N_7792);
nand U14076 (N_14076,N_7762,N_7943);
nand U14077 (N_14077,N_9311,N_7364);
and U14078 (N_14078,N_5108,N_6924);
or U14079 (N_14079,N_9981,N_6312);
or U14080 (N_14080,N_9481,N_5158);
nand U14081 (N_14081,N_8457,N_5698);
nand U14082 (N_14082,N_8504,N_8952);
or U14083 (N_14083,N_7966,N_7271);
nand U14084 (N_14084,N_7123,N_6947);
or U14085 (N_14085,N_7100,N_9303);
nor U14086 (N_14086,N_5397,N_6189);
nor U14087 (N_14087,N_5270,N_8050);
nor U14088 (N_14088,N_9011,N_9261);
and U14089 (N_14089,N_8880,N_7609);
and U14090 (N_14090,N_5674,N_9050);
nand U14091 (N_14091,N_9891,N_5046);
xnor U14092 (N_14092,N_7481,N_8058);
xnor U14093 (N_14093,N_8915,N_5090);
nor U14094 (N_14094,N_5857,N_8357);
nor U14095 (N_14095,N_9231,N_5663);
and U14096 (N_14096,N_7500,N_7005);
nor U14097 (N_14097,N_6688,N_8104);
or U14098 (N_14098,N_5405,N_8637);
nand U14099 (N_14099,N_9586,N_5448);
nor U14100 (N_14100,N_5845,N_7405);
nor U14101 (N_14101,N_6897,N_6622);
nand U14102 (N_14102,N_5913,N_7113);
nor U14103 (N_14103,N_5873,N_5402);
nor U14104 (N_14104,N_9756,N_6780);
nor U14105 (N_14105,N_6118,N_9809);
or U14106 (N_14106,N_8617,N_9752);
nand U14107 (N_14107,N_5070,N_8498);
nor U14108 (N_14108,N_5936,N_9352);
nand U14109 (N_14109,N_5668,N_6625);
xnor U14110 (N_14110,N_6899,N_7393);
nand U14111 (N_14111,N_6164,N_8406);
nor U14112 (N_14112,N_8375,N_6423);
or U14113 (N_14113,N_6202,N_6614);
or U14114 (N_14114,N_8670,N_6924);
or U14115 (N_14115,N_5562,N_7564);
xor U14116 (N_14116,N_9885,N_5731);
nand U14117 (N_14117,N_7107,N_6068);
and U14118 (N_14118,N_8544,N_8992);
nand U14119 (N_14119,N_8214,N_8155);
nor U14120 (N_14120,N_9516,N_6141);
nand U14121 (N_14121,N_6405,N_7120);
and U14122 (N_14122,N_7588,N_7420);
nor U14123 (N_14123,N_9366,N_7563);
and U14124 (N_14124,N_7390,N_9557);
nand U14125 (N_14125,N_8744,N_6829);
or U14126 (N_14126,N_7642,N_7004);
nand U14127 (N_14127,N_8506,N_5225);
or U14128 (N_14128,N_7783,N_8329);
and U14129 (N_14129,N_6908,N_6989);
nor U14130 (N_14130,N_7988,N_9050);
and U14131 (N_14131,N_6087,N_5841);
nand U14132 (N_14132,N_6957,N_5432);
nor U14133 (N_14133,N_8602,N_6876);
nand U14134 (N_14134,N_7971,N_6808);
xor U14135 (N_14135,N_8292,N_8447);
or U14136 (N_14136,N_6815,N_5434);
nand U14137 (N_14137,N_8571,N_6044);
nand U14138 (N_14138,N_7174,N_7613);
and U14139 (N_14139,N_8086,N_9013);
nor U14140 (N_14140,N_5795,N_5509);
and U14141 (N_14141,N_9422,N_8979);
and U14142 (N_14142,N_6389,N_9973);
or U14143 (N_14143,N_8154,N_8745);
nor U14144 (N_14144,N_9608,N_8270);
xnor U14145 (N_14145,N_6937,N_9593);
and U14146 (N_14146,N_8733,N_8050);
or U14147 (N_14147,N_8278,N_7195);
nor U14148 (N_14148,N_7513,N_5200);
or U14149 (N_14149,N_5787,N_5554);
or U14150 (N_14150,N_8356,N_5613);
or U14151 (N_14151,N_8283,N_8529);
and U14152 (N_14152,N_7691,N_7870);
nor U14153 (N_14153,N_5674,N_7051);
nand U14154 (N_14154,N_6023,N_8915);
or U14155 (N_14155,N_7878,N_5078);
or U14156 (N_14156,N_5669,N_8136);
nand U14157 (N_14157,N_7790,N_6577);
nand U14158 (N_14158,N_5944,N_8139);
nand U14159 (N_14159,N_9657,N_5074);
or U14160 (N_14160,N_6303,N_5476);
nand U14161 (N_14161,N_9935,N_8604);
xnor U14162 (N_14162,N_7004,N_9619);
nand U14163 (N_14163,N_7151,N_9804);
nor U14164 (N_14164,N_7521,N_5668);
or U14165 (N_14165,N_7824,N_8338);
or U14166 (N_14166,N_7318,N_7001);
or U14167 (N_14167,N_9806,N_7330);
and U14168 (N_14168,N_8209,N_8228);
or U14169 (N_14169,N_5353,N_7732);
or U14170 (N_14170,N_6170,N_6708);
nor U14171 (N_14171,N_5891,N_5194);
nor U14172 (N_14172,N_5937,N_6784);
nand U14173 (N_14173,N_8631,N_7506);
nor U14174 (N_14174,N_9287,N_6310);
or U14175 (N_14175,N_8633,N_7381);
or U14176 (N_14176,N_7593,N_9317);
nand U14177 (N_14177,N_8154,N_7385);
nor U14178 (N_14178,N_9193,N_9668);
and U14179 (N_14179,N_6428,N_8272);
and U14180 (N_14180,N_6128,N_8841);
and U14181 (N_14181,N_8812,N_8374);
or U14182 (N_14182,N_9549,N_6219);
or U14183 (N_14183,N_9036,N_9590);
and U14184 (N_14184,N_5374,N_9064);
nand U14185 (N_14185,N_7785,N_5418);
nand U14186 (N_14186,N_7083,N_6595);
nand U14187 (N_14187,N_8483,N_6245);
nand U14188 (N_14188,N_7465,N_6604);
and U14189 (N_14189,N_7523,N_6638);
nand U14190 (N_14190,N_5459,N_7410);
and U14191 (N_14191,N_8058,N_8221);
xnor U14192 (N_14192,N_9176,N_6139);
nor U14193 (N_14193,N_5210,N_7890);
nor U14194 (N_14194,N_5615,N_6067);
nand U14195 (N_14195,N_7212,N_5105);
xnor U14196 (N_14196,N_9637,N_5962);
nor U14197 (N_14197,N_7123,N_8786);
nand U14198 (N_14198,N_7815,N_7004);
nor U14199 (N_14199,N_8043,N_9695);
or U14200 (N_14200,N_7638,N_8289);
nand U14201 (N_14201,N_8915,N_6942);
nor U14202 (N_14202,N_7484,N_8988);
nand U14203 (N_14203,N_6001,N_7343);
nor U14204 (N_14204,N_7513,N_7540);
nor U14205 (N_14205,N_7439,N_7537);
xnor U14206 (N_14206,N_7556,N_7014);
nor U14207 (N_14207,N_6526,N_8613);
nand U14208 (N_14208,N_5252,N_9562);
nand U14209 (N_14209,N_9271,N_8472);
or U14210 (N_14210,N_6516,N_7102);
and U14211 (N_14211,N_6215,N_9208);
or U14212 (N_14212,N_7328,N_7729);
xor U14213 (N_14213,N_8745,N_6778);
nor U14214 (N_14214,N_6779,N_9369);
and U14215 (N_14215,N_5301,N_9087);
xor U14216 (N_14216,N_7841,N_7847);
or U14217 (N_14217,N_9573,N_9437);
nor U14218 (N_14218,N_9169,N_5653);
and U14219 (N_14219,N_5888,N_6724);
and U14220 (N_14220,N_7788,N_9892);
and U14221 (N_14221,N_6802,N_8681);
nand U14222 (N_14222,N_8720,N_5662);
or U14223 (N_14223,N_7492,N_6714);
nor U14224 (N_14224,N_6866,N_9636);
nand U14225 (N_14225,N_9407,N_5444);
nand U14226 (N_14226,N_8631,N_9039);
nand U14227 (N_14227,N_9623,N_9665);
xnor U14228 (N_14228,N_9257,N_9697);
and U14229 (N_14229,N_7082,N_6625);
nor U14230 (N_14230,N_9431,N_6315);
or U14231 (N_14231,N_7426,N_7796);
nor U14232 (N_14232,N_8866,N_9154);
nor U14233 (N_14233,N_8901,N_5595);
nor U14234 (N_14234,N_6288,N_6171);
or U14235 (N_14235,N_8641,N_7834);
nor U14236 (N_14236,N_9770,N_9919);
or U14237 (N_14237,N_9418,N_9976);
nor U14238 (N_14238,N_5503,N_5562);
nor U14239 (N_14239,N_5304,N_8489);
and U14240 (N_14240,N_7400,N_9578);
or U14241 (N_14241,N_6414,N_9107);
nor U14242 (N_14242,N_7127,N_8396);
and U14243 (N_14243,N_6750,N_6120);
nor U14244 (N_14244,N_6466,N_9301);
and U14245 (N_14245,N_9290,N_6888);
nor U14246 (N_14246,N_5036,N_5060);
xnor U14247 (N_14247,N_7115,N_8205);
nand U14248 (N_14248,N_8129,N_6992);
or U14249 (N_14249,N_5688,N_6305);
nor U14250 (N_14250,N_7683,N_6215);
and U14251 (N_14251,N_6071,N_9734);
nor U14252 (N_14252,N_6125,N_9895);
nor U14253 (N_14253,N_5679,N_7524);
nand U14254 (N_14254,N_5435,N_8628);
and U14255 (N_14255,N_6045,N_5509);
nand U14256 (N_14256,N_5681,N_6071);
or U14257 (N_14257,N_7377,N_9091);
and U14258 (N_14258,N_7895,N_9225);
and U14259 (N_14259,N_5354,N_7977);
and U14260 (N_14260,N_6311,N_9052);
nor U14261 (N_14261,N_9020,N_8612);
and U14262 (N_14262,N_8261,N_7914);
nand U14263 (N_14263,N_5581,N_5703);
xor U14264 (N_14264,N_8212,N_7090);
xor U14265 (N_14265,N_9068,N_5732);
nand U14266 (N_14266,N_9921,N_6452);
and U14267 (N_14267,N_7625,N_5871);
and U14268 (N_14268,N_5733,N_7945);
nand U14269 (N_14269,N_7360,N_9002);
xnor U14270 (N_14270,N_6191,N_6481);
and U14271 (N_14271,N_7747,N_5404);
xor U14272 (N_14272,N_7606,N_7248);
or U14273 (N_14273,N_7859,N_7423);
nand U14274 (N_14274,N_9955,N_9825);
xor U14275 (N_14275,N_7720,N_9015);
nor U14276 (N_14276,N_5985,N_5681);
nor U14277 (N_14277,N_6809,N_8170);
or U14278 (N_14278,N_7487,N_5812);
or U14279 (N_14279,N_7086,N_9401);
or U14280 (N_14280,N_5552,N_5650);
or U14281 (N_14281,N_5472,N_7251);
or U14282 (N_14282,N_5042,N_5643);
nor U14283 (N_14283,N_7194,N_6894);
and U14284 (N_14284,N_8068,N_8647);
nor U14285 (N_14285,N_5796,N_5992);
and U14286 (N_14286,N_5588,N_8636);
xor U14287 (N_14287,N_7959,N_7841);
xor U14288 (N_14288,N_5086,N_5635);
xor U14289 (N_14289,N_6520,N_9082);
or U14290 (N_14290,N_8293,N_9227);
and U14291 (N_14291,N_5842,N_7676);
and U14292 (N_14292,N_9103,N_8601);
or U14293 (N_14293,N_7356,N_7093);
or U14294 (N_14294,N_7034,N_5900);
nand U14295 (N_14295,N_9323,N_6314);
and U14296 (N_14296,N_6720,N_7444);
or U14297 (N_14297,N_7320,N_8618);
and U14298 (N_14298,N_6025,N_8982);
xnor U14299 (N_14299,N_5060,N_6310);
nor U14300 (N_14300,N_5248,N_9397);
and U14301 (N_14301,N_6715,N_5821);
or U14302 (N_14302,N_8540,N_9427);
and U14303 (N_14303,N_8671,N_8530);
or U14304 (N_14304,N_7620,N_9178);
and U14305 (N_14305,N_9670,N_9634);
and U14306 (N_14306,N_9536,N_6878);
or U14307 (N_14307,N_8279,N_9674);
or U14308 (N_14308,N_7533,N_8854);
or U14309 (N_14309,N_7797,N_8689);
nor U14310 (N_14310,N_6688,N_6315);
nor U14311 (N_14311,N_8691,N_7794);
nand U14312 (N_14312,N_6025,N_9477);
nand U14313 (N_14313,N_7746,N_9022);
and U14314 (N_14314,N_6207,N_5272);
nor U14315 (N_14315,N_7046,N_9058);
nor U14316 (N_14316,N_7447,N_8842);
nor U14317 (N_14317,N_5398,N_7221);
or U14318 (N_14318,N_9294,N_9354);
or U14319 (N_14319,N_7848,N_8242);
nor U14320 (N_14320,N_7406,N_6480);
xnor U14321 (N_14321,N_7575,N_7704);
xnor U14322 (N_14322,N_8049,N_6576);
and U14323 (N_14323,N_8248,N_8559);
nand U14324 (N_14324,N_5461,N_5285);
nand U14325 (N_14325,N_6281,N_9128);
xor U14326 (N_14326,N_5610,N_9413);
or U14327 (N_14327,N_6996,N_9127);
or U14328 (N_14328,N_5245,N_6468);
or U14329 (N_14329,N_8606,N_8475);
xor U14330 (N_14330,N_5461,N_5345);
and U14331 (N_14331,N_6911,N_8655);
nand U14332 (N_14332,N_9570,N_9755);
xor U14333 (N_14333,N_7619,N_7570);
or U14334 (N_14334,N_8111,N_6363);
nand U14335 (N_14335,N_8613,N_5564);
or U14336 (N_14336,N_5329,N_7166);
and U14337 (N_14337,N_5169,N_5565);
nor U14338 (N_14338,N_6151,N_7336);
nand U14339 (N_14339,N_6720,N_9422);
nor U14340 (N_14340,N_9919,N_5067);
and U14341 (N_14341,N_9813,N_6930);
and U14342 (N_14342,N_8607,N_5263);
nand U14343 (N_14343,N_6072,N_5506);
nand U14344 (N_14344,N_9108,N_8682);
xnor U14345 (N_14345,N_5380,N_8634);
and U14346 (N_14346,N_7050,N_6266);
nand U14347 (N_14347,N_9952,N_5172);
or U14348 (N_14348,N_9668,N_7705);
and U14349 (N_14349,N_6019,N_5477);
or U14350 (N_14350,N_6054,N_9657);
or U14351 (N_14351,N_7417,N_5357);
and U14352 (N_14352,N_6302,N_5515);
and U14353 (N_14353,N_7365,N_5765);
and U14354 (N_14354,N_5482,N_7246);
or U14355 (N_14355,N_7255,N_8712);
or U14356 (N_14356,N_6020,N_7812);
nor U14357 (N_14357,N_9910,N_7200);
and U14358 (N_14358,N_7253,N_5956);
nand U14359 (N_14359,N_9120,N_7004);
nand U14360 (N_14360,N_6273,N_6255);
nor U14361 (N_14361,N_9674,N_6083);
xor U14362 (N_14362,N_7110,N_7951);
and U14363 (N_14363,N_8663,N_9037);
nand U14364 (N_14364,N_5139,N_6943);
and U14365 (N_14365,N_8867,N_8106);
nor U14366 (N_14366,N_9369,N_6146);
or U14367 (N_14367,N_5987,N_5258);
or U14368 (N_14368,N_5527,N_9539);
nand U14369 (N_14369,N_6450,N_5721);
and U14370 (N_14370,N_7547,N_6008);
xnor U14371 (N_14371,N_7731,N_5312);
nand U14372 (N_14372,N_9922,N_7516);
or U14373 (N_14373,N_6145,N_5618);
and U14374 (N_14374,N_6296,N_5460);
nand U14375 (N_14375,N_9377,N_7272);
and U14376 (N_14376,N_7266,N_8528);
or U14377 (N_14377,N_9011,N_9935);
or U14378 (N_14378,N_5904,N_5159);
nor U14379 (N_14379,N_8001,N_6621);
nand U14380 (N_14380,N_5449,N_7634);
nor U14381 (N_14381,N_5918,N_5519);
and U14382 (N_14382,N_8796,N_6210);
or U14383 (N_14383,N_8753,N_7178);
or U14384 (N_14384,N_5590,N_8006);
xor U14385 (N_14385,N_5687,N_8342);
nor U14386 (N_14386,N_6393,N_5818);
nor U14387 (N_14387,N_8715,N_9380);
and U14388 (N_14388,N_7681,N_9701);
and U14389 (N_14389,N_5220,N_8022);
or U14390 (N_14390,N_5990,N_9812);
xnor U14391 (N_14391,N_7323,N_5842);
or U14392 (N_14392,N_9549,N_6393);
nand U14393 (N_14393,N_9172,N_6772);
and U14394 (N_14394,N_9315,N_6894);
nand U14395 (N_14395,N_5215,N_9853);
nand U14396 (N_14396,N_8948,N_9819);
and U14397 (N_14397,N_8634,N_5386);
or U14398 (N_14398,N_6657,N_7051);
or U14399 (N_14399,N_8979,N_9592);
nor U14400 (N_14400,N_8699,N_7954);
and U14401 (N_14401,N_9929,N_7477);
nor U14402 (N_14402,N_8012,N_7299);
xnor U14403 (N_14403,N_5565,N_8295);
xnor U14404 (N_14404,N_6970,N_7924);
nor U14405 (N_14405,N_9663,N_6331);
xnor U14406 (N_14406,N_7758,N_5484);
nor U14407 (N_14407,N_7201,N_8037);
nand U14408 (N_14408,N_5099,N_7253);
nor U14409 (N_14409,N_8441,N_9827);
or U14410 (N_14410,N_9640,N_6447);
or U14411 (N_14411,N_8064,N_7217);
nand U14412 (N_14412,N_9962,N_8004);
xnor U14413 (N_14413,N_6416,N_5618);
or U14414 (N_14414,N_9217,N_9042);
and U14415 (N_14415,N_6737,N_9985);
nor U14416 (N_14416,N_9099,N_6437);
or U14417 (N_14417,N_7049,N_9814);
and U14418 (N_14418,N_5035,N_8158);
xor U14419 (N_14419,N_7625,N_7252);
nand U14420 (N_14420,N_7192,N_9840);
nor U14421 (N_14421,N_5888,N_6035);
or U14422 (N_14422,N_8257,N_7726);
or U14423 (N_14423,N_9272,N_6596);
nor U14424 (N_14424,N_8825,N_8361);
or U14425 (N_14425,N_8454,N_7440);
nor U14426 (N_14426,N_9045,N_6155);
and U14427 (N_14427,N_7331,N_7615);
nor U14428 (N_14428,N_8231,N_5740);
xnor U14429 (N_14429,N_8791,N_7010);
nand U14430 (N_14430,N_8340,N_5912);
nor U14431 (N_14431,N_6646,N_9966);
and U14432 (N_14432,N_6860,N_8087);
xnor U14433 (N_14433,N_8424,N_7967);
nor U14434 (N_14434,N_9195,N_5292);
or U14435 (N_14435,N_5187,N_8800);
nor U14436 (N_14436,N_8476,N_7608);
and U14437 (N_14437,N_7976,N_9278);
nor U14438 (N_14438,N_5451,N_8591);
nand U14439 (N_14439,N_9001,N_6898);
nand U14440 (N_14440,N_5860,N_8846);
nand U14441 (N_14441,N_6140,N_6744);
or U14442 (N_14442,N_7161,N_6579);
nand U14443 (N_14443,N_7345,N_5673);
or U14444 (N_14444,N_8349,N_5869);
and U14445 (N_14445,N_7734,N_5285);
xor U14446 (N_14446,N_5922,N_9011);
nor U14447 (N_14447,N_9053,N_6883);
xnor U14448 (N_14448,N_8102,N_7662);
nand U14449 (N_14449,N_8557,N_8778);
nand U14450 (N_14450,N_7667,N_8284);
or U14451 (N_14451,N_8992,N_8822);
or U14452 (N_14452,N_8056,N_5659);
nor U14453 (N_14453,N_8453,N_6185);
nand U14454 (N_14454,N_5890,N_7606);
or U14455 (N_14455,N_5703,N_7343);
nand U14456 (N_14456,N_6590,N_6505);
and U14457 (N_14457,N_5377,N_5679);
and U14458 (N_14458,N_7897,N_8249);
or U14459 (N_14459,N_7333,N_9361);
xor U14460 (N_14460,N_6434,N_7949);
or U14461 (N_14461,N_9300,N_7590);
or U14462 (N_14462,N_6099,N_8231);
nand U14463 (N_14463,N_6136,N_6517);
nand U14464 (N_14464,N_5808,N_7385);
nor U14465 (N_14465,N_7613,N_6067);
nand U14466 (N_14466,N_9853,N_9091);
nor U14467 (N_14467,N_5935,N_8989);
and U14468 (N_14468,N_7187,N_8263);
nand U14469 (N_14469,N_5035,N_9855);
and U14470 (N_14470,N_5849,N_7777);
nand U14471 (N_14471,N_5348,N_7743);
or U14472 (N_14472,N_6010,N_5418);
nor U14473 (N_14473,N_5726,N_9600);
nand U14474 (N_14474,N_8646,N_9591);
and U14475 (N_14475,N_8147,N_5482);
or U14476 (N_14476,N_7681,N_8376);
and U14477 (N_14477,N_6472,N_6527);
or U14478 (N_14478,N_6876,N_9052);
xor U14479 (N_14479,N_6118,N_9697);
or U14480 (N_14480,N_8072,N_6320);
xnor U14481 (N_14481,N_8151,N_7221);
nor U14482 (N_14482,N_8864,N_5649);
and U14483 (N_14483,N_9104,N_6910);
and U14484 (N_14484,N_9606,N_9105);
nand U14485 (N_14485,N_6760,N_8572);
or U14486 (N_14486,N_8894,N_7859);
or U14487 (N_14487,N_6164,N_8752);
nand U14488 (N_14488,N_6525,N_7292);
nand U14489 (N_14489,N_7380,N_5695);
or U14490 (N_14490,N_5938,N_8357);
or U14491 (N_14491,N_6784,N_6032);
nand U14492 (N_14492,N_6373,N_7749);
or U14493 (N_14493,N_8933,N_6472);
and U14494 (N_14494,N_7553,N_7833);
or U14495 (N_14495,N_6001,N_5895);
or U14496 (N_14496,N_6356,N_5886);
nand U14497 (N_14497,N_6208,N_5701);
and U14498 (N_14498,N_7186,N_8148);
nor U14499 (N_14499,N_7495,N_5892);
nand U14500 (N_14500,N_8290,N_7166);
and U14501 (N_14501,N_5220,N_9169);
or U14502 (N_14502,N_6989,N_9821);
nor U14503 (N_14503,N_5508,N_7733);
nor U14504 (N_14504,N_6357,N_9521);
and U14505 (N_14505,N_9524,N_9403);
and U14506 (N_14506,N_5615,N_6302);
or U14507 (N_14507,N_8228,N_8705);
nand U14508 (N_14508,N_9949,N_6153);
nand U14509 (N_14509,N_6844,N_9923);
and U14510 (N_14510,N_8773,N_8238);
nor U14511 (N_14511,N_9133,N_6718);
or U14512 (N_14512,N_8454,N_9884);
nand U14513 (N_14513,N_5061,N_5044);
and U14514 (N_14514,N_7541,N_6983);
and U14515 (N_14515,N_8194,N_6482);
nand U14516 (N_14516,N_7235,N_8179);
and U14517 (N_14517,N_7027,N_8316);
nand U14518 (N_14518,N_5441,N_5832);
nor U14519 (N_14519,N_6457,N_5840);
and U14520 (N_14520,N_6892,N_5646);
nand U14521 (N_14521,N_6634,N_8427);
nand U14522 (N_14522,N_8472,N_7568);
nor U14523 (N_14523,N_5309,N_7271);
and U14524 (N_14524,N_7353,N_6695);
nor U14525 (N_14525,N_8548,N_8030);
or U14526 (N_14526,N_6383,N_8118);
nor U14527 (N_14527,N_6365,N_8251);
xnor U14528 (N_14528,N_7673,N_5787);
nand U14529 (N_14529,N_6426,N_5649);
xor U14530 (N_14530,N_6208,N_6247);
and U14531 (N_14531,N_5684,N_7424);
or U14532 (N_14532,N_5627,N_7238);
and U14533 (N_14533,N_7293,N_6220);
nor U14534 (N_14534,N_6932,N_9805);
or U14535 (N_14535,N_6490,N_8330);
nor U14536 (N_14536,N_5160,N_6717);
or U14537 (N_14537,N_7456,N_8136);
and U14538 (N_14538,N_9404,N_5884);
or U14539 (N_14539,N_7308,N_5302);
and U14540 (N_14540,N_9833,N_6074);
nand U14541 (N_14541,N_9099,N_9665);
nand U14542 (N_14542,N_8641,N_5776);
and U14543 (N_14543,N_9204,N_9611);
nor U14544 (N_14544,N_9999,N_6476);
and U14545 (N_14545,N_7841,N_9557);
nand U14546 (N_14546,N_5551,N_9260);
nand U14547 (N_14547,N_8671,N_6463);
or U14548 (N_14548,N_9604,N_7035);
and U14549 (N_14549,N_9329,N_5090);
nand U14550 (N_14550,N_5356,N_7973);
nor U14551 (N_14551,N_7318,N_7524);
and U14552 (N_14552,N_7841,N_9152);
or U14553 (N_14553,N_9868,N_6852);
and U14554 (N_14554,N_8843,N_8702);
and U14555 (N_14555,N_6779,N_8793);
nand U14556 (N_14556,N_9225,N_6512);
and U14557 (N_14557,N_8312,N_9088);
and U14558 (N_14558,N_6628,N_6255);
nand U14559 (N_14559,N_5655,N_7606);
and U14560 (N_14560,N_9520,N_9580);
nor U14561 (N_14561,N_6325,N_6521);
nor U14562 (N_14562,N_8214,N_6393);
nand U14563 (N_14563,N_7266,N_8443);
nand U14564 (N_14564,N_8982,N_9254);
nand U14565 (N_14565,N_8910,N_8599);
and U14566 (N_14566,N_8621,N_7747);
and U14567 (N_14567,N_6386,N_6290);
or U14568 (N_14568,N_9026,N_6329);
nor U14569 (N_14569,N_8480,N_7262);
nor U14570 (N_14570,N_7804,N_8258);
nor U14571 (N_14571,N_7182,N_8883);
nand U14572 (N_14572,N_6416,N_7453);
or U14573 (N_14573,N_6731,N_6614);
or U14574 (N_14574,N_7139,N_6035);
nor U14575 (N_14575,N_5690,N_8265);
nand U14576 (N_14576,N_8061,N_5661);
nand U14577 (N_14577,N_5970,N_9907);
nand U14578 (N_14578,N_7158,N_5245);
or U14579 (N_14579,N_6334,N_5369);
nand U14580 (N_14580,N_8695,N_8727);
or U14581 (N_14581,N_9953,N_5627);
or U14582 (N_14582,N_5355,N_6464);
nor U14583 (N_14583,N_8900,N_8944);
and U14584 (N_14584,N_5721,N_9165);
and U14585 (N_14585,N_5877,N_9789);
or U14586 (N_14586,N_5555,N_9748);
nor U14587 (N_14587,N_9139,N_8102);
nand U14588 (N_14588,N_6470,N_5301);
nor U14589 (N_14589,N_7634,N_8159);
and U14590 (N_14590,N_7406,N_5092);
nor U14591 (N_14591,N_5275,N_9044);
nand U14592 (N_14592,N_5875,N_5266);
nor U14593 (N_14593,N_7446,N_9260);
and U14594 (N_14594,N_8804,N_9341);
nor U14595 (N_14595,N_5102,N_5965);
nor U14596 (N_14596,N_6899,N_9123);
and U14597 (N_14597,N_5994,N_7932);
nand U14598 (N_14598,N_8652,N_7601);
nor U14599 (N_14599,N_9028,N_7353);
or U14600 (N_14600,N_8829,N_7397);
nor U14601 (N_14601,N_5402,N_9624);
nor U14602 (N_14602,N_5920,N_6788);
or U14603 (N_14603,N_7580,N_5201);
nor U14604 (N_14604,N_9092,N_5735);
xnor U14605 (N_14605,N_6709,N_7867);
or U14606 (N_14606,N_6315,N_8699);
and U14607 (N_14607,N_9407,N_9687);
and U14608 (N_14608,N_7766,N_5918);
or U14609 (N_14609,N_8848,N_6114);
and U14610 (N_14610,N_8730,N_6663);
and U14611 (N_14611,N_5753,N_9522);
nor U14612 (N_14612,N_9878,N_6264);
or U14613 (N_14613,N_6103,N_5481);
nand U14614 (N_14614,N_7677,N_7106);
or U14615 (N_14615,N_9236,N_8795);
nor U14616 (N_14616,N_7014,N_6704);
xor U14617 (N_14617,N_7411,N_6675);
or U14618 (N_14618,N_5758,N_5418);
and U14619 (N_14619,N_5682,N_5575);
and U14620 (N_14620,N_6257,N_5103);
and U14621 (N_14621,N_8670,N_6043);
nor U14622 (N_14622,N_7369,N_7266);
or U14623 (N_14623,N_8332,N_8333);
nor U14624 (N_14624,N_6287,N_7159);
and U14625 (N_14625,N_8323,N_5847);
or U14626 (N_14626,N_8577,N_7402);
or U14627 (N_14627,N_9604,N_9115);
nor U14628 (N_14628,N_8950,N_5780);
and U14629 (N_14629,N_7161,N_7480);
and U14630 (N_14630,N_8081,N_9423);
xor U14631 (N_14631,N_5544,N_8086);
nand U14632 (N_14632,N_6570,N_6207);
nor U14633 (N_14633,N_5185,N_9233);
xor U14634 (N_14634,N_5986,N_5382);
nand U14635 (N_14635,N_6624,N_8966);
nand U14636 (N_14636,N_5301,N_6871);
nor U14637 (N_14637,N_6061,N_8386);
and U14638 (N_14638,N_7459,N_5926);
nand U14639 (N_14639,N_7228,N_9849);
or U14640 (N_14640,N_9347,N_9667);
xnor U14641 (N_14641,N_7368,N_8308);
nor U14642 (N_14642,N_6201,N_7618);
or U14643 (N_14643,N_7737,N_8200);
or U14644 (N_14644,N_6993,N_5427);
nor U14645 (N_14645,N_9321,N_8639);
xnor U14646 (N_14646,N_5601,N_7290);
nor U14647 (N_14647,N_6822,N_7426);
nor U14648 (N_14648,N_8523,N_6046);
xor U14649 (N_14649,N_5386,N_6617);
xnor U14650 (N_14650,N_6932,N_6341);
or U14651 (N_14651,N_8023,N_7057);
and U14652 (N_14652,N_9488,N_6319);
nor U14653 (N_14653,N_7102,N_6362);
or U14654 (N_14654,N_5180,N_5487);
or U14655 (N_14655,N_8272,N_8264);
and U14656 (N_14656,N_6837,N_6156);
and U14657 (N_14657,N_9007,N_5351);
nand U14658 (N_14658,N_5664,N_5546);
xor U14659 (N_14659,N_5068,N_6412);
or U14660 (N_14660,N_6661,N_8696);
or U14661 (N_14661,N_8161,N_9582);
nand U14662 (N_14662,N_8514,N_7320);
nor U14663 (N_14663,N_5583,N_8240);
nand U14664 (N_14664,N_5293,N_5816);
or U14665 (N_14665,N_9644,N_7847);
or U14666 (N_14666,N_5371,N_8244);
and U14667 (N_14667,N_5645,N_9311);
and U14668 (N_14668,N_6047,N_5296);
and U14669 (N_14669,N_7472,N_7160);
and U14670 (N_14670,N_9244,N_9609);
xnor U14671 (N_14671,N_6094,N_8460);
or U14672 (N_14672,N_9659,N_8538);
nand U14673 (N_14673,N_5901,N_5027);
nand U14674 (N_14674,N_5549,N_8248);
and U14675 (N_14675,N_6272,N_6269);
xnor U14676 (N_14676,N_6734,N_6765);
nand U14677 (N_14677,N_5479,N_8474);
and U14678 (N_14678,N_5955,N_6469);
nand U14679 (N_14679,N_9870,N_5871);
and U14680 (N_14680,N_8438,N_8868);
nor U14681 (N_14681,N_8395,N_5116);
xor U14682 (N_14682,N_7008,N_8260);
nor U14683 (N_14683,N_6686,N_7446);
nand U14684 (N_14684,N_6613,N_9659);
nor U14685 (N_14685,N_7242,N_8632);
and U14686 (N_14686,N_7059,N_9375);
nor U14687 (N_14687,N_5236,N_5215);
and U14688 (N_14688,N_9411,N_6013);
nor U14689 (N_14689,N_9161,N_5333);
nand U14690 (N_14690,N_9566,N_6976);
or U14691 (N_14691,N_5232,N_6989);
or U14692 (N_14692,N_5671,N_8932);
or U14693 (N_14693,N_9497,N_5809);
xnor U14694 (N_14694,N_7796,N_5763);
nor U14695 (N_14695,N_7152,N_6570);
nor U14696 (N_14696,N_9049,N_6409);
nand U14697 (N_14697,N_5680,N_9495);
nand U14698 (N_14698,N_5449,N_8740);
nand U14699 (N_14699,N_9499,N_9417);
and U14700 (N_14700,N_5764,N_5680);
nand U14701 (N_14701,N_7973,N_8902);
nand U14702 (N_14702,N_7477,N_6486);
nor U14703 (N_14703,N_8897,N_8244);
and U14704 (N_14704,N_7152,N_9373);
and U14705 (N_14705,N_5168,N_7649);
or U14706 (N_14706,N_7889,N_9096);
xnor U14707 (N_14707,N_6719,N_7495);
or U14708 (N_14708,N_8190,N_5641);
or U14709 (N_14709,N_9642,N_6689);
or U14710 (N_14710,N_9115,N_6560);
nor U14711 (N_14711,N_8105,N_7076);
nand U14712 (N_14712,N_6987,N_8960);
nand U14713 (N_14713,N_7175,N_5597);
xnor U14714 (N_14714,N_9811,N_7803);
nand U14715 (N_14715,N_5784,N_9865);
or U14716 (N_14716,N_7311,N_6627);
nand U14717 (N_14717,N_7319,N_7318);
and U14718 (N_14718,N_9190,N_5381);
or U14719 (N_14719,N_7372,N_8813);
or U14720 (N_14720,N_5660,N_6489);
nor U14721 (N_14721,N_6001,N_8805);
xnor U14722 (N_14722,N_5080,N_7939);
and U14723 (N_14723,N_8965,N_7133);
xnor U14724 (N_14724,N_8455,N_5302);
or U14725 (N_14725,N_8559,N_6325);
nand U14726 (N_14726,N_6979,N_9297);
nand U14727 (N_14727,N_8911,N_6627);
nor U14728 (N_14728,N_8580,N_7298);
and U14729 (N_14729,N_7144,N_6864);
nor U14730 (N_14730,N_7720,N_6225);
nor U14731 (N_14731,N_9646,N_9572);
nand U14732 (N_14732,N_9428,N_8092);
or U14733 (N_14733,N_7198,N_9155);
nand U14734 (N_14734,N_9795,N_6893);
nand U14735 (N_14735,N_9596,N_9234);
xnor U14736 (N_14736,N_8287,N_5834);
or U14737 (N_14737,N_8668,N_5725);
nand U14738 (N_14738,N_5645,N_6115);
nand U14739 (N_14739,N_6507,N_9685);
nand U14740 (N_14740,N_5604,N_6095);
or U14741 (N_14741,N_5231,N_6454);
and U14742 (N_14742,N_5420,N_7149);
nand U14743 (N_14743,N_9548,N_8115);
and U14744 (N_14744,N_5225,N_7654);
xor U14745 (N_14745,N_9253,N_7469);
nand U14746 (N_14746,N_6909,N_9378);
or U14747 (N_14747,N_5675,N_5840);
or U14748 (N_14748,N_8628,N_6806);
and U14749 (N_14749,N_8863,N_7577);
or U14750 (N_14750,N_9089,N_9725);
xor U14751 (N_14751,N_8813,N_6281);
nand U14752 (N_14752,N_9495,N_8798);
nor U14753 (N_14753,N_9003,N_9389);
and U14754 (N_14754,N_7292,N_7881);
and U14755 (N_14755,N_7409,N_5118);
or U14756 (N_14756,N_9213,N_6334);
nor U14757 (N_14757,N_6844,N_7352);
nor U14758 (N_14758,N_5199,N_7234);
xor U14759 (N_14759,N_8612,N_7998);
nand U14760 (N_14760,N_9751,N_8190);
nor U14761 (N_14761,N_7092,N_6951);
or U14762 (N_14762,N_9540,N_7642);
and U14763 (N_14763,N_5117,N_7963);
nor U14764 (N_14764,N_7764,N_6757);
xor U14765 (N_14765,N_9043,N_8340);
nand U14766 (N_14766,N_8543,N_5788);
nor U14767 (N_14767,N_5380,N_7700);
or U14768 (N_14768,N_5764,N_7864);
nand U14769 (N_14769,N_7776,N_7157);
or U14770 (N_14770,N_8733,N_8102);
xor U14771 (N_14771,N_5055,N_5514);
and U14772 (N_14772,N_8601,N_8695);
or U14773 (N_14773,N_9838,N_6205);
and U14774 (N_14774,N_5490,N_8960);
nand U14775 (N_14775,N_5250,N_9011);
xor U14776 (N_14776,N_6722,N_9492);
nand U14777 (N_14777,N_8270,N_9190);
or U14778 (N_14778,N_9203,N_9131);
and U14779 (N_14779,N_5449,N_9083);
nand U14780 (N_14780,N_7138,N_7239);
nand U14781 (N_14781,N_5032,N_9021);
and U14782 (N_14782,N_6967,N_8663);
or U14783 (N_14783,N_8753,N_7246);
nor U14784 (N_14784,N_7801,N_5236);
nor U14785 (N_14785,N_8833,N_7980);
nor U14786 (N_14786,N_5564,N_5228);
nor U14787 (N_14787,N_8821,N_8940);
or U14788 (N_14788,N_5059,N_9008);
nand U14789 (N_14789,N_5821,N_6176);
nand U14790 (N_14790,N_6446,N_5274);
and U14791 (N_14791,N_6819,N_6310);
and U14792 (N_14792,N_6900,N_6096);
nor U14793 (N_14793,N_9605,N_6055);
nor U14794 (N_14794,N_6946,N_9914);
or U14795 (N_14795,N_5674,N_7152);
or U14796 (N_14796,N_8942,N_8468);
nor U14797 (N_14797,N_9463,N_7511);
xnor U14798 (N_14798,N_8730,N_7093);
nand U14799 (N_14799,N_7118,N_8490);
xnor U14800 (N_14800,N_9816,N_8963);
nand U14801 (N_14801,N_8595,N_8255);
nand U14802 (N_14802,N_9757,N_9406);
nand U14803 (N_14803,N_9017,N_9276);
nand U14804 (N_14804,N_9116,N_7584);
nor U14805 (N_14805,N_9349,N_7736);
nor U14806 (N_14806,N_8299,N_5223);
or U14807 (N_14807,N_5428,N_7730);
nand U14808 (N_14808,N_8373,N_9704);
nand U14809 (N_14809,N_6522,N_7208);
and U14810 (N_14810,N_8804,N_6456);
and U14811 (N_14811,N_7924,N_5731);
or U14812 (N_14812,N_6685,N_5207);
or U14813 (N_14813,N_9454,N_5908);
and U14814 (N_14814,N_6850,N_5063);
nor U14815 (N_14815,N_6209,N_6439);
xor U14816 (N_14816,N_7027,N_6533);
and U14817 (N_14817,N_7482,N_6077);
nor U14818 (N_14818,N_5956,N_7614);
nor U14819 (N_14819,N_7723,N_9864);
nand U14820 (N_14820,N_5819,N_8585);
or U14821 (N_14821,N_7367,N_9043);
nand U14822 (N_14822,N_8724,N_5805);
or U14823 (N_14823,N_8472,N_7985);
and U14824 (N_14824,N_8128,N_8819);
nor U14825 (N_14825,N_8673,N_8166);
nor U14826 (N_14826,N_6134,N_9822);
nand U14827 (N_14827,N_9565,N_9298);
nor U14828 (N_14828,N_6036,N_9237);
nor U14829 (N_14829,N_9070,N_7017);
nand U14830 (N_14830,N_9656,N_5228);
nor U14831 (N_14831,N_7575,N_8862);
xnor U14832 (N_14832,N_8796,N_8687);
xnor U14833 (N_14833,N_8626,N_8740);
or U14834 (N_14834,N_9102,N_6345);
xnor U14835 (N_14835,N_8610,N_5876);
and U14836 (N_14836,N_7656,N_9875);
nor U14837 (N_14837,N_7141,N_7794);
and U14838 (N_14838,N_6674,N_9751);
or U14839 (N_14839,N_5320,N_6969);
nand U14840 (N_14840,N_6627,N_9186);
nor U14841 (N_14841,N_6793,N_5332);
or U14842 (N_14842,N_5337,N_8202);
nor U14843 (N_14843,N_7801,N_6844);
nor U14844 (N_14844,N_7728,N_6762);
and U14845 (N_14845,N_8277,N_5665);
nor U14846 (N_14846,N_8185,N_7855);
and U14847 (N_14847,N_6230,N_8712);
and U14848 (N_14848,N_5504,N_8539);
or U14849 (N_14849,N_6369,N_7869);
nor U14850 (N_14850,N_7400,N_7831);
nor U14851 (N_14851,N_7536,N_6184);
xnor U14852 (N_14852,N_7528,N_8175);
nand U14853 (N_14853,N_6699,N_6358);
xor U14854 (N_14854,N_9537,N_5270);
nor U14855 (N_14855,N_5675,N_6164);
nor U14856 (N_14856,N_8062,N_7934);
nand U14857 (N_14857,N_6452,N_9064);
nand U14858 (N_14858,N_7072,N_6099);
nand U14859 (N_14859,N_8598,N_5174);
and U14860 (N_14860,N_9577,N_7368);
or U14861 (N_14861,N_5515,N_5658);
or U14862 (N_14862,N_6255,N_6947);
or U14863 (N_14863,N_9491,N_7420);
nor U14864 (N_14864,N_7313,N_8851);
nor U14865 (N_14865,N_8714,N_7634);
and U14866 (N_14866,N_8131,N_5422);
nor U14867 (N_14867,N_7323,N_8904);
nor U14868 (N_14868,N_7561,N_9422);
and U14869 (N_14869,N_5137,N_5758);
nand U14870 (N_14870,N_9784,N_6743);
nand U14871 (N_14871,N_9187,N_8105);
nand U14872 (N_14872,N_7690,N_7218);
and U14873 (N_14873,N_9147,N_5608);
nor U14874 (N_14874,N_8463,N_5542);
and U14875 (N_14875,N_9243,N_9192);
and U14876 (N_14876,N_7780,N_8390);
nand U14877 (N_14877,N_6187,N_6803);
nand U14878 (N_14878,N_8666,N_8226);
nand U14879 (N_14879,N_9587,N_8902);
nand U14880 (N_14880,N_8368,N_7479);
and U14881 (N_14881,N_8913,N_9402);
xor U14882 (N_14882,N_6348,N_8857);
nand U14883 (N_14883,N_8704,N_9711);
or U14884 (N_14884,N_5911,N_8064);
nor U14885 (N_14885,N_6234,N_8409);
nor U14886 (N_14886,N_6889,N_6045);
nand U14887 (N_14887,N_8086,N_7893);
nor U14888 (N_14888,N_6351,N_9742);
nor U14889 (N_14889,N_8077,N_9781);
nand U14890 (N_14890,N_5213,N_6930);
nor U14891 (N_14891,N_5774,N_6764);
nor U14892 (N_14892,N_8281,N_9757);
xor U14893 (N_14893,N_8087,N_9009);
nor U14894 (N_14894,N_6262,N_7092);
and U14895 (N_14895,N_5915,N_8002);
nor U14896 (N_14896,N_7135,N_9143);
and U14897 (N_14897,N_9665,N_6427);
nor U14898 (N_14898,N_5006,N_5418);
and U14899 (N_14899,N_6901,N_5778);
xor U14900 (N_14900,N_8607,N_9343);
xor U14901 (N_14901,N_7016,N_8689);
nand U14902 (N_14902,N_7767,N_6332);
xnor U14903 (N_14903,N_8527,N_6935);
nor U14904 (N_14904,N_7204,N_9986);
and U14905 (N_14905,N_8778,N_5843);
nand U14906 (N_14906,N_8662,N_7232);
nand U14907 (N_14907,N_5780,N_9779);
or U14908 (N_14908,N_7758,N_5338);
or U14909 (N_14909,N_7382,N_7783);
nand U14910 (N_14910,N_6160,N_9665);
nor U14911 (N_14911,N_5327,N_7913);
or U14912 (N_14912,N_9543,N_8319);
nor U14913 (N_14913,N_9960,N_7874);
and U14914 (N_14914,N_6978,N_7288);
xnor U14915 (N_14915,N_6872,N_6118);
nand U14916 (N_14916,N_6402,N_7065);
nor U14917 (N_14917,N_5257,N_5647);
and U14918 (N_14918,N_9397,N_8646);
xor U14919 (N_14919,N_9226,N_5388);
nor U14920 (N_14920,N_7105,N_6957);
or U14921 (N_14921,N_6995,N_9993);
xor U14922 (N_14922,N_8997,N_7888);
and U14923 (N_14923,N_7733,N_8481);
nand U14924 (N_14924,N_8491,N_8169);
and U14925 (N_14925,N_9020,N_9138);
nor U14926 (N_14926,N_6688,N_9744);
nand U14927 (N_14927,N_7456,N_5926);
xor U14928 (N_14928,N_7922,N_8318);
or U14929 (N_14929,N_8253,N_5390);
nor U14930 (N_14930,N_6581,N_5012);
and U14931 (N_14931,N_7242,N_6604);
and U14932 (N_14932,N_9253,N_8787);
nand U14933 (N_14933,N_8019,N_5547);
and U14934 (N_14934,N_6530,N_5469);
or U14935 (N_14935,N_8242,N_6755);
and U14936 (N_14936,N_9518,N_6676);
nand U14937 (N_14937,N_7577,N_6954);
and U14938 (N_14938,N_9854,N_5836);
nor U14939 (N_14939,N_7576,N_8600);
or U14940 (N_14940,N_7373,N_5699);
nor U14941 (N_14941,N_6082,N_6491);
nand U14942 (N_14942,N_5809,N_5447);
nand U14943 (N_14943,N_7971,N_9853);
nor U14944 (N_14944,N_9833,N_9130);
nand U14945 (N_14945,N_5453,N_5227);
and U14946 (N_14946,N_9492,N_5886);
and U14947 (N_14947,N_7277,N_8994);
or U14948 (N_14948,N_5135,N_7907);
nor U14949 (N_14949,N_9305,N_8006);
or U14950 (N_14950,N_8538,N_7763);
nand U14951 (N_14951,N_8182,N_8055);
or U14952 (N_14952,N_7569,N_6048);
xnor U14953 (N_14953,N_9622,N_6504);
nand U14954 (N_14954,N_9794,N_5218);
and U14955 (N_14955,N_5576,N_5680);
nor U14956 (N_14956,N_7592,N_6586);
nand U14957 (N_14957,N_5310,N_9458);
xor U14958 (N_14958,N_7446,N_7119);
nand U14959 (N_14959,N_6744,N_8942);
nand U14960 (N_14960,N_7774,N_8119);
or U14961 (N_14961,N_7569,N_5527);
or U14962 (N_14962,N_5932,N_9264);
and U14963 (N_14963,N_5606,N_7329);
or U14964 (N_14964,N_8530,N_9213);
nor U14965 (N_14965,N_5099,N_8500);
and U14966 (N_14966,N_9050,N_9744);
nand U14967 (N_14967,N_8036,N_9523);
and U14968 (N_14968,N_8081,N_6674);
or U14969 (N_14969,N_8682,N_8253);
nand U14970 (N_14970,N_6574,N_5354);
xor U14971 (N_14971,N_9178,N_9775);
nor U14972 (N_14972,N_5505,N_9813);
nand U14973 (N_14973,N_5122,N_7991);
or U14974 (N_14974,N_5655,N_9191);
and U14975 (N_14975,N_7806,N_6747);
nor U14976 (N_14976,N_7636,N_8981);
xnor U14977 (N_14977,N_5134,N_8926);
or U14978 (N_14978,N_6663,N_7425);
nand U14979 (N_14979,N_7179,N_9652);
or U14980 (N_14980,N_5280,N_8048);
xor U14981 (N_14981,N_8876,N_9633);
nand U14982 (N_14982,N_8847,N_5675);
or U14983 (N_14983,N_8870,N_7770);
or U14984 (N_14984,N_9304,N_5959);
nand U14985 (N_14985,N_7041,N_9188);
and U14986 (N_14986,N_5538,N_7225);
xor U14987 (N_14987,N_7972,N_7875);
or U14988 (N_14988,N_8027,N_5152);
or U14989 (N_14989,N_5968,N_9031);
nand U14990 (N_14990,N_5999,N_8759);
nor U14991 (N_14991,N_5174,N_7403);
nor U14992 (N_14992,N_5508,N_6975);
nor U14993 (N_14993,N_6436,N_8840);
nand U14994 (N_14994,N_8108,N_6741);
xnor U14995 (N_14995,N_7798,N_9381);
nand U14996 (N_14996,N_8708,N_5529);
nor U14997 (N_14997,N_9052,N_7876);
nand U14998 (N_14998,N_5875,N_5524);
or U14999 (N_14999,N_6936,N_8843);
and UO_0 (O_0,N_14614,N_11912);
nand UO_1 (O_1,N_10897,N_13953);
nand UO_2 (O_2,N_10776,N_12113);
or UO_3 (O_3,N_12127,N_10971);
or UO_4 (O_4,N_14224,N_10644);
nand UO_5 (O_5,N_11847,N_11278);
or UO_6 (O_6,N_13823,N_10909);
or UO_7 (O_7,N_13401,N_13513);
and UO_8 (O_8,N_14307,N_12834);
and UO_9 (O_9,N_11559,N_13882);
or UO_10 (O_10,N_13389,N_11526);
and UO_11 (O_11,N_10052,N_13411);
xnor UO_12 (O_12,N_14930,N_14944);
and UO_13 (O_13,N_10327,N_11984);
and UO_14 (O_14,N_12605,N_13161);
nand UO_15 (O_15,N_10062,N_14085);
nor UO_16 (O_16,N_10175,N_10854);
or UO_17 (O_17,N_11011,N_12081);
and UO_18 (O_18,N_10920,N_13450);
or UO_19 (O_19,N_14851,N_11820);
or UO_20 (O_20,N_11357,N_10713);
nor UO_21 (O_21,N_14675,N_11301);
nor UO_22 (O_22,N_14560,N_13261);
xnor UO_23 (O_23,N_10057,N_12474);
nor UO_24 (O_24,N_14194,N_14423);
nand UO_25 (O_25,N_14990,N_13655);
nand UO_26 (O_26,N_13364,N_10182);
or UO_27 (O_27,N_14342,N_13010);
or UO_28 (O_28,N_14884,N_10682);
nor UO_29 (O_29,N_14980,N_13277);
nor UO_30 (O_30,N_11591,N_11259);
or UO_31 (O_31,N_13665,N_14165);
nand UO_32 (O_32,N_13127,N_11530);
and UO_33 (O_33,N_12946,N_11411);
nor UO_34 (O_34,N_14648,N_12489);
or UO_35 (O_35,N_11106,N_11406);
and UO_36 (O_36,N_12135,N_14511);
nor UO_37 (O_37,N_10792,N_14719);
nor UO_38 (O_38,N_10267,N_12886);
nor UO_39 (O_39,N_14592,N_14200);
nor UO_40 (O_40,N_12402,N_13550);
and UO_41 (O_41,N_11523,N_10159);
nand UO_42 (O_42,N_12646,N_10141);
and UO_43 (O_43,N_10108,N_11175);
or UO_44 (O_44,N_14397,N_14067);
nor UO_45 (O_45,N_11068,N_11260);
and UO_46 (O_46,N_13527,N_10212);
nand UO_47 (O_47,N_10911,N_13256);
and UO_48 (O_48,N_11448,N_12577);
xor UO_49 (O_49,N_10051,N_10979);
and UO_50 (O_50,N_13770,N_11556);
nand UO_51 (O_51,N_10600,N_10518);
or UO_52 (O_52,N_11635,N_10030);
nor UO_53 (O_53,N_13562,N_11241);
xnor UO_54 (O_54,N_10548,N_11945);
nor UO_55 (O_55,N_13821,N_13503);
or UO_56 (O_56,N_10875,N_11898);
nor UO_57 (O_57,N_12374,N_13995);
and UO_58 (O_58,N_12719,N_14618);
nand UO_59 (O_59,N_13881,N_10386);
and UO_60 (O_60,N_14570,N_11949);
or UO_61 (O_61,N_12027,N_11538);
nand UO_62 (O_62,N_11296,N_12410);
and UO_63 (O_63,N_12465,N_14571);
and UO_64 (O_64,N_11210,N_14345);
and UO_65 (O_65,N_11777,N_11476);
and UO_66 (O_66,N_12133,N_14802);
xnor UO_67 (O_67,N_10752,N_10213);
and UO_68 (O_68,N_10705,N_14781);
and UO_69 (O_69,N_11959,N_14244);
and UO_70 (O_70,N_13819,N_13347);
and UO_71 (O_71,N_14514,N_14185);
or UO_72 (O_72,N_13700,N_10860);
or UO_73 (O_73,N_12412,N_14332);
nor UO_74 (O_74,N_10173,N_13789);
and UO_75 (O_75,N_14541,N_13748);
or UO_76 (O_76,N_14487,N_11835);
or UO_77 (O_77,N_10310,N_14764);
and UO_78 (O_78,N_12877,N_12009);
or UO_79 (O_79,N_12989,N_10525);
or UO_80 (O_80,N_12645,N_11824);
nand UO_81 (O_81,N_10719,N_14843);
or UO_82 (O_82,N_10318,N_13738);
nand UO_83 (O_83,N_13293,N_13908);
nor UO_84 (O_84,N_11087,N_12068);
xnor UO_85 (O_85,N_14279,N_13142);
or UO_86 (O_86,N_11300,N_14286);
xor UO_87 (O_87,N_12040,N_14956);
or UO_88 (O_88,N_10599,N_12999);
xnor UO_89 (O_89,N_14892,N_11646);
nor UO_90 (O_90,N_12026,N_11261);
nand UO_91 (O_91,N_13940,N_11943);
xnor UO_92 (O_92,N_13420,N_12682);
and UO_93 (O_93,N_14533,N_14744);
nor UO_94 (O_94,N_13195,N_12840);
and UO_95 (O_95,N_10556,N_14965);
nor UO_96 (O_96,N_13791,N_11527);
xor UO_97 (O_97,N_10199,N_12299);
and UO_98 (O_98,N_11219,N_11931);
and UO_99 (O_99,N_14974,N_10382);
or UO_100 (O_100,N_11314,N_11917);
nor UO_101 (O_101,N_10029,N_12042);
nor UO_102 (O_102,N_13581,N_10769);
or UO_103 (O_103,N_11188,N_14867);
or UO_104 (O_104,N_12253,N_13651);
and UO_105 (O_105,N_14115,N_12643);
or UO_106 (O_106,N_14605,N_12310);
nor UO_107 (O_107,N_12647,N_11829);
nor UO_108 (O_108,N_11404,N_13190);
or UO_109 (O_109,N_13184,N_12820);
and UO_110 (O_110,N_12771,N_10228);
or UO_111 (O_111,N_13152,N_11623);
nand UO_112 (O_112,N_12794,N_10586);
and UO_113 (O_113,N_10862,N_12676);
or UO_114 (O_114,N_10451,N_12243);
nor UO_115 (O_115,N_12229,N_12066);
nand UO_116 (O_116,N_10211,N_14335);
nor UO_117 (O_117,N_10903,N_11833);
or UO_118 (O_118,N_10631,N_14470);
and UO_119 (O_119,N_12504,N_11694);
nand UO_120 (O_120,N_14654,N_11667);
and UO_121 (O_121,N_12260,N_11170);
and UO_122 (O_122,N_11946,N_14769);
nand UO_123 (O_123,N_13658,N_10630);
nand UO_124 (O_124,N_12439,N_13050);
and UO_125 (O_125,N_11294,N_12190);
nand UO_126 (O_126,N_12912,N_13439);
nor UO_127 (O_127,N_10954,N_14117);
or UO_128 (O_128,N_12815,N_13484);
or UO_129 (O_129,N_11209,N_13680);
nand UO_130 (O_130,N_13039,N_11127);
nor UO_131 (O_131,N_14603,N_11579);
nand UO_132 (O_132,N_10594,N_12411);
nor UO_133 (O_133,N_12369,N_14049);
and UO_134 (O_134,N_13017,N_13002);
or UO_135 (O_135,N_10014,N_12514);
nand UO_136 (O_136,N_13070,N_13843);
nand UO_137 (O_137,N_14650,N_13260);
or UO_138 (O_138,N_12881,N_13577);
nor UO_139 (O_139,N_11644,N_14242);
nor UO_140 (O_140,N_13345,N_13631);
nand UO_141 (O_141,N_11135,N_12516);
xnor UO_142 (O_142,N_13165,N_14499);
and UO_143 (O_143,N_11573,N_12657);
or UO_144 (O_144,N_10231,N_14938);
and UO_145 (O_145,N_11168,N_12562);
nand UO_146 (O_146,N_13136,N_14078);
and UO_147 (O_147,N_11304,N_14091);
or UO_148 (O_148,N_12856,N_13031);
or UO_149 (O_149,N_13210,N_13979);
or UO_150 (O_150,N_14072,N_10272);
xnor UO_151 (O_151,N_13699,N_13653);
nand UO_152 (O_152,N_11902,N_13138);
and UO_153 (O_153,N_14850,N_13637);
or UO_154 (O_154,N_14154,N_11090);
or UO_155 (O_155,N_11332,N_13590);
nand UO_156 (O_156,N_12426,N_13842);
and UO_157 (O_157,N_14416,N_10571);
nor UO_158 (O_158,N_14303,N_14446);
xnor UO_159 (O_159,N_13643,N_12298);
nor UO_160 (O_160,N_13755,N_14164);
or UO_161 (O_161,N_14700,N_11504);
nand UO_162 (O_162,N_11725,N_11836);
nand UO_163 (O_163,N_12874,N_11749);
and UO_164 (O_164,N_13857,N_14756);
nand UO_165 (O_165,N_10890,N_13215);
nand UO_166 (O_166,N_10957,N_10237);
nor UO_167 (O_167,N_13774,N_13160);
nand UO_168 (O_168,N_14429,N_11861);
and UO_169 (O_169,N_12028,N_10385);
nor UO_170 (O_170,N_10045,N_11325);
nor UO_171 (O_171,N_10475,N_11617);
or UO_172 (O_172,N_13130,N_13818);
nor UO_173 (O_173,N_11409,N_14052);
and UO_174 (O_174,N_11763,N_13139);
nor UO_175 (O_175,N_12328,N_14858);
and UO_176 (O_176,N_12954,N_11752);
nand UO_177 (O_177,N_10892,N_13758);
and UO_178 (O_178,N_14264,N_11044);
or UO_179 (O_179,N_10483,N_11501);
or UO_180 (O_180,N_14882,N_10239);
and UO_181 (O_181,N_11452,N_12007);
or UO_182 (O_182,N_12166,N_10789);
or UO_183 (O_183,N_13100,N_10166);
and UO_184 (O_184,N_13385,N_12824);
nand UO_185 (O_185,N_10526,N_14494);
nand UO_186 (O_186,N_14210,N_13896);
xnor UO_187 (O_187,N_14056,N_10528);
and UO_188 (O_188,N_10895,N_12837);
nand UO_189 (O_189,N_13088,N_12958);
nor UO_190 (O_190,N_12724,N_14437);
nor UO_191 (O_191,N_10395,N_14540);
or UO_192 (O_192,N_11052,N_11095);
nor UO_193 (O_193,N_13993,N_13131);
or UO_194 (O_194,N_12276,N_13778);
nand UO_195 (O_195,N_11512,N_12383);
nor UO_196 (O_196,N_12671,N_10210);
or UO_197 (O_197,N_14656,N_13098);
and UO_198 (O_198,N_10939,N_13464);
and UO_199 (O_199,N_12071,N_14667);
nor UO_200 (O_200,N_12679,N_14529);
nor UO_201 (O_201,N_14193,N_10338);
nand UO_202 (O_202,N_12231,N_14142);
and UO_203 (O_203,N_12680,N_13853);
or UO_204 (O_204,N_11392,N_13648);
nand UO_205 (O_205,N_12666,N_11568);
and UO_206 (O_206,N_11212,N_14758);
nor UO_207 (O_207,N_10624,N_12628);
or UO_208 (O_208,N_10142,N_14120);
nor UO_209 (O_209,N_13382,N_13056);
and UO_210 (O_210,N_13478,N_11181);
and UO_211 (O_211,N_12911,N_11198);
and UO_212 (O_212,N_13588,N_11930);
and UO_213 (O_213,N_11952,N_11475);
nand UO_214 (O_214,N_12070,N_10236);
nand UO_215 (O_215,N_11654,N_11834);
and UO_216 (O_216,N_12300,N_12313);
nor UO_217 (O_217,N_14737,N_10059);
or UO_218 (O_218,N_14704,N_12082);
nand UO_219 (O_219,N_12897,N_10330);
nor UO_220 (O_220,N_14891,N_13945);
nor UO_221 (O_221,N_14443,N_10986);
nor UO_222 (O_222,N_12960,N_13296);
and UO_223 (O_223,N_13122,N_11904);
and UO_224 (O_224,N_13434,N_13745);
nor UO_225 (O_225,N_14839,N_10956);
nor UO_226 (O_226,N_10540,N_10550);
nand UO_227 (O_227,N_13801,N_10855);
xnor UO_228 (O_228,N_10400,N_13558);
nand UO_229 (O_229,N_13603,N_11603);
nand UO_230 (O_230,N_10521,N_12611);
nor UO_231 (O_231,N_13063,N_10282);
nor UO_232 (O_232,N_12937,N_13222);
nor UO_233 (O_233,N_12029,N_10100);
and UO_234 (O_234,N_12626,N_13423);
nand UO_235 (O_235,N_13390,N_11599);
or UO_236 (O_236,N_12964,N_14204);
or UO_237 (O_237,N_13959,N_10061);
nand UO_238 (O_238,N_11339,N_11905);
nor UO_239 (O_239,N_14819,N_14993);
nand UO_240 (O_240,N_12708,N_13368);
and UO_241 (O_241,N_11581,N_14042);
nor UO_242 (O_242,N_13875,N_14326);
nand UO_243 (O_243,N_12011,N_12161);
nor UO_244 (O_244,N_14348,N_13790);
and UO_245 (O_245,N_10646,N_12706);
nor UO_246 (O_246,N_12675,N_12479);
nor UO_247 (O_247,N_10777,N_10053);
or UO_248 (O_248,N_14738,N_14496);
nand UO_249 (O_249,N_13621,N_12084);
or UO_250 (O_250,N_12574,N_13556);
nand UO_251 (O_251,N_12335,N_10444);
or UO_252 (O_252,N_13013,N_11534);
nor UO_253 (O_253,N_14674,N_12156);
and UO_254 (O_254,N_13114,N_13982);
or UO_255 (O_255,N_13150,N_14623);
or UO_256 (O_256,N_14823,N_14714);
xor UO_257 (O_257,N_12726,N_11896);
or UO_258 (O_258,N_14889,N_13822);
and UO_259 (O_259,N_10465,N_12786);
nor UO_260 (O_260,N_14825,N_14915);
and UO_261 (O_261,N_11852,N_11439);
nor UO_262 (O_262,N_11340,N_11493);
or UO_263 (O_263,N_13447,N_13463);
or UO_264 (O_264,N_10036,N_13416);
or UO_265 (O_265,N_11253,N_10974);
and UO_266 (O_266,N_10454,N_10703);
or UO_267 (O_267,N_11506,N_11808);
or UO_268 (O_268,N_10568,N_11935);
and UO_269 (O_269,N_10573,N_10563);
xnor UO_270 (O_270,N_12755,N_14518);
nor UO_271 (O_271,N_13760,N_11481);
xor UO_272 (O_272,N_13816,N_11310);
nor UO_273 (O_273,N_14246,N_13797);
xor UO_274 (O_274,N_10094,N_14118);
nor UO_275 (O_275,N_13291,N_13584);
and UO_276 (O_276,N_13904,N_13099);
nor UO_277 (O_277,N_14989,N_14346);
nand UO_278 (O_278,N_11708,N_13807);
or UO_279 (O_279,N_12875,N_10641);
or UO_280 (O_280,N_13473,N_13639);
nor UO_281 (O_281,N_11477,N_14163);
nor UO_282 (O_282,N_11350,N_10306);
nor UO_283 (O_283,N_11862,N_12921);
or UO_284 (O_284,N_12406,N_14642);
nand UO_285 (O_285,N_10998,N_10350);
nand UO_286 (O_286,N_10021,N_13043);
xor UO_287 (O_287,N_14096,N_11728);
and UO_288 (O_288,N_14613,N_11462);
and UO_289 (O_289,N_14879,N_10771);
or UO_290 (O_290,N_14316,N_14151);
nand UO_291 (O_291,N_11699,N_11323);
nor UO_292 (O_292,N_12083,N_14372);
or UO_293 (O_293,N_12783,N_12076);
nor UO_294 (O_294,N_14886,N_12491);
xor UO_295 (O_295,N_12423,N_10251);
nand UO_296 (O_296,N_12058,N_13972);
nor UO_297 (O_297,N_10812,N_14698);
and UO_298 (O_298,N_12902,N_12947);
and UO_299 (O_299,N_14266,N_11059);
nor UO_300 (O_300,N_13897,N_10531);
or UO_301 (O_301,N_10613,N_12545);
or UO_302 (O_302,N_11343,N_12022);
and UO_303 (O_303,N_10346,N_10990);
or UO_304 (O_304,N_14475,N_11626);
or UO_305 (O_305,N_11971,N_11919);
nand UO_306 (O_306,N_11213,N_14713);
and UO_307 (O_307,N_10214,N_11584);
nand UO_308 (O_308,N_13985,N_10118);
or UO_309 (O_309,N_12373,N_12388);
nand UO_310 (O_310,N_11562,N_11001);
nor UO_311 (O_311,N_13384,N_12012);
and UO_312 (O_312,N_12554,N_10167);
nand UO_313 (O_313,N_11467,N_11826);
or UO_314 (O_314,N_13788,N_12717);
or UO_315 (O_315,N_11140,N_14816);
nand UO_316 (O_316,N_11792,N_13155);
nand UO_317 (O_317,N_14040,N_13606);
xnor UO_318 (O_318,N_12879,N_14804);
and UO_319 (O_319,N_11064,N_14716);
nand UO_320 (O_320,N_13518,N_12255);
and UO_321 (O_321,N_11753,N_13548);
or UO_322 (O_322,N_14874,N_12334);
or UO_323 (O_323,N_10656,N_10733);
or UO_324 (O_324,N_13943,N_10222);
xor UO_325 (O_325,N_10806,N_11660);
or UO_326 (O_326,N_14114,N_10828);
nand UO_327 (O_327,N_13640,N_12450);
or UO_328 (O_328,N_10435,N_12621);
or UO_329 (O_329,N_10924,N_12641);
nand UO_330 (O_330,N_10022,N_13538);
and UO_331 (O_331,N_11152,N_11857);
nor UO_332 (O_332,N_13027,N_11316);
nand UO_333 (O_333,N_12592,N_13105);
or UO_334 (O_334,N_14350,N_14616);
or UO_335 (O_335,N_12606,N_13274);
or UO_336 (O_336,N_11016,N_13193);
xor UO_337 (O_337,N_11057,N_10690);
nor UO_338 (O_338,N_11262,N_11767);
nor UO_339 (O_339,N_14840,N_14094);
nor UO_340 (O_340,N_10541,N_13486);
xnor UO_341 (O_341,N_14004,N_13804);
and UO_342 (O_342,N_11061,N_12660);
nor UO_343 (O_343,N_10598,N_10050);
nor UO_344 (O_344,N_12435,N_10420);
nor UO_345 (O_345,N_13925,N_10219);
xor UO_346 (O_346,N_11202,N_11208);
nand UO_347 (O_347,N_14864,N_14972);
nor UO_348 (O_348,N_14741,N_12064);
nor UO_349 (O_349,N_14670,N_14920);
nor UO_350 (O_350,N_12387,N_11369);
nor UO_351 (O_351,N_10148,N_14845);
nor UO_352 (O_352,N_10693,N_11056);
and UO_353 (O_353,N_13858,N_14685);
nand UO_354 (O_354,N_10574,N_13634);
or UO_355 (O_355,N_11828,N_13701);
xor UO_356 (O_356,N_12268,N_14373);
or UO_357 (O_357,N_10084,N_12159);
nand UO_358 (O_358,N_10487,N_12976);
and UO_359 (O_359,N_13487,N_14009);
nor UO_360 (O_360,N_12662,N_12443);
or UO_361 (O_361,N_10996,N_13325);
nor UO_362 (O_362,N_10116,N_12106);
and UO_363 (O_363,N_11105,N_12583);
or UO_364 (O_364,N_11410,N_12111);
and UO_365 (O_365,N_13311,N_13137);
xnor UO_366 (O_366,N_14485,N_14452);
and UO_367 (O_367,N_12473,N_14543);
and UO_368 (O_368,N_14601,N_11881);
nor UO_369 (O_369,N_12788,N_12674);
nor UO_370 (O_370,N_12975,N_14299);
or UO_371 (O_371,N_13149,N_14697);
and UO_372 (O_372,N_12468,N_10925);
nand UO_373 (O_373,N_14772,N_14523);
nand UO_374 (O_374,N_13488,N_10344);
nor UO_375 (O_375,N_11220,N_11967);
or UO_376 (O_376,N_11283,N_10028);
xnor UO_377 (O_377,N_14051,N_11096);
or UO_378 (O_378,N_10155,N_11938);
nor UO_379 (O_379,N_14222,N_14537);
nand UO_380 (O_380,N_10750,N_13987);
and UO_381 (O_381,N_11111,N_14073);
nor UO_382 (O_382,N_13042,N_14849);
nor UO_383 (O_383,N_12321,N_13549);
and UO_384 (O_384,N_12077,N_11953);
or UO_385 (O_385,N_14389,N_13712);
nand UO_386 (O_386,N_12032,N_10362);
and UO_387 (O_387,N_11223,N_13044);
nand UO_388 (O_388,N_10217,N_11863);
or UO_389 (O_389,N_12703,N_12134);
and UO_390 (O_390,N_12579,N_11236);
nor UO_391 (O_391,N_14268,N_10151);
nor UO_392 (O_392,N_13598,N_13182);
nor UO_393 (O_393,N_13438,N_14676);
nand UO_394 (O_394,N_14320,N_14739);
or UO_395 (O_395,N_14968,N_10507);
nor UO_396 (O_396,N_12804,N_14167);
nand UO_397 (O_397,N_13301,N_14767);
or UO_398 (O_398,N_13014,N_10720);
xor UO_399 (O_399,N_12700,N_14016);
or UO_400 (O_400,N_10512,N_12205);
and UO_401 (O_401,N_12015,N_13086);
nand UO_402 (O_402,N_14095,N_14219);
nor UO_403 (O_403,N_14856,N_13468);
nand UO_404 (O_404,N_14014,N_10287);
and UO_405 (O_405,N_13624,N_12521);
or UO_406 (O_406,N_14524,N_13188);
and UO_407 (O_407,N_11637,N_10074);
or UO_408 (O_408,N_10423,N_12385);
or UO_409 (O_409,N_10933,N_12586);
nand UO_410 (O_410,N_10683,N_13886);
or UO_411 (O_411,N_13154,N_10826);
or UO_412 (O_412,N_10716,N_12180);
nand UO_413 (O_413,N_13349,N_14206);
or UO_414 (O_414,N_10622,N_11201);
nor UO_415 (O_415,N_13388,N_11718);
and UO_416 (O_416,N_10744,N_14731);
or UO_417 (O_417,N_13749,N_12224);
nor UO_418 (O_418,N_13294,N_12761);
and UO_419 (O_419,N_14566,N_10421);
xor UO_420 (O_420,N_13064,N_11769);
nor UO_421 (O_421,N_12904,N_11832);
xnor UO_422 (O_422,N_10987,N_12456);
nand UO_423 (O_423,N_11146,N_10628);
or UO_424 (O_424,N_14595,N_12930);
or UO_425 (O_425,N_13870,N_12060);
and UO_426 (O_426,N_14636,N_12734);
or UO_427 (O_427,N_12144,N_10808);
or UO_428 (O_428,N_14702,N_12471);
nand UO_429 (O_429,N_11706,N_13900);
nand UO_430 (O_430,N_10853,N_13961);
nand UO_431 (O_431,N_12857,N_13459);
nand UO_432 (O_432,N_10952,N_12668);
xor UO_433 (O_433,N_10603,N_12803);
or UO_434 (O_434,N_11774,N_10227);
or UO_435 (O_435,N_14564,N_11440);
and UO_436 (O_436,N_13009,N_13094);
or UO_437 (O_437,N_10846,N_13794);
nor UO_438 (O_438,N_14929,N_14466);
nor UO_439 (O_439,N_14484,N_13912);
nor UO_440 (O_440,N_14135,N_12951);
and UO_441 (O_441,N_13555,N_10527);
and UO_442 (O_442,N_11229,N_13242);
and UO_443 (O_443,N_12983,N_13183);
or UO_444 (O_444,N_11614,N_11850);
nand UO_445 (O_445,N_11915,N_12017);
nor UO_446 (O_446,N_10662,N_14836);
xor UO_447 (O_447,N_10044,N_14138);
or UO_448 (O_448,N_12594,N_13072);
or UO_449 (O_449,N_10503,N_13844);
nand UO_450 (O_450,N_13828,N_10146);
nand UO_451 (O_451,N_13023,N_13431);
nand UO_452 (O_452,N_12202,N_13626);
and UO_453 (O_453,N_14383,N_12195);
nor UO_454 (O_454,N_13968,N_12116);
and UO_455 (O_455,N_11545,N_13197);
and UO_456 (O_456,N_10005,N_13251);
and UO_457 (O_457,N_10796,N_12050);
nor UO_458 (O_458,N_14183,N_11216);
nand UO_459 (O_459,N_11804,N_13954);
xnor UO_460 (O_460,N_12063,N_10658);
nand UO_461 (O_461,N_10001,N_10611);
or UO_462 (O_462,N_12633,N_10374);
and UO_463 (O_463,N_12532,N_12293);
nand UO_464 (O_464,N_13695,N_12138);
and UO_465 (O_465,N_12528,N_11567);
or UO_466 (O_466,N_14652,N_14983);
nor UO_467 (O_467,N_13557,N_10940);
nor UO_468 (O_468,N_12262,N_14969);
and UO_469 (O_469,N_12740,N_14671);
nand UO_470 (O_470,N_11239,N_11680);
nand UO_471 (O_471,N_14734,N_11600);
and UO_472 (O_472,N_13803,N_12887);
nand UO_473 (O_473,N_10262,N_12955);
nor UO_474 (O_474,N_11782,N_10366);
nor UO_475 (O_475,N_13723,N_10476);
or UO_476 (O_476,N_13834,N_12792);
or UO_477 (O_477,N_13007,N_14593);
nand UO_478 (O_478,N_14630,N_12573);
nor UO_479 (O_479,N_11040,N_12663);
and UO_480 (O_480,N_13033,N_13540);
and UO_481 (O_481,N_14917,N_13799);
or UO_482 (O_482,N_12520,N_12922);
and UO_483 (O_483,N_12120,N_12123);
xnor UO_484 (O_484,N_11653,N_11375);
and UO_485 (O_485,N_11693,N_13359);
and UO_486 (O_486,N_11269,N_12893);
or UO_487 (O_487,N_11793,N_10647);
nand UO_488 (O_488,N_13898,N_13236);
xnor UO_489 (O_489,N_11539,N_14122);
or UO_490 (O_490,N_10835,N_12544);
xor UO_491 (O_491,N_11355,N_13074);
or UO_492 (O_492,N_12670,N_11430);
or UO_493 (O_493,N_13406,N_14597);
and UO_494 (O_494,N_12392,N_14863);
nand UO_495 (O_495,N_11453,N_10840);
nand UO_496 (O_496,N_13232,N_14418);
nor UO_497 (O_497,N_11073,N_12961);
and UO_498 (O_498,N_11727,N_13418);
nor UO_499 (O_499,N_12816,N_13931);
and UO_500 (O_500,N_11317,N_13342);
nor UO_501 (O_501,N_14844,N_11492);
and UO_502 (O_502,N_12838,N_14292);
and UO_503 (O_503,N_10587,N_13906);
or UO_504 (O_504,N_11674,N_12099);
xnor UO_505 (O_505,N_12723,N_13263);
nand UO_506 (O_506,N_13091,N_13874);
nand UO_507 (O_507,N_14202,N_12796);
nand UO_508 (O_508,N_11601,N_11060);
nand UO_509 (O_509,N_13836,N_10448);
nor UO_510 (O_510,N_10016,N_12197);
and UO_511 (O_511,N_11129,N_13353);
nor UO_512 (O_512,N_11385,N_10742);
or UO_513 (O_513,N_14937,N_12873);
nor UO_514 (O_514,N_13271,N_14251);
and UO_515 (O_515,N_13292,N_13737);
or UO_516 (O_516,N_14762,N_13559);
nor UO_517 (O_517,N_10779,N_12010);
or UO_518 (O_518,N_10801,N_10864);
xnor UO_519 (O_519,N_10431,N_11378);
nand UO_520 (O_520,N_11437,N_12536);
or UO_521 (O_521,N_14861,N_13726);
nand UO_522 (O_522,N_11775,N_10495);
xnor UO_523 (O_523,N_14542,N_10802);
and UO_524 (O_524,N_11083,N_12432);
and UO_525 (O_525,N_14786,N_12183);
nand UO_526 (O_526,N_14790,N_12575);
nor UO_527 (O_527,N_14233,N_14637);
nor UO_528 (O_528,N_13209,N_14344);
xor UO_529 (O_529,N_14860,N_13860);
and UO_530 (O_530,N_12326,N_10532);
nand UO_531 (O_531,N_14363,N_12057);
nand UO_532 (O_532,N_11926,N_14057);
and UO_533 (O_533,N_14872,N_13890);
nand UO_534 (O_534,N_14378,N_13732);
and UO_535 (O_535,N_14288,N_13185);
nand UO_536 (O_536,N_12130,N_13851);
nand UO_537 (O_537,N_14712,N_12409);
or UO_538 (O_538,N_12888,N_11276);
nand UO_539 (O_539,N_12351,N_10091);
or UO_540 (O_540,N_10552,N_14551);
or UO_541 (O_541,N_13286,N_12110);
or UO_542 (O_542,N_14512,N_12522);
and UO_543 (O_543,N_13761,N_11705);
or UO_544 (O_544,N_11342,N_14628);
xor UO_545 (O_545,N_10634,N_13047);
or UO_546 (O_546,N_10816,N_14155);
and UO_547 (O_547,N_13395,N_13254);
nor UO_548 (O_548,N_13402,N_10334);
or UO_549 (O_549,N_10446,N_10010);
nand UO_550 (O_550,N_10031,N_14797);
nand UO_551 (O_551,N_11731,N_12476);
nor UO_552 (O_552,N_11399,N_13025);
or UO_553 (O_553,N_11593,N_14620);
nor UO_554 (O_554,N_12323,N_14156);
and UO_555 (O_555,N_11227,N_10560);
nor UO_556 (O_556,N_13586,N_14870);
and UO_557 (O_557,N_14569,N_12806);
or UO_558 (O_558,N_12977,N_12973);
nor UO_559 (O_559,N_13466,N_10186);
nand UO_560 (O_560,N_14759,N_13361);
nand UO_561 (O_561,N_11648,N_11427);
nor UO_562 (O_562,N_10543,N_11622);
and UO_563 (O_563,N_13481,N_14904);
nand UO_564 (O_564,N_11683,N_11737);
or UO_565 (O_565,N_10354,N_12002);
or UO_566 (O_566,N_13902,N_11858);
nor UO_567 (O_567,N_12217,N_12051);
xor UO_568 (O_568,N_14999,N_11373);
xor UO_569 (O_569,N_13646,N_14586);
or UO_570 (O_570,N_11423,N_12750);
nor UO_571 (O_571,N_11704,N_10202);
nor UO_572 (O_572,N_13692,N_13752);
nand UO_573 (O_573,N_14984,N_13206);
nor UO_574 (O_574,N_10831,N_14942);
xnor UO_575 (O_575,N_13281,N_12702);
nor UO_576 (O_576,N_12649,N_12762);
or UO_577 (O_577,N_11882,N_14659);
xnor UO_578 (O_578,N_14510,N_10484);
nand UO_579 (O_579,N_12752,N_12618);
nand UO_580 (O_580,N_14950,N_13849);
and UO_581 (O_581,N_12619,N_11416);
nand UO_582 (O_582,N_13410,N_13196);
nand UO_583 (O_583,N_12927,N_10414);
nand UO_584 (O_584,N_13567,N_14994);
nor UO_585 (O_585,N_10468,N_10201);
nand UO_586 (O_586,N_10313,N_14693);
xor UO_587 (O_587,N_11092,N_13365);
and UO_588 (O_588,N_13265,N_12263);
xor UO_589 (O_589,N_13866,N_14876);
nor UO_590 (O_590,N_10462,N_13536);
and UO_591 (O_591,N_14896,N_12995);
nor UO_592 (O_592,N_13820,N_13612);
nor UO_593 (O_593,N_11756,N_12315);
and UO_594 (O_594,N_10643,N_13950);
and UO_595 (O_595,N_13057,N_14906);
nor UO_596 (O_596,N_14563,N_12769);
nand UO_597 (O_597,N_10732,N_14177);
or UO_598 (O_598,N_12168,N_10559);
or UO_599 (O_599,N_11179,N_12691);
nand UO_600 (O_600,N_10749,N_13641);
and UO_601 (O_601,N_12290,N_13024);
xor UO_602 (O_602,N_10502,N_10880);
nor UO_603 (O_603,N_12230,N_12623);
nor UO_604 (O_604,N_12566,N_11258);
nand UO_605 (O_605,N_11449,N_13255);
nor UO_606 (O_606,N_11702,N_13106);
nor UO_607 (O_607,N_13151,N_11305);
nand UO_608 (O_608,N_11352,N_11267);
or UO_609 (O_609,N_13537,N_12118);
and UO_610 (O_610,N_13337,N_10967);
and UO_611 (O_611,N_12457,N_13073);
xnor UO_612 (O_612,N_14403,N_10642);
or UO_613 (O_613,N_13504,N_14074);
nand UO_614 (O_614,N_14557,N_11356);
nand UO_615 (O_615,N_10357,N_12347);
nor UO_616 (O_616,N_12781,N_13529);
or UO_617 (O_617,N_14159,N_10493);
or UO_618 (O_618,N_12950,N_13202);
and UO_619 (O_619,N_12375,N_11062);
nor UO_620 (O_620,N_10434,N_14761);
or UO_621 (O_621,N_11969,N_12148);
and UO_622 (O_622,N_13735,N_12278);
nand UO_623 (O_623,N_11459,N_12399);
and UO_624 (O_624,N_13706,N_12832);
or UO_625 (O_625,N_14076,N_11972);
nor UO_626 (O_626,N_11907,N_11389);
or UO_627 (O_627,N_13355,N_14647);
or UO_628 (O_628,N_14088,N_11446);
nor UO_629 (O_629,N_11751,N_10973);
or UO_630 (O_630,N_14033,N_12622);
and UO_631 (O_631,N_10604,N_10640);
and UO_632 (O_632,N_10685,N_12226);
or UO_633 (O_633,N_13449,N_13097);
or UO_634 (O_634,N_11575,N_11722);
nor UO_635 (O_635,N_11529,N_11844);
or UO_636 (O_636,N_13519,N_10137);
xnor UO_637 (O_637,N_11266,N_11750);
or UO_638 (O_638,N_13614,N_12087);
nand UO_639 (O_639,N_12265,N_12819);
and UO_640 (O_640,N_11108,N_13032);
nand UO_641 (O_641,N_10891,N_11620);
nor UO_642 (O_642,N_10072,N_11597);
xnor UO_643 (O_643,N_10976,N_14457);
nand UO_644 (O_644,N_14639,N_12305);
nor UO_645 (O_645,N_12153,N_12177);
and UO_646 (O_646,N_12591,N_10601);
nand UO_647 (O_647,N_14402,N_10963);
xor UO_648 (O_648,N_13451,N_11214);
nand UO_649 (O_649,N_10847,N_14388);
nor UO_650 (O_650,N_11205,N_13145);
and UO_651 (O_651,N_10972,N_13990);
or UO_652 (O_652,N_14478,N_11787);
or UO_653 (O_653,N_12045,N_14089);
nor UO_654 (O_654,N_11649,N_12851);
or UO_655 (O_655,N_14658,N_11494);
or UO_656 (O_656,N_14381,N_11590);
nor UO_657 (O_657,N_14123,N_10351);
and UO_658 (O_658,N_10695,N_12339);
xor UO_659 (O_659,N_10964,N_14180);
nand UO_660 (O_660,N_14973,N_10266);
or UO_661 (O_661,N_10244,N_11628);
and UO_662 (O_662,N_14561,N_14489);
nor UO_663 (O_663,N_12685,N_12039);
or UO_664 (O_664,N_14231,N_13994);
or UO_665 (O_665,N_12483,N_10193);
or UO_666 (O_666,N_13442,N_11768);
and UO_667 (O_667,N_11746,N_12981);
nor UO_668 (O_668,N_13030,N_12174);
or UO_669 (O_669,N_14677,N_12557);
or UO_670 (O_670,N_10935,N_13541);
or UO_671 (O_671,N_12756,N_10843);
nor UO_672 (O_672,N_14015,N_12687);
or UO_673 (O_673,N_11438,N_10687);
nor UO_674 (O_674,N_14087,N_14474);
xor UO_675 (O_675,N_10171,N_13784);
nand UO_676 (O_676,N_14784,N_13705);
nor UO_677 (O_677,N_14841,N_12164);
nor UO_678 (O_678,N_10725,N_10549);
nor UO_679 (O_679,N_12333,N_13894);
xnor UO_680 (O_680,N_10004,N_11663);
or UO_681 (O_681,N_10547,N_10706);
xnor UO_682 (O_682,N_10520,N_14258);
and UO_683 (O_683,N_14486,N_11024);
nand UO_684 (O_684,N_14392,N_10260);
and UO_685 (O_685,N_12968,N_10365);
nand UO_686 (O_686,N_11028,N_11687);
or UO_687 (O_687,N_12712,N_14121);
nand UO_688 (O_688,N_11672,N_10436);
or UO_689 (O_689,N_12247,N_11630);
or UO_690 (O_690,N_11341,N_11698);
or UO_691 (O_691,N_10832,N_12737);
nand UO_692 (O_692,N_10721,N_12852);
and UO_693 (O_693,N_10488,N_14412);
and UO_694 (O_694,N_11334,N_10070);
and UO_695 (O_695,N_10983,N_13189);
or UO_696 (O_696,N_14259,N_12239);
and UO_697 (O_697,N_10043,N_12206);
nand UO_698 (O_698,N_14396,N_12648);
and UO_699 (O_699,N_13863,N_12517);
and UO_700 (O_700,N_12301,N_12043);
or UO_701 (O_701,N_10968,N_13205);
or UO_702 (O_702,N_10132,N_14038);
and UO_703 (O_703,N_10965,N_10677);
xnor UO_704 (O_704,N_11131,N_13808);
and UO_705 (O_705,N_13630,N_12590);
and UO_706 (O_706,N_13470,N_14166);
xnor UO_707 (O_707,N_14562,N_12035);
nand UO_708 (O_708,N_13569,N_10168);
nor UO_709 (O_709,N_12836,N_11551);
nand UO_710 (O_710,N_11547,N_13417);
nand UO_711 (O_711,N_10353,N_11272);
nor UO_712 (O_712,N_10349,N_13062);
nand UO_713 (O_713,N_10743,N_12365);
and UO_714 (O_714,N_11845,N_12720);
or UO_715 (O_715,N_12407,N_11465);
and UO_716 (O_716,N_11041,N_11791);
or UO_717 (O_717,N_11187,N_12598);
and UO_718 (O_718,N_13996,N_12386);
or UO_719 (O_719,N_11143,N_14720);
and UO_720 (O_720,N_13662,N_13809);
nand UO_721 (O_721,N_14105,N_11417);
and UO_722 (O_722,N_12154,N_12746);
and UO_723 (O_723,N_10111,N_11933);
and UO_724 (O_724,N_14708,N_14173);
and UO_725 (O_725,N_12482,N_10405);
xnor UO_726 (O_726,N_14473,N_12149);
or UO_727 (O_727,N_14433,N_10407);
or UO_728 (O_728,N_14083,N_11724);
nor UO_729 (O_729,N_10491,N_13445);
nand UO_730 (O_730,N_12546,N_12088);
xor UO_731 (O_731,N_14998,N_14188);
nand UO_732 (O_732,N_12447,N_10852);
nor UO_733 (O_733,N_13578,N_12291);
nor UO_734 (O_734,N_13724,N_13964);
and UO_735 (O_735,N_11684,N_13572);
nor UO_736 (O_736,N_14148,N_14235);
nand UO_737 (O_737,N_14077,N_12768);
nor UO_738 (O_738,N_13733,N_11743);
nand UO_739 (O_739,N_10054,N_11874);
nor UO_740 (O_740,N_11098,N_14376);
or UO_741 (O_741,N_12698,N_13939);
or UO_742 (O_742,N_14498,N_10389);
nand UO_743 (O_743,N_13198,N_14441);
and UO_744 (O_744,N_12141,N_11318);
nand UO_745 (O_745,N_14366,N_14108);
nand UO_746 (O_746,N_13907,N_13244);
nor UO_747 (O_747,N_10791,N_14262);
and UO_748 (O_748,N_14572,N_14622);
xor UO_749 (O_749,N_14216,N_14280);
nor UO_750 (O_750,N_12695,N_13419);
or UO_751 (O_751,N_12258,N_10722);
xnor UO_752 (O_752,N_10089,N_12974);
and UO_753 (O_753,N_12533,N_10384);
nor UO_754 (O_754,N_11790,N_13644);
nor UO_755 (O_755,N_12863,N_10071);
nor UO_756 (O_756,N_14046,N_10390);
nand UO_757 (O_757,N_11894,N_10368);
and UO_758 (O_758,N_13657,N_10918);
nand UO_759 (O_759,N_13949,N_10617);
nor UO_760 (O_760,N_12610,N_13343);
nor UO_761 (O_761,N_14277,N_11366);
nand UO_762 (O_762,N_12540,N_14414);
and UO_763 (O_763,N_14005,N_14451);
xnor UO_764 (O_764,N_11035,N_13262);
nand UO_765 (O_765,N_10782,N_13505);
nor UO_766 (O_766,N_10180,N_10977);
nand UO_767 (O_767,N_13363,N_11518);
nor UO_768 (O_768,N_11125,N_12952);
and UO_769 (O_769,N_12853,N_12397);
and UO_770 (O_770,N_14643,N_13885);
or UO_771 (O_771,N_11403,N_11625);
or UO_772 (O_772,N_14919,N_13273);
and UO_773 (O_773,N_13986,N_12234);
nor UO_774 (O_774,N_12733,N_10342);
nand UO_775 (O_775,N_14589,N_10768);
or UO_776 (O_776,N_13975,N_12890);
or UO_777 (O_777,N_14574,N_14090);
nor UO_778 (O_778,N_12257,N_12731);
nor UO_779 (O_779,N_10786,N_14684);
nor UO_780 (O_780,N_14255,N_14107);
and UO_781 (O_781,N_14554,N_14955);
nand UO_782 (O_782,N_13227,N_10416);
or UO_783 (O_783,N_11508,N_12932);
nand UO_784 (O_784,N_12165,N_13714);
and UO_785 (O_785,N_11650,N_10837);
nor UO_786 (O_786,N_12656,N_14931);
nand UO_787 (O_787,N_13593,N_13045);
and UO_788 (O_788,N_13081,N_12972);
nand UO_789 (O_789,N_11237,N_12469);
and UO_790 (O_790,N_10413,N_13352);
nand UO_791 (O_791,N_13796,N_13877);
nor UO_792 (O_792,N_12359,N_14646);
or UO_793 (O_793,N_11218,N_10017);
or UO_794 (O_794,N_12889,N_14694);
or UO_795 (O_795,N_13085,N_12223);
nor UO_796 (O_796,N_13498,N_12499);
nor UO_797 (O_797,N_12281,N_11928);
or UO_798 (O_798,N_12381,N_11461);
and UO_799 (O_799,N_10739,N_11848);
and UO_800 (O_800,N_12495,N_12140);
xor UO_801 (O_801,N_11813,N_13016);
nand UO_802 (O_802,N_14075,N_14615);
or UO_803 (O_803,N_13642,N_10865);
and UO_804 (O_804,N_10093,N_12349);
nand UO_805 (O_805,N_14908,N_13354);
or UO_806 (O_806,N_10803,N_11729);
nand UO_807 (O_807,N_10068,N_10297);
nand UO_808 (O_808,N_14706,N_12370);
or UO_809 (O_809,N_12021,N_11554);
or UO_810 (O_810,N_12772,N_10321);
or UO_811 (O_811,N_12459,N_14273);
nand UO_812 (O_812,N_10856,N_11524);
nor UO_813 (O_813,N_10758,N_10815);
or UO_814 (O_814,N_12547,N_13302);
or UO_815 (O_815,N_13125,N_14028);
and UO_816 (O_816,N_11451,N_14295);
or UO_817 (O_817,N_13523,N_13055);
nor UO_818 (O_818,N_14838,N_13269);
nand UO_819 (O_819,N_14338,N_13454);
nand UO_820 (O_820,N_10754,N_14689);
xor UO_821 (O_821,N_11689,N_10221);
or UO_822 (O_822,N_11760,N_11569);
nor UO_823 (O_823,N_14873,N_13663);
nand UO_824 (O_824,N_12843,N_13422);
nand UO_825 (O_825,N_10930,N_12470);
and UO_826 (O_826,N_10433,N_13576);
nand UO_827 (O_827,N_13698,N_13702);
or UO_828 (O_828,N_13192,N_14869);
nand UO_829 (O_829,N_10781,N_14347);
or UO_830 (O_830,N_13156,N_13717);
or UO_831 (O_831,N_10388,N_11031);
nor UO_832 (O_832,N_14359,N_12894);
xor UO_833 (O_833,N_13707,N_12207);
nand UO_834 (O_834,N_11231,N_14198);
nand UO_835 (O_835,N_10467,N_12721);
nor UO_836 (O_836,N_12689,N_10308);
or UO_837 (O_837,N_13123,N_12196);
nand UO_838 (O_838,N_14490,N_12526);
and UO_839 (O_839,N_10265,N_11050);
and UO_840 (O_840,N_11932,N_12235);
nand UO_841 (O_841,N_11772,N_12049);
nand UO_842 (O_842,N_14055,N_10341);
xnor UO_843 (O_843,N_12510,N_10098);
or UO_844 (O_844,N_11701,N_11299);
nor UO_845 (O_845,N_12037,N_11747);
and UO_846 (O_846,N_11901,N_11849);
and UO_847 (O_847,N_12061,N_14945);
and UO_848 (O_848,N_13729,N_12751);
and UO_849 (O_849,N_12003,N_10921);
and UO_850 (O_850,N_11157,N_14161);
and UO_851 (O_851,N_12286,N_11981);
xnor UO_852 (O_852,N_10567,N_10887);
nor UO_853 (O_853,N_13587,N_10412);
and UO_854 (O_854,N_10049,N_13040);
or UO_855 (O_855,N_10944,N_12074);
and UO_856 (O_856,N_11347,N_11588);
xor UO_857 (O_857,N_10204,N_10296);
nand UO_858 (O_858,N_14898,N_10629);
or UO_859 (O_859,N_10443,N_10147);
or UO_860 (O_860,N_12861,N_13946);
nor UO_861 (O_861,N_10470,N_10387);
nand UO_862 (O_862,N_12396,N_14099);
nor UO_863 (O_863,N_10788,N_10938);
and UO_864 (O_864,N_14290,N_13595);
or UO_865 (O_865,N_12210,N_12194);
nand UO_866 (O_866,N_11837,N_14261);
and UO_867 (O_867,N_13691,N_14946);
or UO_868 (O_868,N_14024,N_12529);
or UO_869 (O_869,N_13109,N_10810);
or UO_870 (O_870,N_12355,N_12117);
nor UO_871 (O_871,N_10899,N_11621);
nor UO_872 (O_872,N_13756,N_12914);
or UO_873 (O_873,N_11113,N_14567);
nand UO_874 (O_874,N_14456,N_10838);
xnor UO_875 (O_875,N_14820,N_10867);
nand UO_876 (O_876,N_14426,N_10663);
or UO_877 (O_877,N_13178,N_10120);
nand UO_878 (O_878,N_11225,N_11442);
and UO_879 (O_879,N_13479,N_12371);
xor UO_880 (O_880,N_10233,N_10316);
nor UO_881 (O_881,N_12075,N_14411);
and UO_882 (O_882,N_11159,N_14782);
xor UO_883 (O_883,N_10474,N_11063);
xor UO_884 (O_884,N_12523,N_11914);
nor UO_885 (O_885,N_14141,N_13090);
nor UO_886 (O_886,N_14846,N_11696);
xnor UO_887 (O_887,N_12745,N_14149);
xor UO_888 (O_888,N_10650,N_10822);
or UO_889 (O_889,N_11732,N_14997);
xor UO_890 (O_890,N_14673,N_10255);
nand UO_891 (O_891,N_14250,N_12336);
nor UO_892 (O_892,N_11380,N_11652);
or UO_893 (O_893,N_13393,N_11434);
or UO_894 (O_894,N_13455,N_14783);
and UO_895 (O_895,N_13407,N_14187);
nor UO_896 (O_896,N_11532,N_14296);
nand UO_897 (O_897,N_13276,N_10409);
and UO_898 (O_898,N_10391,N_12693);
nor UO_899 (O_899,N_14110,N_11864);
and UO_900 (O_900,N_11311,N_14472);
xnor UO_901 (O_901,N_10612,N_12360);
nand UO_902 (O_902,N_11514,N_11631);
nor UO_903 (O_903,N_11485,N_12858);
nand UO_904 (O_904,N_12172,N_11456);
nor UO_905 (O_905,N_12801,N_11585);
or UO_906 (O_906,N_12569,N_12595);
nor UO_907 (O_907,N_13357,N_13604);
nor UO_908 (O_908,N_13742,N_12446);
and UO_909 (O_909,N_12160,N_11985);
nor UO_910 (O_910,N_13530,N_13335);
nand UO_911 (O_911,N_13666,N_10129);
and UO_912 (O_912,N_11633,N_12617);
or UO_913 (O_913,N_12324,N_13688);
nor UO_914 (O_914,N_11735,N_13824);
nand UO_915 (O_915,N_11293,N_13921);
nor UO_916 (O_916,N_12451,N_12747);
or UO_917 (O_917,N_13825,N_10648);
nor UO_918 (O_918,N_14535,N_13471);
or UO_919 (O_919,N_12092,N_13128);
or UO_920 (O_920,N_14722,N_10773);
and UO_921 (O_921,N_13397,N_12085);
and UO_922 (O_922,N_11823,N_11137);
and UO_923 (O_923,N_10932,N_12631);
nor UO_924 (O_924,N_12025,N_13372);
nand UO_925 (O_925,N_13677,N_10295);
or UO_926 (O_926,N_13862,N_13403);
and UO_927 (O_927,N_13597,N_11466);
nor UO_928 (O_928,N_13887,N_12478);
nand UO_929 (O_929,N_11666,N_12115);
or UO_930 (O_930,N_13672,N_14390);
nor UO_931 (O_931,N_11245,N_14237);
or UO_932 (O_932,N_14415,N_11079);
or UO_933 (O_933,N_12101,N_14097);
nand UO_934 (O_934,N_14463,N_14668);
nand UO_935 (O_935,N_14365,N_13884);
nor UO_936 (O_936,N_14550,N_10085);
or UO_937 (O_937,N_13427,N_12222);
nand UO_938 (O_938,N_12956,N_11773);
or UO_939 (O_939,N_11548,N_14692);
and UO_940 (O_940,N_12855,N_14186);
or UO_941 (O_941,N_12132,N_11963);
nor UO_942 (O_942,N_10198,N_13444);
and UO_943 (O_943,N_13927,N_12609);
or UO_944 (O_944,N_10919,N_10893);
nand UO_945 (O_945,N_11022,N_11616);
or UO_946 (O_946,N_11934,N_13075);
and UO_947 (O_947,N_10206,N_11838);
or UO_948 (O_948,N_13771,N_10539);
nor UO_949 (O_949,N_12442,N_14147);
nand UO_950 (O_950,N_14967,N_14298);
nor UO_951 (O_951,N_13873,N_13275);
nand UO_952 (O_952,N_14360,N_12650);
nand UO_953 (O_953,N_13366,N_10273);
nor UO_954 (O_954,N_14393,N_12139);
xnor UO_955 (O_955,N_12325,N_10702);
or UO_956 (O_956,N_10544,N_11574);
xor UO_957 (O_957,N_13344,N_11719);
or UO_958 (O_958,N_11873,N_12891);
nand UO_959 (O_959,N_10302,N_10717);
nor UO_960 (O_960,N_13240,N_10197);
xnor UO_961 (O_961,N_13708,N_12965);
or UO_962 (O_962,N_10842,N_14763);
or UO_963 (O_963,N_14454,N_11155);
nor UO_964 (O_964,N_13048,N_10113);
nand UO_965 (O_965,N_13573,N_14172);
nand UO_966 (O_966,N_13001,N_11664);
nand UO_967 (O_967,N_10649,N_10286);
xnor UO_968 (O_968,N_10811,N_11609);
nand UO_969 (O_969,N_12108,N_12093);
nand UO_970 (O_970,N_14760,N_10460);
or UO_971 (O_971,N_14284,N_10764);
nand UO_972 (O_972,N_14894,N_10418);
nand UO_973 (O_973,N_14531,N_12391);
and UO_974 (O_974,N_10913,N_11431);
nand UO_975 (O_975,N_10406,N_10904);
nor UO_976 (O_976,N_14021,N_14625);
nand UO_977 (O_977,N_13711,N_14913);
nor UO_978 (O_978,N_10680,N_10438);
or UO_979 (O_979,N_10595,N_10257);
or UO_980 (O_980,N_11923,N_11742);
nand UO_981 (O_981,N_10114,N_11879);
nor UO_982 (O_982,N_11428,N_14522);
nand UO_983 (O_983,N_13214,N_13525);
xnor UO_984 (O_984,N_12340,N_13845);
nor UO_985 (O_985,N_10929,N_12636);
and UO_986 (O_986,N_13058,N_11089);
nand UO_987 (O_987,N_12434,N_12272);
and UO_988 (O_988,N_13494,N_12714);
nand UO_989 (O_989,N_12279,N_13485);
or UO_990 (O_990,N_10960,N_13230);
and UO_991 (O_991,N_12137,N_10735);
and UO_992 (O_992,N_11618,N_12030);
nor UO_993 (O_993,N_13600,N_12729);
or UO_994 (O_994,N_14662,N_11419);
nor UO_995 (O_995,N_14638,N_13457);
or UO_996 (O_996,N_11128,N_11275);
or UO_997 (O_997,N_10699,N_13266);
nand UO_998 (O_998,N_11700,N_10379);
nand UO_999 (O_999,N_10107,N_13472);
nor UO_1000 (O_1000,N_14408,N_13703);
nor UO_1001 (O_1001,N_13533,N_10894);
and UO_1002 (O_1002,N_11101,N_14368);
nand UO_1003 (O_1003,N_11759,N_11232);
or UO_1004 (O_1004,N_10675,N_12332);
nor UO_1005 (O_1005,N_14125,N_14060);
nor UO_1006 (O_1006,N_11484,N_10827);
nor UO_1007 (O_1007,N_14380,N_11036);
and UO_1008 (O_1008,N_12632,N_10799);
xor UO_1009 (O_1009,N_11328,N_10660);
or UO_1010 (O_1010,N_14963,N_11080);
or UO_1011 (O_1011,N_10726,N_11019);
nor UO_1012 (O_1012,N_13141,N_11961);
nand UO_1013 (O_1013,N_10746,N_14828);
nor UO_1014 (O_1014,N_10651,N_12681);
nor UO_1015 (O_1015,N_14022,N_10298);
or UO_1016 (O_1016,N_10326,N_13580);
xnor UO_1017 (O_1017,N_11002,N_14297);
and UO_1018 (O_1018,N_13446,N_12380);
nand UO_1019 (O_1019,N_10018,N_13913);
or UO_1020 (O_1020,N_14978,N_10902);
xor UO_1021 (O_1021,N_12966,N_13633);
or UO_1022 (O_1022,N_12320,N_12993);
nor UO_1023 (O_1023,N_14627,N_14318);
xnor UO_1024 (O_1024,N_13546,N_10347);
and UO_1025 (O_1025,N_11114,N_13199);
and UO_1026 (O_1026,N_10664,N_13369);
nand UO_1027 (O_1027,N_12248,N_13841);
nand UO_1028 (O_1028,N_11271,N_13903);
and UO_1029 (O_1029,N_14384,N_12472);
nand UO_1030 (O_1030,N_10194,N_10632);
xnor UO_1031 (O_1031,N_13810,N_14354);
or UO_1032 (O_1032,N_10970,N_11851);
nand UO_1033 (O_1033,N_10745,N_12484);
or UO_1034 (O_1034,N_13243,N_10319);
and UO_1035 (O_1035,N_12097,N_10969);
nor UO_1036 (O_1036,N_10396,N_14996);
nand UO_1037 (O_1037,N_11843,N_11546);
xor UO_1038 (O_1038,N_12348,N_11993);
or UO_1039 (O_1039,N_10482,N_14619);
nor UO_1040 (O_1040,N_14267,N_14100);
nand UO_1041 (O_1041,N_12006,N_14045);
or UO_1042 (O_1042,N_12765,N_10403);
and UO_1043 (O_1043,N_13476,N_11803);
or UO_1044 (O_1044,N_11612,N_11639);
xnor UO_1045 (O_1045,N_11185,N_10839);
nand UO_1046 (O_1046,N_14182,N_12020);
nor UO_1047 (O_1047,N_10140,N_12233);
nand UO_1048 (O_1048,N_11206,N_11368);
nor UO_1049 (O_1049,N_14208,N_12245);
nand UO_1050 (O_1050,N_13356,N_12543);
or UO_1051 (O_1051,N_14407,N_13060);
or UO_1052 (O_1052,N_10836,N_12377);
nor UO_1053 (O_1053,N_10619,N_12424);
or UO_1054 (O_1054,N_10095,N_10498);
and UO_1055 (O_1055,N_14302,N_10626);
nor UO_1056 (O_1056,N_11498,N_11394);
nor UO_1057 (O_1057,N_12612,N_12053);
or UO_1058 (O_1058,N_14621,N_10506);
and UO_1059 (O_1059,N_10728,N_13367);
or UO_1060 (O_1060,N_10937,N_13988);
and UO_1061 (O_1061,N_14493,N_10243);
xnor UO_1062 (O_1062,N_13306,N_14488);
and UO_1063 (O_1063,N_12096,N_14481);
nor UO_1064 (O_1064,N_11884,N_13326);
or UO_1065 (O_1065,N_12735,N_10399);
nand UO_1066 (O_1066,N_10235,N_11207);
nor UO_1067 (O_1067,N_14477,N_11327);
and UO_1068 (O_1068,N_13005,N_11887);
and UO_1069 (O_1069,N_13336,N_10122);
or UO_1070 (O_1070,N_14006,N_10485);
and UO_1071 (O_1071,N_13547,N_13645);
and UO_1072 (O_1072,N_10218,N_12103);
xor UO_1073 (O_1073,N_14711,N_11365);
nand UO_1074 (O_1074,N_13579,N_13971);
or UO_1075 (O_1075,N_10982,N_14479);
nor UO_1076 (O_1076,N_12357,N_11306);
xnor UO_1077 (O_1077,N_13095,N_14035);
nor UO_1078 (O_1078,N_10614,N_14826);
or UO_1079 (O_1079,N_14467,N_13041);
and UO_1080 (O_1080,N_14184,N_11571);
and UO_1081 (O_1081,N_13375,N_12213);
nand UO_1082 (O_1082,N_10411,N_13228);
nand UO_1083 (O_1083,N_14923,N_12338);
nand UO_1084 (O_1084,N_13101,N_11075);
and UO_1085 (O_1085,N_10009,N_12924);
and UO_1086 (O_1086,N_12031,N_13969);
nor UO_1087 (O_1087,N_11457,N_13008);
nor UO_1088 (O_1088,N_10670,N_14213);
nor UO_1089 (O_1089,N_13916,N_12283);
nor UO_1090 (O_1090,N_12630,N_11273);
nor UO_1091 (O_1091,N_14026,N_11697);
xor UO_1092 (O_1092,N_13776,N_14672);
nor UO_1093 (O_1093,N_13966,N_11138);
and UO_1094 (O_1094,N_12778,N_14534);
and UO_1095 (O_1095,N_10580,N_14103);
nand UO_1096 (O_1096,N_12664,N_12898);
nor UO_1097 (O_1097,N_14803,N_14092);
nor UO_1098 (O_1098,N_12269,N_11082);
or UO_1099 (O_1099,N_12331,N_11572);
or UO_1100 (O_1100,N_13249,N_10553);
and UO_1101 (O_1101,N_14951,N_11000);
and UO_1102 (O_1102,N_14583,N_14549);
or UO_1103 (O_1103,N_13867,N_14835);
or UO_1104 (O_1104,N_12524,N_12112);
and UO_1105 (O_1105,N_12589,N_10356);
nand UO_1106 (O_1106,N_12684,N_14515);
xor UO_1107 (O_1107,N_10710,N_10790);
or UO_1108 (O_1108,N_11661,N_10271);
xnor UO_1109 (O_1109,N_10562,N_11023);
nor UO_1110 (O_1110,N_13528,N_11383);
nor UO_1111 (O_1111,N_14336,N_10082);
xnor UO_1112 (O_1112,N_13129,N_13753);
nand UO_1113 (O_1113,N_14313,N_11720);
nand UO_1114 (O_1114,N_14160,N_14806);
or UO_1115 (O_1115,N_11243,N_10163);
nand UO_1116 (O_1116,N_14238,N_10157);
xor UO_1117 (O_1117,N_14323,N_14687);
or UO_1118 (O_1118,N_12184,N_12883);
nand UO_1119 (O_1119,N_12046,N_10729);
and UO_1120 (O_1120,N_10339,N_13909);
nand UO_1121 (O_1121,N_10795,N_13891);
nor UO_1122 (O_1122,N_10731,N_12805);
and UO_1123 (O_1123,N_14361,N_14265);
or UO_1124 (O_1124,N_10676,N_13035);
nand UO_1125 (O_1125,N_10055,N_12818);
nor UO_1126 (O_1126,N_10694,N_11348);
and UO_1127 (O_1127,N_13831,N_14281);
xnor UO_1128 (O_1128,N_11978,N_13607);
or UO_1129 (O_1129,N_12710,N_11676);
or UO_1130 (O_1130,N_14269,N_10027);
nor UO_1131 (O_1131,N_11091,N_14608);
nand UO_1132 (O_1132,N_13436,N_13084);
or UO_1133 (O_1133,N_12044,N_11797);
xnor UO_1134 (O_1134,N_12421,N_11391);
nor UO_1135 (O_1135,N_10352,N_14176);
xor UO_1136 (O_1136,N_10426,N_13314);
or UO_1137 (O_1137,N_11867,N_10691);
nand UO_1138 (O_1138,N_10134,N_10709);
nor UO_1139 (O_1139,N_11801,N_13984);
nor UO_1140 (O_1140,N_13787,N_11541);
nand UO_1141 (O_1141,N_10370,N_10112);
nor UO_1142 (O_1142,N_11865,N_10951);
nand UO_1143 (O_1143,N_13443,N_13467);
and UO_1144 (O_1144,N_11396,N_12537);
and UO_1145 (O_1145,N_12455,N_12067);
or UO_1146 (O_1146,N_10727,N_11288);
nand UO_1147 (O_1147,N_14069,N_12748);
nor UO_1148 (O_1148,N_13676,N_10185);
xnor UO_1149 (O_1149,N_11469,N_14226);
and UO_1150 (O_1150,N_12054,N_14439);
xor UO_1151 (O_1151,N_10410,N_10160);
nor UO_1152 (O_1152,N_10569,N_11286);
xnor UO_1153 (O_1153,N_14773,N_13795);
xor UO_1154 (O_1154,N_11714,N_14821);
and UO_1155 (O_1155,N_11986,N_13295);
nand UO_1156 (O_1156,N_14230,N_11167);
nor UO_1157 (O_1157,N_10187,N_11265);
nor UO_1158 (O_1158,N_14771,N_13782);
and UO_1159 (O_1159,N_14750,N_14733);
nor UO_1160 (O_1160,N_11084,N_11796);
nor UO_1161 (O_1161,N_14174,N_13671);
and UO_1162 (O_1162,N_10578,N_12008);
nor UO_1163 (O_1163,N_11051,N_12220);
nand UO_1164 (O_1164,N_12953,N_13177);
and UO_1165 (O_1165,N_10269,N_12361);
and UO_1166 (O_1166,N_14893,N_11692);
nand UO_1167 (O_1167,N_12214,N_10824);
and UO_1168 (O_1168,N_12169,N_11890);
xor UO_1169 (O_1169,N_10280,N_10961);
nor UO_1170 (O_1170,N_13111,N_13895);
and UO_1171 (O_1171,N_10581,N_11730);
or UO_1172 (O_1172,N_14526,N_13020);
and UO_1173 (O_1173,N_10714,N_11414);
nor UO_1174 (O_1174,N_12627,N_10523);
or UO_1175 (O_1175,N_12433,N_13892);
or UO_1176 (O_1176,N_14153,N_13620);
and UO_1177 (O_1177,N_10404,N_11292);
nor UO_1178 (O_1178,N_10590,N_14539);
or UO_1179 (O_1179,N_12867,N_11120);
or UO_1180 (O_1180,N_14805,N_13998);
and UO_1181 (O_1181,N_13490,N_13901);
or UO_1182 (O_1182,N_14236,N_14399);
and UO_1183 (O_1183,N_12502,N_13802);
or UO_1184 (O_1184,N_11610,N_14398);
and UO_1185 (O_1185,N_12500,N_11379);
and UO_1186 (O_1186,N_13004,N_10380);
xor UO_1187 (O_1187,N_12560,N_11596);
xnor UO_1188 (O_1188,N_10329,N_11418);
and UO_1189 (O_1189,N_12302,N_11911);
and UO_1190 (O_1190,N_10708,N_12835);
or UO_1191 (O_1191,N_12460,N_14131);
and UO_1192 (O_1192,N_11710,N_11712);
nand UO_1193 (O_1193,N_14641,N_11789);
nand UO_1194 (O_1194,N_14240,N_10442);
nor UO_1195 (O_1195,N_12422,N_12507);
nand UO_1196 (O_1196,N_13693,N_13224);
nand UO_1197 (O_1197,N_14364,N_13772);
nand UO_1198 (O_1198,N_14678,N_14578);
or UO_1199 (O_1199,N_12019,N_11454);
nor UO_1200 (O_1200,N_10874,N_13911);
xor UO_1201 (O_1201,N_12452,N_10325);
nand UO_1202 (O_1202,N_10358,N_10439);
or UO_1203 (O_1203,N_14768,N_12170);
nor UO_1204 (O_1204,N_13305,N_10343);
or UO_1205 (O_1205,N_10978,N_14465);
and UO_1206 (O_1206,N_11889,N_14272);
and UO_1207 (O_1207,N_10674,N_10494);
nand UO_1208 (O_1208,N_14285,N_14847);
nor UO_1209 (O_1209,N_14143,N_12795);
and UO_1210 (O_1210,N_11678,N_13116);
and UO_1211 (O_1211,N_12145,N_10554);
or UO_1212 (O_1212,N_10597,N_11362);
nand UO_1213 (O_1213,N_11049,N_12034);
nand UO_1214 (O_1214,N_13563,N_10305);
or UO_1215 (O_1215,N_14599,N_13037);
nor UO_1216 (O_1216,N_14109,N_13387);
or UO_1217 (O_1217,N_12651,N_10825);
or UO_1218 (O_1218,N_12842,N_13798);
and UO_1219 (O_1219,N_10481,N_11384);
xor UO_1220 (O_1220,N_10991,N_14011);
or UO_1221 (O_1221,N_14749,N_12267);
and UO_1222 (O_1222,N_10751,N_14220);
nor UO_1223 (O_1223,N_13465,N_10497);
nand UO_1224 (O_1224,N_11346,N_13107);
nor UO_1225 (O_1225,N_12652,N_12982);
or UO_1226 (O_1226,N_13203,N_14765);
nor UO_1227 (O_1227,N_11855,N_10020);
or UO_1228 (O_1228,N_13461,N_11289);
nor UO_1229 (O_1229,N_11013,N_14221);
nand UO_1230 (O_1230,N_11558,N_10718);
or UO_1231 (O_1231,N_14104,N_13856);
or UO_1232 (O_1232,N_10184,N_14343);
nor UO_1233 (O_1233,N_14301,N_12764);
and UO_1234 (O_1234,N_12831,N_13613);
nor UO_1235 (O_1235,N_12018,N_12823);
or UO_1236 (O_1236,N_11398,N_14661);
and UO_1237 (O_1237,N_13340,N_13250);
and UO_1238 (O_1238,N_12284,N_12732);
or UO_1239 (O_1239,N_10117,N_10536);
or UO_1240 (O_1240,N_11240,N_12738);
nor UO_1241 (O_1241,N_11037,N_12107);
or UO_1242 (O_1242,N_12716,N_13204);
nor UO_1243 (O_1243,N_13594,N_12929);
nand UO_1244 (O_1244,N_11359,N_12800);
or UO_1245 (O_1245,N_14421,N_13687);
nand UO_1246 (O_1246,N_11405,N_13679);
nand UO_1247 (O_1247,N_10131,N_10254);
xor UO_1248 (O_1248,N_13709,N_13076);
and UO_1249 (O_1249,N_14949,N_12957);
xnor UO_1250 (O_1250,N_11162,N_12688);
or UO_1251 (O_1251,N_11651,N_12561);
and UO_1252 (O_1252,N_14371,N_10736);
and UO_1253 (O_1253,N_10275,N_10576);
or UO_1254 (O_1254,N_14519,N_13012);
nand UO_1255 (O_1255,N_14229,N_14189);
xnor UO_1256 (O_1256,N_12062,N_14940);
nand UO_1257 (O_1257,N_11875,N_11764);
nor UO_1258 (O_1258,N_13148,N_12987);
nand UO_1259 (O_1259,N_11636,N_13739);
nor UO_1260 (O_1260,N_10360,N_11594);
or UO_1261 (O_1261,N_13619,N_10457);
nand UO_1262 (O_1262,N_10311,N_13526);
nor UO_1263 (O_1263,N_11395,N_14726);
and UO_1264 (O_1264,N_12306,N_11464);
nor UO_1265 (O_1265,N_14755,N_11134);
and UO_1266 (O_1266,N_10033,N_10079);
nor UO_1267 (O_1267,N_10994,N_14241);
nor UO_1268 (O_1268,N_13922,N_10741);
and UO_1269 (O_1269,N_11263,N_12715);
nor UO_1270 (O_1270,N_10627,N_14513);
xnor UO_1271 (O_1271,N_12200,N_11130);
xor UO_1272 (O_1272,N_10588,N_10417);
and UO_1273 (O_1273,N_11509,N_13110);
xor UO_1274 (O_1274,N_12122,N_13428);
nor UO_1275 (O_1275,N_10756,N_10767);
nand UO_1276 (O_1276,N_14587,N_10900);
xor UO_1277 (O_1277,N_11827,N_13158);
or UO_1278 (O_1278,N_14112,N_11613);
or UO_1279 (O_1279,N_10364,N_14947);
nand UO_1280 (O_1280,N_13146,N_11429);
nand UO_1281 (O_1281,N_10335,N_14199);
or UO_1282 (O_1282,N_14328,N_11377);
nand UO_1283 (O_1283,N_11112,N_10783);
xnor UO_1284 (O_1284,N_14505,N_12404);
or UO_1285 (O_1285,N_12713,N_12920);
nor UO_1286 (O_1286,N_14880,N_13029);
nand UO_1287 (O_1287,N_14239,N_11755);
and UO_1288 (O_1288,N_13173,N_13694);
nor UO_1289 (O_1289,N_12352,N_11247);
and UO_1290 (O_1290,N_11007,N_13974);
and UO_1291 (O_1291,N_14552,N_11994);
xnor UO_1292 (O_1292,N_11337,N_11815);
xnor UO_1293 (O_1293,N_11513,N_10770);
nor UO_1294 (O_1294,N_13399,N_14362);
nor UO_1295 (O_1295,N_14400,N_13750);
xor UO_1296 (O_1296,N_13021,N_13304);
xor UO_1297 (O_1297,N_12188,N_10469);
nand UO_1298 (O_1298,N_11973,N_14145);
xnor UO_1299 (O_1299,N_10177,N_10858);
nand UO_1300 (O_1300,N_11172,N_14669);
and UO_1301 (O_1301,N_11153,N_11748);
xnor UO_1302 (O_1302,N_12445,N_13632);
nand UO_1303 (O_1303,N_12665,N_14725);
or UO_1304 (O_1304,N_12790,N_10582);
nand UO_1305 (O_1305,N_12944,N_11053);
or UO_1306 (O_1306,N_14469,N_14939);
nand UO_1307 (O_1307,N_14282,N_12882);
nand UO_1308 (O_1308,N_11988,N_13469);
or UO_1309 (O_1309,N_10164,N_13452);
nor UO_1310 (O_1310,N_14140,N_11948);
or UO_1311 (O_1311,N_14832,N_11121);
nor UO_1312 (O_1312,N_11627,N_12065);
nand UO_1313 (O_1313,N_14061,N_12942);
and UO_1314 (O_1314,N_11645,N_10323);
nor UO_1315 (O_1315,N_14442,N_14943);
xor UO_1316 (O_1316,N_14936,N_14953);
or UO_1317 (O_1317,N_11376,N_13848);
and UO_1318 (O_1318,N_11133,N_12862);
or UO_1319 (O_1319,N_12901,N_11983);
or UO_1320 (O_1320,N_11047,N_10013);
and UO_1321 (O_1321,N_10299,N_14101);
and UO_1322 (O_1322,N_12105,N_14690);
and UO_1323 (O_1323,N_14321,N_13229);
or UO_1324 (O_1324,N_11682,N_13690);
or UO_1325 (O_1325,N_10669,N_13282);
nor UO_1326 (O_1326,N_13322,N_12694);
and UO_1327 (O_1327,N_13298,N_11543);
nand UO_1328 (O_1328,N_11954,N_14082);
or UO_1329 (O_1329,N_14008,N_10143);
nand UO_1330 (O_1330,N_10432,N_14425);
nor UO_1331 (O_1331,N_11470,N_10427);
and UO_1332 (O_1332,N_14907,N_12461);
nor UO_1333 (O_1333,N_11432,N_10333);
nand UO_1334 (O_1334,N_13743,N_12419);
nor UO_1335 (O_1335,N_13348,N_10449);
nand UO_1336 (O_1336,N_12615,N_10546);
xor UO_1337 (O_1337,N_14367,N_12441);
and UO_1338 (O_1338,N_10152,N_10424);
and UO_1339 (O_1339,N_11372,N_11812);
nand UO_1340 (O_1340,N_10196,N_14317);
nand UO_1341 (O_1341,N_14329,N_14245);
nor UO_1342 (O_1342,N_13917,N_14196);
and UO_1343 (O_1343,N_11222,N_12440);
and UO_1344 (O_1344,N_14705,N_14508);
and UO_1345 (O_1345,N_13914,N_12318);
nand UO_1346 (O_1346,N_14885,N_13623);
and UO_1347 (O_1347,N_10156,N_10659);
nand UO_1348 (O_1348,N_10946,N_13826);
nand UO_1349 (O_1349,N_13477,N_13248);
nand UO_1350 (O_1350,N_13783,N_11413);
nor UO_1351 (O_1351,N_11944,N_10813);
and UO_1352 (O_1352,N_12449,N_11156);
and UO_1353 (O_1353,N_13575,N_10402);
xor UO_1354 (O_1354,N_12487,N_13200);
and UO_1355 (O_1355,N_12552,N_13736);
nand UO_1356 (O_1356,N_12211,N_12136);
or UO_1357 (O_1357,N_11880,N_13565);
xnor UO_1358 (O_1358,N_10304,N_11126);
nor UO_1359 (O_1359,N_13278,N_13006);
and UO_1360 (O_1360,N_11822,N_10884);
and UO_1361 (O_1361,N_11038,N_13667);
or UO_1362 (O_1362,N_14723,N_11147);
and UO_1363 (O_1363,N_13038,N_14445);
and UO_1364 (O_1364,N_13570,N_14232);
nand UO_1365 (O_1365,N_10277,N_14436);
or UO_1366 (O_1366,N_13731,N_14912);
xor UO_1367 (O_1367,N_12186,N_10139);
or UO_1368 (O_1368,N_10238,N_13234);
and UO_1369 (O_1369,N_11922,N_13910);
nor UO_1370 (O_1370,N_10090,N_14976);
and UO_1371 (O_1371,N_10678,N_14168);
xor UO_1372 (O_1372,N_12024,N_11421);
nor UO_1373 (O_1373,N_10508,N_10575);
xor UO_1374 (O_1374,N_13532,N_13120);
xor UO_1375 (O_1375,N_11783,N_14401);
and UO_1376 (O_1376,N_11681,N_14468);
or UO_1377 (O_1377,N_11071,N_11415);
or UO_1378 (O_1378,N_11280,N_12189);
nor UO_1379 (O_1379,N_14799,N_12865);
and UO_1380 (O_1380,N_10378,N_13303);
and UO_1381 (O_1381,N_11761,N_11754);
nand UO_1382 (O_1382,N_13589,N_12438);
nand UO_1383 (O_1383,N_13948,N_10450);
nand UO_1384 (O_1384,N_14043,N_12201);
or UO_1385 (O_1385,N_14150,N_12653);
nor UO_1386 (O_1386,N_13585,N_11516);
nor UO_1387 (O_1387,N_11669,N_10615);
or UO_1388 (O_1388,N_14611,N_10591);
xnor UO_1389 (O_1389,N_12129,N_13635);
nor UO_1390 (O_1390,N_10372,N_10538);
xor UO_1391 (O_1391,N_13500,N_11736);
or UO_1392 (O_1392,N_10577,N_12530);
nor UO_1393 (O_1393,N_14665,N_11805);
nor UO_1394 (O_1394,N_12892,N_12498);
and UO_1395 (O_1395,N_10376,N_12142);
nand UO_1396 (O_1396,N_10962,N_12599);
nand UO_1397 (O_1397,N_10056,N_10882);
nand UO_1398 (O_1398,N_13935,N_11408);
or UO_1399 (O_1399,N_12244,N_13670);
and UO_1400 (O_1400,N_14883,N_10256);
nor UO_1401 (O_1401,N_11888,N_13115);
and UO_1402 (O_1402,N_11758,N_12970);
or UO_1403 (O_1403,N_13919,N_11976);
and UO_1404 (O_1404,N_12366,N_11785);
nor UO_1405 (O_1405,N_14252,N_10819);
and UO_1406 (O_1406,N_14027,N_12098);
nor UO_1407 (O_1407,N_13521,N_13409);
and UO_1408 (O_1408,N_12329,N_14766);
nand UO_1409 (O_1409,N_11741,N_13941);
nor UO_1410 (O_1410,N_11191,N_12337);
xnor UO_1411 (O_1411,N_12000,N_10857);
nand UO_1412 (O_1412,N_10514,N_11006);
nand UO_1413 (O_1413,N_10928,N_11675);
nand UO_1414 (O_1414,N_12686,N_13223);
nand UO_1415 (O_1415,N_12555,N_11998);
and UO_1416 (O_1416,N_11307,N_13245);
or UO_1417 (O_1417,N_14724,N_10492);
xnor UO_1418 (O_1418,N_10314,N_14192);
and UO_1419 (O_1419,N_12570,N_11029);
or UO_1420 (O_1420,N_14902,N_12711);
and UO_1421 (O_1421,N_12467,N_13426);
and UO_1422 (O_1422,N_14553,N_13015);
xnor UO_1423 (O_1423,N_14093,N_10099);
nand UO_1424 (O_1424,N_11962,N_14903);
nor UO_1425 (O_1425,N_11811,N_14491);
nand UO_1426 (O_1426,N_10337,N_12979);
nand UO_1427 (O_1427,N_11242,N_12672);
or UO_1428 (O_1428,N_11184,N_11274);
and UO_1429 (O_1429,N_11883,N_11141);
and UO_1430 (O_1430,N_13686,N_14394);
nor UO_1431 (O_1431,N_11163,N_13153);
and UO_1432 (O_1432,N_11315,N_12308);
and UO_1433 (O_1433,N_10355,N_14987);
nor UO_1434 (O_1434,N_11668,N_13520);
and UO_1435 (O_1435,N_13817,N_14975);
nand UO_1436 (O_1436,N_12548,N_10381);
and UO_1437 (O_1437,N_14545,N_10579);
or UO_1438 (O_1438,N_14501,N_12551);
and UO_1439 (O_1439,N_12225,N_10889);
nand UO_1440 (O_1440,N_12564,N_11331);
or UO_1441 (O_1441,N_12933,N_12870);
xnor UO_1442 (O_1442,N_12812,N_10065);
and UO_1443 (O_1443,N_11515,N_11441);
xor UO_1444 (O_1444,N_14126,N_14036);
or UO_1445 (O_1445,N_14314,N_10914);
and UO_1446 (O_1446,N_10761,N_14339);
and UO_1447 (O_1447,N_13053,N_13768);
nand UO_1448 (O_1448,N_11281,N_10288);
nor UO_1449 (O_1449,N_10097,N_12978);
nor UO_1450 (O_1450,N_14736,N_14770);
or UO_1451 (O_1451,N_11066,N_14822);
nand UO_1452 (O_1452,N_14503,N_14283);
xor UO_1453 (O_1453,N_10270,N_10473);
nand UO_1454 (O_1454,N_13811,N_13838);
nand UO_1455 (O_1455,N_11381,N_10555);
xnor UO_1456 (O_1456,N_11321,N_10075);
nand UO_1457 (O_1457,N_12527,N_10153);
or UO_1458 (O_1458,N_11480,N_11956);
and UO_1459 (O_1459,N_12041,N_13068);
xnor UO_1460 (O_1460,N_11165,N_12287);
nand UO_1461 (O_1461,N_11656,N_10178);
nand UO_1462 (O_1462,N_14576,N_10060);
nor UO_1463 (O_1463,N_10076,N_13511);
and UO_1464 (O_1464,N_14207,N_12341);
nand UO_1465 (O_1465,N_14375,N_11784);
nor UO_1466 (O_1466,N_14502,N_11991);
and UO_1467 (O_1467,N_11995,N_11957);
nand UO_1468 (O_1468,N_13069,N_13785);
and UO_1469 (O_1469,N_10332,N_10102);
and UO_1470 (O_1470,N_12327,N_10639);
nor UO_1471 (O_1471,N_10780,N_11795);
or UO_1472 (O_1472,N_13315,N_13133);
or UO_1473 (O_1473,N_11074,N_11496);
xor UO_1474 (O_1474,N_14787,N_14178);
or UO_1475 (O_1475,N_11479,N_12249);
nand UO_1476 (O_1476,N_14887,N_13320);
or UO_1477 (O_1477,N_10127,N_11221);
nor UO_1478 (O_1478,N_13233,N_11624);
and UO_1479 (O_1479,N_14504,N_12519);
xnor UO_1480 (O_1480,N_13915,N_14596);
nand UO_1481 (O_1481,N_13617,N_10144);
or UO_1482 (O_1482,N_10224,N_10215);
or UO_1483 (O_1483,N_11695,N_10661);
or UO_1484 (O_1484,N_13764,N_12845);
or UO_1485 (O_1485,N_14895,N_12839);
nand UO_1486 (O_1486,N_14260,N_13951);
or UO_1487 (O_1487,N_14776,N_13124);
or UO_1488 (O_1488,N_13430,N_14877);
or UO_1489 (O_1489,N_12114,N_14679);
or UO_1490 (O_1490,N_12453,N_13967);
nand UO_1491 (O_1491,N_14054,N_14905);
or UO_1492 (O_1492,N_13019,N_12252);
or UO_1493 (O_1493,N_10734,N_12971);
nand UO_1494 (O_1494,N_14664,N_13247);
and UO_1495 (O_1495,N_13319,N_10529);
or UO_1496 (O_1496,N_10188,N_10309);
nand UO_1497 (O_1497,N_14696,N_13207);
nand UO_1498 (O_1498,N_10636,N_14699);
or UO_1499 (O_1499,N_13358,N_11333);
nand UO_1500 (O_1500,N_10023,N_14217);
nor UO_1501 (O_1501,N_14139,N_13308);
and UO_1502 (O_1502,N_13373,N_12846);
nand UO_1503 (O_1503,N_13169,N_13253);
nand UO_1504 (O_1504,N_12926,N_13049);
or UO_1505 (O_1505,N_11608,N_14119);
nand UO_1506 (O_1506,N_10565,N_10516);
nand UO_1507 (O_1507,N_13394,N_11282);
xnor UO_1508 (O_1508,N_13947,N_11564);
and UO_1509 (O_1509,N_11407,N_11659);
nand UO_1510 (O_1510,N_11685,N_12055);
nor UO_1511 (O_1511,N_13609,N_13079);
and UO_1512 (O_1512,N_11673,N_12109);
and UO_1513 (O_1513,N_10688,N_11570);
nand UO_1514 (O_1514,N_11367,N_10711);
and UO_1515 (O_1515,N_14315,N_13524);
and UO_1516 (O_1516,N_12817,N_14124);
nor UO_1517 (O_1517,N_10105,N_13871);
or UO_1518 (O_1518,N_12173,N_13596);
xnor UO_1519 (O_1519,N_13383,N_12849);
xor UO_1520 (O_1520,N_13093,N_11450);
or UO_1521 (O_1521,N_14146,N_12931);
nor UO_1522 (O_1522,N_11054,N_10686);
and UO_1523 (O_1523,N_12394,N_14914);
nor UO_1524 (O_1524,N_11606,N_12364);
nand UO_1525 (O_1525,N_11151,N_12481);
nor UO_1526 (O_1526,N_12620,N_10229);
and UO_1527 (O_1527,N_13618,N_10138);
and UO_1528 (O_1528,N_14337,N_14910);
and UO_1529 (O_1529,N_14034,N_11422);
xnor UO_1530 (O_1530,N_14565,N_13793);
nand UO_1531 (O_1531,N_11215,N_14453);
nand UO_1532 (O_1532,N_14449,N_14982);
nand UO_1533 (O_1533,N_11598,N_13003);
or UO_1534 (O_1534,N_12475,N_12616);
and UO_1535 (O_1535,N_11382,N_10747);
nor UO_1536 (O_1536,N_13333,N_13883);
nand UO_1537 (O_1537,N_13201,N_12884);
nand UO_1538 (O_1538,N_10274,N_13054);
xnor UO_1539 (O_1539,N_13564,N_14356);
or UO_1540 (O_1540,N_10863,N_12854);
and UO_1541 (O_1541,N_12949,N_12934);
nand UO_1542 (O_1542,N_10225,N_13458);
or UO_1543 (O_1543,N_14807,N_11313);
nor UO_1544 (O_1544,N_11478,N_12654);
nor UO_1545 (O_1545,N_10471,N_14102);
or UO_1546 (O_1546,N_10557,N_11999);
and UO_1547 (O_1547,N_13280,N_11816);
or UO_1548 (O_1548,N_13332,N_12730);
and UO_1549 (O_1549,N_12872,N_10109);
and UO_1550 (O_1550,N_11319,N_14927);
or UO_1551 (O_1551,N_14528,N_11160);
and UO_1552 (O_1552,N_14683,N_10623);
and UO_1553 (O_1553,N_12635,N_14195);
nor UO_1554 (O_1554,N_13341,N_11565);
nand UO_1555 (O_1555,N_10126,N_14158);
nand UO_1556 (O_1556,N_10245,N_12625);
xnor UO_1557 (O_1557,N_13963,N_14068);
nor UO_1558 (O_1558,N_11026,N_11345);
and UO_1559 (O_1559,N_12317,N_12992);
and UO_1560 (O_1560,N_11580,N_12271);
nand UO_1561 (O_1561,N_14532,N_10246);
nor UO_1562 (O_1562,N_10910,N_13571);
or UO_1563 (O_1563,N_14681,N_10907);
nand UO_1564 (O_1564,N_11005,N_14853);
xnor UO_1565 (O_1565,N_12869,N_12354);
and UO_1566 (O_1566,N_12350,N_11195);
nor UO_1567 (O_1567,N_11642,N_14911);
xor UO_1568 (O_1568,N_13956,N_11780);
and UO_1569 (O_1569,N_10208,N_13284);
or UO_1570 (O_1570,N_11629,N_13722);
nor UO_1571 (O_1571,N_13241,N_10564);
nor UO_1572 (O_1572,N_13379,N_13592);
or UO_1573 (O_1573,N_14031,N_11297);
nand UO_1574 (O_1574,N_10558,N_11110);
and UO_1575 (O_1575,N_11193,N_10817);
and UO_1576 (O_1576,N_11964,N_11204);
or UO_1577 (O_1577,N_10007,N_10988);
nor UO_1578 (O_1578,N_11576,N_12069);
nand UO_1579 (O_1579,N_10833,N_12744);
and UO_1580 (O_1580,N_13957,N_12701);
nand UO_1581 (O_1581,N_13412,N_11940);
and UO_1582 (O_1582,N_11338,N_14455);
nor UO_1583 (O_1583,N_10006,N_10697);
or UO_1584 (O_1584,N_12866,N_13113);
nand UO_1585 (O_1585,N_12868,N_13918);
xnor UO_1586 (O_1586,N_14023,N_13629);
nor UO_1587 (O_1587,N_10517,N_10814);
or UO_1588 (O_1588,N_10252,N_10258);
and UO_1589 (O_1589,N_11899,N_12885);
nor UO_1590 (O_1590,N_11638,N_11721);
or UO_1591 (O_1591,N_14962,N_12004);
or UO_1592 (O_1592,N_12400,N_12639);
xor UO_1593 (O_1593,N_11500,N_12629);
nand UO_1594 (O_1594,N_14127,N_11686);
and UO_1595 (O_1595,N_13163,N_12760);
nand UO_1596 (O_1596,N_11197,N_14789);
nand UO_1597 (O_1597,N_13501,N_13181);
nand UO_1598 (O_1598,N_12124,N_11840);
nand UO_1599 (O_1599,N_11248,N_14129);
nand UO_1600 (O_1600,N_10602,N_11671);
or UO_1601 (O_1601,N_13414,N_13876);
nand UO_1602 (O_1602,N_14745,N_12131);
or UO_1603 (O_1603,N_14404,N_10737);
nand UO_1604 (O_1604,N_11716,N_11148);
and UO_1605 (O_1605,N_11230,N_14136);
nor UO_1606 (O_1606,N_12052,N_10320);
nand UO_1607 (O_1607,N_13854,N_11176);
nand UO_1608 (O_1608,N_14521,N_14958);
nand UO_1609 (O_1609,N_10877,N_10486);
or UO_1610 (O_1610,N_11401,N_12941);
nand UO_1611 (O_1611,N_11587,N_14050);
nor UO_1612 (O_1612,N_11186,N_11776);
nand UO_1613 (O_1613,N_10250,N_10715);
or UO_1614 (O_1614,N_14800,N_12603);
or UO_1615 (O_1615,N_14417,N_10915);
and UO_1616 (O_1616,N_10941,N_10844);
and UO_1617 (O_1617,N_14691,N_10441);
and UO_1618 (O_1618,N_11942,N_14573);
or UO_1619 (O_1619,N_13330,N_11891);
and UO_1620 (O_1620,N_11119,N_10609);
and UO_1621 (O_1621,N_10704,N_13754);
nand UO_1622 (O_1622,N_14509,N_11872);
nand UO_1623 (O_1623,N_11142,N_11521);
and UO_1624 (O_1624,N_13746,N_14379);
xnor UO_1625 (O_1625,N_13078,N_11136);
or UO_1626 (O_1626,N_14961,N_13924);
nor UO_1627 (O_1627,N_14308,N_10931);
nor UO_1628 (O_1628,N_11182,N_12191);
nor UO_1629 (O_1629,N_14604,N_14718);
nand UO_1630 (O_1630,N_14536,N_14959);
nand UO_1631 (O_1631,N_13929,N_14134);
nand UO_1632 (O_1632,N_14709,N_12295);
or UO_1633 (O_1633,N_14017,N_12568);
xnor UO_1634 (O_1634,N_13852,N_10293);
nor UO_1635 (O_1635,N_11235,N_12496);
nor UO_1636 (O_1636,N_13805,N_14334);
nor UO_1637 (O_1637,N_10519,N_12395);
or UO_1638 (O_1638,N_14214,N_11445);
and UO_1639 (O_1639,N_11929,N_13448);
and UO_1640 (O_1640,N_12311,N_12073);
and UO_1641 (O_1641,N_14310,N_10530);
or UO_1642 (O_1642,N_11909,N_11950);
nor UO_1643 (O_1643,N_13339,N_10024);
nor UO_1644 (O_1644,N_10542,N_14865);
xor UO_1645 (O_1645,N_10162,N_11335);
nand UO_1646 (O_1646,N_13507,N_11903);
or UO_1647 (O_1647,N_13800,N_11118);
and UO_1648 (O_1648,N_12918,N_10985);
nand UO_1649 (O_1649,N_11102,N_13172);
nand UO_1650 (O_1650,N_10128,N_11018);
xnor UO_1651 (O_1651,N_10885,N_11412);
nand UO_1652 (O_1652,N_14830,N_11886);
nor UO_1653 (O_1653,N_14113,N_14833);
xnor UO_1654 (O_1654,N_12658,N_14868);
xnor UO_1655 (O_1655,N_12204,N_12294);
and UO_1656 (O_1656,N_14248,N_11390);
and UO_1657 (O_1657,N_12725,N_11088);
or UO_1658 (O_1658,N_10625,N_13660);
nor UO_1659 (O_1659,N_11097,N_10700);
or UO_1660 (O_1660,N_11150,N_11109);
xor UO_1661 (O_1661,N_13252,N_13678);
nor UO_1662 (O_1662,N_10189,N_13378);
or UO_1663 (O_1663,N_13827,N_13942);
xor UO_1664 (O_1664,N_13159,N_14406);
nor UO_1665 (O_1665,N_11990,N_12089);
or UO_1666 (O_1666,N_12903,N_11171);
or UO_1667 (O_1667,N_14727,N_10367);
nand UO_1668 (O_1668,N_14432,N_10805);
nor UO_1669 (O_1669,N_10279,N_10589);
nand UO_1670 (O_1670,N_14066,N_14507);
nand UO_1671 (O_1671,N_12429,N_11885);
and UO_1672 (O_1672,N_13958,N_10593);
or UO_1673 (O_1673,N_12494,N_11979);
nand UO_1674 (O_1674,N_13279,N_12967);
xnor UO_1675 (O_1675,N_13934,N_14079);
nor UO_1676 (O_1676,N_14041,N_10645);
nor UO_1677 (O_1677,N_10765,N_11471);
nand UO_1678 (O_1678,N_11364,N_14001);
nor UO_1679 (O_1679,N_11703,N_12634);
nand UO_1680 (O_1680,N_12833,N_11825);
and UO_1681 (O_1681,N_10248,N_11549);
and UO_1682 (O_1682,N_11158,N_13036);
nor UO_1683 (O_1683,N_11055,N_11924);
xor UO_1684 (O_1684,N_14926,N_10452);
nor UO_1685 (O_1685,N_12415,N_14970);
nor UO_1686 (O_1686,N_11298,N_11854);
or UO_1687 (O_1687,N_12319,N_12033);
nor UO_1688 (O_1688,N_12997,N_12828);
nand UO_1689 (O_1689,N_10534,N_12250);
nor UO_1690 (O_1690,N_13937,N_10019);
or UO_1691 (O_1691,N_12023,N_11595);
nand UO_1692 (O_1692,N_11004,N_12556);
nand UO_1693 (O_1693,N_14058,N_13119);
nor UO_1694 (O_1694,N_12916,N_12163);
nand UO_1695 (O_1695,N_14918,N_13777);
nand UO_1696 (O_1696,N_12013,N_10730);
and UO_1697 (O_1697,N_11178,N_13267);
nand UO_1698 (O_1698,N_10778,N_12696);
nor UO_1699 (O_1699,N_14340,N_11435);
nand UO_1700 (O_1700,N_12185,N_12940);
nor UO_1701 (O_1701,N_10453,N_11799);
and UO_1702 (O_1702,N_11099,N_11771);
nand UO_1703 (O_1703,N_11302,N_10328);
and UO_1704 (O_1704,N_10294,N_10345);
nor UO_1705 (O_1705,N_10463,N_14304);
or UO_1706 (O_1706,N_10845,N_10809);
nor UO_1707 (O_1707,N_13194,N_14319);
or UO_1708 (O_1708,N_14495,N_14721);
nand UO_1709 (O_1709,N_10220,N_13779);
and UO_1710 (O_1710,N_10509,N_13211);
nor UO_1711 (O_1711,N_12808,N_14979);
nor UO_1712 (O_1712,N_14130,N_14606);
and UO_1713 (O_1713,N_12988,N_10572);
nor UO_1714 (O_1714,N_12739,N_11226);
nand UO_1715 (O_1715,N_12638,N_13514);
and UO_1716 (O_1716,N_11081,N_13018);
and UO_1717 (O_1717,N_13591,N_13307);
nor UO_1718 (O_1718,N_11015,N_12342);
and UO_1719 (O_1719,N_10035,N_14447);
xnor UO_1720 (O_1720,N_11360,N_12608);
nand UO_1721 (O_1721,N_12307,N_10997);
nand UO_1722 (O_1722,N_10533,N_12518);
nor UO_1723 (O_1723,N_11420,N_11966);
or UO_1724 (O_1724,N_11893,N_10637);
nor UO_1725 (O_1725,N_11256,N_12486);
nor UO_1726 (O_1726,N_11284,N_13460);
or UO_1727 (O_1727,N_11974,N_13545);
nor UO_1728 (O_1728,N_11604,N_13983);
and UO_1729 (O_1729,N_12362,N_12876);
or UO_1730 (O_1730,N_13135,N_11374);
and UO_1731 (O_1731,N_10394,N_14274);
nor UO_1732 (O_1732,N_11510,N_11502);
or UO_1733 (O_1733,N_12847,N_11691);
or UO_1734 (O_1734,N_11303,N_13697);
and UO_1735 (O_1735,N_10759,N_14897);
nand UO_1736 (O_1736,N_12353,N_10610);
or UO_1737 (O_1737,N_14888,N_13652);
or UO_1738 (O_1738,N_10121,N_12428);
or UO_1739 (O_1739,N_11144,N_13608);
nor UO_1740 (O_1740,N_11279,N_13289);
or UO_1741 (O_1741,N_13492,N_13170);
nand UO_1742 (O_1742,N_12907,N_12936);
nand UO_1743 (O_1743,N_12330,N_10103);
nand UO_1744 (O_1744,N_12661,N_13077);
or UO_1745 (O_1745,N_12513,N_12463);
nand UO_1746 (O_1746,N_11444,N_10429);
or UO_1747 (O_1747,N_14086,N_12829);
nor UO_1748 (O_1748,N_14525,N_14710);
or UO_1749 (O_1749,N_12288,N_11657);
or UO_1750 (O_1750,N_12758,N_10268);
or UO_1751 (O_1751,N_12699,N_12827);
or UO_1752 (O_1752,N_13928,N_13728);
nand UO_1753 (O_1753,N_11472,N_14353);
nor UO_1754 (O_1754,N_12219,N_10596);
or UO_1755 (O_1755,N_13704,N_10515);
nand UO_1756 (O_1756,N_14435,N_13574);
or UO_1757 (O_1757,N_14387,N_10917);
xor UO_1758 (O_1758,N_14497,N_10067);
nor UO_1759 (O_1759,N_12980,N_13300);
and UO_1760 (O_1760,N_10415,N_13221);
or UO_1761 (O_1761,N_12984,N_14377);
or UO_1762 (O_1762,N_11841,N_13508);
nor UO_1763 (O_1763,N_10037,N_12895);
or UO_1764 (O_1764,N_13212,N_10861);
nor UO_1765 (O_1765,N_12176,N_11566);
or UO_1766 (O_1766,N_13191,N_10348);
or UO_1767 (O_1767,N_13681,N_12218);
nand UO_1768 (O_1768,N_10223,N_12773);
or UO_1769 (O_1769,N_10869,N_10240);
or UO_1770 (O_1770,N_13059,N_13976);
nand UO_1771 (O_1771,N_10226,N_12707);
nor UO_1772 (O_1772,N_12613,N_13441);
and UO_1773 (O_1773,N_12844,N_12822);
and UO_1774 (O_1774,N_12962,N_10999);
nor UO_1775 (O_1775,N_14420,N_13865);
nor UO_1776 (O_1776,N_13566,N_11003);
nor UO_1777 (O_1777,N_14062,N_11738);
and UO_1778 (O_1778,N_14612,N_12935);
or UO_1779 (O_1779,N_12587,N_13730);
nor UO_1780 (O_1780,N_12588,N_12346);
or UO_1781 (O_1781,N_12690,N_14409);
nand UO_1782 (O_1782,N_11169,N_13815);
or UO_1783 (O_1783,N_13905,N_11781);
nand UO_1784 (O_1784,N_13052,N_11196);
and UO_1785 (O_1785,N_10087,N_14063);
nand UO_1786 (O_1786,N_11277,N_14254);
nor UO_1787 (O_1787,N_11711,N_11192);
and UO_1788 (O_1788,N_14294,N_10104);
nor UO_1789 (O_1789,N_11817,N_14988);
or UO_1790 (O_1790,N_12151,N_13377);
nand UO_1791 (O_1791,N_11103,N_11046);
xnor UO_1792 (O_1792,N_12275,N_14438);
or UO_1793 (O_1793,N_11077,N_11309);
and UO_1794 (O_1794,N_12909,N_12203);
nor UO_1795 (O_1795,N_10012,N_11536);
nand UO_1796 (O_1796,N_14932,N_10284);
nor UO_1797 (O_1797,N_14581,N_11048);
nand UO_1798 (O_1798,N_12506,N_12413);
nand UO_1799 (O_1799,N_12477,N_13000);
nand UO_1800 (O_1800,N_12379,N_12372);
and UO_1801 (O_1801,N_10888,N_11778);
nor UO_1802 (O_1802,N_13179,N_12789);
nand UO_1803 (O_1803,N_13553,N_13238);
and UO_1804 (O_1804,N_13832,N_11800);
nor UO_1805 (O_1805,N_11388,N_11351);
nand UO_1806 (O_1806,N_10738,N_12811);
or UO_1807 (O_1807,N_12462,N_12384);
or UO_1808 (O_1808,N_14257,N_13837);
or UO_1809 (O_1809,N_14170,N_14548);
and UO_1810 (O_1810,N_11295,N_11164);
and UO_1811 (O_1811,N_10984,N_13166);
nand UO_1812 (O_1812,N_10873,N_13846);
nor UO_1813 (O_1813,N_13213,N_13220);
and UO_1814 (O_1814,N_14582,N_13944);
or UO_1815 (O_1815,N_13162,N_10896);
nand UO_1816 (O_1816,N_13605,N_11619);
and UO_1817 (O_1817,N_10455,N_13258);
and UO_1818 (O_1818,N_12959,N_14243);
nand UO_1819 (O_1819,N_13938,N_14293);
and UO_1820 (O_1820,N_12086,N_11977);
and UO_1821 (O_1821,N_13328,N_10478);
nor UO_1822 (O_1822,N_13496,N_10136);
nor UO_1823 (O_1823,N_13991,N_12094);
or UO_1824 (O_1824,N_14754,N_10397);
and UO_1825 (O_1825,N_11679,N_10621);
and UO_1826 (O_1826,N_10283,N_14653);
and UO_1827 (O_1827,N_10301,N_10681);
nand UO_1828 (O_1828,N_10499,N_11033);
nor UO_1829 (O_1829,N_12787,N_14966);
nand UO_1830 (O_1830,N_14928,N_10866);
xor UO_1831 (O_1831,N_10684,N_10980);
and UO_1832 (O_1832,N_13627,N_11228);
and UO_1833 (O_1833,N_12767,N_10760);
and UO_1834 (O_1834,N_13290,N_13685);
and UO_1835 (O_1835,N_14922,N_10259);
and UO_1836 (O_1836,N_12538,N_11734);
nor UO_1837 (O_1837,N_11533,N_11540);
or UO_1838 (O_1838,N_11027,N_11358);
or UO_1839 (O_1839,N_13813,N_12550);
nor UO_1840 (O_1840,N_10249,N_14598);
nor UO_1841 (O_1841,N_10377,N_13104);
or UO_1842 (O_1842,N_14933,N_12531);
nor UO_1843 (O_1843,N_12238,N_11076);
xnor UO_1844 (O_1844,N_14059,N_14568);
or UO_1845 (O_1845,N_11116,N_12162);
nor UO_1846 (O_1846,N_13552,N_14538);
nand UO_1847 (O_1847,N_13362,N_11997);
nand UO_1848 (O_1848,N_13741,N_10032);
and UO_1849 (O_1849,N_12669,N_14580);
and UO_1850 (O_1850,N_14977,N_13544);
and UO_1851 (O_1851,N_12221,N_12779);
and UO_1852 (O_1852,N_10841,N_13531);
xor UO_1853 (O_1853,N_12963,N_11308);
nand UO_1854 (O_1854,N_10537,N_12722);
or UO_1855 (O_1855,N_10766,N_13515);
or UO_1856 (O_1856,N_11939,N_13350);
nor UO_1857 (O_1857,N_13374,N_14657);
xor UO_1858 (O_1858,N_14322,N_12525);
xnor UO_1859 (O_1859,N_11349,N_12192);
and UO_1860 (O_1860,N_11180,N_11139);
or UO_1861 (O_1861,N_14645,N_11447);
and UO_1862 (O_1862,N_12198,N_13398);
nand UO_1863 (O_1863,N_10652,N_11870);
nor UO_1864 (O_1864,N_10242,N_13175);
or UO_1865 (O_1865,N_13654,N_11788);
or UO_1866 (O_1866,N_10524,N_12915);
or UO_1867 (O_1867,N_12464,N_10665);
or UO_1868 (O_1868,N_12488,N_12048);
or UO_1869 (O_1869,N_11647,N_11145);
nor UO_1870 (O_1870,N_12490,N_10993);
nand UO_1871 (O_1871,N_10317,N_14516);
or UO_1872 (O_1872,N_12774,N_11900);
or UO_1873 (O_1873,N_13144,N_10154);
nand UO_1874 (O_1874,N_13147,N_14591);
nor UO_1875 (O_1875,N_12572,N_14144);
nor UO_1876 (O_1876,N_11014,N_10848);
or UO_1877 (O_1877,N_11030,N_14954);
and UO_1878 (O_1878,N_12056,N_10876);
xor UO_1879 (O_1879,N_11330,N_11641);
and UO_1880 (O_1880,N_13981,N_11528);
nand UO_1881 (O_1881,N_14957,N_14588);
and UO_1882 (O_1882,N_12604,N_13134);
nand UO_1883 (O_1883,N_14175,N_10472);
or UO_1884 (O_1884,N_13720,N_11807);
nand UO_1885 (O_1885,N_14003,N_10905);
nor UO_1886 (O_1886,N_10002,N_12565);
or UO_1887 (O_1887,N_12683,N_12240);
or UO_1888 (O_1888,N_13257,N_14419);
nand UO_1889 (O_1889,N_11970,N_11802);
or UO_1890 (O_1890,N_12913,N_12431);
or UO_1891 (O_1891,N_14848,N_11329);
nor UO_1892 (O_1892,N_12938,N_12727);
xnor UO_1893 (O_1893,N_11503,N_12559);
xnor UO_1894 (O_1894,N_11238,N_11065);
xnor UO_1895 (O_1895,N_10638,N_12312);
and UO_1896 (O_1896,N_14663,N_13601);
xor UO_1897 (O_1897,N_11779,N_13675);
nor UO_1898 (O_1898,N_10209,N_10995);
nor UO_1899 (O_1899,N_10948,N_11250);
or UO_1900 (O_1900,N_12378,N_11605);
or UO_1901 (O_1901,N_13425,N_12777);
nand UO_1902 (O_1902,N_14644,N_11611);
nand UO_1903 (O_1903,N_11897,N_14624);
nor UO_1904 (O_1904,N_14866,N_10285);
or UO_1905 (O_1905,N_13583,N_13180);
xnor UO_1906 (O_1906,N_12259,N_13453);
or UO_1907 (O_1907,N_13264,N_12512);
or UO_1908 (O_1908,N_14635,N_11344);
or UO_1909 (O_1909,N_10671,N_10291);
and UO_1910 (O_1910,N_14181,N_13839);
nor UO_1911 (O_1911,N_13775,N_10383);
nor UO_1912 (O_1912,N_13386,N_13327);
and UO_1913 (O_1913,N_11203,N_10881);
and UO_1914 (O_1914,N_10740,N_10419);
or UO_1915 (O_1915,N_13568,N_10679);
nor UO_1916 (O_1916,N_14461,N_10821);
nor UO_1917 (O_1917,N_11072,N_10692);
or UO_1918 (O_1918,N_13669,N_14909);
and UO_1919 (O_1919,N_10698,N_10762);
and UO_1920 (O_1920,N_13806,N_13926);
nor UO_1921 (O_1921,N_13757,N_11257);
nand UO_1922 (O_1922,N_12216,N_14333);
and UO_1923 (O_1923,N_14209,N_11115);
nand UO_1924 (O_1924,N_14735,N_10785);
nor UO_1925 (O_1925,N_14289,N_12119);
nand UO_1926 (O_1926,N_13309,N_11542);
or UO_1927 (O_1927,N_13028,N_14609);
and UO_1928 (O_1928,N_10425,N_10174);
nor UO_1929 (O_1929,N_13780,N_10798);
or UO_1930 (O_1930,N_14171,N_14827);
nand UO_1931 (O_1931,N_11069,N_12578);
nor UO_1932 (O_1932,N_12228,N_10566);
nand UO_1933 (O_1933,N_14351,N_10551);
nor UO_1934 (O_1934,N_10607,N_14584);
and UO_1935 (O_1935,N_10496,N_12314);
nand UO_1936 (O_1936,N_14358,N_12102);
nand UO_1937 (O_1937,N_10608,N_11798);
nand UO_1938 (O_1938,N_14459,N_12511);
xnor UO_1939 (O_1939,N_10046,N_13329);
nand UO_1940 (O_1940,N_10086,N_12155);
nand UO_1941 (O_1941,N_14680,N_12208);
and UO_1942 (O_1942,N_11511,N_14785);
or UO_1943 (O_1943,N_12405,N_13747);
nand UO_1944 (O_1944,N_13659,N_13235);
and UO_1945 (O_1945,N_12358,N_13187);
and UO_1946 (O_1946,N_12437,N_13080);
or UO_1947 (O_1947,N_13535,N_11602);
nand UO_1948 (O_1948,N_14462,N_10261);
nand UO_1949 (O_1949,N_10080,N_13560);
or UO_1950 (O_1950,N_12782,N_14325);
and UO_1951 (O_1951,N_11517,N_10672);
nand UO_1952 (O_1952,N_11460,N_12427);
or UO_1953 (O_1953,N_12503,N_14324);
xor UO_1954 (O_1954,N_14476,N_11537);
xnor UO_1955 (O_1955,N_14530,N_10207);
xor UO_1956 (O_1956,N_12563,N_10047);
or UO_1957 (O_1957,N_12906,N_14309);
nor UO_1958 (O_1958,N_13432,N_11842);
or UO_1959 (O_1959,N_10110,N_11488);
or UO_1960 (O_1960,N_14044,N_10135);
and UO_1961 (O_1961,N_10950,N_13715);
or UO_1962 (O_1962,N_11989,N_14862);
or UO_1963 (O_1963,N_10657,N_13396);
or UO_1964 (O_1964,N_10130,N_11473);
nor UO_1965 (O_1965,N_12878,N_14740);
and UO_1966 (O_1966,N_10456,N_14287);
xnor UO_1967 (O_1967,N_11895,N_14128);
nand UO_1968 (O_1968,N_13684,N_11583);
nand UO_1969 (O_1969,N_11285,N_12596);
xnor UO_1970 (O_1970,N_14448,N_12212);
or UO_1971 (O_1971,N_11925,N_12181);
nor UO_1972 (O_1972,N_14211,N_10011);
nand UO_1973 (O_1973,N_13786,N_14941);
nand UO_1974 (O_1974,N_12539,N_14617);
and UO_1975 (O_1975,N_12444,N_13168);
or UO_1976 (O_1976,N_10015,N_14703);
and UO_1977 (O_1977,N_10000,N_13859);
or UO_1978 (O_1978,N_12784,N_14349);
and UO_1979 (O_1979,N_14037,N_11324);
nand UO_1980 (O_1980,N_11497,N_14464);
or UO_1981 (O_1981,N_14746,N_10479);
or UO_1982 (O_1982,N_10322,N_10955);
xor UO_1983 (O_1983,N_12741,N_14585);
or UO_1984 (O_1984,N_11632,N_13616);
xnor UO_1985 (O_1985,N_13889,N_10654);
or UO_1986 (O_1986,N_13219,N_14899);
or UO_1987 (O_1987,N_14311,N_13483);
nor UO_1988 (O_1988,N_11234,N_11009);
or UO_1989 (O_1989,N_13610,N_14271);
or UO_1990 (O_1990,N_10234,N_11892);
and UO_1991 (O_1991,N_12809,N_12430);
and UO_1992 (O_1992,N_11723,N_14013);
nor UO_1993 (O_1993,N_10172,N_12793);
nand UO_1994 (O_1994,N_11557,N_10092);
and UO_1995 (O_1995,N_14070,N_12848);
nor UO_1996 (O_1996,N_14575,N_13833);
and UO_1997 (O_1997,N_11563,N_14460);
nor UO_1998 (O_1998,N_11194,N_11397);
or UO_1999 (O_1999,N_12289,N_14253);
endmodule