module basic_1500_15000_2000_120_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1217,In_277);
nor U1 (N_1,In_1353,In_1439);
or U2 (N_2,In_228,In_543);
or U3 (N_3,In_780,In_500);
or U4 (N_4,In_1462,In_342);
nor U5 (N_5,In_1345,In_866);
nand U6 (N_6,In_529,In_258);
nand U7 (N_7,In_658,In_626);
nand U8 (N_8,In_1493,In_252);
and U9 (N_9,In_883,In_900);
nand U10 (N_10,In_396,In_956);
nor U11 (N_11,In_466,In_1383);
nor U12 (N_12,In_905,In_236);
nand U13 (N_13,In_457,In_765);
or U14 (N_14,In_1275,In_701);
or U15 (N_15,In_738,In_672);
nand U16 (N_16,In_1074,In_328);
nor U17 (N_17,In_56,In_407);
nand U18 (N_18,In_948,In_633);
nand U19 (N_19,In_1129,In_1330);
xnor U20 (N_20,In_359,In_747);
or U21 (N_21,In_1201,In_7);
or U22 (N_22,In_212,In_1005);
and U23 (N_23,In_611,In_895);
or U24 (N_24,In_355,In_1393);
or U25 (N_25,In_1496,In_570);
nor U26 (N_26,In_1009,In_518);
and U27 (N_27,In_48,In_422);
or U28 (N_28,In_566,In_931);
or U29 (N_29,In_1309,In_1279);
nor U30 (N_30,In_970,In_975);
nor U31 (N_31,In_1165,In_698);
nor U32 (N_32,In_247,In_446);
nand U33 (N_33,In_794,In_1347);
and U34 (N_34,In_1448,In_485);
or U35 (N_35,In_408,In_1116);
nand U36 (N_36,In_49,In_312);
nand U37 (N_37,In_650,In_332);
and U38 (N_38,In_234,In_631);
nor U39 (N_39,In_730,In_1293);
nand U40 (N_40,In_1106,In_143);
or U41 (N_41,In_1160,In_642);
nand U42 (N_42,In_280,In_654);
or U43 (N_43,In_782,In_879);
and U44 (N_44,In_267,In_481);
and U45 (N_45,In_1028,In_237);
or U46 (N_46,In_74,In_996);
and U47 (N_47,In_612,In_1412);
nor U48 (N_48,In_785,In_580);
or U49 (N_49,In_824,In_6);
or U50 (N_50,In_474,In_475);
nor U51 (N_51,In_551,In_75);
nand U52 (N_52,In_1428,In_515);
nand U53 (N_53,In_510,In_1410);
or U54 (N_54,In_856,In_655);
and U55 (N_55,In_1359,In_185);
nand U56 (N_56,In_1220,In_773);
or U57 (N_57,In_641,In_189);
nor U58 (N_58,In_852,In_853);
nand U59 (N_59,In_604,In_674);
nand U60 (N_60,In_958,In_851);
nor U61 (N_61,In_1468,In_424);
nand U62 (N_62,In_1012,In_1270);
nand U63 (N_63,In_445,In_837);
and U64 (N_64,In_1102,In_315);
nand U65 (N_65,In_386,In_357);
nand U66 (N_66,In_1022,In_66);
xnor U67 (N_67,In_346,In_1017);
nor U68 (N_68,In_819,In_1046);
and U69 (N_69,In_1172,In_540);
and U70 (N_70,In_243,In_881);
or U71 (N_71,In_1485,In_547);
and U72 (N_72,In_141,In_462);
or U73 (N_73,In_439,In_1039);
or U74 (N_74,In_1161,In_8);
nor U75 (N_75,In_1465,In_902);
and U76 (N_76,In_1049,In_1027);
or U77 (N_77,In_1284,In_99);
and U78 (N_78,In_345,In_942);
or U79 (N_79,In_1195,In_398);
nand U80 (N_80,In_1385,In_925);
or U81 (N_81,In_192,In_1148);
nand U82 (N_82,In_1119,In_331);
and U83 (N_83,In_1072,In_53);
or U84 (N_84,In_982,In_193);
or U85 (N_85,In_65,In_860);
xor U86 (N_86,In_1218,In_1114);
nor U87 (N_87,In_104,In_1137);
and U88 (N_88,In_1300,In_148);
nand U89 (N_89,In_945,In_708);
nor U90 (N_90,In_400,In_1475);
xor U91 (N_91,In_1288,In_1324);
xnor U92 (N_92,In_1036,In_714);
nand U93 (N_93,In_1372,In_303);
nor U94 (N_94,In_629,In_419);
nand U95 (N_95,In_1232,In_335);
nor U96 (N_96,In_1344,In_1379);
and U97 (N_97,In_806,In_906);
nor U98 (N_98,In_517,In_197);
and U99 (N_99,In_1040,In_125);
and U100 (N_100,In_669,In_717);
xnor U101 (N_101,In_1269,In_1223);
nor U102 (N_102,In_84,In_711);
or U103 (N_103,In_157,In_416);
and U104 (N_104,In_645,In_39);
nor U105 (N_105,In_1489,In_82);
nand U106 (N_106,In_1250,In_204);
or U107 (N_107,In_1084,In_1378);
and U108 (N_108,In_751,In_493);
nor U109 (N_109,In_435,In_1305);
nand U110 (N_110,In_401,In_1308);
nor U111 (N_111,In_735,In_534);
nor U112 (N_112,In_89,In_377);
or U113 (N_113,In_271,In_387);
nor U114 (N_114,In_993,In_987);
nand U115 (N_115,In_671,In_1155);
and U116 (N_116,In_1041,In_1000);
and U117 (N_117,In_702,In_1138);
nand U118 (N_118,In_791,In_308);
nor U119 (N_119,In_1268,In_423);
nand U120 (N_120,In_1229,In_553);
nor U121 (N_121,In_829,In_1093);
nor U122 (N_122,In_362,In_184);
nor U123 (N_123,In_709,In_318);
and U124 (N_124,In_167,In_873);
and U125 (N_125,In_743,In_992);
nand U126 (N_126,In_924,In_297);
nor U127 (N_127,In_1086,In_1149);
nor U128 (N_128,In_241,N_104);
nor U129 (N_129,N_1,In_678);
and U130 (N_130,In_284,N_15);
or U131 (N_131,In_1101,In_634);
nand U132 (N_132,In_1486,In_968);
nand U133 (N_133,In_898,N_29);
xnor U134 (N_134,In_150,In_1488);
or U135 (N_135,In_1450,In_131);
or U136 (N_136,In_820,In_734);
or U137 (N_137,In_1170,In_295);
nor U138 (N_138,In_657,N_73);
or U139 (N_139,In_821,In_1388);
or U140 (N_140,In_144,In_27);
and U141 (N_141,In_1076,In_661);
nand U142 (N_142,In_390,In_927);
nand U143 (N_143,In_206,In_953);
nor U144 (N_144,In_1211,In_878);
nor U145 (N_145,In_684,In_1168);
or U146 (N_146,In_899,N_99);
and U147 (N_147,In_1209,In_615);
nor U148 (N_148,In_499,In_1071);
nand U149 (N_149,In_618,In_863);
nand U150 (N_150,In_1479,In_771);
nor U151 (N_151,In_1253,In_313);
nor U152 (N_152,In_699,In_0);
and U153 (N_153,In_1145,In_855);
nor U154 (N_154,In_746,In_1113);
nand U155 (N_155,In_1011,In_859);
or U156 (N_156,In_1075,In_455);
nand U157 (N_157,In_244,N_114);
nor U158 (N_158,In_757,In_1206);
nor U159 (N_159,In_1451,In_456);
nand U160 (N_160,N_94,In_978);
or U161 (N_161,In_512,In_1440);
or U162 (N_162,In_882,In_323);
xor U163 (N_163,In_1096,In_681);
or U164 (N_164,In_767,In_1497);
xnor U165 (N_165,In_999,In_181);
or U166 (N_166,In_546,In_223);
nand U167 (N_167,In_253,In_894);
or U168 (N_168,In_1391,In_364);
or U169 (N_169,In_316,In_660);
and U170 (N_170,In_1291,In_1081);
nor U171 (N_171,In_1136,In_1010);
and U172 (N_172,In_179,In_1097);
nand U173 (N_173,In_245,In_716);
and U174 (N_174,In_838,In_868);
nand U175 (N_175,N_119,In_38);
or U176 (N_176,N_117,In_380);
nor U177 (N_177,In_1225,In_1277);
and U178 (N_178,In_298,N_102);
nor U179 (N_179,N_23,In_915);
and U180 (N_180,In_501,In_375);
or U181 (N_181,In_688,In_473);
nor U182 (N_182,In_614,In_1342);
nor U183 (N_183,In_412,In_1243);
or U184 (N_184,In_101,In_935);
and U185 (N_185,In_726,In_610);
or U186 (N_186,In_1200,In_112);
nand U187 (N_187,In_922,In_1408);
and U188 (N_188,In_3,In_1435);
and U189 (N_189,In_1152,In_847);
and U190 (N_190,N_88,In_46);
or U191 (N_191,In_1397,In_1013);
xnor U192 (N_192,In_100,In_431);
xnor U193 (N_193,In_957,In_536);
or U194 (N_194,In_1228,In_57);
xnor U195 (N_195,In_651,In_1058);
nor U196 (N_196,In_590,N_79);
and U197 (N_197,In_124,In_81);
or U198 (N_198,In_279,In_995);
and U199 (N_199,In_1216,In_918);
nand U200 (N_200,In_222,In_903);
nor U201 (N_201,In_938,In_487);
or U202 (N_202,In_344,N_103);
or U203 (N_203,In_1381,In_319);
nor U204 (N_204,In_613,N_50);
nand U205 (N_205,In_797,In_102);
or U206 (N_206,In_453,In_1060);
nand U207 (N_207,In_256,In_349);
nand U208 (N_208,In_353,N_31);
nand U209 (N_209,In_1219,In_673);
and U210 (N_210,In_1331,In_4);
nand U211 (N_211,In_1190,In_617);
nor U212 (N_212,In_558,N_63);
nor U213 (N_213,In_1470,In_1240);
or U214 (N_214,In_320,In_530);
nand U215 (N_215,In_1455,In_827);
or U216 (N_216,In_1377,In_1251);
or U217 (N_217,In_814,In_168);
xnor U218 (N_218,In_1290,In_1019);
nand U219 (N_219,In_128,In_55);
nand U220 (N_220,In_524,In_1115);
nand U221 (N_221,In_115,In_26);
nor U222 (N_222,In_1373,In_679);
or U223 (N_223,In_561,In_801);
nand U224 (N_224,In_1436,In_5);
and U225 (N_225,In_923,In_800);
nand U226 (N_226,In_766,In_35);
nand U227 (N_227,In_707,In_1057);
or U228 (N_228,In_273,In_378);
xnor U229 (N_229,In_763,In_194);
and U230 (N_230,In_973,In_748);
xnor U231 (N_231,In_263,In_976);
and U232 (N_232,In_1338,In_966);
nand U233 (N_233,In_638,In_219);
and U234 (N_234,In_1360,In_960);
and U235 (N_235,In_1431,In_984);
and U236 (N_236,In_625,In_781);
nor U237 (N_237,In_506,In_725);
and U238 (N_238,In_176,In_393);
and U239 (N_239,In_1454,In_33);
and U240 (N_240,In_483,In_283);
nor U241 (N_241,In_261,In_595);
and U242 (N_242,N_52,In_1303);
xor U243 (N_243,In_593,In_77);
nand U244 (N_244,In_1273,In_62);
and U245 (N_245,In_94,In_1258);
nand U246 (N_246,In_199,In_1307);
and U247 (N_247,In_1214,In_209);
and U248 (N_248,In_370,In_208);
and U249 (N_249,In_229,In_405);
nor U250 (N_250,In_1355,In_1108);
nor U251 (N_251,In_1314,In_663);
nor U252 (N_252,In_1018,In_490);
nand U253 (N_253,In_685,In_255);
xnor U254 (N_254,In_498,N_34);
nor U255 (N_255,In_695,In_913);
nand U256 (N_256,In_1318,In_565);
xor U257 (N_257,In_1380,In_107);
nand U258 (N_258,In_962,In_884);
and U259 (N_259,In_582,In_290);
nor U260 (N_260,N_35,In_1052);
nor U261 (N_261,N_158,In_527);
and U262 (N_262,N_231,In_731);
nand U263 (N_263,In_1133,In_542);
nor U264 (N_264,In_299,In_823);
xnor U265 (N_265,In_268,In_1267);
nand U266 (N_266,N_134,In_1083);
nor U267 (N_267,In_1491,In_694);
or U268 (N_268,In_1490,In_514);
and U269 (N_269,In_594,In_103);
nand U270 (N_270,In_307,In_843);
and U271 (N_271,In_581,In_225);
nor U272 (N_272,In_394,In_213);
nor U273 (N_273,In_979,In_1241);
or U274 (N_274,In_86,In_682);
and U275 (N_275,In_154,N_54);
nand U276 (N_276,N_135,In_1182);
nand U277 (N_277,In_1463,In_1237);
nor U278 (N_278,In_1098,In_1069);
nand U279 (N_279,N_74,In_1064);
xor U280 (N_280,In_722,In_1321);
nand U281 (N_281,In_272,In_1316);
or U282 (N_282,In_949,In_488);
nor U283 (N_283,N_217,N_200);
and U284 (N_284,In_1419,In_1498);
nor U285 (N_285,In_482,In_37);
nor U286 (N_286,In_788,In_933);
nor U287 (N_287,In_1474,In_72);
nand U288 (N_288,N_132,N_5);
nor U289 (N_289,N_46,In_519);
or U290 (N_290,In_539,N_221);
or U291 (N_291,In_152,In_108);
and U292 (N_292,In_248,N_246);
and U293 (N_293,In_1274,In_1325);
and U294 (N_294,In_1319,In_58);
xnor U295 (N_295,In_494,In_178);
and U296 (N_296,In_778,In_693);
nor U297 (N_297,In_207,N_97);
nor U298 (N_298,In_959,N_98);
or U299 (N_299,In_952,In_1346);
and U300 (N_300,In_1197,In_1204);
or U301 (N_301,In_239,In_156);
or U302 (N_302,In_162,In_220);
or U303 (N_303,In_784,In_1394);
or U304 (N_304,In_1352,In_950);
nor U305 (N_305,N_78,N_65);
xor U306 (N_306,In_232,N_118);
nand U307 (N_307,In_361,In_338);
nand U308 (N_308,In_1401,N_109);
nor U309 (N_309,In_919,In_1128);
nor U310 (N_310,In_381,In_1443);
or U311 (N_311,In_18,In_1449);
nor U312 (N_312,In_1429,In_1295);
nand U313 (N_313,In_1007,In_1174);
and U314 (N_314,In_779,In_656);
nand U315 (N_315,In_591,In_532);
nand U316 (N_316,In_955,In_1016);
nand U317 (N_317,In_341,In_755);
nor U318 (N_318,In_1476,In_1301);
and U319 (N_319,In_1374,In_1226);
nor U320 (N_320,N_211,In_121);
xnor U321 (N_321,In_789,N_18);
nor U322 (N_322,N_185,In_160);
and U323 (N_323,In_704,In_226);
and U324 (N_324,In_598,In_1326);
xnor U325 (N_325,In_795,In_861);
and U326 (N_326,In_1315,In_436);
nor U327 (N_327,In_1208,In_577);
nand U328 (N_328,N_47,In_1079);
nand U329 (N_329,In_1131,In_434);
nand U330 (N_330,In_1185,In_23);
and U331 (N_331,N_176,N_170);
and U332 (N_332,In_1409,In_1398);
nor U333 (N_333,In_1164,In_721);
xnor U334 (N_334,N_168,In_841);
or U335 (N_335,In_1162,In_662);
nand U336 (N_336,N_129,In_1447);
nor U337 (N_337,N_230,N_96);
and U338 (N_338,In_418,In_109);
nand U339 (N_339,In_274,In_737);
or U340 (N_340,In_281,In_259);
and U341 (N_341,In_496,N_186);
and U342 (N_342,In_1461,N_207);
and U343 (N_343,In_276,N_142);
nand U344 (N_344,In_217,In_584);
or U345 (N_345,In_1065,N_49);
or U346 (N_346,N_241,In_1323);
and U347 (N_347,In_745,In_1175);
xnor U348 (N_348,In_291,N_147);
and U349 (N_349,In_145,In_211);
nor U350 (N_350,In_605,In_568);
or U351 (N_351,In_10,N_16);
and U352 (N_352,In_550,In_51);
nand U353 (N_353,In_1406,In_1051);
nor U354 (N_354,In_1213,N_90);
nor U355 (N_355,In_1395,In_822);
nor U356 (N_356,In_1441,N_166);
and U357 (N_357,In_1091,N_174);
nand U358 (N_358,In_87,In_653);
and U359 (N_359,In_1422,In_659);
xor U360 (N_360,In_1239,In_1361);
nand U361 (N_361,In_151,N_228);
and U362 (N_362,N_243,N_111);
or U363 (N_363,In_224,In_203);
and U364 (N_364,N_220,In_599);
xor U365 (N_365,In_1003,N_108);
and U366 (N_366,In_420,N_245);
nor U367 (N_367,In_14,In_586);
xnor U368 (N_368,In_454,N_69);
or U369 (N_369,In_376,In_831);
nor U370 (N_370,In_729,In_535);
and U371 (N_371,N_187,In_1231);
nand U372 (N_372,In_1387,In_1357);
nand U373 (N_373,In_43,In_783);
or U374 (N_374,N_6,In_1246);
nor U375 (N_375,In_842,In_44);
and U376 (N_376,In_1358,In_114);
nor U377 (N_377,In_1212,N_195);
or U378 (N_378,In_1222,In_122);
or U379 (N_379,In_428,In_1163);
nor U380 (N_380,N_274,In_639);
or U381 (N_381,In_119,In_1034);
or U382 (N_382,N_91,In_1276);
or U383 (N_383,In_1283,In_609);
and U384 (N_384,In_1442,In_667);
nor U385 (N_385,In_1281,In_523);
nor U386 (N_386,N_234,N_307);
nor U387 (N_387,In_1337,In_1023);
nor U388 (N_388,In_804,In_834);
or U389 (N_389,In_1280,In_1238);
or U390 (N_390,In_2,N_115);
nand U391 (N_391,In_1469,In_603);
nor U392 (N_392,N_339,In_628);
xnor U393 (N_393,N_139,N_36);
nor U394 (N_394,In_668,N_335);
nand U395 (N_395,In_972,N_271);
and U396 (N_396,In_665,In_286);
nor U397 (N_397,In_867,N_337);
or U398 (N_398,In_620,In_468);
or U399 (N_399,In_240,In_813);
nor U400 (N_400,N_2,In_1193);
and U401 (N_401,N_279,In_606);
nor U402 (N_402,In_977,In_505);
nor U403 (N_403,N_58,N_38);
and U404 (N_404,In_1473,N_363);
and U405 (N_405,In_1085,N_165);
nand U406 (N_406,N_329,In_1176);
xor U407 (N_407,In_816,In_30);
and U408 (N_408,N_260,In_643);
and U409 (N_409,In_11,N_67);
and U410 (N_410,N_44,In_300);
xnor U411 (N_411,In_644,In_1370);
or U412 (N_412,In_875,N_323);
and U413 (N_413,N_302,In_917);
and U414 (N_414,In_525,In_1188);
or U415 (N_415,In_1433,N_161);
nand U416 (N_416,In_441,In_1066);
nand U417 (N_417,In_202,In_417);
nor U418 (N_418,N_296,In_1404);
or U419 (N_419,In_1260,In_742);
nand U420 (N_420,In_397,In_368);
nand U421 (N_421,In_980,In_502);
and U422 (N_422,In_173,In_880);
nor U423 (N_423,In_1282,In_559);
or U424 (N_424,In_1339,In_385);
and U425 (N_425,In_817,In_845);
nor U426 (N_426,In_1171,N_303);
or U427 (N_427,In_1014,In_583);
nand U428 (N_428,In_458,In_713);
nor U429 (N_429,In_994,In_835);
nand U430 (N_430,In_164,In_340);
or U431 (N_431,N_250,In_1221);
or U432 (N_432,In_1090,In_775);
xnor U433 (N_433,N_287,In_607);
nor U434 (N_434,In_932,N_19);
nand U435 (N_435,In_1499,In_451);
or U436 (N_436,In_1392,In_862);
nor U437 (N_437,In_744,In_139);
and U438 (N_438,In_588,N_189);
nand U439 (N_439,In_438,N_202);
or U440 (N_440,N_4,In_552);
and U441 (N_441,In_34,In_974);
nor U442 (N_442,In_233,N_24);
or U443 (N_443,In_537,In_712);
nor U444 (N_444,In_1460,N_225);
or U445 (N_445,In_1198,N_190);
xor U446 (N_446,In_632,In_1317);
nand U447 (N_447,N_0,In_1);
nor U448 (N_448,In_753,N_86);
nor U449 (N_449,In_491,In_928);
or U450 (N_450,In_1367,In_137);
nand U451 (N_451,In_251,N_237);
or U452 (N_452,In_560,In_929);
xor U453 (N_453,N_235,In_1169);
nor U454 (N_454,N_22,In_1426);
or U455 (N_455,In_1127,N_100);
nand U456 (N_456,In_373,N_136);
nor U457 (N_457,In_413,In_69);
or U458 (N_458,N_191,In_324);
nor U459 (N_459,In_117,In_443);
and U460 (N_460,In_1363,N_128);
nor U461 (N_461,In_20,N_286);
nor U462 (N_462,In_1088,In_1118);
or U463 (N_463,N_360,In_521);
or U464 (N_464,In_325,In_705);
nand U465 (N_465,In_288,N_272);
or U466 (N_466,N_373,In_1297);
nand U467 (N_467,In_149,In_1159);
nor U468 (N_468,In_624,In_250);
and U469 (N_469,In_116,N_155);
nor U470 (N_470,In_374,In_1207);
or U471 (N_471,In_1061,In_334);
nand U472 (N_472,N_162,In_1492);
and U473 (N_473,In_772,In_1224);
nor U474 (N_474,In_637,In_88);
nand U475 (N_475,N_248,In_776);
nand U476 (N_476,N_257,In_360);
nand U477 (N_477,N_332,N_361);
and U478 (N_478,In_1037,In_664);
and U479 (N_479,In_965,In_182);
nand U480 (N_480,In_759,In_191);
nor U481 (N_481,In_1153,In_365);
nand U482 (N_482,In_347,N_180);
or U483 (N_483,In_1247,In_936);
xnor U484 (N_484,In_1077,In_739);
nor U485 (N_485,In_574,N_345);
nand U486 (N_486,N_334,In_1230);
nor U487 (N_487,In_1092,In_1340);
nor U488 (N_488,N_148,In_478);
nand U489 (N_489,N_290,N_70);
and U490 (N_490,In_1456,N_89);
xnor U491 (N_491,N_194,In_1144);
nand U492 (N_492,In_1026,In_442);
nor U493 (N_493,In_322,In_1110);
and U494 (N_494,N_359,N_258);
nand U495 (N_495,In_123,N_85);
xor U496 (N_496,N_41,In_246);
nand U497 (N_497,In_538,In_554);
nor U498 (N_498,In_1215,In_939);
nor U499 (N_499,In_602,N_9);
nor U500 (N_500,In_1452,In_120);
or U501 (N_501,In_670,N_351);
or U502 (N_502,N_33,In_61);
nand U503 (N_503,In_1329,In_1272);
nand U504 (N_504,In_840,In_1327);
nor U505 (N_505,In_1365,In_1453);
and U506 (N_506,N_140,In_200);
xnor U507 (N_507,In_770,N_285);
xor U508 (N_508,In_616,In_142);
nor U509 (N_509,In_1389,N_43);
xnor U510 (N_510,In_444,N_472);
and U511 (N_511,N_397,N_163);
nand U512 (N_512,In_410,In_68);
xor U513 (N_513,N_427,In_1055);
nand U514 (N_514,In_1117,In_293);
nor U515 (N_515,In_25,N_413);
or U516 (N_516,N_293,In_1302);
or U517 (N_517,N_379,N_459);
nor U518 (N_518,N_381,In_528);
nor U519 (N_519,In_460,In_177);
or U520 (N_520,In_850,N_160);
nand U521 (N_521,N_196,In_480);
nor U522 (N_522,In_1254,N_138);
nor U523 (N_523,In_235,In_1348);
and U524 (N_524,N_364,In_1477);
xnor U525 (N_525,In_1471,In_596);
or U526 (N_526,In_1350,In_476);
and U527 (N_527,In_282,In_808);
or U528 (N_528,In_391,In_306);
and U529 (N_529,In_1021,In_91);
nand U530 (N_530,In_343,In_1286);
nor U531 (N_531,In_1199,In_576);
xnor U532 (N_532,N_410,N_490);
or U533 (N_533,N_365,N_324);
nor U534 (N_534,In_946,In_1033);
nor U535 (N_535,In_384,In_135);
nor U536 (N_536,In_269,In_469);
nor U537 (N_537,In_872,In_1167);
xor U538 (N_538,N_450,In_1423);
or U539 (N_539,In_1006,In_1062);
or U540 (N_540,In_1244,In_1032);
and U541 (N_541,In_1313,N_122);
or U542 (N_542,In_28,In_161);
nand U543 (N_543,In_1407,In_326);
nand U544 (N_544,In_1362,N_295);
nand U545 (N_545,In_511,In_1140);
and U546 (N_546,In_155,In_221);
and U547 (N_547,N_484,In_991);
nor U548 (N_548,N_382,In_1142);
nand U549 (N_549,In_934,In_85);
and U550 (N_550,In_686,In_409);
nor U551 (N_551,N_242,In_635);
xnor U552 (N_552,N_238,N_188);
or U553 (N_553,In_429,In_230);
and U554 (N_554,In_587,N_437);
xnor U555 (N_555,In_1483,In_118);
xor U556 (N_556,N_21,N_292);
and U557 (N_557,In_196,In_1178);
nor U558 (N_558,In_908,N_197);
xnor U559 (N_559,In_1434,In_1264);
xor U560 (N_560,N_439,N_254);
and U561 (N_561,N_66,N_396);
and U562 (N_562,In_758,N_62);
or U563 (N_563,N_488,N_214);
nor U564 (N_564,In_652,In_833);
or U565 (N_565,In_1002,In_1487);
nand U566 (N_566,N_282,In_47);
nand U567 (N_567,N_487,In_21);
and U568 (N_568,N_204,N_362);
or U569 (N_569,In_1432,In_1143);
or U570 (N_570,In_495,In_304);
nor U571 (N_571,In_40,In_174);
nand U572 (N_572,In_1048,In_126);
nand U573 (N_573,N_256,In_544);
and U574 (N_574,In_777,In_1015);
and U575 (N_575,In_1405,In_358);
nand U576 (N_576,In_697,In_64);
nand U577 (N_577,In_12,In_388);
or U578 (N_578,N_486,N_55);
and U579 (N_579,In_509,N_480);
and U580 (N_580,In_1335,In_383);
nor U581 (N_581,In_836,In_470);
and U582 (N_582,In_136,N_239);
or U583 (N_583,In_869,N_398);
nor U584 (N_584,In_1139,In_440);
or U585 (N_585,In_1044,In_1256);
nand U586 (N_586,N_431,In_50);
nand U587 (N_587,In_1296,N_298);
or U588 (N_588,In_1146,In_914);
nor U589 (N_589,In_1415,In_1437);
or U590 (N_590,In_1100,N_312);
or U591 (N_591,In_1369,N_144);
nand U592 (N_592,N_319,N_283);
nor U593 (N_593,In_165,In_1482);
and U594 (N_594,In_1078,N_224);
or U595 (N_595,In_787,N_92);
and U596 (N_596,In_807,In_1425);
or U597 (N_597,In_548,N_356);
or U598 (N_598,In_623,N_278);
nor U599 (N_599,In_1166,In_706);
nor U600 (N_600,In_736,N_61);
or U601 (N_601,In_1126,In_1236);
nand U602 (N_602,In_921,In_330);
nor U603 (N_603,In_1177,N_412);
nor U604 (N_604,In_459,In_98);
nand U605 (N_605,In_22,N_268);
nor U606 (N_606,In_1234,In_826);
nand U607 (N_607,In_180,In_1262);
and U608 (N_608,In_916,N_26);
and U609 (N_609,N_222,N_84);
and U610 (N_610,In_60,In_1371);
nor U611 (N_611,In_815,In_1063);
nand U612 (N_612,In_309,In_1306);
nand U613 (N_613,In_489,In_1386);
nor U614 (N_614,In_564,N_227);
or U615 (N_615,In_472,In_1125);
nor U616 (N_616,In_1376,In_336);
nand U617 (N_617,In_727,In_877);
xor U618 (N_618,N_416,N_56);
nor U619 (N_619,In_406,N_493);
nor U620 (N_620,N_3,N_14);
and U621 (N_621,N_421,In_555);
and U622 (N_622,N_232,N_327);
or U623 (N_623,N_358,In_1008);
or U624 (N_624,In_71,N_451);
nor U625 (N_625,In_885,N_206);
nor U626 (N_626,N_582,N_213);
nor U627 (N_627,In_1123,N_265);
nand U628 (N_628,N_591,N_247);
nand U629 (N_629,In_1259,In_1024);
nor U630 (N_630,In_187,N_306);
xnor U631 (N_631,N_476,N_516);
or U632 (N_632,In_19,In_463);
or U633 (N_633,In_503,In_52);
xnor U634 (N_634,In_1478,N_328);
xor U635 (N_635,N_473,N_175);
nor U636 (N_636,In_163,N_309);
nand U637 (N_637,In_1047,In_1157);
and U638 (N_638,N_299,N_218);
nor U639 (N_639,In_1271,In_1147);
nand U640 (N_640,N_394,N_420);
or U641 (N_641,In_369,In_1043);
or U642 (N_642,In_990,N_375);
or U643 (N_643,In_79,In_687);
nor U644 (N_644,N_512,N_39);
and U645 (N_645,N_372,N_284);
nand U646 (N_646,In_961,In_311);
xnor U647 (N_647,In_969,In_159);
or U648 (N_648,N_124,N_45);
or U649 (N_649,In_427,In_106);
or U650 (N_650,In_1444,In_967);
nor U651 (N_651,N_407,N_561);
and U652 (N_652,N_349,In_943);
and U653 (N_653,In_573,In_1186);
nor U654 (N_654,N_322,In_1400);
nand U655 (N_655,In_153,N_320);
and U656 (N_656,In_985,In_31);
nand U657 (N_657,N_475,In_569);
or U658 (N_658,N_146,N_542);
or U659 (N_659,N_553,In_983);
nand U660 (N_660,N_496,N_380);
and U661 (N_661,In_1495,In_1067);
xnor U662 (N_662,N_357,In_1333);
nand U663 (N_663,In_414,N_311);
and U664 (N_664,In_433,N_40);
nand U665 (N_665,N_266,In_830);
nand U666 (N_666,In_1311,N_580);
nand U667 (N_667,N_192,N_527);
nand U668 (N_668,N_106,N_318);
nor U669 (N_669,N_354,N_419);
and U670 (N_670,N_203,In_147);
or U671 (N_671,N_442,N_544);
and U672 (N_672,N_560,In_1354);
nand U673 (N_673,In_1349,In_1249);
nor U674 (N_674,In_216,In_392);
or U675 (N_675,In_981,In_278);
nor U676 (N_676,In_29,N_606);
nand U677 (N_677,N_201,N_367);
nand U678 (N_678,In_80,In_762);
nand U679 (N_679,In_526,In_238);
and U680 (N_680,N_548,In_522);
nor U681 (N_681,N_593,N_338);
xnor U682 (N_682,N_471,In_205);
nand U683 (N_683,N_617,N_383);
nand U684 (N_684,N_369,N_313);
or U685 (N_685,In_556,In_809);
nand U686 (N_686,N_489,In_1257);
nand U687 (N_687,N_178,In_887);
nor U688 (N_688,In_812,In_798);
nor U689 (N_689,In_864,N_558);
and U690 (N_690,In_1203,N_12);
and U691 (N_691,N_432,N_482);
or U692 (N_692,In_54,In_910);
nor U693 (N_693,N_251,In_16);
or U694 (N_694,N_552,N_281);
xnor U695 (N_695,In_254,In_871);
nor U696 (N_696,N_308,In_676);
or U697 (N_697,In_1341,N_198);
nor U698 (N_698,In_1094,In_1445);
or U699 (N_699,N_401,N_470);
nor U700 (N_700,N_156,In_649);
and U701 (N_701,In_421,In_911);
and U702 (N_702,In_354,In_17);
nor U703 (N_703,In_1130,In_260);
xnor U704 (N_704,In_858,In_113);
nand U705 (N_705,N_599,N_193);
and U706 (N_706,In_1089,N_112);
or U707 (N_707,N_151,In_1187);
and U708 (N_708,N_434,In_262);
nor U709 (N_709,N_453,N_422);
nor U710 (N_710,In_622,In_266);
and U711 (N_711,In_350,In_1427);
or U712 (N_712,In_1480,In_1059);
or U713 (N_713,In_732,In_1266);
or U714 (N_714,In_426,In_1252);
nand U715 (N_715,In_1466,N_504);
nand U716 (N_716,In_504,In_811);
nand U717 (N_717,In_720,In_865);
nor U718 (N_718,In_1320,N_399);
nand U719 (N_719,In_1134,N_574);
nand U720 (N_720,In_1481,In_96);
nor U721 (N_721,N_481,In_723);
and U722 (N_722,N_425,N_621);
or U723 (N_723,In_411,In_310);
and U724 (N_724,In_36,N_169);
or U725 (N_725,In_404,In_367);
or U726 (N_726,N_521,N_406);
nand U727 (N_727,N_572,In_1227);
nor U728 (N_728,In_321,N_13);
or U729 (N_729,N_154,In_465);
and U730 (N_730,In_828,In_752);
or U731 (N_731,N_595,N_137);
nor U732 (N_732,N_321,N_377);
nand U733 (N_733,N_261,In_944);
nor U734 (N_734,N_598,In_854);
and U735 (N_735,In_111,N_457);
or U736 (N_736,N_609,In_1356);
nand U737 (N_737,N_275,In_680);
nor U738 (N_738,In_1375,N_565);
or U739 (N_739,N_182,N_353);
nand U740 (N_740,In_719,In_848);
and U741 (N_741,In_769,In_371);
and U742 (N_742,N_263,N_557);
nand U743 (N_743,N_348,N_436);
xnor U744 (N_744,In_105,N_164);
nand U745 (N_745,N_607,N_441);
and U746 (N_746,N_8,N_536);
or U747 (N_747,In_621,In_792);
nand U748 (N_748,N_264,In_399);
nor U749 (N_749,N_215,In_301);
and U750 (N_750,In_287,In_718);
or U751 (N_751,N_386,In_1390);
xnor U752 (N_752,In_507,In_1310);
or U753 (N_753,N_559,In_636);
nor U754 (N_754,N_705,In_619);
or U755 (N_755,In_448,N_549);
and U756 (N_756,In_1073,N_693);
and U757 (N_757,N_662,In_1438);
nand U758 (N_758,N_414,N_710);
or U759 (N_759,N_589,N_625);
nor U760 (N_760,N_586,In_585);
nor U761 (N_761,N_7,N_42);
nor U762 (N_762,N_682,In_1038);
nor U763 (N_763,N_474,N_656);
nand U764 (N_764,In_802,In_1068);
nor U765 (N_765,In_1494,In_32);
nor U766 (N_766,N_498,In_1210);
and U767 (N_767,In_270,N_466);
xor U768 (N_768,In_1111,N_10);
or U769 (N_769,In_1261,N_212);
or U770 (N_770,N_640,N_240);
and U771 (N_771,In_600,In_1179);
nand U772 (N_772,In_907,In_889);
nand U773 (N_773,In_846,N_703);
nor U774 (N_774,In_1351,In_186);
and U775 (N_775,N_667,N_87);
nand U776 (N_776,N_430,N_433);
or U777 (N_777,In_964,N_276);
and U778 (N_778,N_644,N_456);
nand U779 (N_779,In_986,N_208);
xor U780 (N_780,N_605,N_262);
nor U781 (N_781,N_60,N_393);
and U782 (N_782,In_479,In_796);
nor U783 (N_783,N_127,N_83);
nand U784 (N_784,In_183,N_624);
nand U785 (N_785,N_502,N_684);
xor U786 (N_786,N_378,N_579);
and U787 (N_787,N_152,N_657);
nor U788 (N_788,In_1156,N_340);
nor U789 (N_789,In_897,In_447);
xor U790 (N_790,In_520,N_28);
or U791 (N_791,N_653,N_655);
and U792 (N_792,N_301,N_458);
nand U793 (N_793,In_1180,In_1020);
and U794 (N_794,N_526,N_330);
nand U795 (N_795,In_352,In_1150);
or U796 (N_796,In_541,N_706);
nand U797 (N_797,N_739,N_347);
nor U798 (N_798,In_740,N_642);
nand U799 (N_799,N_563,N_101);
and U800 (N_800,N_460,In_90);
and U801 (N_801,N_632,In_285);
nor U802 (N_802,In_134,In_1173);
nand U803 (N_803,N_691,N_355);
nor U804 (N_804,N_229,N_637);
and U805 (N_805,In_1312,N_269);
or U806 (N_806,N_491,N_708);
xnor U807 (N_807,In_562,N_415);
nor U808 (N_808,N_686,In_579);
nor U809 (N_809,N_726,N_447);
and U810 (N_810,In_1285,N_209);
nand U811 (N_811,N_25,N_539);
nand U812 (N_812,In_329,N_395);
nand U813 (N_813,In_333,In_1053);
or U814 (N_814,N_503,N_692);
and U815 (N_815,In_382,In_1472);
or U816 (N_816,In_1082,In_997);
or U817 (N_817,N_342,N_478);
or U818 (N_818,In_857,N_627);
or U819 (N_819,N_408,In_1151);
nand U820 (N_820,N_143,In_513);
and U821 (N_821,In_1099,In_1154);
or U822 (N_822,N_64,N_573);
and U823 (N_823,N_123,N_288);
or U824 (N_824,N_145,N_405);
or U825 (N_825,In_557,In_567);
and U826 (N_826,N_730,N_623);
nand U827 (N_827,In_1484,In_690);
or U828 (N_828,In_1384,N_674);
xnor U829 (N_829,In_339,N_371);
nor U830 (N_830,In_1459,N_153);
nand U831 (N_831,N_80,N_464);
and U832 (N_832,N_718,N_551);
xor U833 (N_833,In_764,In_988);
xor U834 (N_834,In_292,In_190);
and U835 (N_835,In_1263,In_1402);
nand U836 (N_836,In_761,In_59);
and U837 (N_837,In_305,In_327);
and U838 (N_838,N_743,N_325);
nor U839 (N_839,N_619,N_280);
or U840 (N_840,In_998,In_1414);
nand U841 (N_841,N_159,In_1382);
and U842 (N_842,N_304,N_455);
or U843 (N_843,In_1194,In_337);
or U844 (N_844,In_13,N_75);
and U845 (N_845,In_1458,In_563);
nor U846 (N_846,In_129,N_443);
or U847 (N_847,N_392,N_244);
nand U848 (N_848,N_518,N_157);
and U849 (N_849,In_450,N_59);
nand U850 (N_850,In_954,In_1464);
nor U851 (N_851,N_594,N_505);
nand U852 (N_852,N_352,N_661);
nand U853 (N_853,N_696,In_432);
nor U854 (N_854,In_351,N_603);
nand U855 (N_855,In_810,In_93);
nand U856 (N_856,In_849,N_446);
nor U857 (N_857,N_629,In_132);
xor U858 (N_858,In_1196,N_616);
or U859 (N_859,N_133,In_589);
nor U860 (N_860,N_564,In_1056);
or U861 (N_861,N_444,N_291);
and U862 (N_862,N_183,N_734);
and U863 (N_863,In_597,In_133);
nand U864 (N_864,In_1004,N_658);
and U865 (N_865,In_127,In_640);
xor U866 (N_866,N_748,N_742);
nor U867 (N_867,In_1042,In_372);
nor U868 (N_868,N_341,In_1421);
nor U869 (N_869,N_715,In_215);
xnor U870 (N_870,N_477,In_296);
nor U871 (N_871,N_650,N_520);
or U872 (N_872,In_492,N_618);
nand U873 (N_873,In_1158,N_631);
and U874 (N_874,N_601,N_116);
and U875 (N_875,In_601,N_666);
nand U876 (N_876,N_836,N_403);
and U877 (N_877,N_807,In_904);
and U878 (N_878,N_862,In_1184);
nor U879 (N_879,N_20,In_832);
or U880 (N_880,N_837,N_671);
and U881 (N_881,In_188,N_30);
and U882 (N_882,In_1045,In_169);
or U883 (N_883,N_590,In_733);
nor U884 (N_884,N_779,N_829);
and U885 (N_885,N_600,N_825);
nand U886 (N_886,N_838,N_823);
or U887 (N_887,N_806,N_778);
or U888 (N_888,N_716,In_1235);
xor U889 (N_889,N_721,N_150);
xnor U890 (N_890,N_664,In_166);
or U891 (N_891,N_612,N_562);
and U892 (N_892,In_516,N_314);
and U893 (N_893,N_113,N_508);
and U894 (N_894,N_294,N_643);
and U895 (N_895,N_376,N_528);
and U896 (N_896,N_525,In_691);
and U897 (N_897,In_545,N_809);
nand U898 (N_898,N_177,In_901);
xor U899 (N_899,N_787,N_857);
and U900 (N_900,N_82,N_610);
nand U901 (N_901,N_717,N_732);
and U902 (N_902,N_756,N_523);
nand U903 (N_903,In_891,In_175);
nand U904 (N_904,In_793,In_1242);
xnor U905 (N_905,N_592,N_448);
xnor U906 (N_906,N_492,N_479);
or U907 (N_907,In_1054,In_1255);
xor U908 (N_908,N_711,N_411);
or U909 (N_909,In_870,In_728);
and U910 (N_910,In_749,N_681);
nand U911 (N_911,In_1248,In_508);
nand U912 (N_912,N_704,In_41);
nor U913 (N_913,N_566,In_1299);
nor U914 (N_914,N_833,N_723);
or U915 (N_915,In_930,In_1416);
nand U916 (N_916,N_860,N_506);
or U917 (N_917,In_1430,N_724);
xor U918 (N_918,N_741,N_343);
xnor U919 (N_919,N_344,In_9);
nand U920 (N_920,N_751,N_93);
and U921 (N_921,N_277,N_390);
nand U922 (N_922,N_828,N_370);
nor U923 (N_923,N_267,In_1087);
and U924 (N_924,In_1107,N_848);
nor U925 (N_925,N_389,N_797);
or U926 (N_926,In_464,N_760);
or U927 (N_927,N_831,N_648);
nand U928 (N_928,N_863,N_861);
or U929 (N_929,In_1031,N_532);
nand U930 (N_930,N_540,N_844);
and U931 (N_931,In_317,N_819);
nor U932 (N_932,N_550,N_873);
and U933 (N_933,N_350,N_556);
xnor U934 (N_934,N_763,In_909);
nor U935 (N_935,N_729,In_790);
and U936 (N_936,N_497,N_712);
or U937 (N_937,In_45,In_896);
nor U938 (N_938,N_864,N_821);
or U939 (N_939,N_694,N_402);
nor U940 (N_940,In_95,In_467);
nand U941 (N_941,In_760,In_395);
and U942 (N_942,N_252,N_683);
or U943 (N_943,In_1132,N_297);
and U944 (N_944,N_738,N_641);
nand U945 (N_945,N_850,In_549);
nand U946 (N_946,N_317,N_81);
nor U947 (N_947,N_181,N_289);
and U948 (N_948,In_768,In_1328);
nor U949 (N_949,N_791,N_820);
nand U950 (N_950,N_513,In_140);
or U951 (N_951,N_462,N_628);
nand U952 (N_952,N_842,N_530);
and U953 (N_953,N_105,In_42);
and U954 (N_954,In_1332,N_588);
nand U955 (N_955,In_1265,N_205);
xnor U956 (N_956,N_346,N_639);
nor U957 (N_957,N_749,N_587);
nand U958 (N_958,N_514,In_70);
nor U959 (N_959,N_668,N_652);
nor U960 (N_960,N_576,In_1446);
and U961 (N_961,N_400,N_141);
nand U962 (N_962,N_812,N_184);
and U963 (N_963,In_170,In_363);
nand U964 (N_964,N_571,N_131);
xnor U965 (N_965,N_469,N_804);
or U966 (N_966,In_1025,N_773);
xnor U967 (N_967,N_223,N_780);
nor U968 (N_968,N_845,N_173);
or U969 (N_969,In_750,In_893);
xor U970 (N_970,N_541,N_300);
nor U971 (N_971,In_572,N_509);
nand U972 (N_972,N_216,N_660);
and U973 (N_973,In_1322,In_1122);
nor U974 (N_974,N_326,N_775);
or U975 (N_975,N_404,In_710);
nor U976 (N_976,N_866,N_867);
nand U977 (N_977,N_37,N_388);
nand U978 (N_978,N_614,In_171);
and U979 (N_979,N_125,In_1418);
and U980 (N_980,In_1399,In_1202);
and U981 (N_981,N_391,In_231);
nand U982 (N_982,In_227,In_1289);
xor U983 (N_983,N_507,N_71);
xor U984 (N_984,N_107,N_126);
xor U985 (N_985,N_429,N_834);
and U986 (N_986,N_537,N_435);
or U987 (N_987,N_495,N_856);
xor U988 (N_988,In_73,N_417);
or U989 (N_989,In_1298,N_698);
or U990 (N_990,In_886,N_733);
and U991 (N_991,N_622,N_798);
nor U992 (N_992,N_810,N_646);
and U993 (N_993,N_501,In_275);
and U994 (N_994,In_1413,N_555);
nor U995 (N_995,N_688,N_315);
nor U996 (N_996,N_785,N_452);
or U997 (N_997,In_195,N_449);
or U998 (N_998,In_630,In_1343);
nand U999 (N_999,In_844,In_1467);
nor U1000 (N_1000,N_336,N_149);
and U1001 (N_1001,N_27,In_289);
or U1002 (N_1002,N_949,N_604);
or U1003 (N_1003,N_11,N_554);
and U1004 (N_1004,N_649,N_947);
nand U1005 (N_1005,N_870,N_700);
nand U1006 (N_1006,N_953,In_575);
and U1007 (N_1007,N_110,N_633);
and U1008 (N_1008,N_762,N_920);
xor U1009 (N_1009,N_894,In_696);
nand U1010 (N_1010,In_971,N_596);
nand U1011 (N_1011,In_1183,In_786);
and U1012 (N_1012,N_529,In_947);
or U1013 (N_1013,In_926,N_57);
and U1014 (N_1014,N_904,N_961);
or U1015 (N_1015,N_774,N_270);
or U1016 (N_1016,N_900,N_835);
and U1017 (N_1017,N_517,N_832);
or U1018 (N_1018,N_385,N_745);
nand U1019 (N_1019,N_305,N_687);
or U1020 (N_1020,In_892,N_720);
and U1021 (N_1021,N_991,N_423);
nor U1022 (N_1022,N_368,In_920);
and U1023 (N_1023,N_915,In_689);
nand U1024 (N_1024,N_750,N_731);
nand U1025 (N_1025,In_571,In_666);
nor U1026 (N_1026,N_792,In_1095);
nand U1027 (N_1027,In_314,N_766);
nor U1028 (N_1028,N_48,N_974);
nor U1029 (N_1029,N_972,N_818);
xor U1030 (N_1030,N_199,N_626);
nand U1031 (N_1031,N_962,In_1001);
nor U1032 (N_1032,N_925,N_950);
nand U1033 (N_1033,N_602,In_379);
or U1034 (N_1034,N_875,N_77);
nor U1035 (N_1035,N_17,N_869);
nand U1036 (N_1036,N_120,In_452);
or U1037 (N_1037,In_437,In_941);
and U1038 (N_1038,N_901,N_535);
nor U1039 (N_1039,N_483,N_824);
or U1040 (N_1040,In_1205,In_675);
or U1041 (N_1041,N_651,N_467);
xor U1042 (N_1042,In_97,N_914);
and U1043 (N_1043,In_692,N_800);
nand U1044 (N_1044,N_440,N_795);
xnor U1045 (N_1045,N_273,N_53);
or U1046 (N_1046,N_996,In_1278);
or U1047 (N_1047,N_813,N_801);
or U1048 (N_1048,N_685,N_233);
and U1049 (N_1049,N_783,N_445);
nor U1050 (N_1050,N_999,N_975);
or U1051 (N_1051,N_752,N_980);
and U1052 (N_1052,N_937,N_968);
nor U1053 (N_1053,In_608,N_570);
nand U1054 (N_1054,N_796,N_882);
nand U1055 (N_1055,N_454,N_675);
or U1056 (N_1056,N_965,N_852);
nand U1057 (N_1057,N_898,In_592);
or U1058 (N_1058,N_815,N_922);
nor U1059 (N_1059,N_567,N_906);
and U1060 (N_1060,In_646,N_995);
and U1061 (N_1061,N_735,In_210);
nand U1062 (N_1062,N_597,N_816);
or U1063 (N_1063,N_615,N_547);
nor U1064 (N_1064,In_415,N_485);
nor U1065 (N_1065,N_888,N_772);
and U1066 (N_1066,N_881,N_545);
nand U1067 (N_1067,N_533,In_1366);
nand U1068 (N_1068,In_1030,N_927);
nor U1069 (N_1069,N_753,In_774);
or U1070 (N_1070,N_630,In_951);
xnor U1071 (N_1071,In_756,N_957);
nand U1072 (N_1072,N_868,N_581);
or U1073 (N_1073,N_670,N_911);
nand U1074 (N_1074,N_855,N_921);
and U1075 (N_1075,In_805,N_895);
and U1076 (N_1076,N_886,N_585);
or U1077 (N_1077,N_967,In_78);
or U1078 (N_1078,In_402,In_1080);
and U1079 (N_1079,In_218,N_959);
or U1080 (N_1080,N_707,N_941);
nand U1081 (N_1081,N_677,N_977);
nand U1082 (N_1082,N_702,In_1294);
nand U1083 (N_1083,N_931,N_989);
nor U1084 (N_1084,N_167,In_484);
and U1085 (N_1085,N_635,N_534);
nand U1086 (N_1086,N_814,N_878);
nand U1087 (N_1087,In_1192,N_993);
and U1088 (N_1088,In_24,N_988);
nor U1089 (N_1089,N_893,N_874);
nor U1090 (N_1090,In_67,N_569);
and U1091 (N_1091,N_672,In_940);
and U1092 (N_1092,N_531,N_500);
nand U1093 (N_1093,In_1233,N_255);
and U1094 (N_1094,In_888,N_638);
nand U1095 (N_1095,In_803,In_1420);
or U1096 (N_1096,In_1124,N_669);
and U1097 (N_1097,N_697,In_461);
nor U1098 (N_1098,N_956,N_689);
or U1099 (N_1099,N_511,N_316);
xor U1100 (N_1100,N_384,N_746);
and U1101 (N_1101,N_902,In_1304);
and U1102 (N_1102,In_110,In_214);
and U1103 (N_1103,N_872,N_912);
nor U1104 (N_1104,In_874,N_923);
nor U1105 (N_1105,N_973,In_366);
nand U1106 (N_1106,In_1109,N_822);
or U1107 (N_1107,N_847,N_935);
nor U1108 (N_1108,N_95,N_727);
xor U1109 (N_1109,In_76,N_522);
or U1110 (N_1110,N_620,N_426);
or U1111 (N_1111,N_659,N_871);
nand U1112 (N_1112,N_952,N_757);
xnor U1113 (N_1113,N_771,In_1135);
or U1114 (N_1114,N_676,N_728);
nand U1115 (N_1115,In_1181,N_584);
or U1116 (N_1116,N_865,In_937);
or U1117 (N_1117,N_709,N_701);
or U1118 (N_1118,In_1103,N_958);
nand U1119 (N_1119,N_976,N_963);
nand U1120 (N_1120,N_846,N_418);
nand U1121 (N_1121,In_198,N_978);
and U1122 (N_1122,N_946,In_754);
and U1123 (N_1123,N_253,In_158);
and U1124 (N_1124,In_425,N_903);
nand U1125 (N_1125,In_1070,N_1042);
or U1126 (N_1126,N_428,In_683);
nor U1127 (N_1127,N_782,N_887);
or U1128 (N_1128,N_575,N_1081);
nand U1129 (N_1129,N_1003,N_1014);
nor U1130 (N_1130,N_924,N_1106);
and U1131 (N_1131,N_1007,N_905);
and U1132 (N_1132,N_634,N_910);
nor U1133 (N_1133,N_1072,N_72);
or U1134 (N_1134,N_1085,N_461);
or U1135 (N_1135,N_1068,N_789);
nand U1136 (N_1136,N_424,N_979);
or U1137 (N_1137,N_1046,N_1101);
and U1138 (N_1138,N_768,N_1112);
xor U1139 (N_1139,N_249,N_538);
nand U1140 (N_1140,N_608,N_1122);
or U1141 (N_1141,N_543,N_964);
nor U1142 (N_1142,N_333,In_1336);
nor U1143 (N_1143,N_1011,In_449);
or U1144 (N_1144,N_896,N_1082);
and U1145 (N_1145,In_1189,In_715);
nand U1146 (N_1146,In_92,In_264);
and U1147 (N_1147,In_201,N_817);
nor U1148 (N_1148,N_969,N_932);
nand U1149 (N_1149,N_1049,N_1096);
nand U1150 (N_1150,In_648,N_1079);
nor U1151 (N_1151,N_1094,N_843);
or U1152 (N_1152,In_677,N_1097);
or U1153 (N_1153,N_1031,In_1035);
or U1154 (N_1154,N_908,N_519);
and U1155 (N_1155,N_1039,In_1403);
xor U1156 (N_1156,N_788,N_943);
and U1157 (N_1157,N_468,N_546);
nand U1158 (N_1158,In_627,N_744);
and U1159 (N_1159,N_877,N_1018);
or U1160 (N_1160,N_1008,N_1078);
nor U1161 (N_1161,N_690,N_1073);
nand U1162 (N_1162,N_695,N_839);
or U1163 (N_1163,In_477,N_1120);
nand U1164 (N_1164,N_892,N_858);
or U1165 (N_1165,N_1110,N_944);
nor U1166 (N_1166,N_1069,N_1123);
and U1167 (N_1167,N_754,N_51);
nand U1168 (N_1168,N_121,In_1364);
nor U1169 (N_1169,In_1396,N_1026);
and U1170 (N_1170,N_755,N_1117);
or U1171 (N_1171,N_611,N_1002);
or U1172 (N_1172,N_1016,N_981);
nand U1173 (N_1173,In_1245,In_799);
nor U1174 (N_1174,In_356,In_876);
nor U1175 (N_1175,N_1107,N_1027);
xnor U1176 (N_1176,N_1013,N_983);
and U1177 (N_1177,In_486,N_1051);
nand U1178 (N_1178,In_1120,N_933);
or U1179 (N_1179,In_302,N_719);
and U1180 (N_1180,N_699,N_758);
or U1181 (N_1181,N_954,N_374);
and U1182 (N_1182,In_130,N_1065);
and U1183 (N_1183,N_808,In_1029);
or U1184 (N_1184,In_741,N_1090);
nand U1185 (N_1185,N_1124,N_1091);
nand U1186 (N_1186,N_1084,N_1109);
nor U1187 (N_1187,N_987,N_803);
xnor U1188 (N_1188,N_1076,N_1098);
or U1189 (N_1189,N_1113,N_1035);
and U1190 (N_1190,N_851,N_1061);
xnor U1191 (N_1191,N_1055,N_1052);
or U1192 (N_1192,In_1417,N_647);
and U1193 (N_1193,In_146,N_577);
nand U1194 (N_1194,N_722,N_1075);
and U1195 (N_1195,N_1038,N_1001);
nor U1196 (N_1196,N_409,N_1034);
nor U1197 (N_1197,N_890,N_997);
nand U1198 (N_1198,In_703,N_1036);
nor U1199 (N_1199,In_531,N_1115);
or U1200 (N_1200,N_613,N_1058);
xor U1201 (N_1201,In_1104,N_438);
nor U1202 (N_1202,N_883,N_1095);
nor U1203 (N_1203,N_984,In_1191);
and U1204 (N_1204,N_1071,N_1104);
or U1205 (N_1205,N_942,N_1028);
nand U1206 (N_1206,N_1020,N_1006);
xnor U1207 (N_1207,In_1292,N_827);
or U1208 (N_1208,N_645,N_811);
nand U1209 (N_1209,In_1121,N_1041);
nor U1210 (N_1210,N_936,N_907);
xor U1211 (N_1211,N_982,N_714);
and U1212 (N_1212,N_1064,N_1121);
nor U1213 (N_1213,In_1368,N_1012);
nand U1214 (N_1214,In_839,N_171);
nand U1215 (N_1215,N_994,In_700);
nor U1216 (N_1216,N_1103,N_926);
nand U1217 (N_1217,N_948,N_784);
nand U1218 (N_1218,In_63,N_465);
and U1219 (N_1219,N_1108,N_1070);
and U1220 (N_1220,N_970,N_876);
and U1221 (N_1221,N_219,N_853);
nor U1222 (N_1222,N_1086,In_257);
nand U1223 (N_1223,N_1043,N_880);
or U1224 (N_1224,N_793,N_1015);
nand U1225 (N_1225,N_179,N_1010);
xor U1226 (N_1226,N_678,N_794);
nor U1227 (N_1227,N_1074,N_891);
or U1228 (N_1228,N_1111,In_389);
or U1229 (N_1229,N_665,N_673);
and U1230 (N_1230,N_805,N_884);
and U1231 (N_1231,N_1102,N_1066);
and U1232 (N_1232,In_1105,N_840);
nor U1233 (N_1233,N_986,In_430);
and U1234 (N_1234,N_1025,N_1100);
nor U1235 (N_1235,N_1044,N_799);
or U1236 (N_1236,N_826,N_1083);
or U1237 (N_1237,N_1093,N_1059);
and U1238 (N_1238,N_765,In_1112);
nor U1239 (N_1239,N_515,N_1088);
nor U1240 (N_1240,N_918,N_928);
nand U1241 (N_1241,N_259,N_663);
nor U1242 (N_1242,N_1105,N_1087);
nand U1243 (N_1243,N_510,N_680);
nand U1244 (N_1244,N_310,N_1062);
and U1245 (N_1245,N_1089,N_747);
and U1246 (N_1246,N_1023,N_945);
nand U1247 (N_1247,N_1056,N_1029);
nand U1248 (N_1248,N_583,N_725);
or U1249 (N_1249,N_1048,N_919);
nand U1250 (N_1250,In_249,N_1205);
nor U1251 (N_1251,N_1143,N_1183);
or U1252 (N_1252,N_494,N_1067);
nor U1253 (N_1253,N_1129,N_929);
xor U1254 (N_1254,In_265,N_776);
and U1255 (N_1255,In_138,N_1126);
nand U1256 (N_1256,N_1057,N_1024);
or U1257 (N_1257,N_1125,N_1173);
and U1258 (N_1258,N_1226,N_1246);
nand U1259 (N_1259,N_1045,N_955);
xor U1260 (N_1260,N_1222,N_1238);
or U1261 (N_1261,N_985,N_1150);
nand U1262 (N_1262,N_1148,N_854);
nor U1263 (N_1263,N_1128,N_1155);
nand U1264 (N_1264,N_1141,In_912);
nand U1265 (N_1265,N_210,N_1127);
and U1266 (N_1266,N_1131,N_992);
and U1267 (N_1267,N_1227,N_916);
or U1268 (N_1268,N_899,In_647);
nor U1269 (N_1269,N_1140,N_897);
or U1270 (N_1270,N_1170,In_1457);
nor U1271 (N_1271,N_1139,N_740);
and U1272 (N_1272,N_998,N_1217);
nand U1273 (N_1273,N_913,N_1221);
and U1274 (N_1274,N_1216,In_1334);
nor U1275 (N_1275,N_1239,N_1144);
and U1276 (N_1276,N_960,N_761);
nand U1277 (N_1277,N_1208,N_1050);
nor U1278 (N_1278,N_802,N_1158);
nand U1279 (N_1279,N_172,N_1168);
and U1280 (N_1280,N_130,N_830);
and U1281 (N_1281,N_1218,N_1130);
nand U1282 (N_1282,N_1193,In_471);
nor U1283 (N_1283,N_1153,N_1040);
nor U1284 (N_1284,N_1176,N_1021);
nand U1285 (N_1285,N_387,N_1243);
nor U1286 (N_1286,N_1195,N_1197);
and U1287 (N_1287,N_236,N_1149);
nor U1288 (N_1288,N_1116,In_825);
and U1289 (N_1289,N_1152,N_938);
and U1290 (N_1290,N_781,In_1424);
and U1291 (N_1291,N_578,In_172);
nor U1292 (N_1292,In_403,N_226);
nand U1293 (N_1293,N_1199,N_777);
nand U1294 (N_1294,In_963,N_1200);
nor U1295 (N_1295,N_1194,N_1249);
and U1296 (N_1296,N_1206,N_1017);
nand U1297 (N_1297,N_1171,N_1215);
nor U1298 (N_1298,N_1186,N_939);
or U1299 (N_1299,N_930,N_971);
and U1300 (N_1300,N_1241,In_83);
and U1301 (N_1301,N_1047,In_989);
or U1302 (N_1302,N_1165,N_1005);
nand U1303 (N_1303,N_1092,N_1177);
xor U1304 (N_1304,N_1234,In_294);
nand U1305 (N_1305,In_497,N_1191);
nand U1306 (N_1306,N_1202,N_1204);
and U1307 (N_1307,N_1209,In_890);
nand U1308 (N_1308,N_859,N_1138);
nand U1309 (N_1309,N_1030,N_1147);
or U1310 (N_1310,N_1185,N_1118);
or U1311 (N_1311,N_1223,N_1054);
or U1312 (N_1312,N_1154,N_1099);
and U1313 (N_1313,N_1210,N_889);
xor U1314 (N_1314,N_1000,N_1211);
nor U1315 (N_1315,N_32,N_366);
nor U1316 (N_1316,N_1151,N_1004);
nor U1317 (N_1317,In_578,N_1231);
nor U1318 (N_1318,N_1159,N_1037);
nand U1319 (N_1319,N_1203,N_1220);
xnor U1320 (N_1320,N_1196,N_769);
nand U1321 (N_1321,N_1033,N_1229);
and U1322 (N_1322,N_1184,N_1180);
and U1323 (N_1323,N_849,N_1187);
xor U1324 (N_1324,N_879,In_1050);
and U1325 (N_1325,N_1233,N_1189);
or U1326 (N_1326,N_1135,In_818);
nor U1327 (N_1327,N_1162,N_770);
nor U1328 (N_1328,N_934,N_1244);
nand U1329 (N_1329,N_1132,N_966);
or U1330 (N_1330,N_940,N_1207);
xnor U1331 (N_1331,N_1167,N_1164);
and U1332 (N_1332,N_654,N_1225);
xnor U1333 (N_1333,N_1219,N_790);
and U1334 (N_1334,N_1146,N_1198);
xnor U1335 (N_1335,N_1009,N_1174);
and U1336 (N_1336,N_331,N_1156);
or U1337 (N_1337,N_1063,N_764);
and U1338 (N_1338,In_1141,N_1188);
nand U1339 (N_1339,N_1134,N_1060);
and U1340 (N_1340,N_1142,In_15);
nor U1341 (N_1341,N_1172,N_636);
nor U1342 (N_1342,In_1287,N_1248);
nand U1343 (N_1343,N_1182,N_759);
and U1344 (N_1344,N_1181,In_724);
and U1345 (N_1345,N_1192,N_1232);
nand U1346 (N_1346,In_1411,N_1212);
and U1347 (N_1347,N_713,N_1114);
and U1348 (N_1348,N_736,N_1213);
and U1349 (N_1349,N_1137,N_909);
or U1350 (N_1350,In_242,N_1160);
or U1351 (N_1351,N_1032,N_767);
nor U1352 (N_1352,N_1022,N_1175);
nand U1353 (N_1353,N_463,N_1235);
or U1354 (N_1354,N_1080,N_737);
nor U1355 (N_1355,N_1157,N_1214);
or U1356 (N_1356,N_1179,N_1228);
nor U1357 (N_1357,N_786,N_679);
nor U1358 (N_1358,N_1163,N_951);
and U1359 (N_1359,N_885,N_1136);
or U1360 (N_1360,N_1236,N_990);
nor U1361 (N_1361,N_1053,N_1245);
and U1362 (N_1362,N_499,N_1169);
or U1363 (N_1363,N_1178,N_1145);
nor U1364 (N_1364,N_841,N_1247);
and U1365 (N_1365,N_1224,N_1166);
or U1366 (N_1366,N_1119,N_1133);
or U1367 (N_1367,N_1237,N_524);
or U1368 (N_1368,In_348,N_76);
and U1369 (N_1369,N_1242,N_68);
and U1370 (N_1370,N_1240,N_1201);
nand U1371 (N_1371,In_533,N_1230);
nor U1372 (N_1372,N_1190,N_1019);
nand U1373 (N_1373,N_917,N_1077);
or U1374 (N_1374,N_1161,N_568);
nand U1375 (N_1375,N_1254,N_1255);
nor U1376 (N_1376,N_1309,N_1351);
and U1377 (N_1377,N_1346,N_1277);
and U1378 (N_1378,N_1316,N_1334);
or U1379 (N_1379,N_1260,N_1335);
nand U1380 (N_1380,N_1327,N_1374);
nor U1381 (N_1381,N_1315,N_1293);
and U1382 (N_1382,N_1333,N_1266);
nor U1383 (N_1383,N_1285,N_1312);
nor U1384 (N_1384,N_1345,N_1303);
xor U1385 (N_1385,N_1368,N_1300);
nand U1386 (N_1386,N_1325,N_1269);
nor U1387 (N_1387,N_1298,N_1367);
or U1388 (N_1388,N_1363,N_1295);
or U1389 (N_1389,N_1328,N_1353);
nand U1390 (N_1390,N_1318,N_1355);
nor U1391 (N_1391,N_1258,N_1263);
and U1392 (N_1392,N_1292,N_1343);
nor U1393 (N_1393,N_1329,N_1305);
or U1394 (N_1394,N_1336,N_1360);
nand U1395 (N_1395,N_1284,N_1253);
and U1396 (N_1396,N_1313,N_1307);
or U1397 (N_1397,N_1371,N_1339);
nand U1398 (N_1398,N_1342,N_1281);
and U1399 (N_1399,N_1296,N_1352);
xnor U1400 (N_1400,N_1319,N_1340);
nand U1401 (N_1401,N_1369,N_1347);
and U1402 (N_1402,N_1301,N_1267);
and U1403 (N_1403,N_1370,N_1272);
xor U1404 (N_1404,N_1306,N_1287);
nand U1405 (N_1405,N_1270,N_1297);
or U1406 (N_1406,N_1275,N_1299);
nor U1407 (N_1407,N_1256,N_1252);
nor U1408 (N_1408,N_1289,N_1321);
or U1409 (N_1409,N_1291,N_1273);
nand U1410 (N_1410,N_1259,N_1311);
and U1411 (N_1411,N_1286,N_1276);
nand U1412 (N_1412,N_1331,N_1302);
xor U1413 (N_1413,N_1358,N_1326);
nor U1414 (N_1414,N_1357,N_1337);
nand U1415 (N_1415,N_1271,N_1251);
or U1416 (N_1416,N_1372,N_1317);
and U1417 (N_1417,N_1341,N_1283);
or U1418 (N_1418,N_1322,N_1310);
nand U1419 (N_1419,N_1354,N_1265);
nand U1420 (N_1420,N_1338,N_1274);
nand U1421 (N_1421,N_1350,N_1356);
nand U1422 (N_1422,N_1264,N_1373);
or U1423 (N_1423,N_1250,N_1279);
nand U1424 (N_1424,N_1294,N_1348);
nand U1425 (N_1425,N_1362,N_1330);
xor U1426 (N_1426,N_1261,N_1257);
or U1427 (N_1427,N_1288,N_1359);
or U1428 (N_1428,N_1323,N_1365);
nand U1429 (N_1429,N_1349,N_1282);
and U1430 (N_1430,N_1280,N_1361);
and U1431 (N_1431,N_1314,N_1268);
nand U1432 (N_1432,N_1304,N_1278);
and U1433 (N_1433,N_1344,N_1366);
xor U1434 (N_1434,N_1290,N_1364);
or U1435 (N_1435,N_1320,N_1324);
or U1436 (N_1436,N_1332,N_1262);
xnor U1437 (N_1437,N_1308,N_1347);
or U1438 (N_1438,N_1297,N_1341);
nand U1439 (N_1439,N_1356,N_1346);
and U1440 (N_1440,N_1306,N_1257);
nand U1441 (N_1441,N_1297,N_1346);
nand U1442 (N_1442,N_1260,N_1317);
nor U1443 (N_1443,N_1293,N_1336);
and U1444 (N_1444,N_1346,N_1337);
xnor U1445 (N_1445,N_1321,N_1263);
or U1446 (N_1446,N_1315,N_1326);
nor U1447 (N_1447,N_1257,N_1255);
and U1448 (N_1448,N_1355,N_1357);
nor U1449 (N_1449,N_1254,N_1311);
nand U1450 (N_1450,N_1295,N_1293);
and U1451 (N_1451,N_1354,N_1374);
xor U1452 (N_1452,N_1285,N_1299);
xor U1453 (N_1453,N_1355,N_1324);
and U1454 (N_1454,N_1358,N_1312);
and U1455 (N_1455,N_1310,N_1268);
and U1456 (N_1456,N_1346,N_1327);
nand U1457 (N_1457,N_1308,N_1259);
nand U1458 (N_1458,N_1279,N_1278);
and U1459 (N_1459,N_1280,N_1346);
and U1460 (N_1460,N_1282,N_1321);
or U1461 (N_1461,N_1323,N_1345);
and U1462 (N_1462,N_1307,N_1358);
nand U1463 (N_1463,N_1322,N_1266);
or U1464 (N_1464,N_1270,N_1326);
or U1465 (N_1465,N_1271,N_1253);
or U1466 (N_1466,N_1314,N_1340);
and U1467 (N_1467,N_1330,N_1339);
and U1468 (N_1468,N_1329,N_1279);
or U1469 (N_1469,N_1277,N_1329);
and U1470 (N_1470,N_1287,N_1363);
nand U1471 (N_1471,N_1364,N_1317);
or U1472 (N_1472,N_1357,N_1304);
and U1473 (N_1473,N_1260,N_1297);
and U1474 (N_1474,N_1251,N_1283);
nor U1475 (N_1475,N_1299,N_1250);
or U1476 (N_1476,N_1363,N_1367);
and U1477 (N_1477,N_1341,N_1357);
and U1478 (N_1478,N_1262,N_1306);
nor U1479 (N_1479,N_1337,N_1269);
nor U1480 (N_1480,N_1352,N_1318);
nor U1481 (N_1481,N_1317,N_1320);
nor U1482 (N_1482,N_1364,N_1335);
xor U1483 (N_1483,N_1354,N_1252);
nand U1484 (N_1484,N_1281,N_1340);
and U1485 (N_1485,N_1267,N_1319);
nand U1486 (N_1486,N_1265,N_1294);
and U1487 (N_1487,N_1316,N_1254);
nor U1488 (N_1488,N_1272,N_1363);
nand U1489 (N_1489,N_1295,N_1273);
xnor U1490 (N_1490,N_1299,N_1308);
nand U1491 (N_1491,N_1300,N_1254);
nor U1492 (N_1492,N_1347,N_1355);
nor U1493 (N_1493,N_1358,N_1362);
or U1494 (N_1494,N_1368,N_1342);
nand U1495 (N_1495,N_1259,N_1306);
nand U1496 (N_1496,N_1270,N_1356);
nor U1497 (N_1497,N_1288,N_1310);
nand U1498 (N_1498,N_1280,N_1334);
or U1499 (N_1499,N_1367,N_1253);
xor U1500 (N_1500,N_1462,N_1432);
xor U1501 (N_1501,N_1485,N_1456);
and U1502 (N_1502,N_1460,N_1409);
and U1503 (N_1503,N_1393,N_1429);
nor U1504 (N_1504,N_1375,N_1384);
xnor U1505 (N_1505,N_1491,N_1417);
and U1506 (N_1506,N_1401,N_1469);
nor U1507 (N_1507,N_1472,N_1470);
nor U1508 (N_1508,N_1413,N_1404);
and U1509 (N_1509,N_1488,N_1453);
nor U1510 (N_1510,N_1438,N_1451);
nor U1511 (N_1511,N_1497,N_1459);
nand U1512 (N_1512,N_1471,N_1475);
nor U1513 (N_1513,N_1406,N_1474);
nor U1514 (N_1514,N_1435,N_1444);
nor U1515 (N_1515,N_1418,N_1467);
nand U1516 (N_1516,N_1378,N_1416);
nor U1517 (N_1517,N_1377,N_1392);
nand U1518 (N_1518,N_1463,N_1380);
xor U1519 (N_1519,N_1419,N_1395);
or U1520 (N_1520,N_1387,N_1396);
or U1521 (N_1521,N_1480,N_1496);
nor U1522 (N_1522,N_1481,N_1415);
nor U1523 (N_1523,N_1422,N_1457);
or U1524 (N_1524,N_1383,N_1490);
or U1525 (N_1525,N_1414,N_1428);
or U1526 (N_1526,N_1478,N_1449);
nand U1527 (N_1527,N_1477,N_1446);
or U1528 (N_1528,N_1399,N_1426);
or U1529 (N_1529,N_1464,N_1398);
nand U1530 (N_1530,N_1483,N_1389);
and U1531 (N_1531,N_1468,N_1388);
xnor U1532 (N_1532,N_1376,N_1394);
or U1533 (N_1533,N_1447,N_1454);
or U1534 (N_1534,N_1430,N_1420);
nand U1535 (N_1535,N_1482,N_1407);
nor U1536 (N_1536,N_1455,N_1433);
or U1537 (N_1537,N_1499,N_1443);
nand U1538 (N_1538,N_1466,N_1410);
and U1539 (N_1539,N_1476,N_1473);
and U1540 (N_1540,N_1437,N_1411);
and U1541 (N_1541,N_1494,N_1452);
or U1542 (N_1542,N_1458,N_1423);
nor U1543 (N_1543,N_1440,N_1445);
xor U1544 (N_1544,N_1434,N_1431);
nand U1545 (N_1545,N_1425,N_1379);
nor U1546 (N_1546,N_1421,N_1439);
or U1547 (N_1547,N_1390,N_1441);
nand U1548 (N_1548,N_1489,N_1484);
or U1549 (N_1549,N_1486,N_1487);
or U1550 (N_1550,N_1465,N_1448);
nand U1551 (N_1551,N_1400,N_1479);
or U1552 (N_1552,N_1402,N_1442);
and U1553 (N_1553,N_1495,N_1461);
xor U1554 (N_1554,N_1424,N_1405);
nor U1555 (N_1555,N_1403,N_1412);
xor U1556 (N_1556,N_1427,N_1397);
nand U1557 (N_1557,N_1498,N_1408);
or U1558 (N_1558,N_1391,N_1436);
and U1559 (N_1559,N_1382,N_1385);
nand U1560 (N_1560,N_1386,N_1492);
nand U1561 (N_1561,N_1493,N_1450);
and U1562 (N_1562,N_1381,N_1482);
or U1563 (N_1563,N_1401,N_1388);
nand U1564 (N_1564,N_1397,N_1422);
nor U1565 (N_1565,N_1378,N_1398);
and U1566 (N_1566,N_1458,N_1399);
nor U1567 (N_1567,N_1492,N_1442);
or U1568 (N_1568,N_1404,N_1489);
nand U1569 (N_1569,N_1441,N_1422);
nand U1570 (N_1570,N_1383,N_1485);
or U1571 (N_1571,N_1428,N_1426);
and U1572 (N_1572,N_1406,N_1419);
and U1573 (N_1573,N_1457,N_1425);
and U1574 (N_1574,N_1378,N_1476);
nand U1575 (N_1575,N_1381,N_1471);
and U1576 (N_1576,N_1486,N_1391);
and U1577 (N_1577,N_1451,N_1399);
or U1578 (N_1578,N_1482,N_1415);
and U1579 (N_1579,N_1438,N_1420);
nor U1580 (N_1580,N_1418,N_1416);
nor U1581 (N_1581,N_1398,N_1417);
nor U1582 (N_1582,N_1492,N_1424);
nor U1583 (N_1583,N_1446,N_1457);
nor U1584 (N_1584,N_1487,N_1460);
and U1585 (N_1585,N_1432,N_1434);
nor U1586 (N_1586,N_1409,N_1382);
and U1587 (N_1587,N_1399,N_1496);
nor U1588 (N_1588,N_1496,N_1452);
nor U1589 (N_1589,N_1415,N_1420);
and U1590 (N_1590,N_1466,N_1398);
or U1591 (N_1591,N_1401,N_1426);
nand U1592 (N_1592,N_1492,N_1497);
and U1593 (N_1593,N_1396,N_1410);
xor U1594 (N_1594,N_1475,N_1493);
nor U1595 (N_1595,N_1417,N_1397);
or U1596 (N_1596,N_1462,N_1385);
nor U1597 (N_1597,N_1442,N_1398);
nor U1598 (N_1598,N_1442,N_1444);
and U1599 (N_1599,N_1458,N_1494);
or U1600 (N_1600,N_1437,N_1443);
nand U1601 (N_1601,N_1489,N_1433);
nor U1602 (N_1602,N_1402,N_1462);
or U1603 (N_1603,N_1474,N_1473);
and U1604 (N_1604,N_1386,N_1397);
or U1605 (N_1605,N_1400,N_1444);
and U1606 (N_1606,N_1489,N_1403);
and U1607 (N_1607,N_1408,N_1403);
or U1608 (N_1608,N_1381,N_1464);
nor U1609 (N_1609,N_1475,N_1392);
xnor U1610 (N_1610,N_1432,N_1459);
nor U1611 (N_1611,N_1419,N_1430);
nor U1612 (N_1612,N_1406,N_1481);
and U1613 (N_1613,N_1490,N_1423);
and U1614 (N_1614,N_1481,N_1489);
nor U1615 (N_1615,N_1419,N_1494);
nand U1616 (N_1616,N_1398,N_1379);
or U1617 (N_1617,N_1375,N_1444);
nand U1618 (N_1618,N_1418,N_1393);
nand U1619 (N_1619,N_1479,N_1405);
and U1620 (N_1620,N_1382,N_1475);
or U1621 (N_1621,N_1480,N_1388);
or U1622 (N_1622,N_1383,N_1421);
nor U1623 (N_1623,N_1483,N_1447);
nor U1624 (N_1624,N_1398,N_1387);
nand U1625 (N_1625,N_1563,N_1614);
nand U1626 (N_1626,N_1531,N_1560);
xor U1627 (N_1627,N_1525,N_1543);
nand U1628 (N_1628,N_1598,N_1597);
xnor U1629 (N_1629,N_1613,N_1565);
or U1630 (N_1630,N_1576,N_1617);
nor U1631 (N_1631,N_1610,N_1522);
and U1632 (N_1632,N_1594,N_1545);
nor U1633 (N_1633,N_1514,N_1524);
or U1634 (N_1634,N_1502,N_1546);
and U1635 (N_1635,N_1612,N_1507);
or U1636 (N_1636,N_1585,N_1537);
or U1637 (N_1637,N_1515,N_1535);
and U1638 (N_1638,N_1561,N_1554);
nor U1639 (N_1639,N_1582,N_1508);
or U1640 (N_1640,N_1606,N_1574);
nand U1641 (N_1641,N_1590,N_1505);
or U1642 (N_1642,N_1622,N_1602);
and U1643 (N_1643,N_1564,N_1586);
and U1644 (N_1644,N_1618,N_1609);
nor U1645 (N_1645,N_1501,N_1527);
or U1646 (N_1646,N_1542,N_1549);
nor U1647 (N_1647,N_1568,N_1605);
and U1648 (N_1648,N_1575,N_1550);
nor U1649 (N_1649,N_1601,N_1553);
xnor U1650 (N_1650,N_1552,N_1504);
and U1651 (N_1651,N_1623,N_1581);
or U1652 (N_1652,N_1580,N_1562);
and U1653 (N_1653,N_1556,N_1533);
nand U1654 (N_1654,N_1595,N_1513);
and U1655 (N_1655,N_1578,N_1607);
and U1656 (N_1656,N_1512,N_1587);
or U1657 (N_1657,N_1511,N_1567);
xor U1658 (N_1658,N_1571,N_1534);
and U1659 (N_1659,N_1620,N_1583);
or U1660 (N_1660,N_1555,N_1519);
xor U1661 (N_1661,N_1593,N_1570);
or U1662 (N_1662,N_1608,N_1538);
and U1663 (N_1663,N_1516,N_1624);
nor U1664 (N_1664,N_1604,N_1569);
or U1665 (N_1665,N_1579,N_1592);
xor U1666 (N_1666,N_1599,N_1559);
or U1667 (N_1667,N_1573,N_1572);
nor U1668 (N_1668,N_1577,N_1521);
nand U1669 (N_1669,N_1621,N_1544);
nand U1670 (N_1670,N_1503,N_1541);
xnor U1671 (N_1671,N_1603,N_1520);
nand U1672 (N_1672,N_1529,N_1540);
or U1673 (N_1673,N_1532,N_1528);
and U1674 (N_1674,N_1539,N_1551);
nand U1675 (N_1675,N_1548,N_1500);
or U1676 (N_1676,N_1518,N_1530);
and U1677 (N_1677,N_1619,N_1616);
nand U1678 (N_1678,N_1557,N_1510);
nor U1679 (N_1679,N_1509,N_1589);
nand U1680 (N_1680,N_1523,N_1596);
nor U1681 (N_1681,N_1517,N_1506);
and U1682 (N_1682,N_1547,N_1526);
nor U1683 (N_1683,N_1611,N_1584);
or U1684 (N_1684,N_1566,N_1536);
nor U1685 (N_1685,N_1600,N_1615);
xor U1686 (N_1686,N_1558,N_1588);
nor U1687 (N_1687,N_1591,N_1584);
and U1688 (N_1688,N_1546,N_1607);
or U1689 (N_1689,N_1562,N_1518);
and U1690 (N_1690,N_1501,N_1604);
xnor U1691 (N_1691,N_1536,N_1543);
and U1692 (N_1692,N_1537,N_1618);
xnor U1693 (N_1693,N_1597,N_1518);
and U1694 (N_1694,N_1511,N_1542);
and U1695 (N_1695,N_1582,N_1600);
or U1696 (N_1696,N_1564,N_1502);
or U1697 (N_1697,N_1617,N_1572);
nand U1698 (N_1698,N_1549,N_1594);
or U1699 (N_1699,N_1623,N_1593);
and U1700 (N_1700,N_1551,N_1544);
or U1701 (N_1701,N_1604,N_1530);
and U1702 (N_1702,N_1542,N_1624);
and U1703 (N_1703,N_1563,N_1580);
nor U1704 (N_1704,N_1550,N_1610);
and U1705 (N_1705,N_1541,N_1612);
or U1706 (N_1706,N_1613,N_1588);
nand U1707 (N_1707,N_1620,N_1586);
or U1708 (N_1708,N_1560,N_1500);
nor U1709 (N_1709,N_1562,N_1552);
and U1710 (N_1710,N_1605,N_1511);
and U1711 (N_1711,N_1548,N_1503);
nand U1712 (N_1712,N_1528,N_1597);
or U1713 (N_1713,N_1616,N_1585);
and U1714 (N_1714,N_1574,N_1601);
nor U1715 (N_1715,N_1612,N_1611);
or U1716 (N_1716,N_1566,N_1558);
xnor U1717 (N_1717,N_1503,N_1578);
or U1718 (N_1718,N_1542,N_1600);
nand U1719 (N_1719,N_1578,N_1564);
nor U1720 (N_1720,N_1606,N_1557);
or U1721 (N_1721,N_1567,N_1580);
nor U1722 (N_1722,N_1586,N_1552);
xor U1723 (N_1723,N_1605,N_1514);
nand U1724 (N_1724,N_1541,N_1531);
or U1725 (N_1725,N_1618,N_1527);
nor U1726 (N_1726,N_1589,N_1605);
and U1727 (N_1727,N_1620,N_1615);
and U1728 (N_1728,N_1556,N_1576);
or U1729 (N_1729,N_1531,N_1610);
nor U1730 (N_1730,N_1524,N_1523);
or U1731 (N_1731,N_1616,N_1500);
xor U1732 (N_1732,N_1510,N_1623);
nor U1733 (N_1733,N_1564,N_1613);
nand U1734 (N_1734,N_1537,N_1619);
nor U1735 (N_1735,N_1584,N_1565);
or U1736 (N_1736,N_1545,N_1535);
and U1737 (N_1737,N_1512,N_1563);
or U1738 (N_1738,N_1539,N_1575);
xor U1739 (N_1739,N_1531,N_1512);
xor U1740 (N_1740,N_1604,N_1514);
nor U1741 (N_1741,N_1592,N_1536);
nand U1742 (N_1742,N_1546,N_1612);
nor U1743 (N_1743,N_1618,N_1608);
nand U1744 (N_1744,N_1541,N_1581);
and U1745 (N_1745,N_1550,N_1572);
xnor U1746 (N_1746,N_1514,N_1547);
nand U1747 (N_1747,N_1589,N_1526);
and U1748 (N_1748,N_1551,N_1565);
and U1749 (N_1749,N_1520,N_1539);
and U1750 (N_1750,N_1701,N_1684);
xor U1751 (N_1751,N_1717,N_1669);
nor U1752 (N_1752,N_1631,N_1689);
nand U1753 (N_1753,N_1737,N_1748);
and U1754 (N_1754,N_1749,N_1735);
or U1755 (N_1755,N_1636,N_1667);
nand U1756 (N_1756,N_1736,N_1661);
xor U1757 (N_1757,N_1668,N_1708);
nor U1758 (N_1758,N_1681,N_1706);
or U1759 (N_1759,N_1633,N_1743);
and U1760 (N_1760,N_1628,N_1682);
nor U1761 (N_1761,N_1625,N_1647);
and U1762 (N_1762,N_1665,N_1699);
nor U1763 (N_1763,N_1732,N_1675);
and U1764 (N_1764,N_1722,N_1634);
and U1765 (N_1765,N_1658,N_1719);
nor U1766 (N_1766,N_1640,N_1710);
or U1767 (N_1767,N_1679,N_1729);
and U1768 (N_1768,N_1680,N_1704);
or U1769 (N_1769,N_1730,N_1683);
nor U1770 (N_1770,N_1738,N_1645);
and U1771 (N_1771,N_1635,N_1663);
or U1772 (N_1772,N_1688,N_1739);
nand U1773 (N_1773,N_1692,N_1639);
nand U1774 (N_1774,N_1711,N_1662);
or U1775 (N_1775,N_1659,N_1698);
and U1776 (N_1776,N_1642,N_1672);
and U1777 (N_1777,N_1673,N_1720);
and U1778 (N_1778,N_1724,N_1670);
nor U1779 (N_1779,N_1686,N_1726);
and U1780 (N_1780,N_1745,N_1637);
nand U1781 (N_1781,N_1644,N_1705);
nor U1782 (N_1782,N_1653,N_1687);
and U1783 (N_1783,N_1742,N_1696);
nand U1784 (N_1784,N_1649,N_1676);
and U1785 (N_1785,N_1666,N_1660);
nor U1786 (N_1786,N_1733,N_1657);
nor U1787 (N_1787,N_1664,N_1626);
nand U1788 (N_1788,N_1671,N_1654);
nand U1789 (N_1789,N_1685,N_1655);
nand U1790 (N_1790,N_1656,N_1650);
and U1791 (N_1791,N_1648,N_1652);
and U1792 (N_1792,N_1721,N_1714);
or U1793 (N_1793,N_1646,N_1746);
nor U1794 (N_1794,N_1627,N_1695);
xnor U1795 (N_1795,N_1630,N_1641);
nand U1796 (N_1796,N_1740,N_1744);
nand U1797 (N_1797,N_1651,N_1747);
nor U1798 (N_1798,N_1638,N_1703);
nor U1799 (N_1799,N_1674,N_1731);
nand U1800 (N_1800,N_1713,N_1691);
xnor U1801 (N_1801,N_1728,N_1643);
xor U1802 (N_1802,N_1693,N_1694);
or U1803 (N_1803,N_1702,N_1718);
nand U1804 (N_1804,N_1677,N_1709);
or U1805 (N_1805,N_1723,N_1712);
nand U1806 (N_1806,N_1700,N_1632);
and U1807 (N_1807,N_1725,N_1715);
nor U1808 (N_1808,N_1690,N_1707);
nand U1809 (N_1809,N_1716,N_1734);
and U1810 (N_1810,N_1697,N_1727);
nor U1811 (N_1811,N_1629,N_1741);
nor U1812 (N_1812,N_1678,N_1744);
nand U1813 (N_1813,N_1674,N_1707);
xor U1814 (N_1814,N_1688,N_1655);
and U1815 (N_1815,N_1686,N_1707);
nand U1816 (N_1816,N_1652,N_1691);
nand U1817 (N_1817,N_1719,N_1727);
nor U1818 (N_1818,N_1723,N_1651);
or U1819 (N_1819,N_1738,N_1747);
nor U1820 (N_1820,N_1709,N_1743);
and U1821 (N_1821,N_1638,N_1636);
or U1822 (N_1822,N_1645,N_1713);
or U1823 (N_1823,N_1748,N_1717);
xor U1824 (N_1824,N_1668,N_1663);
or U1825 (N_1825,N_1746,N_1685);
or U1826 (N_1826,N_1734,N_1696);
and U1827 (N_1827,N_1717,N_1666);
and U1828 (N_1828,N_1692,N_1698);
nor U1829 (N_1829,N_1675,N_1701);
or U1830 (N_1830,N_1638,N_1732);
nand U1831 (N_1831,N_1726,N_1709);
and U1832 (N_1832,N_1633,N_1720);
nor U1833 (N_1833,N_1685,N_1635);
and U1834 (N_1834,N_1715,N_1640);
nor U1835 (N_1835,N_1681,N_1741);
nor U1836 (N_1836,N_1714,N_1671);
nand U1837 (N_1837,N_1659,N_1643);
and U1838 (N_1838,N_1674,N_1630);
and U1839 (N_1839,N_1742,N_1711);
and U1840 (N_1840,N_1668,N_1680);
nor U1841 (N_1841,N_1631,N_1741);
nor U1842 (N_1842,N_1736,N_1630);
or U1843 (N_1843,N_1688,N_1705);
or U1844 (N_1844,N_1649,N_1626);
nand U1845 (N_1845,N_1726,N_1646);
and U1846 (N_1846,N_1727,N_1637);
or U1847 (N_1847,N_1742,N_1743);
or U1848 (N_1848,N_1707,N_1654);
or U1849 (N_1849,N_1649,N_1682);
nor U1850 (N_1850,N_1694,N_1745);
and U1851 (N_1851,N_1668,N_1657);
nand U1852 (N_1852,N_1710,N_1656);
nor U1853 (N_1853,N_1732,N_1722);
or U1854 (N_1854,N_1736,N_1737);
and U1855 (N_1855,N_1709,N_1729);
or U1856 (N_1856,N_1659,N_1628);
and U1857 (N_1857,N_1742,N_1703);
nor U1858 (N_1858,N_1717,N_1625);
and U1859 (N_1859,N_1712,N_1675);
nor U1860 (N_1860,N_1713,N_1670);
or U1861 (N_1861,N_1670,N_1710);
nor U1862 (N_1862,N_1680,N_1689);
nor U1863 (N_1863,N_1692,N_1709);
nor U1864 (N_1864,N_1646,N_1714);
and U1865 (N_1865,N_1709,N_1686);
nor U1866 (N_1866,N_1733,N_1743);
xnor U1867 (N_1867,N_1631,N_1642);
or U1868 (N_1868,N_1629,N_1714);
or U1869 (N_1869,N_1714,N_1694);
or U1870 (N_1870,N_1673,N_1700);
or U1871 (N_1871,N_1720,N_1689);
and U1872 (N_1872,N_1737,N_1706);
and U1873 (N_1873,N_1681,N_1684);
nor U1874 (N_1874,N_1733,N_1727);
nor U1875 (N_1875,N_1841,N_1777);
nand U1876 (N_1876,N_1766,N_1773);
or U1877 (N_1877,N_1852,N_1823);
xor U1878 (N_1878,N_1849,N_1838);
and U1879 (N_1879,N_1847,N_1784);
or U1880 (N_1880,N_1820,N_1833);
nor U1881 (N_1881,N_1768,N_1753);
or U1882 (N_1882,N_1857,N_1850);
nor U1883 (N_1883,N_1756,N_1818);
or U1884 (N_1884,N_1815,N_1826);
nor U1885 (N_1885,N_1785,N_1861);
xnor U1886 (N_1886,N_1757,N_1835);
and U1887 (N_1887,N_1804,N_1810);
and U1888 (N_1888,N_1869,N_1872);
nand U1889 (N_1889,N_1811,N_1814);
and U1890 (N_1890,N_1769,N_1798);
and U1891 (N_1891,N_1870,N_1824);
or U1892 (N_1892,N_1863,N_1802);
or U1893 (N_1893,N_1764,N_1755);
nor U1894 (N_1894,N_1817,N_1827);
nor U1895 (N_1895,N_1874,N_1873);
or U1896 (N_1896,N_1828,N_1867);
nor U1897 (N_1897,N_1792,N_1839);
nor U1898 (N_1898,N_1853,N_1801);
and U1899 (N_1899,N_1866,N_1845);
or U1900 (N_1900,N_1796,N_1805);
and U1901 (N_1901,N_1779,N_1859);
nand U1902 (N_1902,N_1761,N_1786);
and U1903 (N_1903,N_1812,N_1807);
xor U1904 (N_1904,N_1832,N_1770);
nand U1905 (N_1905,N_1758,N_1848);
nor U1906 (N_1906,N_1809,N_1836);
or U1907 (N_1907,N_1868,N_1825);
nor U1908 (N_1908,N_1771,N_1821);
nand U1909 (N_1909,N_1808,N_1787);
nand U1910 (N_1910,N_1799,N_1762);
xor U1911 (N_1911,N_1759,N_1772);
nor U1912 (N_1912,N_1760,N_1765);
nand U1913 (N_1913,N_1837,N_1862);
nand U1914 (N_1914,N_1819,N_1822);
and U1915 (N_1915,N_1803,N_1842);
and U1916 (N_1916,N_1781,N_1795);
and U1917 (N_1917,N_1754,N_1794);
and U1918 (N_1918,N_1865,N_1791);
or U1919 (N_1919,N_1855,N_1783);
nor U1920 (N_1920,N_1752,N_1846);
or U1921 (N_1921,N_1830,N_1864);
or U1922 (N_1922,N_1816,N_1840);
nand U1923 (N_1923,N_1793,N_1750);
nor U1924 (N_1924,N_1790,N_1797);
nor U1925 (N_1925,N_1789,N_1788);
or U1926 (N_1926,N_1780,N_1858);
and U1927 (N_1927,N_1813,N_1856);
nand U1928 (N_1928,N_1776,N_1782);
or U1929 (N_1929,N_1854,N_1763);
nor U1930 (N_1930,N_1843,N_1844);
nand U1931 (N_1931,N_1751,N_1774);
nor U1932 (N_1932,N_1775,N_1851);
and U1933 (N_1933,N_1800,N_1806);
nor U1934 (N_1934,N_1860,N_1829);
nor U1935 (N_1935,N_1831,N_1834);
nor U1936 (N_1936,N_1778,N_1871);
nand U1937 (N_1937,N_1767,N_1831);
nand U1938 (N_1938,N_1762,N_1848);
and U1939 (N_1939,N_1870,N_1809);
or U1940 (N_1940,N_1803,N_1772);
and U1941 (N_1941,N_1799,N_1760);
and U1942 (N_1942,N_1817,N_1799);
nor U1943 (N_1943,N_1790,N_1805);
nor U1944 (N_1944,N_1760,N_1843);
nand U1945 (N_1945,N_1854,N_1791);
nand U1946 (N_1946,N_1784,N_1785);
and U1947 (N_1947,N_1771,N_1853);
or U1948 (N_1948,N_1811,N_1783);
xnor U1949 (N_1949,N_1769,N_1791);
nand U1950 (N_1950,N_1817,N_1824);
nand U1951 (N_1951,N_1831,N_1865);
nor U1952 (N_1952,N_1774,N_1771);
nor U1953 (N_1953,N_1757,N_1759);
nor U1954 (N_1954,N_1820,N_1769);
nand U1955 (N_1955,N_1840,N_1828);
nand U1956 (N_1956,N_1787,N_1845);
nand U1957 (N_1957,N_1751,N_1856);
and U1958 (N_1958,N_1779,N_1870);
xor U1959 (N_1959,N_1783,N_1750);
nand U1960 (N_1960,N_1803,N_1831);
nand U1961 (N_1961,N_1776,N_1751);
nand U1962 (N_1962,N_1822,N_1804);
or U1963 (N_1963,N_1851,N_1872);
and U1964 (N_1964,N_1792,N_1794);
nor U1965 (N_1965,N_1802,N_1853);
nand U1966 (N_1966,N_1808,N_1798);
and U1967 (N_1967,N_1796,N_1819);
nor U1968 (N_1968,N_1802,N_1858);
or U1969 (N_1969,N_1822,N_1871);
nor U1970 (N_1970,N_1857,N_1782);
and U1971 (N_1971,N_1799,N_1826);
nor U1972 (N_1972,N_1843,N_1804);
nor U1973 (N_1973,N_1772,N_1829);
or U1974 (N_1974,N_1823,N_1798);
and U1975 (N_1975,N_1762,N_1871);
xnor U1976 (N_1976,N_1787,N_1779);
or U1977 (N_1977,N_1850,N_1860);
and U1978 (N_1978,N_1750,N_1839);
nand U1979 (N_1979,N_1865,N_1769);
or U1980 (N_1980,N_1836,N_1863);
nand U1981 (N_1981,N_1783,N_1804);
nand U1982 (N_1982,N_1756,N_1826);
nor U1983 (N_1983,N_1828,N_1796);
nor U1984 (N_1984,N_1855,N_1823);
nor U1985 (N_1985,N_1809,N_1768);
nor U1986 (N_1986,N_1776,N_1852);
nand U1987 (N_1987,N_1820,N_1797);
xor U1988 (N_1988,N_1853,N_1752);
nand U1989 (N_1989,N_1847,N_1825);
and U1990 (N_1990,N_1764,N_1765);
nand U1991 (N_1991,N_1832,N_1836);
and U1992 (N_1992,N_1854,N_1817);
and U1993 (N_1993,N_1869,N_1785);
xnor U1994 (N_1994,N_1802,N_1867);
and U1995 (N_1995,N_1793,N_1784);
or U1996 (N_1996,N_1812,N_1771);
nand U1997 (N_1997,N_1857,N_1767);
nor U1998 (N_1998,N_1846,N_1833);
and U1999 (N_1999,N_1858,N_1778);
and U2000 (N_2000,N_1895,N_1980);
nand U2001 (N_2001,N_1961,N_1940);
or U2002 (N_2002,N_1970,N_1936);
nor U2003 (N_2003,N_1950,N_1998);
and U2004 (N_2004,N_1900,N_1888);
and U2005 (N_2005,N_1886,N_1892);
or U2006 (N_2006,N_1987,N_1994);
nand U2007 (N_2007,N_1880,N_1971);
xor U2008 (N_2008,N_1929,N_1930);
and U2009 (N_2009,N_1915,N_1974);
xor U2010 (N_2010,N_1899,N_1889);
nor U2011 (N_2011,N_1938,N_1965);
and U2012 (N_2012,N_1977,N_1964);
nand U2013 (N_2013,N_1944,N_1924);
nand U2014 (N_2014,N_1932,N_1942);
or U2015 (N_2015,N_1920,N_1887);
or U2016 (N_2016,N_1962,N_1960);
nor U2017 (N_2017,N_1957,N_1991);
xor U2018 (N_2018,N_1934,N_1947);
nor U2019 (N_2019,N_1952,N_1933);
or U2020 (N_2020,N_1926,N_1875);
or U2021 (N_2021,N_1969,N_1978);
and U2022 (N_2022,N_1959,N_1877);
nor U2023 (N_2023,N_1979,N_1997);
or U2024 (N_2024,N_1999,N_1975);
or U2025 (N_2025,N_1984,N_1927);
nand U2026 (N_2026,N_1911,N_1966);
or U2027 (N_2027,N_1990,N_1890);
and U2028 (N_2028,N_1909,N_1879);
nor U2029 (N_2029,N_1878,N_1919);
nand U2030 (N_2030,N_1925,N_1935);
nand U2031 (N_2031,N_1923,N_1901);
and U2032 (N_2032,N_1913,N_1954);
or U2033 (N_2033,N_1943,N_1955);
nor U2034 (N_2034,N_1912,N_1983);
and U2035 (N_2035,N_1956,N_1885);
nor U2036 (N_2036,N_1905,N_1906);
or U2037 (N_2037,N_1893,N_1985);
xor U2038 (N_2038,N_1894,N_1949);
or U2039 (N_2039,N_1903,N_1946);
and U2040 (N_2040,N_1988,N_1918);
xnor U2041 (N_2041,N_1881,N_1972);
xor U2042 (N_2042,N_1922,N_1907);
xor U2043 (N_2043,N_1883,N_1921);
or U2044 (N_2044,N_1882,N_1916);
nor U2045 (N_2045,N_1902,N_1884);
or U2046 (N_2046,N_1891,N_1897);
or U2047 (N_2047,N_1995,N_1993);
or U2048 (N_2048,N_1973,N_1982);
and U2049 (N_2049,N_1996,N_1908);
nor U2050 (N_2050,N_1928,N_1931);
xor U2051 (N_2051,N_1986,N_1941);
or U2052 (N_2052,N_1898,N_1989);
nand U2053 (N_2053,N_1963,N_1896);
nand U2054 (N_2054,N_1917,N_1937);
nand U2055 (N_2055,N_1904,N_1981);
xor U2056 (N_2056,N_1945,N_1914);
nand U2057 (N_2057,N_1992,N_1958);
nor U2058 (N_2058,N_1968,N_1976);
nand U2059 (N_2059,N_1939,N_1967);
or U2060 (N_2060,N_1953,N_1951);
or U2061 (N_2061,N_1948,N_1910);
and U2062 (N_2062,N_1876,N_1958);
nor U2063 (N_2063,N_1984,N_1985);
nor U2064 (N_2064,N_1887,N_1907);
nand U2065 (N_2065,N_1904,N_1940);
and U2066 (N_2066,N_1904,N_1971);
or U2067 (N_2067,N_1995,N_1964);
xnor U2068 (N_2068,N_1955,N_1909);
nor U2069 (N_2069,N_1975,N_1955);
and U2070 (N_2070,N_1988,N_1909);
nor U2071 (N_2071,N_1950,N_1894);
nor U2072 (N_2072,N_1875,N_1924);
or U2073 (N_2073,N_1935,N_1978);
nor U2074 (N_2074,N_1881,N_1923);
and U2075 (N_2075,N_1975,N_1881);
nor U2076 (N_2076,N_1991,N_1968);
nand U2077 (N_2077,N_1894,N_1996);
and U2078 (N_2078,N_1888,N_1988);
or U2079 (N_2079,N_1947,N_1893);
nand U2080 (N_2080,N_1898,N_1923);
and U2081 (N_2081,N_1950,N_1976);
nand U2082 (N_2082,N_1889,N_1929);
nor U2083 (N_2083,N_1931,N_1998);
nand U2084 (N_2084,N_1924,N_1999);
nor U2085 (N_2085,N_1953,N_1893);
or U2086 (N_2086,N_1899,N_1977);
and U2087 (N_2087,N_1944,N_1967);
xor U2088 (N_2088,N_1938,N_1916);
and U2089 (N_2089,N_1911,N_1961);
nand U2090 (N_2090,N_1914,N_1935);
nand U2091 (N_2091,N_1941,N_1935);
nand U2092 (N_2092,N_1942,N_1893);
xnor U2093 (N_2093,N_1930,N_1907);
or U2094 (N_2094,N_1891,N_1947);
and U2095 (N_2095,N_1957,N_1955);
nand U2096 (N_2096,N_1989,N_1998);
nand U2097 (N_2097,N_1876,N_1964);
xor U2098 (N_2098,N_1926,N_1895);
and U2099 (N_2099,N_1944,N_1936);
xnor U2100 (N_2100,N_1948,N_1884);
nand U2101 (N_2101,N_1950,N_1992);
nor U2102 (N_2102,N_1889,N_1911);
or U2103 (N_2103,N_1962,N_1879);
and U2104 (N_2104,N_1886,N_1913);
nor U2105 (N_2105,N_1919,N_1891);
or U2106 (N_2106,N_1973,N_1954);
and U2107 (N_2107,N_1909,N_1941);
and U2108 (N_2108,N_1990,N_1994);
nand U2109 (N_2109,N_1949,N_1954);
or U2110 (N_2110,N_1876,N_1931);
and U2111 (N_2111,N_1930,N_1944);
or U2112 (N_2112,N_1935,N_1880);
or U2113 (N_2113,N_1963,N_1937);
nand U2114 (N_2114,N_1893,N_1936);
and U2115 (N_2115,N_1896,N_1990);
xor U2116 (N_2116,N_1991,N_1958);
or U2117 (N_2117,N_1947,N_1909);
and U2118 (N_2118,N_1978,N_1900);
and U2119 (N_2119,N_1995,N_1952);
nand U2120 (N_2120,N_1993,N_1911);
xnor U2121 (N_2121,N_1924,N_1910);
or U2122 (N_2122,N_1888,N_1921);
nor U2123 (N_2123,N_1967,N_1884);
nand U2124 (N_2124,N_1946,N_1935);
nor U2125 (N_2125,N_2075,N_2085);
and U2126 (N_2126,N_2053,N_2081);
and U2127 (N_2127,N_2003,N_2076);
or U2128 (N_2128,N_2035,N_2115);
nor U2129 (N_2129,N_2088,N_2110);
nor U2130 (N_2130,N_2008,N_2052);
and U2131 (N_2131,N_2106,N_2108);
xnor U2132 (N_2132,N_2020,N_2036);
and U2133 (N_2133,N_2065,N_2119);
nor U2134 (N_2134,N_2014,N_2006);
nand U2135 (N_2135,N_2021,N_2074);
nor U2136 (N_2136,N_2078,N_2120);
nor U2137 (N_2137,N_2079,N_2044);
nor U2138 (N_2138,N_2045,N_2117);
nor U2139 (N_2139,N_2093,N_2097);
and U2140 (N_2140,N_2041,N_2051);
nor U2141 (N_2141,N_2090,N_2011);
nand U2142 (N_2142,N_2094,N_2015);
or U2143 (N_2143,N_2038,N_2025);
or U2144 (N_2144,N_2103,N_2019);
and U2145 (N_2145,N_2027,N_2050);
and U2146 (N_2146,N_2064,N_2067);
nand U2147 (N_2147,N_2086,N_2016);
or U2148 (N_2148,N_2084,N_2013);
nor U2149 (N_2149,N_2005,N_2105);
nor U2150 (N_2150,N_2091,N_2007);
nor U2151 (N_2151,N_2055,N_2037);
xnor U2152 (N_2152,N_2002,N_2107);
or U2153 (N_2153,N_2089,N_2073);
nand U2154 (N_2154,N_2111,N_2069);
and U2155 (N_2155,N_2121,N_2012);
and U2156 (N_2156,N_2054,N_2018);
nand U2157 (N_2157,N_2048,N_2062);
nand U2158 (N_2158,N_2063,N_2001);
nor U2159 (N_2159,N_2118,N_2109);
or U2160 (N_2160,N_2095,N_2028);
nand U2161 (N_2161,N_2010,N_2026);
nor U2162 (N_2162,N_2022,N_2082);
or U2163 (N_2163,N_2043,N_2100);
and U2164 (N_2164,N_2123,N_2057);
nand U2165 (N_2165,N_2059,N_2099);
and U2166 (N_2166,N_2004,N_2080);
nor U2167 (N_2167,N_2000,N_2077);
and U2168 (N_2168,N_2071,N_2058);
xor U2169 (N_2169,N_2070,N_2046);
and U2170 (N_2170,N_2009,N_2124);
or U2171 (N_2171,N_2092,N_2061);
or U2172 (N_2172,N_2031,N_2042);
nor U2173 (N_2173,N_2024,N_2032);
and U2174 (N_2174,N_2096,N_2114);
or U2175 (N_2175,N_2029,N_2034);
nor U2176 (N_2176,N_2102,N_2056);
nand U2177 (N_2177,N_2030,N_2116);
and U2178 (N_2178,N_2072,N_2098);
nand U2179 (N_2179,N_2033,N_2060);
or U2180 (N_2180,N_2047,N_2066);
and U2181 (N_2181,N_2112,N_2083);
or U2182 (N_2182,N_2040,N_2039);
or U2183 (N_2183,N_2101,N_2104);
or U2184 (N_2184,N_2113,N_2122);
nand U2185 (N_2185,N_2087,N_2017);
and U2186 (N_2186,N_2023,N_2049);
nor U2187 (N_2187,N_2068,N_2033);
and U2188 (N_2188,N_2067,N_2028);
and U2189 (N_2189,N_2027,N_2007);
and U2190 (N_2190,N_2067,N_2059);
xnor U2191 (N_2191,N_2050,N_2065);
xor U2192 (N_2192,N_2120,N_2094);
nor U2193 (N_2193,N_2056,N_2064);
xnor U2194 (N_2194,N_2061,N_2068);
nand U2195 (N_2195,N_2120,N_2095);
or U2196 (N_2196,N_2085,N_2097);
nor U2197 (N_2197,N_2123,N_2016);
nand U2198 (N_2198,N_2022,N_2119);
nor U2199 (N_2199,N_2080,N_2051);
nand U2200 (N_2200,N_2106,N_2050);
nor U2201 (N_2201,N_2034,N_2099);
or U2202 (N_2202,N_2053,N_2099);
nor U2203 (N_2203,N_2081,N_2004);
or U2204 (N_2204,N_2029,N_2103);
or U2205 (N_2205,N_2052,N_2001);
and U2206 (N_2206,N_2086,N_2077);
and U2207 (N_2207,N_2095,N_2043);
or U2208 (N_2208,N_2025,N_2059);
and U2209 (N_2209,N_2087,N_2051);
xnor U2210 (N_2210,N_2010,N_2017);
or U2211 (N_2211,N_2033,N_2047);
and U2212 (N_2212,N_2000,N_2043);
nor U2213 (N_2213,N_2017,N_2015);
nor U2214 (N_2214,N_2089,N_2045);
nand U2215 (N_2215,N_2097,N_2059);
nand U2216 (N_2216,N_2044,N_2093);
nand U2217 (N_2217,N_2076,N_2024);
nand U2218 (N_2218,N_2018,N_2010);
nor U2219 (N_2219,N_2055,N_2025);
nand U2220 (N_2220,N_2062,N_2023);
or U2221 (N_2221,N_2083,N_2040);
or U2222 (N_2222,N_2080,N_2045);
nor U2223 (N_2223,N_2045,N_2099);
nand U2224 (N_2224,N_2088,N_2059);
nor U2225 (N_2225,N_2078,N_2053);
and U2226 (N_2226,N_2012,N_2124);
xnor U2227 (N_2227,N_2004,N_2002);
and U2228 (N_2228,N_2046,N_2105);
nor U2229 (N_2229,N_2066,N_2059);
or U2230 (N_2230,N_2110,N_2109);
xnor U2231 (N_2231,N_2058,N_2036);
nor U2232 (N_2232,N_2004,N_2069);
and U2233 (N_2233,N_2026,N_2110);
and U2234 (N_2234,N_2113,N_2082);
and U2235 (N_2235,N_2122,N_2029);
and U2236 (N_2236,N_2085,N_2021);
and U2237 (N_2237,N_2055,N_2058);
and U2238 (N_2238,N_2033,N_2086);
nor U2239 (N_2239,N_2113,N_2107);
nand U2240 (N_2240,N_2001,N_2058);
nand U2241 (N_2241,N_2124,N_2085);
nand U2242 (N_2242,N_2065,N_2115);
and U2243 (N_2243,N_2116,N_2086);
and U2244 (N_2244,N_2096,N_2001);
or U2245 (N_2245,N_2055,N_2002);
nor U2246 (N_2246,N_2048,N_2099);
nor U2247 (N_2247,N_2110,N_2047);
xnor U2248 (N_2248,N_2105,N_2010);
xor U2249 (N_2249,N_2046,N_2085);
xnor U2250 (N_2250,N_2187,N_2180);
or U2251 (N_2251,N_2179,N_2155);
nor U2252 (N_2252,N_2161,N_2197);
nor U2253 (N_2253,N_2243,N_2219);
xnor U2254 (N_2254,N_2249,N_2218);
nand U2255 (N_2255,N_2138,N_2184);
and U2256 (N_2256,N_2168,N_2225);
and U2257 (N_2257,N_2231,N_2191);
or U2258 (N_2258,N_2166,N_2227);
nand U2259 (N_2259,N_2143,N_2229);
and U2260 (N_2260,N_2212,N_2159);
or U2261 (N_2261,N_2128,N_2148);
or U2262 (N_2262,N_2190,N_2196);
xnor U2263 (N_2263,N_2223,N_2172);
nor U2264 (N_2264,N_2162,N_2156);
nor U2265 (N_2265,N_2239,N_2169);
nand U2266 (N_2266,N_2207,N_2137);
and U2267 (N_2267,N_2226,N_2240);
or U2268 (N_2268,N_2147,N_2228);
nand U2269 (N_2269,N_2130,N_2200);
and U2270 (N_2270,N_2189,N_2158);
or U2271 (N_2271,N_2176,N_2213);
xor U2272 (N_2272,N_2133,N_2193);
xor U2273 (N_2273,N_2188,N_2224);
nand U2274 (N_2274,N_2167,N_2208);
nand U2275 (N_2275,N_2248,N_2242);
or U2276 (N_2276,N_2203,N_2237);
and U2277 (N_2277,N_2163,N_2150);
nor U2278 (N_2278,N_2129,N_2205);
nor U2279 (N_2279,N_2173,N_2145);
nand U2280 (N_2280,N_2195,N_2233);
or U2281 (N_2281,N_2181,N_2211);
nand U2282 (N_2282,N_2135,N_2127);
and U2283 (N_2283,N_2220,N_2178);
xor U2284 (N_2284,N_2154,N_2132);
nand U2285 (N_2285,N_2182,N_2202);
nor U2286 (N_2286,N_2183,N_2194);
or U2287 (N_2287,N_2185,N_2140);
xor U2288 (N_2288,N_2215,N_2192);
xnor U2289 (N_2289,N_2198,N_2216);
and U2290 (N_2290,N_2247,N_2165);
or U2291 (N_2291,N_2238,N_2142);
nor U2292 (N_2292,N_2139,N_2186);
and U2293 (N_2293,N_2199,N_2146);
nor U2294 (N_2294,N_2234,N_2149);
or U2295 (N_2295,N_2210,N_2126);
nand U2296 (N_2296,N_2235,N_2209);
or U2297 (N_2297,N_2170,N_2125);
nand U2298 (N_2298,N_2204,N_2206);
and U2299 (N_2299,N_2232,N_2144);
xnor U2300 (N_2300,N_2153,N_2236);
nand U2301 (N_2301,N_2134,N_2244);
or U2302 (N_2302,N_2136,N_2141);
nand U2303 (N_2303,N_2230,N_2151);
nand U2304 (N_2304,N_2152,N_2177);
nor U2305 (N_2305,N_2171,N_2214);
xor U2306 (N_2306,N_2131,N_2164);
or U2307 (N_2307,N_2222,N_2217);
or U2308 (N_2308,N_2221,N_2246);
or U2309 (N_2309,N_2157,N_2174);
and U2310 (N_2310,N_2245,N_2241);
nand U2311 (N_2311,N_2175,N_2160);
or U2312 (N_2312,N_2201,N_2200);
nor U2313 (N_2313,N_2177,N_2226);
or U2314 (N_2314,N_2175,N_2194);
and U2315 (N_2315,N_2168,N_2161);
nand U2316 (N_2316,N_2172,N_2128);
nand U2317 (N_2317,N_2210,N_2186);
nor U2318 (N_2318,N_2183,N_2205);
nor U2319 (N_2319,N_2243,N_2173);
and U2320 (N_2320,N_2183,N_2228);
and U2321 (N_2321,N_2187,N_2175);
nand U2322 (N_2322,N_2172,N_2247);
and U2323 (N_2323,N_2169,N_2182);
nand U2324 (N_2324,N_2142,N_2209);
or U2325 (N_2325,N_2181,N_2232);
xnor U2326 (N_2326,N_2242,N_2197);
or U2327 (N_2327,N_2177,N_2244);
nand U2328 (N_2328,N_2178,N_2217);
or U2329 (N_2329,N_2156,N_2207);
and U2330 (N_2330,N_2215,N_2156);
or U2331 (N_2331,N_2233,N_2215);
xor U2332 (N_2332,N_2177,N_2141);
and U2333 (N_2333,N_2220,N_2168);
nand U2334 (N_2334,N_2158,N_2202);
nand U2335 (N_2335,N_2184,N_2243);
nor U2336 (N_2336,N_2152,N_2190);
or U2337 (N_2337,N_2156,N_2238);
xnor U2338 (N_2338,N_2169,N_2200);
or U2339 (N_2339,N_2133,N_2228);
nor U2340 (N_2340,N_2163,N_2131);
nor U2341 (N_2341,N_2181,N_2152);
xnor U2342 (N_2342,N_2177,N_2236);
nand U2343 (N_2343,N_2236,N_2150);
or U2344 (N_2344,N_2169,N_2130);
nor U2345 (N_2345,N_2196,N_2153);
nand U2346 (N_2346,N_2239,N_2225);
nand U2347 (N_2347,N_2158,N_2171);
or U2348 (N_2348,N_2198,N_2215);
and U2349 (N_2349,N_2235,N_2143);
or U2350 (N_2350,N_2149,N_2247);
and U2351 (N_2351,N_2180,N_2204);
and U2352 (N_2352,N_2173,N_2170);
and U2353 (N_2353,N_2134,N_2213);
nor U2354 (N_2354,N_2148,N_2212);
nor U2355 (N_2355,N_2216,N_2127);
and U2356 (N_2356,N_2174,N_2201);
nor U2357 (N_2357,N_2170,N_2242);
or U2358 (N_2358,N_2155,N_2173);
nor U2359 (N_2359,N_2206,N_2184);
xor U2360 (N_2360,N_2149,N_2171);
or U2361 (N_2361,N_2129,N_2151);
nand U2362 (N_2362,N_2125,N_2245);
nor U2363 (N_2363,N_2138,N_2196);
nor U2364 (N_2364,N_2150,N_2134);
or U2365 (N_2365,N_2223,N_2165);
nor U2366 (N_2366,N_2196,N_2167);
or U2367 (N_2367,N_2141,N_2154);
nand U2368 (N_2368,N_2130,N_2199);
xnor U2369 (N_2369,N_2240,N_2146);
or U2370 (N_2370,N_2155,N_2163);
and U2371 (N_2371,N_2203,N_2161);
nor U2372 (N_2372,N_2184,N_2146);
or U2373 (N_2373,N_2191,N_2214);
nand U2374 (N_2374,N_2164,N_2241);
and U2375 (N_2375,N_2334,N_2303);
or U2376 (N_2376,N_2317,N_2263);
and U2377 (N_2377,N_2286,N_2278);
xnor U2378 (N_2378,N_2321,N_2257);
or U2379 (N_2379,N_2366,N_2345);
nand U2380 (N_2380,N_2277,N_2298);
nor U2381 (N_2381,N_2273,N_2337);
or U2382 (N_2382,N_2361,N_2287);
nor U2383 (N_2383,N_2368,N_2349);
and U2384 (N_2384,N_2346,N_2312);
and U2385 (N_2385,N_2323,N_2355);
nor U2386 (N_2386,N_2367,N_2300);
nand U2387 (N_2387,N_2324,N_2270);
nand U2388 (N_2388,N_2284,N_2262);
and U2389 (N_2389,N_2302,N_2306);
nor U2390 (N_2390,N_2338,N_2353);
nor U2391 (N_2391,N_2370,N_2255);
and U2392 (N_2392,N_2319,N_2327);
nor U2393 (N_2393,N_2374,N_2314);
and U2394 (N_2394,N_2343,N_2329);
or U2395 (N_2395,N_2351,N_2264);
xnor U2396 (N_2396,N_2362,N_2364);
or U2397 (N_2397,N_2259,N_2254);
nor U2398 (N_2398,N_2354,N_2363);
nand U2399 (N_2399,N_2357,N_2251);
or U2400 (N_2400,N_2299,N_2325);
nor U2401 (N_2401,N_2289,N_2365);
or U2402 (N_2402,N_2292,N_2272);
nor U2403 (N_2403,N_2297,N_2274);
and U2404 (N_2404,N_2256,N_2332);
and U2405 (N_2405,N_2252,N_2341);
nand U2406 (N_2406,N_2347,N_2280);
nor U2407 (N_2407,N_2307,N_2369);
or U2408 (N_2408,N_2328,N_2311);
xor U2409 (N_2409,N_2275,N_2265);
xnor U2410 (N_2410,N_2283,N_2339);
and U2411 (N_2411,N_2293,N_2282);
nand U2412 (N_2412,N_2269,N_2371);
nor U2413 (N_2413,N_2288,N_2291);
nand U2414 (N_2414,N_2342,N_2261);
nor U2415 (N_2415,N_2304,N_2320);
nand U2416 (N_2416,N_2352,N_2335);
nor U2417 (N_2417,N_2268,N_2336);
and U2418 (N_2418,N_2344,N_2310);
or U2419 (N_2419,N_2326,N_2308);
and U2420 (N_2420,N_2276,N_2260);
and U2421 (N_2421,N_2356,N_2316);
nand U2422 (N_2422,N_2331,N_2350);
nor U2423 (N_2423,N_2322,N_2294);
nor U2424 (N_2424,N_2281,N_2313);
or U2425 (N_2425,N_2305,N_2360);
nor U2426 (N_2426,N_2340,N_2330);
and U2427 (N_2427,N_2318,N_2253);
nand U2428 (N_2428,N_2290,N_2359);
or U2429 (N_2429,N_2372,N_2358);
nor U2430 (N_2430,N_2296,N_2295);
and U2431 (N_2431,N_2267,N_2315);
and U2432 (N_2432,N_2285,N_2301);
and U2433 (N_2433,N_2266,N_2333);
or U2434 (N_2434,N_2250,N_2258);
and U2435 (N_2435,N_2309,N_2373);
and U2436 (N_2436,N_2348,N_2279);
nor U2437 (N_2437,N_2271,N_2316);
nor U2438 (N_2438,N_2285,N_2357);
or U2439 (N_2439,N_2317,N_2259);
or U2440 (N_2440,N_2302,N_2301);
or U2441 (N_2441,N_2250,N_2291);
and U2442 (N_2442,N_2319,N_2370);
nor U2443 (N_2443,N_2355,N_2370);
nor U2444 (N_2444,N_2283,N_2349);
nand U2445 (N_2445,N_2284,N_2296);
nor U2446 (N_2446,N_2325,N_2366);
nand U2447 (N_2447,N_2311,N_2359);
and U2448 (N_2448,N_2257,N_2282);
nand U2449 (N_2449,N_2337,N_2312);
or U2450 (N_2450,N_2315,N_2349);
or U2451 (N_2451,N_2345,N_2298);
and U2452 (N_2452,N_2332,N_2372);
and U2453 (N_2453,N_2365,N_2350);
or U2454 (N_2454,N_2345,N_2291);
nor U2455 (N_2455,N_2372,N_2299);
nor U2456 (N_2456,N_2346,N_2356);
and U2457 (N_2457,N_2358,N_2272);
nand U2458 (N_2458,N_2297,N_2316);
and U2459 (N_2459,N_2328,N_2349);
and U2460 (N_2460,N_2342,N_2289);
nand U2461 (N_2461,N_2291,N_2303);
or U2462 (N_2462,N_2323,N_2276);
nor U2463 (N_2463,N_2256,N_2324);
and U2464 (N_2464,N_2341,N_2250);
nor U2465 (N_2465,N_2261,N_2263);
or U2466 (N_2466,N_2354,N_2348);
nand U2467 (N_2467,N_2260,N_2259);
nand U2468 (N_2468,N_2347,N_2363);
nand U2469 (N_2469,N_2316,N_2285);
nor U2470 (N_2470,N_2290,N_2250);
or U2471 (N_2471,N_2255,N_2299);
nor U2472 (N_2472,N_2262,N_2362);
or U2473 (N_2473,N_2368,N_2319);
xor U2474 (N_2474,N_2369,N_2279);
and U2475 (N_2475,N_2250,N_2322);
or U2476 (N_2476,N_2369,N_2341);
nor U2477 (N_2477,N_2370,N_2361);
and U2478 (N_2478,N_2364,N_2371);
or U2479 (N_2479,N_2319,N_2270);
xnor U2480 (N_2480,N_2335,N_2299);
nor U2481 (N_2481,N_2347,N_2292);
and U2482 (N_2482,N_2250,N_2277);
and U2483 (N_2483,N_2266,N_2302);
or U2484 (N_2484,N_2260,N_2292);
and U2485 (N_2485,N_2281,N_2312);
and U2486 (N_2486,N_2272,N_2312);
nand U2487 (N_2487,N_2273,N_2268);
and U2488 (N_2488,N_2370,N_2352);
xor U2489 (N_2489,N_2287,N_2351);
and U2490 (N_2490,N_2297,N_2284);
and U2491 (N_2491,N_2341,N_2256);
or U2492 (N_2492,N_2261,N_2317);
nor U2493 (N_2493,N_2304,N_2291);
or U2494 (N_2494,N_2320,N_2271);
nand U2495 (N_2495,N_2314,N_2372);
or U2496 (N_2496,N_2282,N_2367);
and U2497 (N_2497,N_2323,N_2339);
or U2498 (N_2498,N_2338,N_2307);
or U2499 (N_2499,N_2319,N_2357);
or U2500 (N_2500,N_2413,N_2434);
or U2501 (N_2501,N_2378,N_2443);
or U2502 (N_2502,N_2410,N_2420);
nand U2503 (N_2503,N_2498,N_2439);
nand U2504 (N_2504,N_2464,N_2472);
or U2505 (N_2505,N_2415,N_2444);
or U2506 (N_2506,N_2389,N_2426);
or U2507 (N_2507,N_2463,N_2465);
nor U2508 (N_2508,N_2491,N_2496);
xor U2509 (N_2509,N_2447,N_2401);
nand U2510 (N_2510,N_2397,N_2459);
and U2511 (N_2511,N_2417,N_2375);
or U2512 (N_2512,N_2475,N_2411);
or U2513 (N_2513,N_2428,N_2381);
xnor U2514 (N_2514,N_2469,N_2432);
and U2515 (N_2515,N_2430,N_2458);
nand U2516 (N_2516,N_2400,N_2488);
nor U2517 (N_2517,N_2487,N_2454);
and U2518 (N_2518,N_2408,N_2385);
nor U2519 (N_2519,N_2479,N_2451);
xnor U2520 (N_2520,N_2497,N_2421);
nand U2521 (N_2521,N_2448,N_2404);
and U2522 (N_2522,N_2399,N_2483);
nand U2523 (N_2523,N_2419,N_2480);
or U2524 (N_2524,N_2412,N_2435);
or U2525 (N_2525,N_2394,N_2481);
nor U2526 (N_2526,N_2393,N_2431);
nand U2527 (N_2527,N_2468,N_2455);
nand U2528 (N_2528,N_2422,N_2494);
xor U2529 (N_2529,N_2405,N_2407);
xnor U2530 (N_2530,N_2427,N_2438);
nor U2531 (N_2531,N_2392,N_2380);
nor U2532 (N_2532,N_2442,N_2376);
or U2533 (N_2533,N_2484,N_2388);
and U2534 (N_2534,N_2489,N_2470);
and U2535 (N_2535,N_2476,N_2424);
or U2536 (N_2536,N_2482,N_2377);
nor U2537 (N_2537,N_2477,N_2403);
or U2538 (N_2538,N_2423,N_2402);
or U2539 (N_2539,N_2466,N_2457);
or U2540 (N_2540,N_2391,N_2437);
nor U2541 (N_2541,N_2445,N_2406);
and U2542 (N_2542,N_2471,N_2433);
nand U2543 (N_2543,N_2386,N_2474);
nor U2544 (N_2544,N_2499,N_2452);
or U2545 (N_2545,N_2478,N_2449);
and U2546 (N_2546,N_2436,N_2450);
and U2547 (N_2547,N_2429,N_2461);
and U2548 (N_2548,N_2383,N_2418);
nand U2549 (N_2549,N_2495,N_2460);
or U2550 (N_2550,N_2486,N_2490);
and U2551 (N_2551,N_2382,N_2440);
xnor U2552 (N_2552,N_2395,N_2416);
nor U2553 (N_2553,N_2485,N_2398);
xnor U2554 (N_2554,N_2493,N_2456);
xor U2555 (N_2555,N_2425,N_2473);
and U2556 (N_2556,N_2462,N_2379);
or U2557 (N_2557,N_2414,N_2390);
xnor U2558 (N_2558,N_2387,N_2467);
nand U2559 (N_2559,N_2441,N_2453);
or U2560 (N_2560,N_2492,N_2409);
or U2561 (N_2561,N_2396,N_2446);
and U2562 (N_2562,N_2384,N_2420);
and U2563 (N_2563,N_2434,N_2384);
or U2564 (N_2564,N_2379,N_2405);
nor U2565 (N_2565,N_2380,N_2402);
or U2566 (N_2566,N_2458,N_2419);
xor U2567 (N_2567,N_2478,N_2411);
or U2568 (N_2568,N_2459,N_2375);
or U2569 (N_2569,N_2384,N_2455);
nand U2570 (N_2570,N_2469,N_2423);
or U2571 (N_2571,N_2412,N_2447);
nand U2572 (N_2572,N_2472,N_2389);
or U2573 (N_2573,N_2427,N_2464);
and U2574 (N_2574,N_2467,N_2444);
xnor U2575 (N_2575,N_2424,N_2430);
or U2576 (N_2576,N_2398,N_2498);
and U2577 (N_2577,N_2493,N_2492);
nor U2578 (N_2578,N_2498,N_2472);
and U2579 (N_2579,N_2488,N_2485);
nand U2580 (N_2580,N_2433,N_2459);
nand U2581 (N_2581,N_2471,N_2458);
nor U2582 (N_2582,N_2481,N_2446);
and U2583 (N_2583,N_2423,N_2396);
nand U2584 (N_2584,N_2484,N_2432);
nor U2585 (N_2585,N_2463,N_2436);
xor U2586 (N_2586,N_2393,N_2473);
or U2587 (N_2587,N_2497,N_2447);
or U2588 (N_2588,N_2464,N_2477);
nand U2589 (N_2589,N_2432,N_2471);
or U2590 (N_2590,N_2458,N_2482);
and U2591 (N_2591,N_2432,N_2377);
nand U2592 (N_2592,N_2487,N_2423);
xor U2593 (N_2593,N_2417,N_2402);
nor U2594 (N_2594,N_2455,N_2382);
and U2595 (N_2595,N_2452,N_2399);
nor U2596 (N_2596,N_2407,N_2487);
nand U2597 (N_2597,N_2468,N_2463);
xor U2598 (N_2598,N_2463,N_2487);
and U2599 (N_2599,N_2415,N_2439);
and U2600 (N_2600,N_2490,N_2424);
nor U2601 (N_2601,N_2475,N_2468);
nand U2602 (N_2602,N_2483,N_2438);
xor U2603 (N_2603,N_2396,N_2483);
xnor U2604 (N_2604,N_2475,N_2456);
and U2605 (N_2605,N_2464,N_2405);
nor U2606 (N_2606,N_2499,N_2487);
nor U2607 (N_2607,N_2486,N_2376);
or U2608 (N_2608,N_2498,N_2496);
nand U2609 (N_2609,N_2416,N_2424);
nor U2610 (N_2610,N_2409,N_2486);
xor U2611 (N_2611,N_2376,N_2408);
xor U2612 (N_2612,N_2498,N_2433);
or U2613 (N_2613,N_2400,N_2468);
and U2614 (N_2614,N_2483,N_2493);
nand U2615 (N_2615,N_2476,N_2485);
or U2616 (N_2616,N_2411,N_2492);
nand U2617 (N_2617,N_2456,N_2482);
or U2618 (N_2618,N_2428,N_2492);
nand U2619 (N_2619,N_2412,N_2414);
nor U2620 (N_2620,N_2386,N_2411);
xor U2621 (N_2621,N_2404,N_2437);
or U2622 (N_2622,N_2388,N_2434);
or U2623 (N_2623,N_2416,N_2420);
nor U2624 (N_2624,N_2485,N_2423);
nor U2625 (N_2625,N_2541,N_2543);
or U2626 (N_2626,N_2616,N_2528);
or U2627 (N_2627,N_2596,N_2614);
nand U2628 (N_2628,N_2604,N_2571);
nand U2629 (N_2629,N_2519,N_2609);
or U2630 (N_2630,N_2589,N_2577);
or U2631 (N_2631,N_2581,N_2569);
and U2632 (N_2632,N_2606,N_2503);
nand U2633 (N_2633,N_2527,N_2561);
nor U2634 (N_2634,N_2542,N_2580);
nand U2635 (N_2635,N_2521,N_2514);
and U2636 (N_2636,N_2555,N_2592);
and U2637 (N_2637,N_2545,N_2520);
and U2638 (N_2638,N_2535,N_2564);
and U2639 (N_2639,N_2598,N_2557);
xnor U2640 (N_2640,N_2530,N_2526);
and U2641 (N_2641,N_2517,N_2550);
nor U2642 (N_2642,N_2576,N_2536);
xnor U2643 (N_2643,N_2591,N_2575);
or U2644 (N_2644,N_2534,N_2508);
or U2645 (N_2645,N_2599,N_2607);
and U2646 (N_2646,N_2584,N_2579);
nor U2647 (N_2647,N_2502,N_2523);
and U2648 (N_2648,N_2568,N_2620);
nand U2649 (N_2649,N_2509,N_2556);
nor U2650 (N_2650,N_2613,N_2501);
or U2651 (N_2651,N_2621,N_2537);
nand U2652 (N_2652,N_2539,N_2611);
nor U2653 (N_2653,N_2574,N_2583);
and U2654 (N_2654,N_2552,N_2553);
nor U2655 (N_2655,N_2540,N_2524);
nor U2656 (N_2656,N_2525,N_2565);
nor U2657 (N_2657,N_2572,N_2544);
and U2658 (N_2658,N_2608,N_2563);
nand U2659 (N_2659,N_2531,N_2617);
or U2660 (N_2660,N_2624,N_2512);
or U2661 (N_2661,N_2618,N_2622);
nor U2662 (N_2662,N_2619,N_2510);
nand U2663 (N_2663,N_2547,N_2600);
xnor U2664 (N_2664,N_2546,N_2533);
or U2665 (N_2665,N_2594,N_2610);
nor U2666 (N_2666,N_2603,N_2570);
nand U2667 (N_2667,N_2507,N_2567);
and U2668 (N_2668,N_2562,N_2585);
or U2669 (N_2669,N_2590,N_2518);
and U2670 (N_2670,N_2548,N_2506);
nor U2671 (N_2671,N_2602,N_2612);
or U2672 (N_2672,N_2558,N_2586);
nor U2673 (N_2673,N_2623,N_2559);
or U2674 (N_2674,N_2511,N_2601);
nand U2675 (N_2675,N_2578,N_2532);
nor U2676 (N_2676,N_2560,N_2582);
nor U2677 (N_2677,N_2504,N_2529);
and U2678 (N_2678,N_2593,N_2551);
nand U2679 (N_2679,N_2538,N_2573);
and U2680 (N_2680,N_2566,N_2515);
nand U2681 (N_2681,N_2505,N_2605);
nor U2682 (N_2682,N_2597,N_2587);
and U2683 (N_2683,N_2615,N_2516);
xnor U2684 (N_2684,N_2500,N_2595);
or U2685 (N_2685,N_2522,N_2549);
xor U2686 (N_2686,N_2554,N_2513);
nand U2687 (N_2687,N_2588,N_2600);
xnor U2688 (N_2688,N_2597,N_2555);
nor U2689 (N_2689,N_2573,N_2519);
or U2690 (N_2690,N_2606,N_2589);
xor U2691 (N_2691,N_2523,N_2530);
or U2692 (N_2692,N_2610,N_2506);
nor U2693 (N_2693,N_2612,N_2524);
nand U2694 (N_2694,N_2526,N_2540);
nor U2695 (N_2695,N_2536,N_2558);
nor U2696 (N_2696,N_2576,N_2505);
and U2697 (N_2697,N_2609,N_2582);
nand U2698 (N_2698,N_2538,N_2525);
or U2699 (N_2699,N_2613,N_2542);
or U2700 (N_2700,N_2589,N_2603);
or U2701 (N_2701,N_2621,N_2505);
nand U2702 (N_2702,N_2616,N_2606);
and U2703 (N_2703,N_2608,N_2567);
or U2704 (N_2704,N_2530,N_2606);
and U2705 (N_2705,N_2559,N_2531);
nor U2706 (N_2706,N_2611,N_2527);
nand U2707 (N_2707,N_2536,N_2545);
nand U2708 (N_2708,N_2523,N_2547);
nand U2709 (N_2709,N_2530,N_2543);
nor U2710 (N_2710,N_2517,N_2597);
nand U2711 (N_2711,N_2601,N_2619);
and U2712 (N_2712,N_2520,N_2517);
and U2713 (N_2713,N_2584,N_2514);
nor U2714 (N_2714,N_2553,N_2609);
and U2715 (N_2715,N_2608,N_2620);
nand U2716 (N_2716,N_2604,N_2503);
or U2717 (N_2717,N_2604,N_2615);
nand U2718 (N_2718,N_2618,N_2613);
nor U2719 (N_2719,N_2522,N_2619);
nor U2720 (N_2720,N_2543,N_2595);
and U2721 (N_2721,N_2549,N_2592);
and U2722 (N_2722,N_2563,N_2622);
nand U2723 (N_2723,N_2599,N_2617);
nor U2724 (N_2724,N_2578,N_2507);
nand U2725 (N_2725,N_2600,N_2572);
or U2726 (N_2726,N_2597,N_2538);
and U2727 (N_2727,N_2525,N_2540);
nor U2728 (N_2728,N_2554,N_2601);
and U2729 (N_2729,N_2547,N_2603);
and U2730 (N_2730,N_2539,N_2610);
and U2731 (N_2731,N_2539,N_2592);
xnor U2732 (N_2732,N_2530,N_2553);
nor U2733 (N_2733,N_2606,N_2521);
or U2734 (N_2734,N_2539,N_2588);
or U2735 (N_2735,N_2576,N_2535);
or U2736 (N_2736,N_2552,N_2579);
and U2737 (N_2737,N_2511,N_2569);
nor U2738 (N_2738,N_2543,N_2583);
nor U2739 (N_2739,N_2530,N_2622);
nand U2740 (N_2740,N_2587,N_2534);
or U2741 (N_2741,N_2524,N_2582);
or U2742 (N_2742,N_2560,N_2566);
and U2743 (N_2743,N_2540,N_2507);
nand U2744 (N_2744,N_2565,N_2530);
nand U2745 (N_2745,N_2581,N_2598);
or U2746 (N_2746,N_2598,N_2616);
and U2747 (N_2747,N_2587,N_2618);
nor U2748 (N_2748,N_2548,N_2534);
nor U2749 (N_2749,N_2560,N_2523);
nor U2750 (N_2750,N_2707,N_2692);
nand U2751 (N_2751,N_2645,N_2651);
nand U2752 (N_2752,N_2650,N_2742);
or U2753 (N_2753,N_2681,N_2697);
nand U2754 (N_2754,N_2685,N_2660);
nor U2755 (N_2755,N_2733,N_2731);
nand U2756 (N_2756,N_2643,N_2698);
xnor U2757 (N_2757,N_2673,N_2631);
and U2758 (N_2758,N_2687,N_2748);
nor U2759 (N_2759,N_2696,N_2663);
or U2760 (N_2760,N_2722,N_2633);
and U2761 (N_2761,N_2716,N_2745);
and U2762 (N_2762,N_2732,N_2720);
or U2763 (N_2763,N_2737,N_2672);
and U2764 (N_2764,N_2647,N_2657);
nand U2765 (N_2765,N_2709,N_2702);
nand U2766 (N_2766,N_2678,N_2646);
nand U2767 (N_2767,N_2718,N_2634);
nand U2768 (N_2768,N_2717,N_2669);
and U2769 (N_2769,N_2724,N_2635);
nor U2770 (N_2770,N_2629,N_2701);
nor U2771 (N_2771,N_2668,N_2726);
and U2772 (N_2772,N_2695,N_2677);
nand U2773 (N_2773,N_2747,N_2704);
and U2774 (N_2774,N_2712,N_2705);
or U2775 (N_2775,N_2727,N_2725);
or U2776 (N_2776,N_2632,N_2734);
nor U2777 (N_2777,N_2699,N_2665);
and U2778 (N_2778,N_2684,N_2653);
nor U2779 (N_2779,N_2743,N_2627);
and U2780 (N_2780,N_2739,N_2679);
nor U2781 (N_2781,N_2723,N_2670);
nor U2782 (N_2782,N_2648,N_2659);
nand U2783 (N_2783,N_2680,N_2736);
nand U2784 (N_2784,N_2719,N_2714);
nor U2785 (N_2785,N_2700,N_2664);
and U2786 (N_2786,N_2649,N_2706);
or U2787 (N_2787,N_2729,N_2626);
xor U2788 (N_2788,N_2638,N_2658);
nand U2789 (N_2789,N_2671,N_2667);
and U2790 (N_2790,N_2628,N_2654);
nand U2791 (N_2791,N_2730,N_2708);
nand U2792 (N_2792,N_2642,N_2625);
nand U2793 (N_2793,N_2728,N_2694);
or U2794 (N_2794,N_2746,N_2666);
nor U2795 (N_2795,N_2688,N_2655);
or U2796 (N_2796,N_2644,N_2662);
and U2797 (N_2797,N_2711,N_2721);
nor U2798 (N_2798,N_2744,N_2630);
xnor U2799 (N_2799,N_2675,N_2710);
and U2800 (N_2800,N_2661,N_2652);
or U2801 (N_2801,N_2641,N_2676);
nand U2802 (N_2802,N_2693,N_2636);
nor U2803 (N_2803,N_2689,N_2639);
xor U2804 (N_2804,N_2637,N_2740);
and U2805 (N_2805,N_2703,N_2741);
nor U2806 (N_2806,N_2715,N_2713);
or U2807 (N_2807,N_2749,N_2686);
and U2808 (N_2808,N_2640,N_2735);
nor U2809 (N_2809,N_2690,N_2656);
xor U2810 (N_2810,N_2682,N_2674);
and U2811 (N_2811,N_2691,N_2683);
nand U2812 (N_2812,N_2738,N_2711);
xor U2813 (N_2813,N_2669,N_2626);
nand U2814 (N_2814,N_2676,N_2717);
and U2815 (N_2815,N_2659,N_2727);
nor U2816 (N_2816,N_2664,N_2715);
xor U2817 (N_2817,N_2658,N_2705);
nand U2818 (N_2818,N_2641,N_2741);
or U2819 (N_2819,N_2628,N_2704);
nor U2820 (N_2820,N_2734,N_2685);
nor U2821 (N_2821,N_2625,N_2700);
nor U2822 (N_2822,N_2715,N_2655);
and U2823 (N_2823,N_2709,N_2634);
nand U2824 (N_2824,N_2686,N_2728);
nor U2825 (N_2825,N_2663,N_2639);
xnor U2826 (N_2826,N_2704,N_2748);
and U2827 (N_2827,N_2691,N_2716);
xnor U2828 (N_2828,N_2741,N_2640);
and U2829 (N_2829,N_2736,N_2626);
and U2830 (N_2830,N_2633,N_2732);
nor U2831 (N_2831,N_2736,N_2731);
nor U2832 (N_2832,N_2638,N_2749);
and U2833 (N_2833,N_2726,N_2681);
nor U2834 (N_2834,N_2743,N_2737);
nand U2835 (N_2835,N_2672,N_2683);
nand U2836 (N_2836,N_2685,N_2648);
nand U2837 (N_2837,N_2745,N_2695);
nand U2838 (N_2838,N_2720,N_2660);
nor U2839 (N_2839,N_2730,N_2670);
and U2840 (N_2840,N_2721,N_2637);
nand U2841 (N_2841,N_2641,N_2734);
or U2842 (N_2842,N_2696,N_2707);
and U2843 (N_2843,N_2708,N_2725);
nor U2844 (N_2844,N_2720,N_2671);
or U2845 (N_2845,N_2689,N_2695);
nor U2846 (N_2846,N_2652,N_2668);
and U2847 (N_2847,N_2713,N_2692);
or U2848 (N_2848,N_2718,N_2657);
or U2849 (N_2849,N_2734,N_2647);
or U2850 (N_2850,N_2724,N_2674);
or U2851 (N_2851,N_2668,N_2712);
or U2852 (N_2852,N_2630,N_2726);
or U2853 (N_2853,N_2729,N_2651);
or U2854 (N_2854,N_2672,N_2736);
or U2855 (N_2855,N_2639,N_2636);
and U2856 (N_2856,N_2714,N_2638);
and U2857 (N_2857,N_2735,N_2676);
or U2858 (N_2858,N_2724,N_2659);
and U2859 (N_2859,N_2665,N_2653);
nor U2860 (N_2860,N_2730,N_2658);
nand U2861 (N_2861,N_2731,N_2656);
and U2862 (N_2862,N_2712,N_2729);
nand U2863 (N_2863,N_2630,N_2682);
and U2864 (N_2864,N_2655,N_2700);
and U2865 (N_2865,N_2650,N_2709);
xnor U2866 (N_2866,N_2674,N_2657);
or U2867 (N_2867,N_2632,N_2707);
or U2868 (N_2868,N_2659,N_2707);
nor U2869 (N_2869,N_2705,N_2704);
nor U2870 (N_2870,N_2635,N_2680);
nor U2871 (N_2871,N_2672,N_2639);
or U2872 (N_2872,N_2743,N_2651);
nand U2873 (N_2873,N_2651,N_2701);
nand U2874 (N_2874,N_2748,N_2669);
nor U2875 (N_2875,N_2767,N_2856);
and U2876 (N_2876,N_2851,N_2796);
and U2877 (N_2877,N_2853,N_2834);
or U2878 (N_2878,N_2775,N_2792);
or U2879 (N_2879,N_2799,N_2759);
or U2880 (N_2880,N_2824,N_2863);
or U2881 (N_2881,N_2750,N_2755);
or U2882 (N_2882,N_2860,N_2810);
or U2883 (N_2883,N_2812,N_2869);
xor U2884 (N_2884,N_2785,N_2854);
nor U2885 (N_2885,N_2770,N_2873);
nor U2886 (N_2886,N_2776,N_2818);
nor U2887 (N_2887,N_2866,N_2845);
nor U2888 (N_2888,N_2781,N_2783);
or U2889 (N_2889,N_2819,N_2805);
xnor U2890 (N_2890,N_2872,N_2757);
nor U2891 (N_2891,N_2849,N_2797);
nor U2892 (N_2892,N_2752,N_2779);
nor U2893 (N_2893,N_2800,N_2861);
nor U2894 (N_2894,N_2764,N_2827);
nor U2895 (N_2895,N_2836,N_2794);
nand U2896 (N_2896,N_2830,N_2820);
nand U2897 (N_2897,N_2772,N_2857);
xor U2898 (N_2898,N_2791,N_2753);
nor U2899 (N_2899,N_2841,N_2874);
or U2900 (N_2900,N_2754,N_2840);
nor U2901 (N_2901,N_2829,N_2807);
nand U2902 (N_2902,N_2825,N_2838);
nor U2903 (N_2903,N_2815,N_2864);
or U2904 (N_2904,N_2788,N_2774);
xor U2905 (N_2905,N_2847,N_2773);
and U2906 (N_2906,N_2833,N_2814);
nand U2907 (N_2907,N_2813,N_2855);
and U2908 (N_2908,N_2811,N_2858);
or U2909 (N_2909,N_2844,N_2843);
or U2910 (N_2910,N_2790,N_2846);
nand U2911 (N_2911,N_2804,N_2839);
nand U2912 (N_2912,N_2762,N_2865);
xor U2913 (N_2913,N_2828,N_2761);
nor U2914 (N_2914,N_2789,N_2766);
nor U2915 (N_2915,N_2803,N_2817);
and U2916 (N_2916,N_2848,N_2859);
nand U2917 (N_2917,N_2867,N_2802);
and U2918 (N_2918,N_2786,N_2801);
or U2919 (N_2919,N_2798,N_2768);
and U2920 (N_2920,N_2868,N_2832);
nand U2921 (N_2921,N_2835,N_2816);
nor U2922 (N_2922,N_2826,N_2871);
and U2923 (N_2923,N_2760,N_2793);
or U2924 (N_2924,N_2806,N_2809);
nand U2925 (N_2925,N_2850,N_2780);
nand U2926 (N_2926,N_2771,N_2795);
nand U2927 (N_2927,N_2778,N_2756);
nor U2928 (N_2928,N_2782,N_2822);
or U2929 (N_2929,N_2870,N_2763);
or U2930 (N_2930,N_2769,N_2784);
xnor U2931 (N_2931,N_2777,N_2837);
xor U2932 (N_2932,N_2821,N_2765);
or U2933 (N_2933,N_2852,N_2831);
nor U2934 (N_2934,N_2758,N_2751);
nor U2935 (N_2935,N_2862,N_2787);
nand U2936 (N_2936,N_2808,N_2823);
or U2937 (N_2937,N_2842,N_2824);
xor U2938 (N_2938,N_2765,N_2808);
nand U2939 (N_2939,N_2795,N_2762);
or U2940 (N_2940,N_2835,N_2870);
and U2941 (N_2941,N_2837,N_2854);
or U2942 (N_2942,N_2752,N_2804);
nor U2943 (N_2943,N_2799,N_2833);
and U2944 (N_2944,N_2799,N_2774);
or U2945 (N_2945,N_2810,N_2849);
nand U2946 (N_2946,N_2776,N_2842);
nand U2947 (N_2947,N_2799,N_2750);
nand U2948 (N_2948,N_2849,N_2786);
nor U2949 (N_2949,N_2874,N_2795);
nor U2950 (N_2950,N_2753,N_2763);
xnor U2951 (N_2951,N_2814,N_2783);
and U2952 (N_2952,N_2822,N_2812);
nand U2953 (N_2953,N_2760,N_2771);
and U2954 (N_2954,N_2784,N_2822);
and U2955 (N_2955,N_2784,N_2763);
or U2956 (N_2956,N_2788,N_2766);
nand U2957 (N_2957,N_2814,N_2855);
nand U2958 (N_2958,N_2801,N_2828);
xnor U2959 (N_2959,N_2825,N_2863);
nand U2960 (N_2960,N_2856,N_2802);
nor U2961 (N_2961,N_2788,N_2758);
xor U2962 (N_2962,N_2750,N_2776);
and U2963 (N_2963,N_2763,N_2823);
or U2964 (N_2964,N_2854,N_2797);
nor U2965 (N_2965,N_2871,N_2860);
nor U2966 (N_2966,N_2803,N_2829);
xnor U2967 (N_2967,N_2766,N_2767);
xor U2968 (N_2968,N_2842,N_2834);
or U2969 (N_2969,N_2831,N_2780);
nor U2970 (N_2970,N_2874,N_2846);
nand U2971 (N_2971,N_2860,N_2824);
nor U2972 (N_2972,N_2777,N_2819);
or U2973 (N_2973,N_2773,N_2837);
or U2974 (N_2974,N_2826,N_2768);
nand U2975 (N_2975,N_2758,N_2844);
or U2976 (N_2976,N_2750,N_2812);
xnor U2977 (N_2977,N_2776,N_2855);
nand U2978 (N_2978,N_2787,N_2815);
xor U2979 (N_2979,N_2870,N_2797);
xor U2980 (N_2980,N_2867,N_2785);
nor U2981 (N_2981,N_2781,N_2762);
nand U2982 (N_2982,N_2759,N_2822);
nor U2983 (N_2983,N_2835,N_2796);
nor U2984 (N_2984,N_2810,N_2863);
nor U2985 (N_2985,N_2853,N_2752);
xnor U2986 (N_2986,N_2829,N_2813);
nor U2987 (N_2987,N_2806,N_2857);
nor U2988 (N_2988,N_2857,N_2767);
or U2989 (N_2989,N_2794,N_2859);
and U2990 (N_2990,N_2798,N_2752);
nand U2991 (N_2991,N_2764,N_2809);
xor U2992 (N_2992,N_2837,N_2863);
or U2993 (N_2993,N_2761,N_2814);
xor U2994 (N_2994,N_2850,N_2846);
nor U2995 (N_2995,N_2758,N_2760);
and U2996 (N_2996,N_2854,N_2841);
nor U2997 (N_2997,N_2784,N_2829);
nor U2998 (N_2998,N_2804,N_2769);
or U2999 (N_2999,N_2855,N_2846);
xor U3000 (N_3000,N_2986,N_2886);
or U3001 (N_3001,N_2927,N_2956);
xnor U3002 (N_3002,N_2938,N_2881);
xnor U3003 (N_3003,N_2924,N_2934);
and U3004 (N_3004,N_2884,N_2912);
nand U3005 (N_3005,N_2932,N_2999);
nand U3006 (N_3006,N_2939,N_2909);
or U3007 (N_3007,N_2906,N_2971);
xor U3008 (N_3008,N_2914,N_2937);
or U3009 (N_3009,N_2976,N_2969);
and U3010 (N_3010,N_2942,N_2964);
xnor U3011 (N_3011,N_2929,N_2952);
or U3012 (N_3012,N_2989,N_2984);
nand U3013 (N_3013,N_2977,N_2879);
or U3014 (N_3014,N_2962,N_2907);
and U3015 (N_3015,N_2970,N_2959);
nand U3016 (N_3016,N_2890,N_2949);
or U3017 (N_3017,N_2901,N_2936);
or U3018 (N_3018,N_2988,N_2995);
nand U3019 (N_3019,N_2987,N_2991);
nor U3020 (N_3020,N_2961,N_2922);
nand U3021 (N_3021,N_2983,N_2877);
or U3022 (N_3022,N_2887,N_2875);
or U3023 (N_3023,N_2946,N_2994);
xor U3024 (N_3024,N_2968,N_2894);
nor U3025 (N_3025,N_2985,N_2917);
nor U3026 (N_3026,N_2950,N_2925);
or U3027 (N_3027,N_2908,N_2990);
nand U3028 (N_3028,N_2960,N_2931);
nand U3029 (N_3029,N_2958,N_2973);
and U3030 (N_3030,N_2933,N_2923);
or U3031 (N_3031,N_2876,N_2882);
and U3032 (N_3032,N_2996,N_2944);
nand U3033 (N_3033,N_2885,N_2911);
nand U3034 (N_3034,N_2903,N_2930);
and U3035 (N_3035,N_2972,N_2948);
or U3036 (N_3036,N_2979,N_2998);
or U3037 (N_3037,N_2880,N_2992);
and U3038 (N_3038,N_2997,N_2919);
and U3039 (N_3039,N_2967,N_2926);
nand U3040 (N_3040,N_2918,N_2974);
or U3041 (N_3041,N_2899,N_2896);
nand U3042 (N_3042,N_2883,N_2955);
and U3043 (N_3043,N_2900,N_2915);
nand U3044 (N_3044,N_2913,N_2963);
nand U3045 (N_3045,N_2910,N_2965);
nand U3046 (N_3046,N_2981,N_2905);
nand U3047 (N_3047,N_2980,N_2954);
xnor U3048 (N_3048,N_2975,N_2928);
nand U3049 (N_3049,N_2904,N_2902);
and U3050 (N_3050,N_2947,N_2878);
nor U3051 (N_3051,N_2966,N_2993);
or U3052 (N_3052,N_2897,N_2893);
nand U3053 (N_3053,N_2953,N_2935);
or U3054 (N_3054,N_2921,N_2888);
nand U3055 (N_3055,N_2940,N_2941);
nand U3056 (N_3056,N_2889,N_2920);
nand U3057 (N_3057,N_2951,N_2978);
or U3058 (N_3058,N_2916,N_2895);
nand U3059 (N_3059,N_2898,N_2945);
nand U3060 (N_3060,N_2957,N_2892);
and U3061 (N_3061,N_2943,N_2982);
and U3062 (N_3062,N_2891,N_2880);
xnor U3063 (N_3063,N_2986,N_2930);
nor U3064 (N_3064,N_2928,N_2938);
and U3065 (N_3065,N_2911,N_2880);
nand U3066 (N_3066,N_2979,N_2977);
or U3067 (N_3067,N_2977,N_2912);
nand U3068 (N_3068,N_2937,N_2920);
nor U3069 (N_3069,N_2918,N_2954);
nand U3070 (N_3070,N_2994,N_2877);
nand U3071 (N_3071,N_2980,N_2890);
and U3072 (N_3072,N_2999,N_2985);
nor U3073 (N_3073,N_2890,N_2990);
or U3074 (N_3074,N_2924,N_2893);
xnor U3075 (N_3075,N_2971,N_2907);
nand U3076 (N_3076,N_2985,N_2974);
or U3077 (N_3077,N_2960,N_2923);
nor U3078 (N_3078,N_2975,N_2895);
or U3079 (N_3079,N_2993,N_2918);
xnor U3080 (N_3080,N_2928,N_2914);
nand U3081 (N_3081,N_2984,N_2919);
nor U3082 (N_3082,N_2985,N_2913);
nand U3083 (N_3083,N_2966,N_2965);
or U3084 (N_3084,N_2988,N_2903);
and U3085 (N_3085,N_2889,N_2881);
nor U3086 (N_3086,N_2951,N_2896);
nor U3087 (N_3087,N_2921,N_2930);
and U3088 (N_3088,N_2942,N_2878);
nand U3089 (N_3089,N_2891,N_2968);
xnor U3090 (N_3090,N_2877,N_2895);
nor U3091 (N_3091,N_2984,N_2901);
or U3092 (N_3092,N_2943,N_2930);
and U3093 (N_3093,N_2975,N_2887);
and U3094 (N_3094,N_2965,N_2963);
or U3095 (N_3095,N_2976,N_2966);
nor U3096 (N_3096,N_2940,N_2927);
xnor U3097 (N_3097,N_2966,N_2989);
nand U3098 (N_3098,N_2908,N_2888);
and U3099 (N_3099,N_2936,N_2986);
nor U3100 (N_3100,N_2995,N_2905);
nor U3101 (N_3101,N_2905,N_2941);
xor U3102 (N_3102,N_2894,N_2875);
or U3103 (N_3103,N_2992,N_2903);
or U3104 (N_3104,N_2967,N_2951);
nand U3105 (N_3105,N_2980,N_2959);
nor U3106 (N_3106,N_2973,N_2922);
and U3107 (N_3107,N_2985,N_2953);
and U3108 (N_3108,N_2920,N_2975);
nand U3109 (N_3109,N_2942,N_2897);
xor U3110 (N_3110,N_2934,N_2986);
nand U3111 (N_3111,N_2905,N_2887);
nand U3112 (N_3112,N_2877,N_2901);
or U3113 (N_3113,N_2943,N_2878);
and U3114 (N_3114,N_2931,N_2990);
and U3115 (N_3115,N_2946,N_2876);
nor U3116 (N_3116,N_2989,N_2926);
nand U3117 (N_3117,N_2975,N_2889);
or U3118 (N_3118,N_2925,N_2935);
nor U3119 (N_3119,N_2953,N_2964);
nand U3120 (N_3120,N_2920,N_2914);
and U3121 (N_3121,N_2946,N_2956);
nand U3122 (N_3122,N_2986,N_2973);
nor U3123 (N_3123,N_2924,N_2903);
nor U3124 (N_3124,N_2985,N_2935);
and U3125 (N_3125,N_3010,N_3067);
nor U3126 (N_3126,N_3057,N_3101);
nand U3127 (N_3127,N_3091,N_3062);
nor U3128 (N_3128,N_3031,N_3109);
or U3129 (N_3129,N_3012,N_3073);
nor U3130 (N_3130,N_3029,N_3047);
nand U3131 (N_3131,N_3065,N_3061);
nor U3132 (N_3132,N_3112,N_3092);
and U3133 (N_3133,N_3028,N_3060);
or U3134 (N_3134,N_3094,N_3068);
or U3135 (N_3135,N_3113,N_3075);
or U3136 (N_3136,N_3093,N_3024);
and U3137 (N_3137,N_3063,N_3049);
xor U3138 (N_3138,N_3116,N_3046);
nor U3139 (N_3139,N_3048,N_3081);
or U3140 (N_3140,N_3018,N_3017);
nand U3141 (N_3141,N_3034,N_3005);
nor U3142 (N_3142,N_3043,N_3124);
nand U3143 (N_3143,N_3069,N_3036);
or U3144 (N_3144,N_3070,N_3102);
or U3145 (N_3145,N_3002,N_3030);
nor U3146 (N_3146,N_3099,N_3110);
nand U3147 (N_3147,N_3019,N_3114);
xor U3148 (N_3148,N_3007,N_3111);
or U3149 (N_3149,N_3071,N_3066);
nor U3150 (N_3150,N_3001,N_3121);
nor U3151 (N_3151,N_3086,N_3050);
or U3152 (N_3152,N_3023,N_3033);
nor U3153 (N_3153,N_3014,N_3096);
xor U3154 (N_3154,N_3082,N_3051);
nand U3155 (N_3155,N_3117,N_3095);
nor U3156 (N_3156,N_3097,N_3003);
nand U3157 (N_3157,N_3058,N_3119);
or U3158 (N_3158,N_3123,N_3016);
xor U3159 (N_3159,N_3000,N_3118);
or U3160 (N_3160,N_3078,N_3104);
nor U3161 (N_3161,N_3079,N_3020);
and U3162 (N_3162,N_3011,N_3006);
nor U3163 (N_3163,N_3009,N_3037);
or U3164 (N_3164,N_3100,N_3077);
and U3165 (N_3165,N_3080,N_3106);
or U3166 (N_3166,N_3022,N_3088);
or U3167 (N_3167,N_3090,N_3035);
or U3168 (N_3168,N_3013,N_3040);
or U3169 (N_3169,N_3059,N_3044);
or U3170 (N_3170,N_3052,N_3089);
and U3171 (N_3171,N_3039,N_3015);
and U3172 (N_3172,N_3072,N_3105);
or U3173 (N_3173,N_3041,N_3098);
or U3174 (N_3174,N_3103,N_3108);
or U3175 (N_3175,N_3107,N_3025);
nor U3176 (N_3176,N_3042,N_3122);
nand U3177 (N_3177,N_3115,N_3004);
nand U3178 (N_3178,N_3076,N_3055);
nor U3179 (N_3179,N_3083,N_3085);
and U3180 (N_3180,N_3008,N_3084);
nor U3181 (N_3181,N_3056,N_3027);
nand U3182 (N_3182,N_3026,N_3053);
xnor U3183 (N_3183,N_3087,N_3054);
or U3184 (N_3184,N_3064,N_3120);
and U3185 (N_3185,N_3038,N_3021);
nand U3186 (N_3186,N_3074,N_3032);
nor U3187 (N_3187,N_3045,N_3020);
nand U3188 (N_3188,N_3060,N_3029);
or U3189 (N_3189,N_3111,N_3104);
nand U3190 (N_3190,N_3115,N_3043);
and U3191 (N_3191,N_3070,N_3029);
nand U3192 (N_3192,N_3051,N_3076);
nor U3193 (N_3193,N_3065,N_3092);
nor U3194 (N_3194,N_3111,N_3084);
and U3195 (N_3195,N_3120,N_3082);
nand U3196 (N_3196,N_3102,N_3116);
and U3197 (N_3197,N_3072,N_3063);
and U3198 (N_3198,N_3064,N_3049);
nand U3199 (N_3199,N_3006,N_3002);
or U3200 (N_3200,N_3115,N_3030);
nand U3201 (N_3201,N_3062,N_3069);
nor U3202 (N_3202,N_3082,N_3008);
xnor U3203 (N_3203,N_3063,N_3031);
xnor U3204 (N_3204,N_3103,N_3005);
or U3205 (N_3205,N_3059,N_3069);
or U3206 (N_3206,N_3060,N_3001);
or U3207 (N_3207,N_3038,N_3057);
or U3208 (N_3208,N_3101,N_3049);
xnor U3209 (N_3209,N_3025,N_3032);
and U3210 (N_3210,N_3104,N_3101);
xor U3211 (N_3211,N_3084,N_3110);
or U3212 (N_3212,N_3093,N_3110);
nor U3213 (N_3213,N_3071,N_3083);
or U3214 (N_3214,N_3103,N_3089);
xor U3215 (N_3215,N_3050,N_3004);
and U3216 (N_3216,N_3046,N_3047);
and U3217 (N_3217,N_3007,N_3047);
or U3218 (N_3218,N_3039,N_3086);
nor U3219 (N_3219,N_3092,N_3051);
and U3220 (N_3220,N_3085,N_3049);
nand U3221 (N_3221,N_3082,N_3000);
or U3222 (N_3222,N_3118,N_3114);
and U3223 (N_3223,N_3060,N_3035);
nor U3224 (N_3224,N_3121,N_3026);
nor U3225 (N_3225,N_3112,N_3116);
and U3226 (N_3226,N_3048,N_3064);
nor U3227 (N_3227,N_3112,N_3106);
and U3228 (N_3228,N_3007,N_3068);
nor U3229 (N_3229,N_3120,N_3093);
nor U3230 (N_3230,N_3073,N_3090);
and U3231 (N_3231,N_3001,N_3089);
nor U3232 (N_3232,N_3069,N_3084);
or U3233 (N_3233,N_3068,N_3091);
and U3234 (N_3234,N_3039,N_3040);
nand U3235 (N_3235,N_3124,N_3060);
nand U3236 (N_3236,N_3029,N_3074);
and U3237 (N_3237,N_3122,N_3049);
nor U3238 (N_3238,N_3087,N_3104);
nor U3239 (N_3239,N_3007,N_3118);
or U3240 (N_3240,N_3068,N_3004);
and U3241 (N_3241,N_3085,N_3043);
xor U3242 (N_3242,N_3113,N_3038);
nor U3243 (N_3243,N_3007,N_3102);
and U3244 (N_3244,N_3087,N_3062);
or U3245 (N_3245,N_3075,N_3021);
nand U3246 (N_3246,N_3069,N_3116);
nand U3247 (N_3247,N_3037,N_3051);
or U3248 (N_3248,N_3068,N_3075);
or U3249 (N_3249,N_3117,N_3064);
nor U3250 (N_3250,N_3154,N_3220);
nor U3251 (N_3251,N_3135,N_3216);
nor U3252 (N_3252,N_3228,N_3198);
nor U3253 (N_3253,N_3171,N_3187);
nor U3254 (N_3254,N_3182,N_3166);
xnor U3255 (N_3255,N_3151,N_3231);
nor U3256 (N_3256,N_3239,N_3132);
nand U3257 (N_3257,N_3212,N_3234);
or U3258 (N_3258,N_3247,N_3142);
nor U3259 (N_3259,N_3176,N_3213);
xor U3260 (N_3260,N_3179,N_3223);
and U3261 (N_3261,N_3169,N_3173);
and U3262 (N_3262,N_3245,N_3221);
nand U3263 (N_3263,N_3195,N_3203);
or U3264 (N_3264,N_3177,N_3188);
or U3265 (N_3265,N_3242,N_3159);
and U3266 (N_3266,N_3134,N_3238);
nand U3267 (N_3267,N_3180,N_3143);
and U3268 (N_3268,N_3225,N_3155);
and U3269 (N_3269,N_3194,N_3127);
nor U3270 (N_3270,N_3219,N_3222);
and U3271 (N_3271,N_3189,N_3207);
nor U3272 (N_3272,N_3125,N_3199);
xor U3273 (N_3273,N_3193,N_3208);
or U3274 (N_3274,N_3235,N_3158);
nand U3275 (N_3275,N_3217,N_3160);
and U3276 (N_3276,N_3241,N_3215);
nor U3277 (N_3277,N_3186,N_3181);
nand U3278 (N_3278,N_3211,N_3196);
nand U3279 (N_3279,N_3229,N_3202);
xnor U3280 (N_3280,N_3145,N_3164);
nand U3281 (N_3281,N_3144,N_3233);
nor U3282 (N_3282,N_3167,N_3126);
and U3283 (N_3283,N_3183,N_3206);
nor U3284 (N_3284,N_3191,N_3204);
or U3285 (N_3285,N_3140,N_3246);
xor U3286 (N_3286,N_3168,N_3190);
nor U3287 (N_3287,N_3165,N_3200);
nor U3288 (N_3288,N_3201,N_3141);
nor U3289 (N_3289,N_3152,N_3192);
nor U3290 (N_3290,N_3131,N_3218);
and U3291 (N_3291,N_3197,N_3138);
nor U3292 (N_3292,N_3137,N_3249);
and U3293 (N_3293,N_3163,N_3184);
nand U3294 (N_3294,N_3148,N_3175);
or U3295 (N_3295,N_3248,N_3156);
and U3296 (N_3296,N_3226,N_3214);
and U3297 (N_3297,N_3174,N_3210);
xor U3298 (N_3298,N_3162,N_3205);
and U3299 (N_3299,N_3240,N_3236);
nand U3300 (N_3300,N_3170,N_3232);
nand U3301 (N_3301,N_3178,N_3185);
xnor U3302 (N_3302,N_3237,N_3133);
and U3303 (N_3303,N_3244,N_3230);
and U3304 (N_3304,N_3209,N_3146);
or U3305 (N_3305,N_3161,N_3172);
nand U3306 (N_3306,N_3157,N_3149);
nor U3307 (N_3307,N_3130,N_3224);
and U3308 (N_3308,N_3147,N_3150);
nor U3309 (N_3309,N_3139,N_3227);
and U3310 (N_3310,N_3128,N_3243);
or U3311 (N_3311,N_3129,N_3136);
xor U3312 (N_3312,N_3153,N_3181);
and U3313 (N_3313,N_3130,N_3135);
nand U3314 (N_3314,N_3196,N_3144);
xor U3315 (N_3315,N_3228,N_3206);
nor U3316 (N_3316,N_3210,N_3190);
nand U3317 (N_3317,N_3137,N_3203);
nand U3318 (N_3318,N_3221,N_3164);
nand U3319 (N_3319,N_3129,N_3203);
xor U3320 (N_3320,N_3207,N_3184);
nor U3321 (N_3321,N_3189,N_3161);
or U3322 (N_3322,N_3225,N_3177);
xor U3323 (N_3323,N_3144,N_3151);
nand U3324 (N_3324,N_3179,N_3215);
or U3325 (N_3325,N_3170,N_3217);
and U3326 (N_3326,N_3230,N_3233);
xnor U3327 (N_3327,N_3202,N_3150);
xor U3328 (N_3328,N_3173,N_3128);
xor U3329 (N_3329,N_3177,N_3156);
and U3330 (N_3330,N_3224,N_3219);
xor U3331 (N_3331,N_3208,N_3213);
or U3332 (N_3332,N_3245,N_3202);
nand U3333 (N_3333,N_3178,N_3204);
or U3334 (N_3334,N_3184,N_3213);
nor U3335 (N_3335,N_3189,N_3205);
nor U3336 (N_3336,N_3125,N_3181);
or U3337 (N_3337,N_3129,N_3237);
and U3338 (N_3338,N_3206,N_3221);
or U3339 (N_3339,N_3197,N_3145);
nand U3340 (N_3340,N_3214,N_3213);
or U3341 (N_3341,N_3224,N_3203);
or U3342 (N_3342,N_3191,N_3221);
nor U3343 (N_3343,N_3147,N_3219);
or U3344 (N_3344,N_3224,N_3194);
and U3345 (N_3345,N_3150,N_3236);
xor U3346 (N_3346,N_3145,N_3210);
and U3347 (N_3347,N_3231,N_3165);
and U3348 (N_3348,N_3237,N_3234);
nor U3349 (N_3349,N_3141,N_3139);
nor U3350 (N_3350,N_3146,N_3145);
or U3351 (N_3351,N_3171,N_3218);
and U3352 (N_3352,N_3145,N_3221);
nor U3353 (N_3353,N_3201,N_3149);
nand U3354 (N_3354,N_3163,N_3202);
or U3355 (N_3355,N_3241,N_3205);
nand U3356 (N_3356,N_3194,N_3150);
xor U3357 (N_3357,N_3187,N_3167);
nor U3358 (N_3358,N_3240,N_3226);
nor U3359 (N_3359,N_3245,N_3223);
nand U3360 (N_3360,N_3125,N_3145);
nor U3361 (N_3361,N_3141,N_3226);
xnor U3362 (N_3362,N_3135,N_3149);
nor U3363 (N_3363,N_3146,N_3176);
nor U3364 (N_3364,N_3169,N_3229);
nand U3365 (N_3365,N_3126,N_3195);
and U3366 (N_3366,N_3221,N_3129);
nand U3367 (N_3367,N_3140,N_3229);
nor U3368 (N_3368,N_3179,N_3133);
nor U3369 (N_3369,N_3190,N_3193);
nand U3370 (N_3370,N_3132,N_3150);
or U3371 (N_3371,N_3224,N_3193);
nor U3372 (N_3372,N_3236,N_3164);
nor U3373 (N_3373,N_3192,N_3163);
nor U3374 (N_3374,N_3130,N_3215);
nor U3375 (N_3375,N_3348,N_3367);
or U3376 (N_3376,N_3360,N_3308);
and U3377 (N_3377,N_3259,N_3301);
nand U3378 (N_3378,N_3276,N_3293);
and U3379 (N_3379,N_3317,N_3289);
nand U3380 (N_3380,N_3334,N_3280);
or U3381 (N_3381,N_3336,N_3267);
and U3382 (N_3382,N_3252,N_3265);
nand U3383 (N_3383,N_3300,N_3342);
and U3384 (N_3384,N_3266,N_3270);
nor U3385 (N_3385,N_3359,N_3304);
or U3386 (N_3386,N_3371,N_3269);
xnor U3387 (N_3387,N_3306,N_3262);
and U3388 (N_3388,N_3286,N_3361);
and U3389 (N_3389,N_3318,N_3330);
or U3390 (N_3390,N_3291,N_3325);
and U3391 (N_3391,N_3366,N_3292);
nand U3392 (N_3392,N_3278,N_3320);
nor U3393 (N_3393,N_3272,N_3290);
or U3394 (N_3394,N_3340,N_3338);
nor U3395 (N_3395,N_3332,N_3327);
and U3396 (N_3396,N_3253,N_3284);
nand U3397 (N_3397,N_3309,N_3322);
nor U3398 (N_3398,N_3313,N_3273);
nand U3399 (N_3399,N_3321,N_3277);
or U3400 (N_3400,N_3365,N_3374);
and U3401 (N_3401,N_3299,N_3261);
nand U3402 (N_3402,N_3312,N_3328);
or U3403 (N_3403,N_3372,N_3370);
nor U3404 (N_3404,N_3307,N_3357);
or U3405 (N_3405,N_3324,N_3294);
nor U3406 (N_3406,N_3285,N_3257);
nand U3407 (N_3407,N_3283,N_3356);
and U3408 (N_3408,N_3369,N_3295);
or U3409 (N_3409,N_3331,N_3274);
xnor U3410 (N_3410,N_3251,N_3329);
nand U3411 (N_3411,N_3279,N_3373);
and U3412 (N_3412,N_3256,N_3275);
xnor U3413 (N_3413,N_3263,N_3260);
or U3414 (N_3414,N_3287,N_3310);
and U3415 (N_3415,N_3302,N_3337);
nand U3416 (N_3416,N_3316,N_3355);
and U3417 (N_3417,N_3323,N_3363);
xor U3418 (N_3418,N_3303,N_3250);
nor U3419 (N_3419,N_3298,N_3345);
or U3420 (N_3420,N_3282,N_3296);
nand U3421 (N_3421,N_3268,N_3254);
or U3422 (N_3422,N_3352,N_3347);
nor U3423 (N_3423,N_3255,N_3305);
xnor U3424 (N_3424,N_3311,N_3351);
and U3425 (N_3425,N_3349,N_3339);
and U3426 (N_3426,N_3288,N_3354);
or U3427 (N_3427,N_3346,N_3362);
and U3428 (N_3428,N_3333,N_3326);
and U3429 (N_3429,N_3353,N_3344);
nand U3430 (N_3430,N_3364,N_3358);
nor U3431 (N_3431,N_3314,N_3264);
and U3432 (N_3432,N_3350,N_3315);
nand U3433 (N_3433,N_3335,N_3343);
or U3434 (N_3434,N_3368,N_3341);
nor U3435 (N_3435,N_3319,N_3281);
and U3436 (N_3436,N_3258,N_3271);
nand U3437 (N_3437,N_3297,N_3277);
or U3438 (N_3438,N_3265,N_3359);
or U3439 (N_3439,N_3261,N_3321);
nor U3440 (N_3440,N_3370,N_3347);
nand U3441 (N_3441,N_3316,N_3321);
nand U3442 (N_3442,N_3295,N_3322);
nand U3443 (N_3443,N_3352,N_3373);
nor U3444 (N_3444,N_3342,N_3314);
nor U3445 (N_3445,N_3361,N_3259);
nand U3446 (N_3446,N_3347,N_3360);
and U3447 (N_3447,N_3313,N_3363);
or U3448 (N_3448,N_3263,N_3372);
nor U3449 (N_3449,N_3374,N_3291);
xor U3450 (N_3450,N_3335,N_3336);
and U3451 (N_3451,N_3342,N_3252);
nor U3452 (N_3452,N_3304,N_3362);
and U3453 (N_3453,N_3250,N_3330);
nor U3454 (N_3454,N_3318,N_3345);
and U3455 (N_3455,N_3364,N_3301);
or U3456 (N_3456,N_3350,N_3339);
and U3457 (N_3457,N_3371,N_3367);
or U3458 (N_3458,N_3323,N_3318);
or U3459 (N_3459,N_3269,N_3363);
nor U3460 (N_3460,N_3344,N_3335);
or U3461 (N_3461,N_3327,N_3259);
or U3462 (N_3462,N_3254,N_3361);
nor U3463 (N_3463,N_3272,N_3373);
nor U3464 (N_3464,N_3307,N_3263);
nand U3465 (N_3465,N_3254,N_3315);
nand U3466 (N_3466,N_3340,N_3347);
or U3467 (N_3467,N_3342,N_3282);
nand U3468 (N_3468,N_3337,N_3301);
and U3469 (N_3469,N_3359,N_3337);
nor U3470 (N_3470,N_3251,N_3370);
nor U3471 (N_3471,N_3329,N_3278);
nor U3472 (N_3472,N_3275,N_3296);
nor U3473 (N_3473,N_3287,N_3309);
and U3474 (N_3474,N_3270,N_3292);
nor U3475 (N_3475,N_3272,N_3277);
nand U3476 (N_3476,N_3267,N_3282);
or U3477 (N_3477,N_3273,N_3256);
and U3478 (N_3478,N_3262,N_3303);
nor U3479 (N_3479,N_3329,N_3274);
nor U3480 (N_3480,N_3277,N_3288);
or U3481 (N_3481,N_3265,N_3268);
xor U3482 (N_3482,N_3330,N_3269);
and U3483 (N_3483,N_3317,N_3336);
nand U3484 (N_3484,N_3304,N_3285);
and U3485 (N_3485,N_3285,N_3298);
nand U3486 (N_3486,N_3297,N_3354);
nor U3487 (N_3487,N_3297,N_3266);
nand U3488 (N_3488,N_3367,N_3333);
and U3489 (N_3489,N_3303,N_3288);
and U3490 (N_3490,N_3355,N_3359);
and U3491 (N_3491,N_3354,N_3316);
nor U3492 (N_3492,N_3296,N_3313);
nand U3493 (N_3493,N_3253,N_3294);
nand U3494 (N_3494,N_3267,N_3330);
xor U3495 (N_3495,N_3259,N_3275);
xor U3496 (N_3496,N_3283,N_3321);
or U3497 (N_3497,N_3269,N_3362);
or U3498 (N_3498,N_3320,N_3356);
nor U3499 (N_3499,N_3365,N_3305);
xor U3500 (N_3500,N_3377,N_3463);
or U3501 (N_3501,N_3401,N_3467);
nand U3502 (N_3502,N_3475,N_3411);
nor U3503 (N_3503,N_3472,N_3464);
nor U3504 (N_3504,N_3445,N_3394);
and U3505 (N_3505,N_3422,N_3421);
nor U3506 (N_3506,N_3444,N_3496);
and U3507 (N_3507,N_3447,N_3451);
nand U3508 (N_3508,N_3487,N_3416);
nand U3509 (N_3509,N_3390,N_3381);
xnor U3510 (N_3510,N_3430,N_3468);
and U3511 (N_3511,N_3406,N_3498);
xnor U3512 (N_3512,N_3458,N_3392);
nor U3513 (N_3513,N_3453,N_3462);
and U3514 (N_3514,N_3480,N_3499);
nor U3515 (N_3515,N_3449,N_3461);
or U3516 (N_3516,N_3409,N_3400);
or U3517 (N_3517,N_3488,N_3443);
or U3518 (N_3518,N_3380,N_3433);
nor U3519 (N_3519,N_3379,N_3479);
or U3520 (N_3520,N_3396,N_3413);
nor U3521 (N_3521,N_3491,N_3484);
and U3522 (N_3522,N_3474,N_3417);
nor U3523 (N_3523,N_3408,N_3442);
xor U3524 (N_3524,N_3375,N_3405);
and U3525 (N_3525,N_3437,N_3399);
nand U3526 (N_3526,N_3391,N_3495);
and U3527 (N_3527,N_3482,N_3448);
xnor U3528 (N_3528,N_3489,N_3469);
or U3529 (N_3529,N_3465,N_3393);
nand U3530 (N_3530,N_3450,N_3497);
nor U3531 (N_3531,N_3492,N_3490);
nand U3532 (N_3532,N_3420,N_3471);
xnor U3533 (N_3533,N_3473,N_3436);
and U3534 (N_3534,N_3425,N_3383);
xor U3535 (N_3535,N_3427,N_3441);
and U3536 (N_3536,N_3477,N_3459);
and U3537 (N_3537,N_3438,N_3423);
xor U3538 (N_3538,N_3429,N_3403);
nand U3539 (N_3539,N_3386,N_3434);
or U3540 (N_3540,N_3428,N_3454);
or U3541 (N_3541,N_3414,N_3440);
xor U3542 (N_3542,N_3395,N_3452);
nor U3543 (N_3543,N_3376,N_3388);
nor U3544 (N_3544,N_3457,N_3446);
nand U3545 (N_3545,N_3424,N_3466);
nand U3546 (N_3546,N_3415,N_3404);
or U3547 (N_3547,N_3456,N_3397);
nor U3548 (N_3548,N_3483,N_3410);
and U3549 (N_3549,N_3432,N_3470);
and U3550 (N_3550,N_3486,N_3485);
and U3551 (N_3551,N_3384,N_3493);
and U3552 (N_3552,N_3478,N_3426);
nand U3553 (N_3553,N_3435,N_3494);
and U3554 (N_3554,N_3387,N_3385);
xnor U3555 (N_3555,N_3431,N_3481);
and U3556 (N_3556,N_3389,N_3402);
and U3557 (N_3557,N_3418,N_3398);
nor U3558 (N_3558,N_3412,N_3378);
nor U3559 (N_3559,N_3455,N_3460);
and U3560 (N_3560,N_3476,N_3419);
and U3561 (N_3561,N_3439,N_3407);
or U3562 (N_3562,N_3382,N_3394);
nor U3563 (N_3563,N_3473,N_3460);
or U3564 (N_3564,N_3483,N_3477);
xor U3565 (N_3565,N_3451,N_3455);
nand U3566 (N_3566,N_3467,N_3475);
and U3567 (N_3567,N_3487,N_3420);
and U3568 (N_3568,N_3379,N_3428);
and U3569 (N_3569,N_3444,N_3413);
nand U3570 (N_3570,N_3462,N_3410);
and U3571 (N_3571,N_3430,N_3420);
and U3572 (N_3572,N_3415,N_3479);
and U3573 (N_3573,N_3496,N_3387);
or U3574 (N_3574,N_3443,N_3436);
nand U3575 (N_3575,N_3389,N_3435);
and U3576 (N_3576,N_3436,N_3438);
and U3577 (N_3577,N_3418,N_3441);
or U3578 (N_3578,N_3438,N_3379);
and U3579 (N_3579,N_3494,N_3434);
or U3580 (N_3580,N_3398,N_3424);
and U3581 (N_3581,N_3383,N_3491);
nand U3582 (N_3582,N_3391,N_3450);
and U3583 (N_3583,N_3442,N_3419);
nor U3584 (N_3584,N_3492,N_3482);
or U3585 (N_3585,N_3392,N_3472);
xnor U3586 (N_3586,N_3395,N_3461);
and U3587 (N_3587,N_3444,N_3425);
nand U3588 (N_3588,N_3440,N_3472);
nand U3589 (N_3589,N_3423,N_3466);
and U3590 (N_3590,N_3376,N_3387);
or U3591 (N_3591,N_3440,N_3486);
nor U3592 (N_3592,N_3376,N_3471);
nand U3593 (N_3593,N_3441,N_3377);
or U3594 (N_3594,N_3461,N_3410);
nand U3595 (N_3595,N_3390,N_3471);
or U3596 (N_3596,N_3441,N_3490);
nor U3597 (N_3597,N_3390,N_3430);
and U3598 (N_3598,N_3442,N_3395);
or U3599 (N_3599,N_3448,N_3434);
or U3600 (N_3600,N_3454,N_3493);
and U3601 (N_3601,N_3399,N_3451);
xor U3602 (N_3602,N_3482,N_3391);
nand U3603 (N_3603,N_3375,N_3389);
nand U3604 (N_3604,N_3390,N_3491);
or U3605 (N_3605,N_3461,N_3432);
nand U3606 (N_3606,N_3469,N_3493);
nor U3607 (N_3607,N_3452,N_3391);
or U3608 (N_3608,N_3451,N_3492);
or U3609 (N_3609,N_3403,N_3443);
nand U3610 (N_3610,N_3412,N_3431);
nor U3611 (N_3611,N_3479,N_3455);
or U3612 (N_3612,N_3424,N_3381);
and U3613 (N_3613,N_3384,N_3392);
or U3614 (N_3614,N_3403,N_3486);
and U3615 (N_3615,N_3457,N_3411);
or U3616 (N_3616,N_3410,N_3491);
and U3617 (N_3617,N_3385,N_3376);
and U3618 (N_3618,N_3417,N_3450);
nand U3619 (N_3619,N_3390,N_3384);
nor U3620 (N_3620,N_3434,N_3495);
or U3621 (N_3621,N_3480,N_3419);
and U3622 (N_3622,N_3376,N_3377);
nand U3623 (N_3623,N_3413,N_3416);
nand U3624 (N_3624,N_3468,N_3400);
and U3625 (N_3625,N_3531,N_3520);
nor U3626 (N_3626,N_3557,N_3552);
or U3627 (N_3627,N_3590,N_3501);
nor U3628 (N_3628,N_3553,N_3570);
nand U3629 (N_3629,N_3514,N_3601);
nand U3630 (N_3630,N_3603,N_3517);
nor U3631 (N_3631,N_3507,N_3618);
or U3632 (N_3632,N_3530,N_3592);
or U3633 (N_3633,N_3577,N_3622);
nor U3634 (N_3634,N_3615,N_3575);
xor U3635 (N_3635,N_3524,N_3582);
nand U3636 (N_3636,N_3594,N_3574);
nor U3637 (N_3637,N_3542,N_3536);
or U3638 (N_3638,N_3543,N_3528);
or U3639 (N_3639,N_3541,N_3579);
nand U3640 (N_3640,N_3581,N_3556);
nand U3641 (N_3641,N_3620,N_3518);
and U3642 (N_3642,N_3521,N_3619);
nor U3643 (N_3643,N_3529,N_3554);
nor U3644 (N_3644,N_3546,N_3578);
or U3645 (N_3645,N_3599,N_3563);
and U3646 (N_3646,N_3540,N_3608);
nor U3647 (N_3647,N_3526,N_3616);
and U3648 (N_3648,N_3564,N_3527);
nand U3649 (N_3649,N_3606,N_3534);
nand U3650 (N_3650,N_3607,N_3509);
xor U3651 (N_3651,N_3600,N_3512);
and U3652 (N_3652,N_3572,N_3547);
nand U3653 (N_3653,N_3614,N_3588);
nand U3654 (N_3654,N_3567,N_3510);
or U3655 (N_3655,N_3576,N_3593);
and U3656 (N_3656,N_3597,N_3612);
nor U3657 (N_3657,N_3555,N_3500);
or U3658 (N_3658,N_3515,N_3605);
and U3659 (N_3659,N_3624,N_3586);
xnor U3660 (N_3660,N_3568,N_3504);
nor U3661 (N_3661,N_3584,N_3589);
nor U3662 (N_3662,N_3511,N_3580);
and U3663 (N_3663,N_3532,N_3573);
and U3664 (N_3664,N_3623,N_3566);
and U3665 (N_3665,N_3559,N_3537);
nor U3666 (N_3666,N_3587,N_3591);
nor U3667 (N_3667,N_3544,N_3551);
nand U3668 (N_3668,N_3583,N_3525);
nor U3669 (N_3669,N_3569,N_3560);
and U3670 (N_3670,N_3558,N_3621);
nor U3671 (N_3671,N_3549,N_3595);
xor U3672 (N_3672,N_3545,N_3611);
xor U3673 (N_3673,N_3503,N_3522);
and U3674 (N_3674,N_3550,N_3596);
nand U3675 (N_3675,N_3535,N_3565);
nor U3676 (N_3676,N_3513,N_3502);
or U3677 (N_3677,N_3617,N_3533);
nand U3678 (N_3678,N_3585,N_3613);
or U3679 (N_3679,N_3562,N_3505);
nand U3680 (N_3680,N_3609,N_3516);
xor U3681 (N_3681,N_3539,N_3610);
or U3682 (N_3682,N_3519,N_3571);
nand U3683 (N_3683,N_3506,N_3602);
and U3684 (N_3684,N_3538,N_3604);
nand U3685 (N_3685,N_3508,N_3523);
or U3686 (N_3686,N_3561,N_3598);
nor U3687 (N_3687,N_3548,N_3559);
nor U3688 (N_3688,N_3565,N_3595);
nor U3689 (N_3689,N_3615,N_3574);
nor U3690 (N_3690,N_3587,N_3564);
nor U3691 (N_3691,N_3557,N_3548);
or U3692 (N_3692,N_3514,N_3607);
or U3693 (N_3693,N_3523,N_3516);
xor U3694 (N_3694,N_3569,N_3540);
xnor U3695 (N_3695,N_3590,N_3612);
and U3696 (N_3696,N_3515,N_3574);
or U3697 (N_3697,N_3509,N_3512);
nand U3698 (N_3698,N_3502,N_3549);
nand U3699 (N_3699,N_3517,N_3508);
or U3700 (N_3700,N_3578,N_3569);
or U3701 (N_3701,N_3567,N_3589);
and U3702 (N_3702,N_3599,N_3533);
or U3703 (N_3703,N_3616,N_3617);
nor U3704 (N_3704,N_3573,N_3517);
nand U3705 (N_3705,N_3602,N_3509);
and U3706 (N_3706,N_3562,N_3514);
or U3707 (N_3707,N_3586,N_3534);
nand U3708 (N_3708,N_3590,N_3619);
or U3709 (N_3709,N_3579,N_3530);
nand U3710 (N_3710,N_3558,N_3508);
xnor U3711 (N_3711,N_3597,N_3594);
and U3712 (N_3712,N_3546,N_3615);
or U3713 (N_3713,N_3502,N_3617);
nand U3714 (N_3714,N_3506,N_3593);
and U3715 (N_3715,N_3616,N_3578);
nand U3716 (N_3716,N_3504,N_3602);
and U3717 (N_3717,N_3562,N_3554);
and U3718 (N_3718,N_3516,N_3533);
or U3719 (N_3719,N_3520,N_3567);
nand U3720 (N_3720,N_3533,N_3527);
or U3721 (N_3721,N_3607,N_3590);
or U3722 (N_3722,N_3548,N_3519);
nand U3723 (N_3723,N_3624,N_3565);
nor U3724 (N_3724,N_3586,N_3610);
or U3725 (N_3725,N_3532,N_3571);
and U3726 (N_3726,N_3545,N_3589);
and U3727 (N_3727,N_3507,N_3512);
nand U3728 (N_3728,N_3521,N_3611);
or U3729 (N_3729,N_3583,N_3599);
nor U3730 (N_3730,N_3600,N_3597);
nor U3731 (N_3731,N_3618,N_3539);
and U3732 (N_3732,N_3599,N_3603);
nor U3733 (N_3733,N_3558,N_3584);
nand U3734 (N_3734,N_3553,N_3563);
or U3735 (N_3735,N_3503,N_3549);
or U3736 (N_3736,N_3519,N_3501);
xnor U3737 (N_3737,N_3552,N_3592);
nand U3738 (N_3738,N_3606,N_3594);
nand U3739 (N_3739,N_3591,N_3615);
xnor U3740 (N_3740,N_3513,N_3620);
or U3741 (N_3741,N_3620,N_3504);
nand U3742 (N_3742,N_3563,N_3524);
or U3743 (N_3743,N_3547,N_3579);
or U3744 (N_3744,N_3603,N_3529);
nor U3745 (N_3745,N_3530,N_3606);
and U3746 (N_3746,N_3597,N_3610);
xor U3747 (N_3747,N_3598,N_3546);
or U3748 (N_3748,N_3559,N_3575);
or U3749 (N_3749,N_3525,N_3599);
and U3750 (N_3750,N_3711,N_3665);
and U3751 (N_3751,N_3745,N_3676);
and U3752 (N_3752,N_3695,N_3741);
or U3753 (N_3753,N_3697,N_3725);
or U3754 (N_3754,N_3634,N_3669);
and U3755 (N_3755,N_3687,N_3718);
xor U3756 (N_3756,N_3650,N_3628);
nand U3757 (N_3757,N_3675,N_3679);
or U3758 (N_3758,N_3668,N_3646);
or U3759 (N_3759,N_3678,N_3660);
or U3760 (N_3760,N_3728,N_3655);
xnor U3761 (N_3761,N_3626,N_3686);
nor U3762 (N_3762,N_3661,N_3713);
nand U3763 (N_3763,N_3719,N_3707);
and U3764 (N_3764,N_3627,N_3690);
or U3765 (N_3765,N_3736,N_3632);
nand U3766 (N_3766,N_3702,N_3699);
or U3767 (N_3767,N_3683,N_3629);
xnor U3768 (N_3768,N_3746,N_3649);
nor U3769 (N_3769,N_3724,N_3656);
nor U3770 (N_3770,N_3696,N_3652);
xor U3771 (N_3771,N_3734,N_3659);
nand U3772 (N_3772,N_3645,N_3743);
or U3773 (N_3773,N_3638,N_3693);
and U3774 (N_3774,N_3643,N_3726);
and U3775 (N_3775,N_3733,N_3653);
and U3776 (N_3776,N_3705,N_3709);
or U3777 (N_3777,N_3747,N_3640);
nand U3778 (N_3778,N_3671,N_3644);
xor U3779 (N_3779,N_3721,N_3714);
nor U3780 (N_3780,N_3636,N_3704);
xor U3781 (N_3781,N_3729,N_3694);
nand U3782 (N_3782,N_3658,N_3674);
nor U3783 (N_3783,N_3685,N_3664);
or U3784 (N_3784,N_3625,N_3737);
or U3785 (N_3785,N_3630,N_3680);
xnor U3786 (N_3786,N_3739,N_3722);
or U3787 (N_3787,N_3723,N_3727);
and U3788 (N_3788,N_3672,N_3700);
nand U3789 (N_3789,N_3716,N_3703);
or U3790 (N_3790,N_3682,N_3712);
or U3791 (N_3791,N_3633,N_3647);
or U3792 (N_3792,N_3648,N_3641);
and U3793 (N_3793,N_3720,N_3730);
nand U3794 (N_3794,N_3662,N_3715);
and U3795 (N_3795,N_3731,N_3701);
nand U3796 (N_3796,N_3684,N_3639);
xor U3797 (N_3797,N_3698,N_3706);
nor U3798 (N_3798,N_3635,N_3748);
nand U3799 (N_3799,N_3689,N_3688);
xnor U3800 (N_3800,N_3657,N_3654);
and U3801 (N_3801,N_3637,N_3663);
or U3802 (N_3802,N_3742,N_3670);
nand U3803 (N_3803,N_3717,N_3740);
or U3804 (N_3804,N_3749,N_3744);
or U3805 (N_3805,N_3677,N_3667);
xnor U3806 (N_3806,N_3631,N_3738);
and U3807 (N_3807,N_3735,N_3673);
or U3808 (N_3808,N_3710,N_3666);
nor U3809 (N_3809,N_3681,N_3642);
nor U3810 (N_3810,N_3692,N_3651);
nor U3811 (N_3811,N_3708,N_3732);
or U3812 (N_3812,N_3691,N_3685);
and U3813 (N_3813,N_3749,N_3699);
nand U3814 (N_3814,N_3732,N_3679);
nor U3815 (N_3815,N_3680,N_3721);
nand U3816 (N_3816,N_3699,N_3627);
or U3817 (N_3817,N_3712,N_3703);
and U3818 (N_3818,N_3704,N_3702);
nor U3819 (N_3819,N_3640,N_3651);
nor U3820 (N_3820,N_3649,N_3626);
nor U3821 (N_3821,N_3727,N_3634);
and U3822 (N_3822,N_3653,N_3658);
and U3823 (N_3823,N_3691,N_3689);
and U3824 (N_3824,N_3738,N_3671);
and U3825 (N_3825,N_3709,N_3642);
or U3826 (N_3826,N_3740,N_3707);
nor U3827 (N_3827,N_3728,N_3647);
nand U3828 (N_3828,N_3633,N_3663);
and U3829 (N_3829,N_3644,N_3735);
nand U3830 (N_3830,N_3643,N_3664);
or U3831 (N_3831,N_3643,N_3708);
nand U3832 (N_3832,N_3633,N_3696);
nor U3833 (N_3833,N_3638,N_3629);
nand U3834 (N_3834,N_3735,N_3705);
nand U3835 (N_3835,N_3668,N_3708);
nand U3836 (N_3836,N_3682,N_3707);
or U3837 (N_3837,N_3748,N_3697);
or U3838 (N_3838,N_3626,N_3655);
nor U3839 (N_3839,N_3634,N_3654);
or U3840 (N_3840,N_3664,N_3675);
nand U3841 (N_3841,N_3673,N_3709);
nor U3842 (N_3842,N_3736,N_3635);
and U3843 (N_3843,N_3713,N_3739);
nand U3844 (N_3844,N_3708,N_3731);
nor U3845 (N_3845,N_3633,N_3690);
and U3846 (N_3846,N_3696,N_3653);
xor U3847 (N_3847,N_3729,N_3718);
xnor U3848 (N_3848,N_3739,N_3648);
nor U3849 (N_3849,N_3685,N_3708);
or U3850 (N_3850,N_3714,N_3738);
or U3851 (N_3851,N_3669,N_3640);
nor U3852 (N_3852,N_3738,N_3696);
nor U3853 (N_3853,N_3747,N_3717);
nor U3854 (N_3854,N_3701,N_3670);
nor U3855 (N_3855,N_3678,N_3718);
or U3856 (N_3856,N_3673,N_3714);
nand U3857 (N_3857,N_3655,N_3644);
nand U3858 (N_3858,N_3658,N_3733);
nor U3859 (N_3859,N_3722,N_3662);
and U3860 (N_3860,N_3683,N_3672);
or U3861 (N_3861,N_3686,N_3724);
and U3862 (N_3862,N_3663,N_3671);
nor U3863 (N_3863,N_3652,N_3659);
and U3864 (N_3864,N_3746,N_3665);
or U3865 (N_3865,N_3676,N_3719);
and U3866 (N_3866,N_3719,N_3657);
nand U3867 (N_3867,N_3646,N_3705);
and U3868 (N_3868,N_3704,N_3694);
and U3869 (N_3869,N_3748,N_3734);
or U3870 (N_3870,N_3654,N_3648);
nor U3871 (N_3871,N_3713,N_3709);
nor U3872 (N_3872,N_3737,N_3746);
or U3873 (N_3873,N_3690,N_3696);
nand U3874 (N_3874,N_3679,N_3741);
and U3875 (N_3875,N_3864,N_3782);
nor U3876 (N_3876,N_3810,N_3779);
nor U3877 (N_3877,N_3768,N_3823);
and U3878 (N_3878,N_3755,N_3840);
or U3879 (N_3879,N_3872,N_3786);
and U3880 (N_3880,N_3844,N_3843);
nand U3881 (N_3881,N_3852,N_3771);
xor U3882 (N_3882,N_3820,N_3776);
or U3883 (N_3883,N_3766,N_3773);
nand U3884 (N_3884,N_3764,N_3870);
and U3885 (N_3885,N_3866,N_3860);
xor U3886 (N_3886,N_3835,N_3759);
or U3887 (N_3887,N_3763,N_3791);
nor U3888 (N_3888,N_3784,N_3853);
nor U3889 (N_3889,N_3774,N_3781);
or U3890 (N_3890,N_3775,N_3858);
or U3891 (N_3891,N_3760,N_3797);
or U3892 (N_3892,N_3854,N_3802);
and U3893 (N_3893,N_3762,N_3809);
nor U3894 (N_3894,N_3777,N_3805);
xor U3895 (N_3895,N_3849,N_3825);
nand U3896 (N_3896,N_3831,N_3850);
or U3897 (N_3897,N_3874,N_3804);
and U3898 (N_3898,N_3796,N_3868);
and U3899 (N_3899,N_3811,N_3756);
nand U3900 (N_3900,N_3750,N_3833);
nand U3901 (N_3901,N_3821,N_3807);
nand U3902 (N_3902,N_3790,N_3846);
nor U3903 (N_3903,N_3818,N_3801);
nor U3904 (N_3904,N_3837,N_3871);
and U3905 (N_3905,N_3867,N_3800);
nor U3906 (N_3906,N_3841,N_3865);
xor U3907 (N_3907,N_3824,N_3753);
or U3908 (N_3908,N_3863,N_3859);
xnor U3909 (N_3909,N_3813,N_3808);
nor U3910 (N_3910,N_3799,N_3803);
or U3911 (N_3911,N_3798,N_3838);
and U3912 (N_3912,N_3847,N_3829);
or U3913 (N_3913,N_3839,N_3778);
nand U3914 (N_3914,N_3752,N_3792);
nand U3915 (N_3915,N_3830,N_3780);
or U3916 (N_3916,N_3817,N_3855);
nor U3917 (N_3917,N_3851,N_3783);
xnor U3918 (N_3918,N_3814,N_3856);
nor U3919 (N_3919,N_3857,N_3861);
nand U3920 (N_3920,N_3765,N_3836);
or U3921 (N_3921,N_3787,N_3826);
nor U3922 (N_3922,N_3751,N_3828);
nand U3923 (N_3923,N_3757,N_3827);
and U3924 (N_3924,N_3832,N_3815);
nor U3925 (N_3925,N_3785,N_3873);
nor U3926 (N_3926,N_3772,N_3812);
xor U3927 (N_3927,N_3789,N_3822);
and U3928 (N_3928,N_3794,N_3761);
xor U3929 (N_3929,N_3819,N_3842);
nand U3930 (N_3930,N_3816,N_3793);
or U3931 (N_3931,N_3806,N_3869);
and U3932 (N_3932,N_3788,N_3795);
nand U3933 (N_3933,N_3758,N_3767);
and U3934 (N_3934,N_3769,N_3834);
xor U3935 (N_3935,N_3862,N_3770);
or U3936 (N_3936,N_3848,N_3845);
xor U3937 (N_3937,N_3754,N_3827);
nand U3938 (N_3938,N_3796,N_3840);
nand U3939 (N_3939,N_3773,N_3820);
or U3940 (N_3940,N_3774,N_3812);
nor U3941 (N_3941,N_3762,N_3834);
or U3942 (N_3942,N_3790,N_3768);
or U3943 (N_3943,N_3834,N_3757);
or U3944 (N_3944,N_3808,N_3802);
and U3945 (N_3945,N_3764,N_3862);
nand U3946 (N_3946,N_3816,N_3768);
or U3947 (N_3947,N_3832,N_3852);
and U3948 (N_3948,N_3858,N_3783);
xor U3949 (N_3949,N_3758,N_3803);
xor U3950 (N_3950,N_3752,N_3784);
or U3951 (N_3951,N_3833,N_3860);
or U3952 (N_3952,N_3783,N_3853);
and U3953 (N_3953,N_3754,N_3857);
and U3954 (N_3954,N_3771,N_3804);
and U3955 (N_3955,N_3771,N_3753);
xnor U3956 (N_3956,N_3763,N_3786);
and U3957 (N_3957,N_3750,N_3817);
or U3958 (N_3958,N_3862,N_3817);
and U3959 (N_3959,N_3824,N_3858);
or U3960 (N_3960,N_3832,N_3861);
and U3961 (N_3961,N_3803,N_3792);
and U3962 (N_3962,N_3827,N_3848);
nor U3963 (N_3963,N_3825,N_3771);
and U3964 (N_3964,N_3857,N_3809);
nor U3965 (N_3965,N_3872,N_3849);
nand U3966 (N_3966,N_3807,N_3812);
and U3967 (N_3967,N_3791,N_3839);
and U3968 (N_3968,N_3789,N_3762);
nand U3969 (N_3969,N_3838,N_3826);
nand U3970 (N_3970,N_3797,N_3778);
and U3971 (N_3971,N_3850,N_3758);
xor U3972 (N_3972,N_3813,N_3860);
and U3973 (N_3973,N_3825,N_3870);
and U3974 (N_3974,N_3798,N_3767);
nand U3975 (N_3975,N_3871,N_3822);
xor U3976 (N_3976,N_3868,N_3816);
xnor U3977 (N_3977,N_3776,N_3794);
and U3978 (N_3978,N_3808,N_3784);
nor U3979 (N_3979,N_3823,N_3794);
and U3980 (N_3980,N_3806,N_3842);
or U3981 (N_3981,N_3831,N_3766);
nand U3982 (N_3982,N_3772,N_3770);
and U3983 (N_3983,N_3797,N_3833);
nand U3984 (N_3984,N_3792,N_3834);
nor U3985 (N_3985,N_3796,N_3821);
nor U3986 (N_3986,N_3831,N_3784);
nor U3987 (N_3987,N_3819,N_3768);
nor U3988 (N_3988,N_3772,N_3824);
nand U3989 (N_3989,N_3810,N_3786);
and U3990 (N_3990,N_3793,N_3810);
nand U3991 (N_3991,N_3776,N_3771);
or U3992 (N_3992,N_3854,N_3853);
nor U3993 (N_3993,N_3774,N_3800);
nand U3994 (N_3994,N_3839,N_3832);
nand U3995 (N_3995,N_3779,N_3845);
nand U3996 (N_3996,N_3813,N_3767);
nand U3997 (N_3997,N_3826,N_3821);
and U3998 (N_3998,N_3769,N_3812);
nor U3999 (N_3999,N_3860,N_3803);
and U4000 (N_4000,N_3916,N_3990);
or U4001 (N_4001,N_3921,N_3949);
and U4002 (N_4002,N_3943,N_3954);
and U4003 (N_4003,N_3937,N_3907);
and U4004 (N_4004,N_3987,N_3945);
nor U4005 (N_4005,N_3974,N_3932);
or U4006 (N_4006,N_3890,N_3884);
nor U4007 (N_4007,N_3982,N_3967);
xnor U4008 (N_4008,N_3924,N_3951);
and U4009 (N_4009,N_3935,N_3956);
and U4010 (N_4010,N_3995,N_3959);
xnor U4011 (N_4011,N_3888,N_3920);
and U4012 (N_4012,N_3986,N_3977);
nor U4013 (N_4013,N_3975,N_3952);
or U4014 (N_4014,N_3904,N_3998);
nor U4015 (N_4015,N_3985,N_3912);
or U4016 (N_4016,N_3882,N_3946);
nor U4017 (N_4017,N_3915,N_3894);
or U4018 (N_4018,N_3942,N_3876);
and U4019 (N_4019,N_3978,N_3941);
nand U4020 (N_4020,N_3897,N_3961);
nand U4021 (N_4021,N_3996,N_3976);
xnor U4022 (N_4022,N_3908,N_3992);
or U4023 (N_4023,N_3925,N_3968);
and U4024 (N_4024,N_3938,N_3940);
or U4025 (N_4025,N_3947,N_3997);
xor U4026 (N_4026,N_3910,N_3944);
nand U4027 (N_4027,N_3896,N_3929);
nor U4028 (N_4028,N_3971,N_3972);
nand U4029 (N_4029,N_3957,N_3955);
and U4030 (N_4030,N_3988,N_3934);
or U4031 (N_4031,N_3983,N_3948);
nor U4032 (N_4032,N_3979,N_3886);
or U4033 (N_4033,N_3991,N_3919);
or U4034 (N_4034,N_3994,N_3928);
and U4035 (N_4035,N_3939,N_3926);
or U4036 (N_4036,N_3981,N_3893);
nand U4037 (N_4037,N_3905,N_3973);
and U4038 (N_4038,N_3962,N_3958);
nand U4039 (N_4039,N_3980,N_3885);
nand U4040 (N_4040,N_3993,N_3898);
or U4041 (N_4041,N_3892,N_3902);
xor U4042 (N_4042,N_3953,N_3984);
nand U4043 (N_4043,N_3989,N_3917);
and U4044 (N_4044,N_3911,N_3965);
nor U4045 (N_4045,N_3963,N_3875);
xor U4046 (N_4046,N_3930,N_3966);
nor U4047 (N_4047,N_3891,N_3901);
nand U4048 (N_4048,N_3881,N_3936);
and U4049 (N_4049,N_3909,N_3900);
nor U4050 (N_4050,N_3931,N_3879);
nand U4051 (N_4051,N_3889,N_3903);
nand U4052 (N_4052,N_3883,N_3877);
or U4053 (N_4053,N_3933,N_3969);
and U4054 (N_4054,N_3914,N_3970);
and U4055 (N_4055,N_3923,N_3895);
and U4056 (N_4056,N_3906,N_3922);
nand U4057 (N_4057,N_3899,N_3950);
and U4058 (N_4058,N_3918,N_3887);
or U4059 (N_4059,N_3960,N_3880);
nand U4060 (N_4060,N_3964,N_3999);
nor U4061 (N_4061,N_3927,N_3913);
nor U4062 (N_4062,N_3878,N_3947);
or U4063 (N_4063,N_3899,N_3895);
nor U4064 (N_4064,N_3997,N_3934);
nand U4065 (N_4065,N_3885,N_3995);
or U4066 (N_4066,N_3878,N_3897);
or U4067 (N_4067,N_3901,N_3953);
or U4068 (N_4068,N_3916,N_3918);
and U4069 (N_4069,N_3881,N_3984);
nor U4070 (N_4070,N_3953,N_3918);
and U4071 (N_4071,N_3933,N_3884);
xnor U4072 (N_4072,N_3904,N_3971);
and U4073 (N_4073,N_3938,N_3875);
or U4074 (N_4074,N_3892,N_3939);
nand U4075 (N_4075,N_3928,N_3905);
or U4076 (N_4076,N_3931,N_3885);
and U4077 (N_4077,N_3920,N_3947);
nand U4078 (N_4078,N_3992,N_3922);
nor U4079 (N_4079,N_3982,N_3894);
xor U4080 (N_4080,N_3930,N_3980);
and U4081 (N_4081,N_3905,N_3994);
or U4082 (N_4082,N_3937,N_3989);
or U4083 (N_4083,N_3952,N_3879);
and U4084 (N_4084,N_3995,N_3894);
or U4085 (N_4085,N_3982,N_3908);
nor U4086 (N_4086,N_3915,N_3969);
nand U4087 (N_4087,N_3894,N_3944);
or U4088 (N_4088,N_3978,N_3975);
nand U4089 (N_4089,N_3975,N_3905);
nand U4090 (N_4090,N_3907,N_3976);
nand U4091 (N_4091,N_3931,N_3975);
and U4092 (N_4092,N_3975,N_3972);
or U4093 (N_4093,N_3947,N_3936);
and U4094 (N_4094,N_3880,N_3990);
or U4095 (N_4095,N_3961,N_3910);
nand U4096 (N_4096,N_3942,N_3976);
nor U4097 (N_4097,N_3910,N_3938);
and U4098 (N_4098,N_3883,N_3986);
or U4099 (N_4099,N_3931,N_3966);
and U4100 (N_4100,N_3875,N_3989);
and U4101 (N_4101,N_3897,N_3942);
or U4102 (N_4102,N_3896,N_3939);
xnor U4103 (N_4103,N_3892,N_3898);
xnor U4104 (N_4104,N_3975,N_3945);
nor U4105 (N_4105,N_3967,N_3906);
or U4106 (N_4106,N_3881,N_3905);
nor U4107 (N_4107,N_3915,N_3892);
and U4108 (N_4108,N_3944,N_3955);
and U4109 (N_4109,N_3923,N_3884);
nor U4110 (N_4110,N_3931,N_3892);
or U4111 (N_4111,N_3906,N_3893);
xnor U4112 (N_4112,N_3899,N_3979);
nand U4113 (N_4113,N_3904,N_3975);
or U4114 (N_4114,N_3961,N_3891);
and U4115 (N_4115,N_3949,N_3993);
nor U4116 (N_4116,N_3937,N_3896);
and U4117 (N_4117,N_3949,N_3956);
or U4118 (N_4118,N_3943,N_3877);
nand U4119 (N_4119,N_3992,N_3930);
nor U4120 (N_4120,N_3943,N_3985);
nor U4121 (N_4121,N_3939,N_3904);
nand U4122 (N_4122,N_3975,N_3878);
nand U4123 (N_4123,N_3939,N_3972);
and U4124 (N_4124,N_3973,N_3896);
nand U4125 (N_4125,N_4086,N_4020);
nand U4126 (N_4126,N_4091,N_4057);
nand U4127 (N_4127,N_4061,N_4118);
and U4128 (N_4128,N_4036,N_4101);
or U4129 (N_4129,N_4046,N_4002);
nand U4130 (N_4130,N_4056,N_4037);
nand U4131 (N_4131,N_4010,N_4021);
nand U4132 (N_4132,N_4060,N_4063);
nor U4133 (N_4133,N_4085,N_4075);
or U4134 (N_4134,N_4108,N_4105);
and U4135 (N_4135,N_4032,N_4041);
or U4136 (N_4136,N_4038,N_4109);
or U4137 (N_4137,N_4117,N_4064);
nor U4138 (N_4138,N_4051,N_4017);
or U4139 (N_4139,N_4080,N_4062);
nand U4140 (N_4140,N_4083,N_4058);
nor U4141 (N_4141,N_4072,N_4115);
and U4142 (N_4142,N_4113,N_4090);
nand U4143 (N_4143,N_4034,N_4013);
nand U4144 (N_4144,N_4102,N_4001);
nand U4145 (N_4145,N_4107,N_4122);
nor U4146 (N_4146,N_4103,N_4049);
and U4147 (N_4147,N_4027,N_4048);
nand U4148 (N_4148,N_4081,N_4093);
and U4149 (N_4149,N_4026,N_4014);
or U4150 (N_4150,N_4025,N_4047);
nand U4151 (N_4151,N_4096,N_4076);
nor U4152 (N_4152,N_4011,N_4069);
or U4153 (N_4153,N_4124,N_4016);
nand U4154 (N_4154,N_4116,N_4029);
and U4155 (N_4155,N_4071,N_4054);
nand U4156 (N_4156,N_4078,N_4007);
or U4157 (N_4157,N_4119,N_4031);
nor U4158 (N_4158,N_4123,N_4092);
or U4159 (N_4159,N_4073,N_4006);
nand U4160 (N_4160,N_4114,N_4094);
nor U4161 (N_4161,N_4023,N_4120);
nand U4162 (N_4162,N_4100,N_4104);
nand U4163 (N_4163,N_4004,N_4084);
and U4164 (N_4164,N_4019,N_4039);
nand U4165 (N_4165,N_4012,N_4077);
and U4166 (N_4166,N_4005,N_4044);
nor U4167 (N_4167,N_4030,N_4098);
and U4168 (N_4168,N_4065,N_4015);
nor U4169 (N_4169,N_4043,N_4035);
xnor U4170 (N_4170,N_4087,N_4045);
xor U4171 (N_4171,N_4070,N_4059);
nand U4172 (N_4172,N_4028,N_4009);
nand U4173 (N_4173,N_4095,N_4111);
nor U4174 (N_4174,N_4121,N_4074);
xnor U4175 (N_4175,N_4112,N_4066);
nor U4176 (N_4176,N_4052,N_4022);
nor U4177 (N_4177,N_4040,N_4089);
nand U4178 (N_4178,N_4008,N_4068);
nor U4179 (N_4179,N_4050,N_4079);
nand U4180 (N_4180,N_4099,N_4055);
and U4181 (N_4181,N_4082,N_4067);
nand U4182 (N_4182,N_4042,N_4000);
and U4183 (N_4183,N_4097,N_4110);
and U4184 (N_4184,N_4106,N_4033);
nor U4185 (N_4185,N_4003,N_4053);
nand U4186 (N_4186,N_4024,N_4018);
or U4187 (N_4187,N_4088,N_4112);
xor U4188 (N_4188,N_4082,N_4091);
nand U4189 (N_4189,N_4062,N_4060);
xnor U4190 (N_4190,N_4108,N_4088);
or U4191 (N_4191,N_4053,N_4074);
nor U4192 (N_4192,N_4094,N_4120);
nand U4193 (N_4193,N_4094,N_4090);
or U4194 (N_4194,N_4003,N_4086);
and U4195 (N_4195,N_4108,N_4122);
xnor U4196 (N_4196,N_4041,N_4091);
nor U4197 (N_4197,N_4063,N_4121);
and U4198 (N_4198,N_4099,N_4053);
nor U4199 (N_4199,N_4120,N_4002);
nand U4200 (N_4200,N_4030,N_4117);
and U4201 (N_4201,N_4004,N_4010);
nor U4202 (N_4202,N_4071,N_4058);
nand U4203 (N_4203,N_4048,N_4066);
nand U4204 (N_4204,N_4105,N_4086);
nand U4205 (N_4205,N_4002,N_4023);
nand U4206 (N_4206,N_4059,N_4083);
xor U4207 (N_4207,N_4053,N_4031);
and U4208 (N_4208,N_4090,N_4088);
nand U4209 (N_4209,N_4086,N_4005);
and U4210 (N_4210,N_4107,N_4086);
and U4211 (N_4211,N_4087,N_4064);
nand U4212 (N_4212,N_4015,N_4036);
and U4213 (N_4213,N_4023,N_4034);
or U4214 (N_4214,N_4067,N_4107);
or U4215 (N_4215,N_4005,N_4124);
or U4216 (N_4216,N_4096,N_4071);
or U4217 (N_4217,N_4078,N_4104);
xnor U4218 (N_4218,N_4115,N_4120);
or U4219 (N_4219,N_4100,N_4076);
or U4220 (N_4220,N_4061,N_4041);
xor U4221 (N_4221,N_4068,N_4011);
and U4222 (N_4222,N_4123,N_4047);
nor U4223 (N_4223,N_4029,N_4089);
and U4224 (N_4224,N_4117,N_4032);
or U4225 (N_4225,N_4061,N_4114);
nor U4226 (N_4226,N_4075,N_4042);
xor U4227 (N_4227,N_4116,N_4093);
nand U4228 (N_4228,N_4079,N_4088);
xor U4229 (N_4229,N_4112,N_4021);
nand U4230 (N_4230,N_4124,N_4002);
xnor U4231 (N_4231,N_4042,N_4106);
xor U4232 (N_4232,N_4052,N_4105);
nand U4233 (N_4233,N_4022,N_4057);
and U4234 (N_4234,N_4030,N_4004);
nand U4235 (N_4235,N_4051,N_4088);
or U4236 (N_4236,N_4079,N_4031);
or U4237 (N_4237,N_4077,N_4009);
or U4238 (N_4238,N_4115,N_4092);
and U4239 (N_4239,N_4011,N_4077);
nor U4240 (N_4240,N_4026,N_4031);
nor U4241 (N_4241,N_4057,N_4012);
or U4242 (N_4242,N_4111,N_4071);
and U4243 (N_4243,N_4063,N_4053);
or U4244 (N_4244,N_4025,N_4076);
or U4245 (N_4245,N_4091,N_4069);
nand U4246 (N_4246,N_4002,N_4081);
and U4247 (N_4247,N_4087,N_4028);
nor U4248 (N_4248,N_4005,N_4087);
nand U4249 (N_4249,N_4103,N_4079);
xnor U4250 (N_4250,N_4175,N_4139);
nand U4251 (N_4251,N_4130,N_4216);
nor U4252 (N_4252,N_4153,N_4164);
or U4253 (N_4253,N_4132,N_4178);
nand U4254 (N_4254,N_4183,N_4241);
nor U4255 (N_4255,N_4235,N_4193);
nor U4256 (N_4256,N_4219,N_4245);
nand U4257 (N_4257,N_4209,N_4232);
nand U4258 (N_4258,N_4190,N_4148);
nor U4259 (N_4259,N_4228,N_4200);
or U4260 (N_4260,N_4156,N_4214);
nand U4261 (N_4261,N_4221,N_4158);
xor U4262 (N_4262,N_4125,N_4237);
nand U4263 (N_4263,N_4233,N_4242);
nand U4264 (N_4264,N_4150,N_4186);
nand U4265 (N_4265,N_4227,N_4247);
xor U4266 (N_4266,N_4191,N_4167);
and U4267 (N_4267,N_4179,N_4220);
nor U4268 (N_4268,N_4218,N_4185);
or U4269 (N_4269,N_4165,N_4163);
or U4270 (N_4270,N_4187,N_4239);
or U4271 (N_4271,N_4238,N_4224);
nor U4272 (N_4272,N_4182,N_4215);
and U4273 (N_4273,N_4181,N_4248);
or U4274 (N_4274,N_4166,N_4230);
or U4275 (N_4275,N_4126,N_4143);
nand U4276 (N_4276,N_4159,N_4160);
nand U4277 (N_4277,N_4134,N_4206);
and U4278 (N_4278,N_4246,N_4203);
nand U4279 (N_4279,N_4210,N_4129);
or U4280 (N_4280,N_4189,N_4229);
and U4281 (N_4281,N_4213,N_4172);
and U4282 (N_4282,N_4205,N_4196);
and U4283 (N_4283,N_4171,N_4127);
nor U4284 (N_4284,N_4202,N_4138);
nand U4285 (N_4285,N_4137,N_4180);
or U4286 (N_4286,N_4152,N_4217);
or U4287 (N_4287,N_4146,N_4194);
nor U4288 (N_4288,N_4195,N_4244);
nor U4289 (N_4289,N_4184,N_4204);
nand U4290 (N_4290,N_4226,N_4149);
xnor U4291 (N_4291,N_4211,N_4198);
and U4292 (N_4292,N_4144,N_4201);
and U4293 (N_4293,N_4225,N_4234);
or U4294 (N_4294,N_4145,N_4157);
or U4295 (N_4295,N_4192,N_4147);
nand U4296 (N_4296,N_4236,N_4222);
nor U4297 (N_4297,N_4131,N_4188);
nand U4298 (N_4298,N_4151,N_4231);
xor U4299 (N_4299,N_4240,N_4249);
and U4300 (N_4300,N_4155,N_4135);
or U4301 (N_4301,N_4162,N_4161);
nand U4302 (N_4302,N_4170,N_4136);
xnor U4303 (N_4303,N_4140,N_4173);
nand U4304 (N_4304,N_4243,N_4141);
xor U4305 (N_4305,N_4174,N_4176);
nor U4306 (N_4306,N_4128,N_4207);
nor U4307 (N_4307,N_4154,N_4168);
nand U4308 (N_4308,N_4169,N_4197);
nor U4309 (N_4309,N_4177,N_4199);
nor U4310 (N_4310,N_4133,N_4223);
nand U4311 (N_4311,N_4142,N_4208);
or U4312 (N_4312,N_4212,N_4185);
and U4313 (N_4313,N_4176,N_4128);
nor U4314 (N_4314,N_4191,N_4143);
or U4315 (N_4315,N_4148,N_4151);
nor U4316 (N_4316,N_4180,N_4201);
and U4317 (N_4317,N_4131,N_4192);
nand U4318 (N_4318,N_4226,N_4139);
nor U4319 (N_4319,N_4227,N_4201);
or U4320 (N_4320,N_4239,N_4161);
nand U4321 (N_4321,N_4128,N_4173);
nand U4322 (N_4322,N_4239,N_4223);
nor U4323 (N_4323,N_4208,N_4186);
and U4324 (N_4324,N_4177,N_4228);
and U4325 (N_4325,N_4183,N_4135);
nor U4326 (N_4326,N_4164,N_4193);
or U4327 (N_4327,N_4222,N_4185);
nand U4328 (N_4328,N_4218,N_4178);
nand U4329 (N_4329,N_4235,N_4166);
and U4330 (N_4330,N_4173,N_4202);
nand U4331 (N_4331,N_4157,N_4189);
xor U4332 (N_4332,N_4134,N_4245);
or U4333 (N_4333,N_4179,N_4217);
nand U4334 (N_4334,N_4194,N_4153);
or U4335 (N_4335,N_4158,N_4244);
and U4336 (N_4336,N_4226,N_4161);
nand U4337 (N_4337,N_4133,N_4178);
xor U4338 (N_4338,N_4247,N_4154);
or U4339 (N_4339,N_4152,N_4188);
xnor U4340 (N_4340,N_4223,N_4226);
or U4341 (N_4341,N_4144,N_4244);
nor U4342 (N_4342,N_4130,N_4214);
nor U4343 (N_4343,N_4195,N_4192);
or U4344 (N_4344,N_4137,N_4217);
or U4345 (N_4345,N_4190,N_4176);
nand U4346 (N_4346,N_4224,N_4189);
or U4347 (N_4347,N_4194,N_4201);
and U4348 (N_4348,N_4132,N_4157);
xor U4349 (N_4349,N_4202,N_4167);
or U4350 (N_4350,N_4205,N_4229);
nor U4351 (N_4351,N_4249,N_4146);
xnor U4352 (N_4352,N_4171,N_4205);
or U4353 (N_4353,N_4197,N_4224);
and U4354 (N_4354,N_4236,N_4213);
or U4355 (N_4355,N_4220,N_4210);
and U4356 (N_4356,N_4129,N_4161);
and U4357 (N_4357,N_4162,N_4184);
xnor U4358 (N_4358,N_4210,N_4228);
nand U4359 (N_4359,N_4161,N_4186);
or U4360 (N_4360,N_4216,N_4241);
nand U4361 (N_4361,N_4153,N_4148);
nor U4362 (N_4362,N_4158,N_4197);
or U4363 (N_4363,N_4153,N_4141);
or U4364 (N_4364,N_4190,N_4151);
nand U4365 (N_4365,N_4234,N_4214);
nor U4366 (N_4366,N_4160,N_4217);
nand U4367 (N_4367,N_4181,N_4204);
nor U4368 (N_4368,N_4248,N_4193);
or U4369 (N_4369,N_4182,N_4209);
nand U4370 (N_4370,N_4215,N_4167);
nand U4371 (N_4371,N_4245,N_4132);
and U4372 (N_4372,N_4176,N_4148);
nor U4373 (N_4373,N_4173,N_4222);
or U4374 (N_4374,N_4247,N_4145);
nand U4375 (N_4375,N_4261,N_4297);
nand U4376 (N_4376,N_4306,N_4257);
and U4377 (N_4377,N_4250,N_4292);
and U4378 (N_4378,N_4328,N_4362);
nor U4379 (N_4379,N_4371,N_4290);
and U4380 (N_4380,N_4293,N_4305);
or U4381 (N_4381,N_4271,N_4255);
and U4382 (N_4382,N_4314,N_4352);
nand U4383 (N_4383,N_4333,N_4368);
and U4384 (N_4384,N_4330,N_4324);
and U4385 (N_4385,N_4321,N_4360);
and U4386 (N_4386,N_4340,N_4253);
nand U4387 (N_4387,N_4345,N_4259);
nand U4388 (N_4388,N_4329,N_4260);
nor U4389 (N_4389,N_4275,N_4318);
and U4390 (N_4390,N_4264,N_4358);
nand U4391 (N_4391,N_4354,N_4254);
and U4392 (N_4392,N_4357,N_4344);
or U4393 (N_4393,N_4336,N_4334);
nor U4394 (N_4394,N_4279,N_4346);
or U4395 (N_4395,N_4313,N_4369);
xnor U4396 (N_4396,N_4288,N_4315);
nand U4397 (N_4397,N_4263,N_4349);
and U4398 (N_4398,N_4301,N_4350);
and U4399 (N_4399,N_4341,N_4326);
and U4400 (N_4400,N_4285,N_4256);
xor U4401 (N_4401,N_4361,N_4342);
or U4402 (N_4402,N_4303,N_4332);
and U4403 (N_4403,N_4356,N_4273);
and U4404 (N_4404,N_4319,N_4278);
nand U4405 (N_4405,N_4309,N_4337);
nand U4406 (N_4406,N_4281,N_4276);
and U4407 (N_4407,N_4373,N_4320);
and U4408 (N_4408,N_4272,N_4353);
or U4409 (N_4409,N_4302,N_4280);
and U4410 (N_4410,N_4258,N_4347);
nand U4411 (N_4411,N_4317,N_4277);
or U4412 (N_4412,N_4283,N_4282);
or U4413 (N_4413,N_4299,N_4323);
and U4414 (N_4414,N_4365,N_4348);
nand U4415 (N_4415,N_4331,N_4372);
nand U4416 (N_4416,N_4251,N_4267);
or U4417 (N_4417,N_4327,N_4300);
or U4418 (N_4418,N_4316,N_4269);
xor U4419 (N_4419,N_4311,N_4307);
xor U4420 (N_4420,N_4265,N_4308);
nor U4421 (N_4421,N_4325,N_4310);
or U4422 (N_4422,N_4363,N_4252);
and U4423 (N_4423,N_4289,N_4268);
nand U4424 (N_4424,N_4351,N_4284);
or U4425 (N_4425,N_4359,N_4298);
xnor U4426 (N_4426,N_4262,N_4335);
or U4427 (N_4427,N_4274,N_4370);
nor U4428 (N_4428,N_4312,N_4291);
nand U4429 (N_4429,N_4266,N_4286);
or U4430 (N_4430,N_4304,N_4364);
nand U4431 (N_4431,N_4270,N_4366);
nand U4432 (N_4432,N_4343,N_4294);
nand U4433 (N_4433,N_4287,N_4322);
or U4434 (N_4434,N_4296,N_4374);
xor U4435 (N_4435,N_4338,N_4355);
and U4436 (N_4436,N_4367,N_4339);
and U4437 (N_4437,N_4295,N_4319);
and U4438 (N_4438,N_4321,N_4349);
and U4439 (N_4439,N_4369,N_4344);
or U4440 (N_4440,N_4358,N_4281);
or U4441 (N_4441,N_4341,N_4298);
and U4442 (N_4442,N_4332,N_4308);
or U4443 (N_4443,N_4269,N_4274);
nand U4444 (N_4444,N_4374,N_4281);
nand U4445 (N_4445,N_4364,N_4328);
nor U4446 (N_4446,N_4314,N_4299);
nor U4447 (N_4447,N_4321,N_4295);
nand U4448 (N_4448,N_4293,N_4295);
nor U4449 (N_4449,N_4267,N_4371);
and U4450 (N_4450,N_4286,N_4305);
nand U4451 (N_4451,N_4302,N_4314);
and U4452 (N_4452,N_4349,N_4283);
and U4453 (N_4453,N_4328,N_4359);
nand U4454 (N_4454,N_4303,N_4322);
nand U4455 (N_4455,N_4356,N_4271);
xor U4456 (N_4456,N_4318,N_4277);
nand U4457 (N_4457,N_4271,N_4280);
and U4458 (N_4458,N_4275,N_4281);
nor U4459 (N_4459,N_4268,N_4364);
or U4460 (N_4460,N_4373,N_4324);
or U4461 (N_4461,N_4367,N_4307);
and U4462 (N_4462,N_4260,N_4318);
or U4463 (N_4463,N_4302,N_4313);
and U4464 (N_4464,N_4369,N_4304);
nor U4465 (N_4465,N_4251,N_4287);
nand U4466 (N_4466,N_4337,N_4304);
nor U4467 (N_4467,N_4277,N_4364);
and U4468 (N_4468,N_4351,N_4361);
or U4469 (N_4469,N_4304,N_4321);
or U4470 (N_4470,N_4302,N_4284);
nand U4471 (N_4471,N_4326,N_4365);
or U4472 (N_4472,N_4297,N_4253);
or U4473 (N_4473,N_4327,N_4305);
nand U4474 (N_4474,N_4339,N_4274);
and U4475 (N_4475,N_4371,N_4348);
and U4476 (N_4476,N_4272,N_4265);
nand U4477 (N_4477,N_4296,N_4266);
nand U4478 (N_4478,N_4269,N_4294);
nor U4479 (N_4479,N_4352,N_4284);
and U4480 (N_4480,N_4336,N_4271);
or U4481 (N_4481,N_4299,N_4311);
nor U4482 (N_4482,N_4293,N_4351);
xor U4483 (N_4483,N_4306,N_4355);
nor U4484 (N_4484,N_4328,N_4257);
nand U4485 (N_4485,N_4313,N_4250);
nand U4486 (N_4486,N_4319,N_4296);
nor U4487 (N_4487,N_4352,N_4325);
and U4488 (N_4488,N_4366,N_4285);
xnor U4489 (N_4489,N_4296,N_4279);
and U4490 (N_4490,N_4356,N_4267);
xnor U4491 (N_4491,N_4312,N_4351);
nand U4492 (N_4492,N_4320,N_4370);
nand U4493 (N_4493,N_4286,N_4363);
nor U4494 (N_4494,N_4360,N_4351);
xor U4495 (N_4495,N_4348,N_4291);
and U4496 (N_4496,N_4334,N_4320);
and U4497 (N_4497,N_4303,N_4335);
nand U4498 (N_4498,N_4368,N_4250);
nor U4499 (N_4499,N_4300,N_4291);
and U4500 (N_4500,N_4465,N_4410);
and U4501 (N_4501,N_4478,N_4420);
or U4502 (N_4502,N_4393,N_4424);
or U4503 (N_4503,N_4455,N_4436);
xnor U4504 (N_4504,N_4386,N_4390);
nor U4505 (N_4505,N_4388,N_4461);
or U4506 (N_4506,N_4376,N_4498);
and U4507 (N_4507,N_4454,N_4432);
nand U4508 (N_4508,N_4458,N_4391);
nor U4509 (N_4509,N_4496,N_4417);
or U4510 (N_4510,N_4405,N_4398);
and U4511 (N_4511,N_4443,N_4479);
or U4512 (N_4512,N_4385,N_4456);
nand U4513 (N_4513,N_4382,N_4430);
and U4514 (N_4514,N_4468,N_4414);
nor U4515 (N_4515,N_4445,N_4435);
and U4516 (N_4516,N_4467,N_4439);
nor U4517 (N_4517,N_4378,N_4448);
and U4518 (N_4518,N_4471,N_4440);
and U4519 (N_4519,N_4476,N_4481);
nor U4520 (N_4520,N_4380,N_4375);
xor U4521 (N_4521,N_4404,N_4377);
nand U4522 (N_4522,N_4412,N_4387);
nand U4523 (N_4523,N_4480,N_4434);
nor U4524 (N_4524,N_4475,N_4482);
nand U4525 (N_4525,N_4407,N_4403);
nor U4526 (N_4526,N_4499,N_4409);
xor U4527 (N_4527,N_4459,N_4497);
and U4528 (N_4528,N_4416,N_4460);
or U4529 (N_4529,N_4477,N_4484);
nand U4530 (N_4530,N_4441,N_4428);
nor U4531 (N_4531,N_4450,N_4495);
nor U4532 (N_4532,N_4457,N_4463);
and U4533 (N_4533,N_4395,N_4383);
nor U4534 (N_4534,N_4408,N_4485);
nand U4535 (N_4535,N_4494,N_4464);
and U4536 (N_4536,N_4397,N_4470);
xnor U4537 (N_4537,N_4406,N_4486);
and U4538 (N_4538,N_4426,N_4490);
and U4539 (N_4539,N_4399,N_4444);
nor U4540 (N_4540,N_4472,N_4453);
nand U4541 (N_4541,N_4401,N_4400);
and U4542 (N_4542,N_4449,N_4469);
or U4543 (N_4543,N_4493,N_4452);
nor U4544 (N_4544,N_4462,N_4433);
or U4545 (N_4545,N_4402,N_4489);
xor U4546 (N_4546,N_4413,N_4423);
and U4547 (N_4547,N_4442,N_4415);
nor U4548 (N_4548,N_4431,N_4381);
and U4549 (N_4549,N_4483,N_4425);
nor U4550 (N_4550,N_4488,N_4418);
nor U4551 (N_4551,N_4411,N_4487);
nand U4552 (N_4552,N_4447,N_4492);
nor U4553 (N_4553,N_4451,N_4392);
or U4554 (N_4554,N_4427,N_4396);
or U4555 (N_4555,N_4474,N_4466);
and U4556 (N_4556,N_4473,N_4429);
and U4557 (N_4557,N_4422,N_4437);
and U4558 (N_4558,N_4394,N_4379);
nand U4559 (N_4559,N_4446,N_4384);
nand U4560 (N_4560,N_4438,N_4421);
and U4561 (N_4561,N_4419,N_4389);
nor U4562 (N_4562,N_4491,N_4421);
xnor U4563 (N_4563,N_4414,N_4454);
nor U4564 (N_4564,N_4444,N_4404);
nand U4565 (N_4565,N_4484,N_4491);
and U4566 (N_4566,N_4431,N_4401);
nand U4567 (N_4567,N_4461,N_4484);
nor U4568 (N_4568,N_4392,N_4390);
nor U4569 (N_4569,N_4390,N_4499);
nand U4570 (N_4570,N_4429,N_4404);
nor U4571 (N_4571,N_4388,N_4419);
and U4572 (N_4572,N_4379,N_4433);
and U4573 (N_4573,N_4441,N_4476);
nor U4574 (N_4574,N_4394,N_4498);
nor U4575 (N_4575,N_4376,N_4403);
xnor U4576 (N_4576,N_4425,N_4495);
nor U4577 (N_4577,N_4429,N_4427);
nand U4578 (N_4578,N_4492,N_4457);
nand U4579 (N_4579,N_4400,N_4453);
and U4580 (N_4580,N_4401,N_4481);
and U4581 (N_4581,N_4380,N_4391);
or U4582 (N_4582,N_4396,N_4474);
nor U4583 (N_4583,N_4462,N_4451);
and U4584 (N_4584,N_4413,N_4394);
and U4585 (N_4585,N_4425,N_4445);
nor U4586 (N_4586,N_4436,N_4396);
or U4587 (N_4587,N_4405,N_4467);
nor U4588 (N_4588,N_4384,N_4418);
and U4589 (N_4589,N_4488,N_4382);
nor U4590 (N_4590,N_4413,N_4481);
or U4591 (N_4591,N_4389,N_4451);
or U4592 (N_4592,N_4422,N_4391);
and U4593 (N_4593,N_4485,N_4452);
or U4594 (N_4594,N_4423,N_4447);
and U4595 (N_4595,N_4394,N_4438);
and U4596 (N_4596,N_4465,N_4415);
nor U4597 (N_4597,N_4387,N_4466);
and U4598 (N_4598,N_4404,N_4406);
nand U4599 (N_4599,N_4448,N_4450);
or U4600 (N_4600,N_4461,N_4407);
nand U4601 (N_4601,N_4497,N_4425);
nor U4602 (N_4602,N_4402,N_4422);
nand U4603 (N_4603,N_4381,N_4419);
or U4604 (N_4604,N_4433,N_4434);
nor U4605 (N_4605,N_4404,N_4437);
xnor U4606 (N_4606,N_4480,N_4403);
nor U4607 (N_4607,N_4406,N_4386);
or U4608 (N_4608,N_4418,N_4431);
xor U4609 (N_4609,N_4485,N_4424);
nand U4610 (N_4610,N_4399,N_4486);
and U4611 (N_4611,N_4464,N_4381);
xor U4612 (N_4612,N_4442,N_4406);
nor U4613 (N_4613,N_4409,N_4394);
nor U4614 (N_4614,N_4388,N_4440);
and U4615 (N_4615,N_4465,N_4489);
and U4616 (N_4616,N_4498,N_4438);
and U4617 (N_4617,N_4421,N_4437);
nand U4618 (N_4618,N_4407,N_4416);
or U4619 (N_4619,N_4496,N_4412);
nor U4620 (N_4620,N_4495,N_4397);
nand U4621 (N_4621,N_4401,N_4428);
nor U4622 (N_4622,N_4464,N_4440);
nand U4623 (N_4623,N_4463,N_4385);
nor U4624 (N_4624,N_4410,N_4426);
nor U4625 (N_4625,N_4587,N_4533);
and U4626 (N_4626,N_4513,N_4554);
xor U4627 (N_4627,N_4519,N_4598);
or U4628 (N_4628,N_4521,N_4616);
nand U4629 (N_4629,N_4534,N_4508);
or U4630 (N_4630,N_4584,N_4602);
and U4631 (N_4631,N_4609,N_4503);
and U4632 (N_4632,N_4590,N_4504);
and U4633 (N_4633,N_4564,N_4618);
xnor U4634 (N_4634,N_4559,N_4550);
nor U4635 (N_4635,N_4577,N_4520);
nand U4636 (N_4636,N_4505,N_4542);
nand U4637 (N_4637,N_4583,N_4604);
nand U4638 (N_4638,N_4573,N_4622);
xnor U4639 (N_4639,N_4506,N_4558);
or U4640 (N_4640,N_4599,N_4620);
and U4641 (N_4641,N_4605,N_4525);
and U4642 (N_4642,N_4565,N_4549);
nand U4643 (N_4643,N_4546,N_4545);
nand U4644 (N_4644,N_4619,N_4518);
and U4645 (N_4645,N_4501,N_4517);
and U4646 (N_4646,N_4553,N_4510);
and U4647 (N_4647,N_4527,N_4566);
nand U4648 (N_4648,N_4529,N_4552);
nor U4649 (N_4649,N_4582,N_4588);
nand U4650 (N_4650,N_4547,N_4574);
nand U4651 (N_4651,N_4624,N_4594);
or U4652 (N_4652,N_4614,N_4569);
and U4653 (N_4653,N_4536,N_4611);
or U4654 (N_4654,N_4580,N_4543);
or U4655 (N_4655,N_4591,N_4528);
or U4656 (N_4656,N_4537,N_4524);
nor U4657 (N_4657,N_4555,N_4568);
nor U4658 (N_4658,N_4586,N_4601);
nand U4659 (N_4659,N_4567,N_4617);
or U4660 (N_4660,N_4606,N_4509);
nor U4661 (N_4661,N_4562,N_4576);
nor U4662 (N_4662,N_4532,N_4538);
nand U4663 (N_4663,N_4593,N_4578);
and U4664 (N_4664,N_4603,N_4544);
nand U4665 (N_4665,N_4522,N_4548);
or U4666 (N_4666,N_4600,N_4539);
or U4667 (N_4667,N_4551,N_4612);
nand U4668 (N_4668,N_4613,N_4608);
nand U4669 (N_4669,N_4563,N_4557);
nor U4670 (N_4670,N_4597,N_4596);
nand U4671 (N_4671,N_4526,N_4531);
xnor U4672 (N_4672,N_4589,N_4585);
nor U4673 (N_4673,N_4579,N_4570);
or U4674 (N_4674,N_4592,N_4621);
or U4675 (N_4675,N_4500,N_4610);
or U4676 (N_4676,N_4541,N_4623);
nand U4677 (N_4677,N_4511,N_4516);
nand U4678 (N_4678,N_4571,N_4561);
nand U4679 (N_4679,N_4535,N_4514);
xor U4680 (N_4680,N_4581,N_4540);
nor U4681 (N_4681,N_4607,N_4515);
and U4682 (N_4682,N_4512,N_4530);
nor U4683 (N_4683,N_4560,N_4595);
and U4684 (N_4684,N_4615,N_4556);
or U4685 (N_4685,N_4507,N_4502);
or U4686 (N_4686,N_4523,N_4575);
nor U4687 (N_4687,N_4572,N_4504);
and U4688 (N_4688,N_4560,N_4544);
and U4689 (N_4689,N_4596,N_4577);
xor U4690 (N_4690,N_4535,N_4608);
and U4691 (N_4691,N_4573,N_4550);
or U4692 (N_4692,N_4601,N_4551);
xor U4693 (N_4693,N_4596,N_4589);
xor U4694 (N_4694,N_4619,N_4550);
nor U4695 (N_4695,N_4525,N_4551);
and U4696 (N_4696,N_4606,N_4588);
nand U4697 (N_4697,N_4522,N_4509);
nand U4698 (N_4698,N_4570,N_4521);
nor U4699 (N_4699,N_4501,N_4566);
or U4700 (N_4700,N_4620,N_4581);
nand U4701 (N_4701,N_4574,N_4500);
nor U4702 (N_4702,N_4573,N_4537);
nand U4703 (N_4703,N_4620,N_4502);
and U4704 (N_4704,N_4593,N_4610);
nor U4705 (N_4705,N_4582,N_4512);
nand U4706 (N_4706,N_4609,N_4541);
nor U4707 (N_4707,N_4509,N_4540);
xor U4708 (N_4708,N_4575,N_4610);
and U4709 (N_4709,N_4588,N_4615);
or U4710 (N_4710,N_4519,N_4615);
nand U4711 (N_4711,N_4581,N_4590);
or U4712 (N_4712,N_4531,N_4587);
nor U4713 (N_4713,N_4501,N_4616);
and U4714 (N_4714,N_4520,N_4504);
nand U4715 (N_4715,N_4579,N_4564);
and U4716 (N_4716,N_4614,N_4563);
nand U4717 (N_4717,N_4567,N_4534);
and U4718 (N_4718,N_4548,N_4534);
nand U4719 (N_4719,N_4536,N_4572);
nand U4720 (N_4720,N_4609,N_4624);
nand U4721 (N_4721,N_4529,N_4576);
nor U4722 (N_4722,N_4581,N_4615);
nor U4723 (N_4723,N_4612,N_4565);
nor U4724 (N_4724,N_4594,N_4590);
nor U4725 (N_4725,N_4589,N_4567);
and U4726 (N_4726,N_4537,N_4575);
xor U4727 (N_4727,N_4521,N_4522);
and U4728 (N_4728,N_4587,N_4548);
and U4729 (N_4729,N_4537,N_4578);
or U4730 (N_4730,N_4596,N_4513);
nand U4731 (N_4731,N_4528,N_4504);
nor U4732 (N_4732,N_4585,N_4525);
or U4733 (N_4733,N_4556,N_4605);
nand U4734 (N_4734,N_4580,N_4579);
or U4735 (N_4735,N_4606,N_4583);
nor U4736 (N_4736,N_4534,N_4509);
nor U4737 (N_4737,N_4554,N_4603);
and U4738 (N_4738,N_4504,N_4609);
and U4739 (N_4739,N_4582,N_4577);
nand U4740 (N_4740,N_4601,N_4584);
and U4741 (N_4741,N_4516,N_4619);
nor U4742 (N_4742,N_4584,N_4505);
nand U4743 (N_4743,N_4602,N_4581);
or U4744 (N_4744,N_4577,N_4521);
nor U4745 (N_4745,N_4605,N_4619);
nor U4746 (N_4746,N_4583,N_4581);
and U4747 (N_4747,N_4536,N_4554);
or U4748 (N_4748,N_4545,N_4566);
nand U4749 (N_4749,N_4589,N_4607);
nor U4750 (N_4750,N_4739,N_4720);
nand U4751 (N_4751,N_4729,N_4717);
nor U4752 (N_4752,N_4730,N_4684);
nand U4753 (N_4753,N_4702,N_4681);
nand U4754 (N_4754,N_4663,N_4643);
nor U4755 (N_4755,N_4733,N_4649);
and U4756 (N_4756,N_4642,N_4716);
and U4757 (N_4757,N_4705,N_4634);
nor U4758 (N_4758,N_4698,N_4660);
nor U4759 (N_4759,N_4695,N_4689);
or U4760 (N_4760,N_4719,N_4671);
or U4761 (N_4761,N_4683,N_4688);
xnor U4762 (N_4762,N_4722,N_4654);
nor U4763 (N_4763,N_4647,N_4666);
or U4764 (N_4764,N_4636,N_4632);
and U4765 (N_4765,N_4718,N_4707);
nor U4766 (N_4766,N_4667,N_4646);
and U4767 (N_4767,N_4664,N_4686);
xor U4768 (N_4768,N_4665,N_4712);
and U4769 (N_4769,N_4697,N_4670);
or U4770 (N_4770,N_4744,N_4680);
or U4771 (N_4771,N_4742,N_4672);
and U4772 (N_4772,N_4737,N_4655);
and U4773 (N_4773,N_4690,N_4662);
and U4774 (N_4774,N_4678,N_4669);
xnor U4775 (N_4775,N_4627,N_4725);
and U4776 (N_4776,N_4743,N_4644);
and U4777 (N_4777,N_4738,N_4652);
or U4778 (N_4778,N_4641,N_4731);
nand U4779 (N_4779,N_4682,N_4701);
nor U4780 (N_4780,N_4704,N_4630);
nor U4781 (N_4781,N_4661,N_4715);
or U4782 (N_4782,N_4721,N_4714);
nor U4783 (N_4783,N_4653,N_4656);
nor U4784 (N_4784,N_4639,N_4710);
and U4785 (N_4785,N_4635,N_4659);
nor U4786 (N_4786,N_4638,N_4708);
or U4787 (N_4787,N_4727,N_4650);
or U4788 (N_4788,N_4749,N_4703);
nand U4789 (N_4789,N_4696,N_4676);
nor U4790 (N_4790,N_4694,N_4626);
or U4791 (N_4791,N_4746,N_4631);
and U4792 (N_4792,N_4693,N_4658);
and U4793 (N_4793,N_4673,N_4726);
nand U4794 (N_4794,N_4711,N_4625);
nor U4795 (N_4795,N_4657,N_4637);
nand U4796 (N_4796,N_4651,N_4723);
nand U4797 (N_4797,N_4629,N_4741);
xnor U4798 (N_4798,N_4674,N_4628);
xor U4799 (N_4799,N_4685,N_4706);
and U4800 (N_4800,N_4724,N_4709);
nand U4801 (N_4801,N_4735,N_4745);
nor U4802 (N_4802,N_4640,N_4692);
and U4803 (N_4803,N_4679,N_4700);
or U4804 (N_4804,N_4648,N_4740);
and U4805 (N_4805,N_4713,N_4747);
and U4806 (N_4806,N_4734,N_4691);
xnor U4807 (N_4807,N_4748,N_4633);
nand U4808 (N_4808,N_4675,N_4728);
nand U4809 (N_4809,N_4699,N_4687);
nand U4810 (N_4810,N_4736,N_4645);
or U4811 (N_4811,N_4677,N_4668);
xor U4812 (N_4812,N_4732,N_4687);
nor U4813 (N_4813,N_4663,N_4700);
nand U4814 (N_4814,N_4726,N_4748);
or U4815 (N_4815,N_4713,N_4629);
or U4816 (N_4816,N_4743,N_4647);
or U4817 (N_4817,N_4731,N_4721);
nor U4818 (N_4818,N_4661,N_4659);
nand U4819 (N_4819,N_4636,N_4726);
nand U4820 (N_4820,N_4705,N_4676);
nand U4821 (N_4821,N_4633,N_4737);
nor U4822 (N_4822,N_4692,N_4735);
nand U4823 (N_4823,N_4681,N_4725);
and U4824 (N_4824,N_4650,N_4633);
and U4825 (N_4825,N_4744,N_4691);
nand U4826 (N_4826,N_4725,N_4709);
and U4827 (N_4827,N_4670,N_4688);
and U4828 (N_4828,N_4724,N_4672);
xor U4829 (N_4829,N_4686,N_4667);
or U4830 (N_4830,N_4742,N_4646);
nand U4831 (N_4831,N_4652,N_4671);
or U4832 (N_4832,N_4687,N_4711);
nand U4833 (N_4833,N_4708,N_4664);
or U4834 (N_4834,N_4671,N_4708);
nand U4835 (N_4835,N_4697,N_4737);
and U4836 (N_4836,N_4708,N_4716);
xor U4837 (N_4837,N_4653,N_4665);
xnor U4838 (N_4838,N_4747,N_4660);
or U4839 (N_4839,N_4699,N_4636);
and U4840 (N_4840,N_4632,N_4693);
or U4841 (N_4841,N_4644,N_4627);
or U4842 (N_4842,N_4715,N_4698);
or U4843 (N_4843,N_4681,N_4671);
and U4844 (N_4844,N_4655,N_4673);
xor U4845 (N_4845,N_4637,N_4726);
nor U4846 (N_4846,N_4654,N_4716);
or U4847 (N_4847,N_4685,N_4724);
or U4848 (N_4848,N_4626,N_4724);
nand U4849 (N_4849,N_4638,N_4641);
nand U4850 (N_4850,N_4674,N_4741);
xor U4851 (N_4851,N_4715,N_4677);
or U4852 (N_4852,N_4731,N_4704);
and U4853 (N_4853,N_4675,N_4633);
xnor U4854 (N_4854,N_4713,N_4702);
nand U4855 (N_4855,N_4678,N_4692);
nor U4856 (N_4856,N_4714,N_4707);
and U4857 (N_4857,N_4739,N_4713);
and U4858 (N_4858,N_4709,N_4634);
and U4859 (N_4859,N_4705,N_4650);
or U4860 (N_4860,N_4653,N_4724);
nor U4861 (N_4861,N_4722,N_4661);
or U4862 (N_4862,N_4649,N_4701);
nand U4863 (N_4863,N_4732,N_4733);
or U4864 (N_4864,N_4673,N_4682);
nor U4865 (N_4865,N_4629,N_4717);
nand U4866 (N_4866,N_4675,N_4662);
or U4867 (N_4867,N_4629,N_4682);
or U4868 (N_4868,N_4653,N_4707);
nand U4869 (N_4869,N_4646,N_4700);
nand U4870 (N_4870,N_4656,N_4673);
nand U4871 (N_4871,N_4689,N_4665);
xor U4872 (N_4872,N_4697,N_4638);
nand U4873 (N_4873,N_4703,N_4723);
nand U4874 (N_4874,N_4741,N_4716);
or U4875 (N_4875,N_4790,N_4783);
or U4876 (N_4876,N_4811,N_4755);
nand U4877 (N_4877,N_4841,N_4864);
or U4878 (N_4878,N_4847,N_4795);
xor U4879 (N_4879,N_4823,N_4861);
or U4880 (N_4880,N_4836,N_4829);
nand U4881 (N_4881,N_4813,N_4846);
or U4882 (N_4882,N_4810,N_4768);
nor U4883 (N_4883,N_4854,N_4817);
nand U4884 (N_4884,N_4848,N_4796);
or U4885 (N_4885,N_4862,N_4759);
nand U4886 (N_4886,N_4870,N_4771);
or U4887 (N_4887,N_4797,N_4816);
or U4888 (N_4888,N_4814,N_4758);
and U4889 (N_4889,N_4837,N_4868);
and U4890 (N_4890,N_4850,N_4859);
or U4891 (N_4891,N_4774,N_4799);
and U4892 (N_4892,N_4853,N_4821);
xnor U4893 (N_4893,N_4826,N_4764);
or U4894 (N_4894,N_4793,N_4751);
or U4895 (N_4895,N_4802,N_4833);
nand U4896 (N_4896,N_4824,N_4867);
nand U4897 (N_4897,N_4825,N_4831);
and U4898 (N_4898,N_4851,N_4762);
and U4899 (N_4899,N_4789,N_4843);
xnor U4900 (N_4900,N_4820,N_4781);
nand U4901 (N_4901,N_4858,N_4775);
or U4902 (N_4902,N_4780,N_4777);
xnor U4903 (N_4903,N_4852,N_4812);
nor U4904 (N_4904,N_4808,N_4828);
and U4905 (N_4905,N_4807,N_4869);
or U4906 (N_4906,N_4779,N_4769);
and U4907 (N_4907,N_4873,N_4801);
nand U4908 (N_4908,N_4806,N_4798);
nand U4909 (N_4909,N_4757,N_4863);
nor U4910 (N_4910,N_4849,N_4756);
or U4911 (N_4911,N_4760,N_4815);
xor U4912 (N_4912,N_4805,N_4822);
nor U4913 (N_4913,N_4844,N_4840);
nor U4914 (N_4914,N_4784,N_4763);
or U4915 (N_4915,N_4818,N_4832);
or U4916 (N_4916,N_4871,N_4872);
and U4917 (N_4917,N_4804,N_4830);
xnor U4918 (N_4918,N_4800,N_4835);
or U4919 (N_4919,N_4791,N_4786);
nand U4920 (N_4920,N_4856,N_4865);
nand U4921 (N_4921,N_4839,N_4838);
and U4922 (N_4922,N_4809,N_4794);
nor U4923 (N_4923,N_4788,N_4787);
nor U4924 (N_4924,N_4866,N_4766);
nand U4925 (N_4925,N_4767,N_4857);
nand U4926 (N_4926,N_4842,N_4752);
nand U4927 (N_4927,N_4765,N_4754);
nand U4928 (N_4928,N_4874,N_4761);
nand U4929 (N_4929,N_4803,N_4770);
nor U4930 (N_4930,N_4792,N_4834);
xor U4931 (N_4931,N_4845,N_4827);
xnor U4932 (N_4932,N_4855,N_4772);
nor U4933 (N_4933,N_4782,N_4860);
xnor U4934 (N_4934,N_4785,N_4753);
nand U4935 (N_4935,N_4819,N_4776);
or U4936 (N_4936,N_4750,N_4778);
nor U4937 (N_4937,N_4773,N_4838);
or U4938 (N_4938,N_4797,N_4827);
or U4939 (N_4939,N_4847,N_4821);
nand U4940 (N_4940,N_4864,N_4865);
or U4941 (N_4941,N_4828,N_4827);
or U4942 (N_4942,N_4759,N_4860);
or U4943 (N_4943,N_4850,N_4818);
and U4944 (N_4944,N_4810,N_4842);
nor U4945 (N_4945,N_4801,N_4836);
nor U4946 (N_4946,N_4840,N_4851);
nand U4947 (N_4947,N_4788,N_4793);
nand U4948 (N_4948,N_4787,N_4784);
nor U4949 (N_4949,N_4822,N_4819);
and U4950 (N_4950,N_4859,N_4866);
nand U4951 (N_4951,N_4773,N_4750);
and U4952 (N_4952,N_4762,N_4810);
nand U4953 (N_4953,N_4841,N_4852);
nor U4954 (N_4954,N_4795,N_4859);
xnor U4955 (N_4955,N_4859,N_4772);
nand U4956 (N_4956,N_4792,N_4791);
nor U4957 (N_4957,N_4765,N_4771);
or U4958 (N_4958,N_4831,N_4819);
or U4959 (N_4959,N_4846,N_4818);
or U4960 (N_4960,N_4870,N_4786);
nor U4961 (N_4961,N_4831,N_4858);
and U4962 (N_4962,N_4808,N_4804);
and U4963 (N_4963,N_4783,N_4810);
and U4964 (N_4964,N_4873,N_4799);
or U4965 (N_4965,N_4793,N_4853);
or U4966 (N_4966,N_4862,N_4772);
or U4967 (N_4967,N_4834,N_4789);
and U4968 (N_4968,N_4802,N_4777);
nor U4969 (N_4969,N_4847,N_4854);
xor U4970 (N_4970,N_4851,N_4873);
nand U4971 (N_4971,N_4826,N_4871);
or U4972 (N_4972,N_4816,N_4785);
and U4973 (N_4973,N_4871,N_4777);
and U4974 (N_4974,N_4842,N_4789);
nand U4975 (N_4975,N_4778,N_4801);
nor U4976 (N_4976,N_4795,N_4786);
nand U4977 (N_4977,N_4839,N_4837);
or U4978 (N_4978,N_4774,N_4838);
and U4979 (N_4979,N_4821,N_4779);
and U4980 (N_4980,N_4817,N_4847);
nor U4981 (N_4981,N_4819,N_4791);
and U4982 (N_4982,N_4768,N_4773);
xnor U4983 (N_4983,N_4845,N_4852);
nand U4984 (N_4984,N_4825,N_4762);
and U4985 (N_4985,N_4860,N_4825);
nor U4986 (N_4986,N_4825,N_4846);
and U4987 (N_4987,N_4833,N_4821);
nor U4988 (N_4988,N_4813,N_4834);
nand U4989 (N_4989,N_4768,N_4843);
nand U4990 (N_4990,N_4867,N_4768);
nor U4991 (N_4991,N_4811,N_4791);
xnor U4992 (N_4992,N_4839,N_4802);
and U4993 (N_4993,N_4827,N_4772);
and U4994 (N_4994,N_4781,N_4841);
or U4995 (N_4995,N_4859,N_4793);
and U4996 (N_4996,N_4750,N_4821);
nor U4997 (N_4997,N_4869,N_4797);
and U4998 (N_4998,N_4840,N_4873);
xor U4999 (N_4999,N_4766,N_4851);
and U5000 (N_5000,N_4999,N_4899);
xnor U5001 (N_5001,N_4916,N_4992);
and U5002 (N_5002,N_4997,N_4971);
nand U5003 (N_5003,N_4988,N_4982);
and U5004 (N_5004,N_4880,N_4879);
and U5005 (N_5005,N_4934,N_4976);
and U5006 (N_5006,N_4968,N_4894);
and U5007 (N_5007,N_4906,N_4957);
nor U5008 (N_5008,N_4943,N_4994);
nand U5009 (N_5009,N_4978,N_4983);
and U5010 (N_5010,N_4949,N_4965);
or U5011 (N_5011,N_4958,N_4951);
nor U5012 (N_5012,N_4977,N_4941);
or U5013 (N_5013,N_4887,N_4919);
xor U5014 (N_5014,N_4929,N_4904);
and U5015 (N_5015,N_4956,N_4960);
nor U5016 (N_5016,N_4938,N_4884);
or U5017 (N_5017,N_4927,N_4970);
nor U5018 (N_5018,N_4913,N_4989);
and U5019 (N_5019,N_4930,N_4935);
and U5020 (N_5020,N_4907,N_4963);
nor U5021 (N_5021,N_4921,N_4952);
and U5022 (N_5022,N_4897,N_4890);
and U5023 (N_5023,N_4990,N_4950);
nor U5024 (N_5024,N_4966,N_4928);
xor U5025 (N_5025,N_4893,N_4912);
and U5026 (N_5026,N_4953,N_4910);
or U5027 (N_5027,N_4892,N_4917);
nor U5028 (N_5028,N_4998,N_4918);
or U5029 (N_5029,N_4885,N_4939);
nand U5030 (N_5030,N_4974,N_4962);
xnor U5031 (N_5031,N_4946,N_4947);
nand U5032 (N_5032,N_4981,N_4920);
nor U5033 (N_5033,N_4984,N_4905);
nand U5034 (N_5034,N_4967,N_4979);
or U5035 (N_5035,N_4902,N_4944);
nand U5036 (N_5036,N_4915,N_4955);
xor U5037 (N_5037,N_4908,N_4940);
and U5038 (N_5038,N_4931,N_4903);
or U5039 (N_5039,N_4896,N_4895);
and U5040 (N_5040,N_4985,N_4942);
or U5041 (N_5041,N_4877,N_4922);
and U5042 (N_5042,N_4986,N_4993);
nor U5043 (N_5043,N_4964,N_4898);
and U5044 (N_5044,N_4980,N_4991);
xnor U5045 (N_5045,N_4945,N_4932);
nand U5046 (N_5046,N_4936,N_4973);
nand U5047 (N_5047,N_4924,N_4948);
or U5048 (N_5048,N_4889,N_4914);
or U5049 (N_5049,N_4901,N_4875);
nand U5050 (N_5050,N_4996,N_4883);
and U5051 (N_5051,N_4911,N_4926);
nor U5052 (N_5052,N_4923,N_4975);
nor U5053 (N_5053,N_4987,N_4886);
nor U5054 (N_5054,N_4878,N_4995);
or U5055 (N_5055,N_4881,N_4972);
or U5056 (N_5056,N_4876,N_4933);
nand U5057 (N_5057,N_4937,N_4900);
or U5058 (N_5058,N_4954,N_4888);
nand U5059 (N_5059,N_4891,N_4909);
and U5060 (N_5060,N_4959,N_4882);
xor U5061 (N_5061,N_4969,N_4925);
nor U5062 (N_5062,N_4961,N_4904);
xor U5063 (N_5063,N_4918,N_4965);
nand U5064 (N_5064,N_4966,N_4890);
nor U5065 (N_5065,N_4875,N_4967);
and U5066 (N_5066,N_4956,N_4922);
or U5067 (N_5067,N_4965,N_4881);
or U5068 (N_5068,N_4892,N_4976);
xor U5069 (N_5069,N_4978,N_4892);
nor U5070 (N_5070,N_4994,N_4892);
and U5071 (N_5071,N_4941,N_4950);
nor U5072 (N_5072,N_4986,N_4955);
xnor U5073 (N_5073,N_4978,N_4882);
nor U5074 (N_5074,N_4880,N_4970);
nand U5075 (N_5075,N_4930,N_4965);
xor U5076 (N_5076,N_4888,N_4988);
nand U5077 (N_5077,N_4919,N_4958);
or U5078 (N_5078,N_4878,N_4935);
nor U5079 (N_5079,N_4927,N_4981);
nor U5080 (N_5080,N_4928,N_4905);
xor U5081 (N_5081,N_4909,N_4926);
and U5082 (N_5082,N_4926,N_4972);
nand U5083 (N_5083,N_4936,N_4932);
and U5084 (N_5084,N_4877,N_4934);
and U5085 (N_5085,N_4925,N_4941);
nand U5086 (N_5086,N_4962,N_4920);
and U5087 (N_5087,N_4911,N_4971);
xor U5088 (N_5088,N_4959,N_4932);
or U5089 (N_5089,N_4912,N_4886);
nor U5090 (N_5090,N_4951,N_4979);
xor U5091 (N_5091,N_4933,N_4927);
nand U5092 (N_5092,N_4962,N_4894);
nor U5093 (N_5093,N_4903,N_4975);
xnor U5094 (N_5094,N_4914,N_4999);
nand U5095 (N_5095,N_4899,N_4931);
or U5096 (N_5096,N_4982,N_4899);
nor U5097 (N_5097,N_4890,N_4937);
nor U5098 (N_5098,N_4886,N_4879);
nor U5099 (N_5099,N_4935,N_4895);
nor U5100 (N_5100,N_4888,N_4920);
xor U5101 (N_5101,N_4884,N_4887);
nand U5102 (N_5102,N_4910,N_4952);
nand U5103 (N_5103,N_4912,N_4946);
nor U5104 (N_5104,N_4976,N_4946);
nand U5105 (N_5105,N_4899,N_4955);
or U5106 (N_5106,N_4997,N_4886);
nor U5107 (N_5107,N_4931,N_4982);
nand U5108 (N_5108,N_4919,N_4948);
nor U5109 (N_5109,N_4975,N_4952);
nand U5110 (N_5110,N_4985,N_4943);
and U5111 (N_5111,N_4922,N_4920);
and U5112 (N_5112,N_4927,N_4909);
or U5113 (N_5113,N_4883,N_4882);
nand U5114 (N_5114,N_4898,N_4917);
xor U5115 (N_5115,N_4966,N_4907);
xnor U5116 (N_5116,N_4919,N_4906);
and U5117 (N_5117,N_4976,N_4882);
nand U5118 (N_5118,N_4915,N_4956);
nand U5119 (N_5119,N_4949,N_4883);
and U5120 (N_5120,N_4952,N_4979);
and U5121 (N_5121,N_4877,N_4928);
nor U5122 (N_5122,N_4882,N_4928);
and U5123 (N_5123,N_4888,N_4966);
nand U5124 (N_5124,N_4918,N_4981);
nor U5125 (N_5125,N_5082,N_5052);
or U5126 (N_5126,N_5038,N_5014);
and U5127 (N_5127,N_5107,N_5048);
nand U5128 (N_5128,N_5000,N_5037);
xnor U5129 (N_5129,N_5102,N_5070);
nand U5130 (N_5130,N_5104,N_5123);
and U5131 (N_5131,N_5055,N_5068);
or U5132 (N_5132,N_5036,N_5023);
nand U5133 (N_5133,N_5039,N_5028);
xnor U5134 (N_5134,N_5080,N_5067);
nand U5135 (N_5135,N_5019,N_5099);
nand U5136 (N_5136,N_5091,N_5010);
nand U5137 (N_5137,N_5121,N_5049);
and U5138 (N_5138,N_5059,N_5018);
xor U5139 (N_5139,N_5017,N_5073);
nor U5140 (N_5140,N_5109,N_5016);
xnor U5141 (N_5141,N_5042,N_5119);
xnor U5142 (N_5142,N_5092,N_5066);
nor U5143 (N_5143,N_5057,N_5097);
nor U5144 (N_5144,N_5120,N_5065);
and U5145 (N_5145,N_5084,N_5124);
nor U5146 (N_5146,N_5112,N_5011);
nand U5147 (N_5147,N_5043,N_5027);
or U5148 (N_5148,N_5034,N_5063);
nand U5149 (N_5149,N_5060,N_5020);
nand U5150 (N_5150,N_5078,N_5013);
nand U5151 (N_5151,N_5108,N_5054);
xor U5152 (N_5152,N_5032,N_5050);
and U5153 (N_5153,N_5100,N_5111);
nor U5154 (N_5154,N_5003,N_5098);
or U5155 (N_5155,N_5022,N_5024);
nor U5156 (N_5156,N_5002,N_5025);
and U5157 (N_5157,N_5005,N_5001);
and U5158 (N_5158,N_5101,N_5105);
or U5159 (N_5159,N_5074,N_5029);
nor U5160 (N_5160,N_5079,N_5095);
or U5161 (N_5161,N_5031,N_5009);
nor U5162 (N_5162,N_5115,N_5106);
or U5163 (N_5163,N_5113,N_5058);
or U5164 (N_5164,N_5040,N_5006);
or U5165 (N_5165,N_5103,N_5096);
or U5166 (N_5166,N_5086,N_5026);
or U5167 (N_5167,N_5041,N_5075);
and U5168 (N_5168,N_5056,N_5030);
or U5169 (N_5169,N_5051,N_5061);
nand U5170 (N_5170,N_5110,N_5089);
and U5171 (N_5171,N_5094,N_5116);
and U5172 (N_5172,N_5008,N_5081);
nand U5173 (N_5173,N_5015,N_5035);
nor U5174 (N_5174,N_5088,N_5053);
nor U5175 (N_5175,N_5076,N_5077);
nor U5176 (N_5176,N_5004,N_5047);
and U5177 (N_5177,N_5072,N_5087);
and U5178 (N_5178,N_5044,N_5033);
nand U5179 (N_5179,N_5085,N_5117);
xor U5180 (N_5180,N_5090,N_5064);
xor U5181 (N_5181,N_5071,N_5083);
or U5182 (N_5182,N_5122,N_5007);
and U5183 (N_5183,N_5118,N_5069);
xnor U5184 (N_5184,N_5045,N_5093);
nand U5185 (N_5185,N_5012,N_5114);
nor U5186 (N_5186,N_5021,N_5046);
and U5187 (N_5187,N_5062,N_5076);
or U5188 (N_5188,N_5074,N_5015);
nor U5189 (N_5189,N_5011,N_5119);
nand U5190 (N_5190,N_5087,N_5068);
or U5191 (N_5191,N_5096,N_5068);
nor U5192 (N_5192,N_5110,N_5061);
nand U5193 (N_5193,N_5018,N_5028);
nor U5194 (N_5194,N_5002,N_5113);
and U5195 (N_5195,N_5124,N_5082);
nor U5196 (N_5196,N_5072,N_5067);
xor U5197 (N_5197,N_5055,N_5117);
nand U5198 (N_5198,N_5077,N_5040);
or U5199 (N_5199,N_5098,N_5124);
or U5200 (N_5200,N_5059,N_5112);
and U5201 (N_5201,N_5014,N_5023);
nor U5202 (N_5202,N_5113,N_5080);
nand U5203 (N_5203,N_5021,N_5113);
nor U5204 (N_5204,N_5064,N_5034);
or U5205 (N_5205,N_5116,N_5108);
or U5206 (N_5206,N_5025,N_5103);
nand U5207 (N_5207,N_5023,N_5086);
and U5208 (N_5208,N_5067,N_5010);
and U5209 (N_5209,N_5027,N_5048);
or U5210 (N_5210,N_5060,N_5120);
nor U5211 (N_5211,N_5035,N_5110);
nor U5212 (N_5212,N_5046,N_5020);
and U5213 (N_5213,N_5009,N_5124);
xor U5214 (N_5214,N_5083,N_5052);
or U5215 (N_5215,N_5042,N_5088);
xnor U5216 (N_5216,N_5095,N_5051);
or U5217 (N_5217,N_5041,N_5097);
xnor U5218 (N_5218,N_5083,N_5085);
nand U5219 (N_5219,N_5035,N_5023);
or U5220 (N_5220,N_5080,N_5124);
nor U5221 (N_5221,N_5079,N_5094);
or U5222 (N_5222,N_5082,N_5083);
nor U5223 (N_5223,N_5068,N_5003);
and U5224 (N_5224,N_5028,N_5116);
nand U5225 (N_5225,N_5028,N_5065);
nor U5226 (N_5226,N_5085,N_5000);
xor U5227 (N_5227,N_5120,N_5009);
and U5228 (N_5228,N_5027,N_5081);
nand U5229 (N_5229,N_5075,N_5044);
and U5230 (N_5230,N_5104,N_5094);
or U5231 (N_5231,N_5041,N_5106);
nor U5232 (N_5232,N_5060,N_5095);
nand U5233 (N_5233,N_5062,N_5089);
nor U5234 (N_5234,N_5007,N_5041);
xnor U5235 (N_5235,N_5042,N_5051);
and U5236 (N_5236,N_5106,N_5071);
or U5237 (N_5237,N_5064,N_5016);
nor U5238 (N_5238,N_5008,N_5031);
nor U5239 (N_5239,N_5075,N_5036);
nand U5240 (N_5240,N_5091,N_5052);
nor U5241 (N_5241,N_5104,N_5084);
or U5242 (N_5242,N_5075,N_5111);
or U5243 (N_5243,N_5098,N_5093);
xnor U5244 (N_5244,N_5083,N_5116);
nor U5245 (N_5245,N_5083,N_5004);
nor U5246 (N_5246,N_5032,N_5011);
and U5247 (N_5247,N_5059,N_5109);
nor U5248 (N_5248,N_5028,N_5001);
xor U5249 (N_5249,N_5034,N_5095);
and U5250 (N_5250,N_5186,N_5210);
nor U5251 (N_5251,N_5177,N_5246);
xnor U5252 (N_5252,N_5166,N_5227);
nor U5253 (N_5253,N_5212,N_5126);
or U5254 (N_5254,N_5248,N_5230);
nand U5255 (N_5255,N_5209,N_5223);
nor U5256 (N_5256,N_5187,N_5217);
and U5257 (N_5257,N_5233,N_5162);
and U5258 (N_5258,N_5127,N_5135);
nand U5259 (N_5259,N_5215,N_5184);
xor U5260 (N_5260,N_5143,N_5152);
or U5261 (N_5261,N_5221,N_5176);
or U5262 (N_5262,N_5200,N_5132);
nor U5263 (N_5263,N_5160,N_5129);
nand U5264 (N_5264,N_5170,N_5128);
nand U5265 (N_5265,N_5157,N_5206);
and U5266 (N_5266,N_5141,N_5150);
nand U5267 (N_5267,N_5218,N_5192);
and U5268 (N_5268,N_5243,N_5174);
or U5269 (N_5269,N_5149,N_5219);
or U5270 (N_5270,N_5216,N_5226);
nand U5271 (N_5271,N_5125,N_5205);
nor U5272 (N_5272,N_5140,N_5146);
and U5273 (N_5273,N_5237,N_5133);
or U5274 (N_5274,N_5231,N_5196);
and U5275 (N_5275,N_5232,N_5181);
xor U5276 (N_5276,N_5175,N_5155);
or U5277 (N_5277,N_5191,N_5151);
or U5278 (N_5278,N_5173,N_5193);
nor U5279 (N_5279,N_5225,N_5249);
or U5280 (N_5280,N_5153,N_5139);
or U5281 (N_5281,N_5165,N_5185);
or U5282 (N_5282,N_5207,N_5229);
nor U5283 (N_5283,N_5220,N_5138);
nor U5284 (N_5284,N_5183,N_5168);
nor U5285 (N_5285,N_5159,N_5178);
xor U5286 (N_5286,N_5194,N_5189);
or U5287 (N_5287,N_5245,N_5213);
nand U5288 (N_5288,N_5147,N_5167);
or U5289 (N_5289,N_5208,N_5241);
or U5290 (N_5290,N_5137,N_5244);
nand U5291 (N_5291,N_5171,N_5239);
nor U5292 (N_5292,N_5188,N_5156);
and U5293 (N_5293,N_5158,N_5164);
nor U5294 (N_5294,N_5148,N_5172);
or U5295 (N_5295,N_5145,N_5203);
xor U5296 (N_5296,N_5136,N_5198);
nand U5297 (N_5297,N_5144,N_5201);
nand U5298 (N_5298,N_5234,N_5169);
nor U5299 (N_5299,N_5142,N_5222);
and U5300 (N_5300,N_5180,N_5202);
or U5301 (N_5301,N_5130,N_5242);
nand U5302 (N_5302,N_5182,N_5235);
nor U5303 (N_5303,N_5154,N_5134);
nand U5304 (N_5304,N_5238,N_5179);
nand U5305 (N_5305,N_5224,N_5236);
and U5306 (N_5306,N_5199,N_5214);
nor U5307 (N_5307,N_5240,N_5197);
and U5308 (N_5308,N_5131,N_5204);
nor U5309 (N_5309,N_5211,N_5228);
or U5310 (N_5310,N_5161,N_5190);
or U5311 (N_5311,N_5195,N_5247);
or U5312 (N_5312,N_5163,N_5211);
or U5313 (N_5313,N_5196,N_5125);
nand U5314 (N_5314,N_5160,N_5172);
or U5315 (N_5315,N_5213,N_5194);
nor U5316 (N_5316,N_5186,N_5157);
nor U5317 (N_5317,N_5214,N_5183);
or U5318 (N_5318,N_5232,N_5129);
or U5319 (N_5319,N_5131,N_5184);
nor U5320 (N_5320,N_5203,N_5149);
nor U5321 (N_5321,N_5127,N_5147);
or U5322 (N_5322,N_5125,N_5214);
nor U5323 (N_5323,N_5178,N_5160);
or U5324 (N_5324,N_5152,N_5140);
xnor U5325 (N_5325,N_5235,N_5246);
nor U5326 (N_5326,N_5234,N_5228);
nor U5327 (N_5327,N_5201,N_5164);
nor U5328 (N_5328,N_5225,N_5126);
nand U5329 (N_5329,N_5157,N_5166);
xnor U5330 (N_5330,N_5228,N_5137);
and U5331 (N_5331,N_5166,N_5204);
or U5332 (N_5332,N_5218,N_5214);
or U5333 (N_5333,N_5206,N_5156);
nand U5334 (N_5334,N_5242,N_5241);
nor U5335 (N_5335,N_5157,N_5143);
xnor U5336 (N_5336,N_5208,N_5247);
and U5337 (N_5337,N_5226,N_5214);
or U5338 (N_5338,N_5246,N_5152);
or U5339 (N_5339,N_5205,N_5157);
or U5340 (N_5340,N_5169,N_5212);
nor U5341 (N_5341,N_5143,N_5160);
or U5342 (N_5342,N_5136,N_5189);
nand U5343 (N_5343,N_5145,N_5173);
nand U5344 (N_5344,N_5145,N_5166);
nor U5345 (N_5345,N_5132,N_5241);
and U5346 (N_5346,N_5215,N_5200);
and U5347 (N_5347,N_5131,N_5191);
nor U5348 (N_5348,N_5171,N_5134);
xor U5349 (N_5349,N_5249,N_5172);
nor U5350 (N_5350,N_5236,N_5177);
nor U5351 (N_5351,N_5137,N_5243);
and U5352 (N_5352,N_5224,N_5215);
nand U5353 (N_5353,N_5245,N_5205);
nor U5354 (N_5354,N_5218,N_5219);
and U5355 (N_5355,N_5176,N_5216);
xnor U5356 (N_5356,N_5196,N_5184);
nor U5357 (N_5357,N_5138,N_5137);
nor U5358 (N_5358,N_5223,N_5145);
nor U5359 (N_5359,N_5213,N_5205);
or U5360 (N_5360,N_5168,N_5205);
xor U5361 (N_5361,N_5127,N_5225);
and U5362 (N_5362,N_5241,N_5181);
and U5363 (N_5363,N_5224,N_5206);
or U5364 (N_5364,N_5198,N_5243);
nor U5365 (N_5365,N_5209,N_5196);
nand U5366 (N_5366,N_5150,N_5178);
and U5367 (N_5367,N_5210,N_5200);
and U5368 (N_5368,N_5226,N_5155);
and U5369 (N_5369,N_5188,N_5216);
or U5370 (N_5370,N_5125,N_5133);
nor U5371 (N_5371,N_5214,N_5241);
and U5372 (N_5372,N_5178,N_5147);
nor U5373 (N_5373,N_5234,N_5151);
nor U5374 (N_5374,N_5200,N_5129);
or U5375 (N_5375,N_5334,N_5262);
nand U5376 (N_5376,N_5351,N_5320);
and U5377 (N_5377,N_5311,N_5353);
xnor U5378 (N_5378,N_5255,N_5319);
nor U5379 (N_5379,N_5363,N_5316);
nand U5380 (N_5380,N_5324,N_5323);
nand U5381 (N_5381,N_5263,N_5297);
xnor U5382 (N_5382,N_5269,N_5322);
nand U5383 (N_5383,N_5283,N_5268);
xor U5384 (N_5384,N_5285,N_5256);
or U5385 (N_5385,N_5371,N_5333);
or U5386 (N_5386,N_5291,N_5264);
and U5387 (N_5387,N_5270,N_5349);
and U5388 (N_5388,N_5354,N_5314);
xnor U5389 (N_5389,N_5317,N_5343);
xnor U5390 (N_5390,N_5366,N_5337);
or U5391 (N_5391,N_5364,N_5276);
and U5392 (N_5392,N_5252,N_5318);
and U5393 (N_5393,N_5294,N_5290);
xnor U5394 (N_5394,N_5310,N_5357);
and U5395 (N_5395,N_5368,N_5288);
xnor U5396 (N_5396,N_5335,N_5309);
or U5397 (N_5397,N_5254,N_5271);
nor U5398 (N_5398,N_5327,N_5273);
or U5399 (N_5399,N_5301,N_5307);
nor U5400 (N_5400,N_5260,N_5257);
and U5401 (N_5401,N_5298,N_5348);
nor U5402 (N_5402,N_5300,N_5286);
nand U5403 (N_5403,N_5299,N_5279);
and U5404 (N_5404,N_5281,N_5274);
nand U5405 (N_5405,N_5284,N_5308);
nor U5406 (N_5406,N_5293,N_5251);
nor U5407 (N_5407,N_5280,N_5369);
nor U5408 (N_5408,N_5272,N_5278);
or U5409 (N_5409,N_5266,N_5342);
and U5410 (N_5410,N_5277,N_5250);
and U5411 (N_5411,N_5315,N_5326);
or U5412 (N_5412,N_5367,N_5352);
nand U5413 (N_5413,N_5355,N_5312);
nor U5414 (N_5414,N_5303,N_5362);
nor U5415 (N_5415,N_5360,N_5295);
nor U5416 (N_5416,N_5338,N_5365);
nor U5417 (N_5417,N_5330,N_5253);
or U5418 (N_5418,N_5332,N_5370);
or U5419 (N_5419,N_5350,N_5374);
nor U5420 (N_5420,N_5359,N_5373);
and U5421 (N_5421,N_5328,N_5292);
nor U5422 (N_5422,N_5361,N_5304);
nand U5423 (N_5423,N_5282,N_5372);
or U5424 (N_5424,N_5340,N_5325);
nand U5425 (N_5425,N_5265,N_5341);
or U5426 (N_5426,N_5344,N_5302);
or U5427 (N_5427,N_5358,N_5267);
nor U5428 (N_5428,N_5287,N_5306);
or U5429 (N_5429,N_5275,N_5345);
nand U5430 (N_5430,N_5331,N_5259);
and U5431 (N_5431,N_5339,N_5296);
and U5432 (N_5432,N_5313,N_5346);
nor U5433 (N_5433,N_5321,N_5258);
and U5434 (N_5434,N_5336,N_5261);
and U5435 (N_5435,N_5347,N_5329);
and U5436 (N_5436,N_5289,N_5305);
xnor U5437 (N_5437,N_5356,N_5276);
xor U5438 (N_5438,N_5292,N_5252);
and U5439 (N_5439,N_5364,N_5334);
nor U5440 (N_5440,N_5374,N_5281);
nor U5441 (N_5441,N_5373,N_5357);
nor U5442 (N_5442,N_5316,N_5257);
or U5443 (N_5443,N_5350,N_5316);
nor U5444 (N_5444,N_5352,N_5310);
and U5445 (N_5445,N_5297,N_5275);
nor U5446 (N_5446,N_5345,N_5305);
and U5447 (N_5447,N_5280,N_5264);
nand U5448 (N_5448,N_5329,N_5278);
xnor U5449 (N_5449,N_5271,N_5302);
nand U5450 (N_5450,N_5313,N_5310);
nand U5451 (N_5451,N_5284,N_5258);
or U5452 (N_5452,N_5305,N_5321);
nand U5453 (N_5453,N_5296,N_5357);
nand U5454 (N_5454,N_5283,N_5302);
and U5455 (N_5455,N_5358,N_5345);
xor U5456 (N_5456,N_5304,N_5268);
and U5457 (N_5457,N_5305,N_5368);
or U5458 (N_5458,N_5302,N_5367);
nor U5459 (N_5459,N_5289,N_5356);
nand U5460 (N_5460,N_5275,N_5253);
or U5461 (N_5461,N_5279,N_5296);
nor U5462 (N_5462,N_5360,N_5373);
nor U5463 (N_5463,N_5328,N_5359);
or U5464 (N_5464,N_5300,N_5280);
and U5465 (N_5465,N_5298,N_5264);
nand U5466 (N_5466,N_5332,N_5286);
nand U5467 (N_5467,N_5262,N_5250);
or U5468 (N_5468,N_5314,N_5286);
nor U5469 (N_5469,N_5351,N_5300);
or U5470 (N_5470,N_5321,N_5301);
and U5471 (N_5471,N_5353,N_5254);
nand U5472 (N_5472,N_5340,N_5354);
and U5473 (N_5473,N_5318,N_5344);
nand U5474 (N_5474,N_5371,N_5277);
and U5475 (N_5475,N_5345,N_5328);
and U5476 (N_5476,N_5269,N_5368);
xnor U5477 (N_5477,N_5273,N_5288);
nand U5478 (N_5478,N_5342,N_5264);
nand U5479 (N_5479,N_5348,N_5270);
or U5480 (N_5480,N_5356,N_5293);
xnor U5481 (N_5481,N_5330,N_5260);
and U5482 (N_5482,N_5253,N_5336);
nor U5483 (N_5483,N_5256,N_5351);
and U5484 (N_5484,N_5370,N_5297);
nor U5485 (N_5485,N_5369,N_5288);
xnor U5486 (N_5486,N_5348,N_5257);
or U5487 (N_5487,N_5268,N_5284);
nand U5488 (N_5488,N_5364,N_5355);
xnor U5489 (N_5489,N_5268,N_5344);
and U5490 (N_5490,N_5336,N_5337);
nor U5491 (N_5491,N_5252,N_5277);
or U5492 (N_5492,N_5288,N_5365);
nor U5493 (N_5493,N_5268,N_5352);
nand U5494 (N_5494,N_5358,N_5265);
and U5495 (N_5495,N_5313,N_5288);
xor U5496 (N_5496,N_5289,N_5267);
nor U5497 (N_5497,N_5366,N_5324);
or U5498 (N_5498,N_5327,N_5284);
and U5499 (N_5499,N_5266,N_5330);
nor U5500 (N_5500,N_5425,N_5456);
nand U5501 (N_5501,N_5437,N_5381);
or U5502 (N_5502,N_5442,N_5390);
nor U5503 (N_5503,N_5448,N_5462);
xnor U5504 (N_5504,N_5479,N_5424);
or U5505 (N_5505,N_5495,N_5393);
or U5506 (N_5506,N_5482,N_5483);
nand U5507 (N_5507,N_5384,N_5465);
nand U5508 (N_5508,N_5414,N_5446);
nor U5509 (N_5509,N_5413,N_5474);
nor U5510 (N_5510,N_5481,N_5440);
and U5511 (N_5511,N_5382,N_5411);
nor U5512 (N_5512,N_5486,N_5380);
nor U5513 (N_5513,N_5439,N_5447);
nand U5514 (N_5514,N_5432,N_5422);
or U5515 (N_5515,N_5431,N_5499);
and U5516 (N_5516,N_5472,N_5410);
or U5517 (N_5517,N_5412,N_5455);
xnor U5518 (N_5518,N_5458,N_5377);
or U5519 (N_5519,N_5405,N_5466);
nand U5520 (N_5520,N_5394,N_5404);
nand U5521 (N_5521,N_5469,N_5493);
nand U5522 (N_5522,N_5489,N_5476);
nor U5523 (N_5523,N_5443,N_5427);
nor U5524 (N_5524,N_5473,N_5397);
or U5525 (N_5525,N_5450,N_5470);
or U5526 (N_5526,N_5441,N_5376);
nand U5527 (N_5527,N_5430,N_5407);
xor U5528 (N_5528,N_5379,N_5385);
nor U5529 (N_5529,N_5484,N_5478);
nor U5530 (N_5530,N_5449,N_5496);
and U5531 (N_5531,N_5464,N_5453);
nor U5532 (N_5532,N_5459,N_5477);
and U5533 (N_5533,N_5378,N_5409);
or U5534 (N_5534,N_5435,N_5436);
nor U5535 (N_5535,N_5399,N_5415);
or U5536 (N_5536,N_5463,N_5406);
or U5537 (N_5537,N_5429,N_5402);
or U5538 (N_5538,N_5480,N_5387);
nor U5539 (N_5539,N_5434,N_5403);
nand U5540 (N_5540,N_5497,N_5457);
or U5541 (N_5541,N_5421,N_5433);
nand U5542 (N_5542,N_5460,N_5418);
or U5543 (N_5543,N_5416,N_5492);
nand U5544 (N_5544,N_5491,N_5426);
nor U5545 (N_5545,N_5452,N_5461);
xnor U5546 (N_5546,N_5398,N_5485);
nor U5547 (N_5547,N_5451,N_5391);
nand U5548 (N_5548,N_5375,N_5396);
nand U5549 (N_5549,N_5475,N_5454);
and U5550 (N_5550,N_5419,N_5498);
or U5551 (N_5551,N_5400,N_5386);
or U5552 (N_5552,N_5488,N_5408);
nor U5553 (N_5553,N_5445,N_5467);
or U5554 (N_5554,N_5389,N_5388);
nand U5555 (N_5555,N_5395,N_5423);
nor U5556 (N_5556,N_5490,N_5428);
nand U5557 (N_5557,N_5487,N_5420);
nand U5558 (N_5558,N_5392,N_5417);
nor U5559 (N_5559,N_5471,N_5401);
nand U5560 (N_5560,N_5438,N_5383);
and U5561 (N_5561,N_5444,N_5494);
and U5562 (N_5562,N_5468,N_5400);
nor U5563 (N_5563,N_5445,N_5419);
nor U5564 (N_5564,N_5385,N_5382);
or U5565 (N_5565,N_5425,N_5396);
and U5566 (N_5566,N_5386,N_5398);
or U5567 (N_5567,N_5493,N_5431);
or U5568 (N_5568,N_5385,N_5461);
or U5569 (N_5569,N_5449,N_5403);
or U5570 (N_5570,N_5424,N_5409);
xor U5571 (N_5571,N_5446,N_5375);
or U5572 (N_5572,N_5479,N_5423);
or U5573 (N_5573,N_5487,N_5469);
nor U5574 (N_5574,N_5449,N_5481);
nor U5575 (N_5575,N_5406,N_5427);
and U5576 (N_5576,N_5394,N_5435);
nand U5577 (N_5577,N_5421,N_5497);
or U5578 (N_5578,N_5378,N_5392);
or U5579 (N_5579,N_5436,N_5421);
xor U5580 (N_5580,N_5381,N_5442);
or U5581 (N_5581,N_5444,N_5463);
xnor U5582 (N_5582,N_5403,N_5439);
nand U5583 (N_5583,N_5401,N_5403);
and U5584 (N_5584,N_5398,N_5492);
or U5585 (N_5585,N_5482,N_5399);
and U5586 (N_5586,N_5483,N_5484);
nand U5587 (N_5587,N_5466,N_5394);
or U5588 (N_5588,N_5496,N_5385);
nand U5589 (N_5589,N_5469,N_5444);
nor U5590 (N_5590,N_5456,N_5484);
nor U5591 (N_5591,N_5384,N_5417);
nand U5592 (N_5592,N_5479,N_5386);
or U5593 (N_5593,N_5483,N_5438);
or U5594 (N_5594,N_5443,N_5465);
nor U5595 (N_5595,N_5456,N_5448);
nor U5596 (N_5596,N_5452,N_5454);
nand U5597 (N_5597,N_5375,N_5398);
or U5598 (N_5598,N_5482,N_5446);
and U5599 (N_5599,N_5440,N_5428);
or U5600 (N_5600,N_5441,N_5410);
nor U5601 (N_5601,N_5478,N_5496);
nand U5602 (N_5602,N_5424,N_5420);
or U5603 (N_5603,N_5390,N_5379);
or U5604 (N_5604,N_5407,N_5408);
nand U5605 (N_5605,N_5417,N_5483);
nor U5606 (N_5606,N_5436,N_5396);
or U5607 (N_5607,N_5495,N_5472);
nand U5608 (N_5608,N_5398,N_5475);
nor U5609 (N_5609,N_5473,N_5430);
nand U5610 (N_5610,N_5410,N_5452);
xor U5611 (N_5611,N_5478,N_5459);
nand U5612 (N_5612,N_5394,N_5456);
xor U5613 (N_5613,N_5472,N_5479);
nand U5614 (N_5614,N_5450,N_5391);
or U5615 (N_5615,N_5405,N_5421);
xnor U5616 (N_5616,N_5477,N_5432);
nor U5617 (N_5617,N_5413,N_5471);
or U5618 (N_5618,N_5429,N_5460);
nand U5619 (N_5619,N_5380,N_5498);
nand U5620 (N_5620,N_5424,N_5416);
nor U5621 (N_5621,N_5387,N_5452);
nand U5622 (N_5622,N_5393,N_5442);
or U5623 (N_5623,N_5469,N_5378);
or U5624 (N_5624,N_5420,N_5380);
xor U5625 (N_5625,N_5593,N_5594);
nor U5626 (N_5626,N_5527,N_5551);
nor U5627 (N_5627,N_5555,N_5612);
nand U5628 (N_5628,N_5600,N_5538);
or U5629 (N_5629,N_5546,N_5614);
nand U5630 (N_5630,N_5563,N_5550);
nor U5631 (N_5631,N_5516,N_5605);
or U5632 (N_5632,N_5558,N_5580);
nand U5633 (N_5633,N_5610,N_5536);
nor U5634 (N_5634,N_5588,N_5541);
or U5635 (N_5635,N_5545,N_5520);
or U5636 (N_5636,N_5519,N_5513);
nand U5637 (N_5637,N_5618,N_5559);
and U5638 (N_5638,N_5508,N_5622);
xnor U5639 (N_5639,N_5624,N_5590);
and U5640 (N_5640,N_5620,N_5599);
or U5641 (N_5641,N_5539,N_5589);
nor U5642 (N_5642,N_5613,N_5530);
and U5643 (N_5643,N_5611,N_5549);
nor U5644 (N_5644,N_5586,N_5578);
or U5645 (N_5645,N_5500,N_5534);
or U5646 (N_5646,N_5596,N_5548);
nand U5647 (N_5647,N_5570,N_5619);
nor U5648 (N_5648,N_5511,N_5606);
nand U5649 (N_5649,N_5526,N_5501);
nand U5650 (N_5650,N_5504,N_5573);
nand U5651 (N_5651,N_5583,N_5609);
or U5652 (N_5652,N_5577,N_5521);
xor U5653 (N_5653,N_5556,N_5517);
nand U5654 (N_5654,N_5544,N_5543);
nor U5655 (N_5655,N_5560,N_5581);
nand U5656 (N_5656,N_5506,N_5522);
and U5657 (N_5657,N_5616,N_5561);
and U5658 (N_5658,N_5557,N_5571);
nand U5659 (N_5659,N_5564,N_5602);
xnor U5660 (N_5660,N_5585,N_5592);
or U5661 (N_5661,N_5512,N_5505);
or U5662 (N_5662,N_5532,N_5572);
nor U5663 (N_5663,N_5607,N_5537);
and U5664 (N_5664,N_5623,N_5582);
and U5665 (N_5665,N_5552,N_5533);
nor U5666 (N_5666,N_5591,N_5601);
xor U5667 (N_5667,N_5617,N_5597);
nand U5668 (N_5668,N_5575,N_5542);
or U5669 (N_5669,N_5568,N_5535);
or U5670 (N_5670,N_5553,N_5562);
nand U5671 (N_5671,N_5604,N_5547);
nand U5672 (N_5672,N_5595,N_5566);
nor U5673 (N_5673,N_5565,N_5603);
and U5674 (N_5674,N_5567,N_5529);
and U5675 (N_5675,N_5523,N_5515);
nand U5676 (N_5676,N_5574,N_5540);
or U5677 (N_5677,N_5510,N_5528);
and U5678 (N_5678,N_5525,N_5621);
nand U5679 (N_5679,N_5518,N_5615);
nand U5680 (N_5680,N_5569,N_5587);
xnor U5681 (N_5681,N_5514,N_5598);
and U5682 (N_5682,N_5502,N_5608);
or U5683 (N_5683,N_5509,N_5507);
or U5684 (N_5684,N_5579,N_5584);
nand U5685 (N_5685,N_5576,N_5554);
or U5686 (N_5686,N_5531,N_5503);
and U5687 (N_5687,N_5524,N_5515);
nand U5688 (N_5688,N_5504,N_5552);
or U5689 (N_5689,N_5613,N_5597);
nand U5690 (N_5690,N_5574,N_5607);
or U5691 (N_5691,N_5526,N_5546);
and U5692 (N_5692,N_5567,N_5560);
and U5693 (N_5693,N_5600,N_5561);
nor U5694 (N_5694,N_5571,N_5549);
nor U5695 (N_5695,N_5578,N_5520);
nand U5696 (N_5696,N_5578,N_5508);
nor U5697 (N_5697,N_5544,N_5586);
and U5698 (N_5698,N_5620,N_5534);
nand U5699 (N_5699,N_5503,N_5581);
nor U5700 (N_5700,N_5508,N_5531);
nand U5701 (N_5701,N_5535,N_5618);
or U5702 (N_5702,N_5567,N_5592);
or U5703 (N_5703,N_5504,N_5610);
or U5704 (N_5704,N_5604,N_5534);
nand U5705 (N_5705,N_5553,N_5576);
and U5706 (N_5706,N_5557,N_5501);
or U5707 (N_5707,N_5523,N_5564);
or U5708 (N_5708,N_5518,N_5506);
or U5709 (N_5709,N_5593,N_5577);
nor U5710 (N_5710,N_5563,N_5534);
or U5711 (N_5711,N_5510,N_5527);
or U5712 (N_5712,N_5620,N_5507);
nand U5713 (N_5713,N_5550,N_5519);
and U5714 (N_5714,N_5611,N_5573);
nand U5715 (N_5715,N_5574,N_5585);
or U5716 (N_5716,N_5590,N_5615);
nor U5717 (N_5717,N_5531,N_5562);
nand U5718 (N_5718,N_5547,N_5579);
or U5719 (N_5719,N_5590,N_5599);
or U5720 (N_5720,N_5505,N_5520);
nor U5721 (N_5721,N_5560,N_5523);
or U5722 (N_5722,N_5558,N_5611);
nand U5723 (N_5723,N_5501,N_5512);
nand U5724 (N_5724,N_5558,N_5616);
xor U5725 (N_5725,N_5588,N_5556);
nor U5726 (N_5726,N_5605,N_5584);
or U5727 (N_5727,N_5520,N_5539);
nor U5728 (N_5728,N_5586,N_5509);
nand U5729 (N_5729,N_5546,N_5567);
nand U5730 (N_5730,N_5590,N_5565);
or U5731 (N_5731,N_5609,N_5550);
or U5732 (N_5732,N_5572,N_5600);
nor U5733 (N_5733,N_5572,N_5612);
and U5734 (N_5734,N_5593,N_5550);
or U5735 (N_5735,N_5530,N_5579);
or U5736 (N_5736,N_5505,N_5618);
nor U5737 (N_5737,N_5502,N_5507);
and U5738 (N_5738,N_5596,N_5593);
or U5739 (N_5739,N_5606,N_5586);
xnor U5740 (N_5740,N_5620,N_5595);
nand U5741 (N_5741,N_5581,N_5559);
or U5742 (N_5742,N_5576,N_5566);
and U5743 (N_5743,N_5607,N_5545);
nor U5744 (N_5744,N_5623,N_5537);
nand U5745 (N_5745,N_5552,N_5602);
or U5746 (N_5746,N_5614,N_5560);
nor U5747 (N_5747,N_5512,N_5593);
xnor U5748 (N_5748,N_5518,N_5572);
nor U5749 (N_5749,N_5592,N_5547);
and U5750 (N_5750,N_5629,N_5665);
nand U5751 (N_5751,N_5714,N_5698);
and U5752 (N_5752,N_5666,N_5638);
or U5753 (N_5753,N_5737,N_5677);
nand U5754 (N_5754,N_5674,N_5676);
nor U5755 (N_5755,N_5745,N_5662);
nor U5756 (N_5756,N_5694,N_5725);
or U5757 (N_5757,N_5693,N_5718);
and U5758 (N_5758,N_5653,N_5733);
and U5759 (N_5759,N_5639,N_5668);
and U5760 (N_5760,N_5731,N_5683);
xnor U5761 (N_5761,N_5735,N_5635);
nand U5762 (N_5762,N_5661,N_5656);
nand U5763 (N_5763,N_5705,N_5711);
nor U5764 (N_5764,N_5691,N_5675);
nand U5765 (N_5765,N_5684,N_5728);
and U5766 (N_5766,N_5647,N_5626);
xnor U5767 (N_5767,N_5658,N_5730);
nor U5768 (N_5768,N_5680,N_5654);
nor U5769 (N_5769,N_5747,N_5736);
and U5770 (N_5770,N_5709,N_5703);
xor U5771 (N_5771,N_5636,N_5710);
nand U5772 (N_5772,N_5744,N_5715);
nand U5773 (N_5773,N_5716,N_5670);
nand U5774 (N_5774,N_5660,N_5679);
nand U5775 (N_5775,N_5672,N_5678);
nor U5776 (N_5776,N_5628,N_5687);
and U5777 (N_5777,N_5739,N_5740);
nor U5778 (N_5778,N_5692,N_5726);
nand U5779 (N_5779,N_5708,N_5651);
or U5780 (N_5780,N_5650,N_5700);
and U5781 (N_5781,N_5640,N_5625);
nor U5782 (N_5782,N_5686,N_5663);
and U5783 (N_5783,N_5720,N_5641);
nor U5784 (N_5784,N_5748,N_5630);
and U5785 (N_5785,N_5706,N_5717);
or U5786 (N_5786,N_5671,N_5637);
nor U5787 (N_5787,N_5741,N_5696);
and U5788 (N_5788,N_5704,N_5734);
nor U5789 (N_5789,N_5657,N_5681);
nand U5790 (N_5790,N_5702,N_5631);
and U5791 (N_5791,N_5646,N_5727);
and U5792 (N_5792,N_5699,N_5669);
or U5793 (N_5793,N_5682,N_5649);
nand U5794 (N_5794,N_5689,N_5749);
nor U5795 (N_5795,N_5690,N_5685);
nand U5796 (N_5796,N_5633,N_5743);
nor U5797 (N_5797,N_5742,N_5673);
or U5798 (N_5798,N_5644,N_5707);
and U5799 (N_5799,N_5724,N_5632);
nand U5800 (N_5800,N_5645,N_5697);
or U5801 (N_5801,N_5738,N_5648);
and U5802 (N_5802,N_5746,N_5721);
nand U5803 (N_5803,N_5667,N_5659);
nand U5804 (N_5804,N_5652,N_5664);
and U5805 (N_5805,N_5712,N_5688);
nand U5806 (N_5806,N_5722,N_5642);
and U5807 (N_5807,N_5732,N_5627);
nor U5808 (N_5808,N_5634,N_5655);
nor U5809 (N_5809,N_5719,N_5713);
or U5810 (N_5810,N_5643,N_5701);
or U5811 (N_5811,N_5695,N_5723);
and U5812 (N_5812,N_5729,N_5709);
and U5813 (N_5813,N_5673,N_5714);
nor U5814 (N_5814,N_5746,N_5729);
xnor U5815 (N_5815,N_5705,N_5635);
and U5816 (N_5816,N_5744,N_5704);
and U5817 (N_5817,N_5733,N_5658);
and U5818 (N_5818,N_5683,N_5668);
and U5819 (N_5819,N_5644,N_5716);
or U5820 (N_5820,N_5666,N_5696);
nand U5821 (N_5821,N_5728,N_5702);
nor U5822 (N_5822,N_5700,N_5626);
and U5823 (N_5823,N_5669,N_5749);
nor U5824 (N_5824,N_5717,N_5628);
or U5825 (N_5825,N_5727,N_5735);
nand U5826 (N_5826,N_5677,N_5747);
and U5827 (N_5827,N_5635,N_5672);
nor U5828 (N_5828,N_5678,N_5641);
xor U5829 (N_5829,N_5635,N_5645);
nand U5830 (N_5830,N_5715,N_5674);
or U5831 (N_5831,N_5703,N_5719);
nand U5832 (N_5832,N_5735,N_5710);
and U5833 (N_5833,N_5702,N_5681);
nor U5834 (N_5834,N_5695,N_5668);
xor U5835 (N_5835,N_5704,N_5676);
or U5836 (N_5836,N_5671,N_5657);
nor U5837 (N_5837,N_5685,N_5740);
and U5838 (N_5838,N_5715,N_5676);
or U5839 (N_5839,N_5729,N_5701);
xnor U5840 (N_5840,N_5721,N_5654);
or U5841 (N_5841,N_5671,N_5727);
nand U5842 (N_5842,N_5680,N_5630);
or U5843 (N_5843,N_5675,N_5645);
nand U5844 (N_5844,N_5702,N_5685);
or U5845 (N_5845,N_5666,N_5702);
nand U5846 (N_5846,N_5678,N_5681);
or U5847 (N_5847,N_5733,N_5699);
or U5848 (N_5848,N_5675,N_5724);
or U5849 (N_5849,N_5672,N_5677);
xor U5850 (N_5850,N_5655,N_5732);
nand U5851 (N_5851,N_5730,N_5675);
nand U5852 (N_5852,N_5708,N_5716);
xor U5853 (N_5853,N_5665,N_5727);
or U5854 (N_5854,N_5728,N_5724);
nor U5855 (N_5855,N_5744,N_5711);
nor U5856 (N_5856,N_5734,N_5695);
nor U5857 (N_5857,N_5734,N_5723);
nand U5858 (N_5858,N_5741,N_5639);
nand U5859 (N_5859,N_5748,N_5665);
nand U5860 (N_5860,N_5727,N_5643);
nor U5861 (N_5861,N_5626,N_5636);
or U5862 (N_5862,N_5633,N_5685);
or U5863 (N_5863,N_5726,N_5699);
nand U5864 (N_5864,N_5721,N_5634);
nor U5865 (N_5865,N_5644,N_5739);
or U5866 (N_5866,N_5663,N_5713);
and U5867 (N_5867,N_5726,N_5651);
nor U5868 (N_5868,N_5711,N_5643);
or U5869 (N_5869,N_5692,N_5716);
and U5870 (N_5870,N_5629,N_5689);
and U5871 (N_5871,N_5716,N_5740);
or U5872 (N_5872,N_5655,N_5741);
or U5873 (N_5873,N_5745,N_5645);
nor U5874 (N_5874,N_5656,N_5696);
xnor U5875 (N_5875,N_5796,N_5852);
xnor U5876 (N_5876,N_5828,N_5836);
or U5877 (N_5877,N_5801,N_5833);
nor U5878 (N_5878,N_5786,N_5814);
or U5879 (N_5879,N_5809,N_5769);
and U5880 (N_5880,N_5874,N_5808);
or U5881 (N_5881,N_5784,N_5851);
nor U5882 (N_5882,N_5843,N_5816);
nor U5883 (N_5883,N_5761,N_5822);
or U5884 (N_5884,N_5758,N_5841);
nand U5885 (N_5885,N_5811,N_5834);
and U5886 (N_5886,N_5792,N_5767);
nand U5887 (N_5887,N_5840,N_5832);
nand U5888 (N_5888,N_5847,N_5760);
and U5889 (N_5889,N_5865,N_5805);
xor U5890 (N_5890,N_5845,N_5863);
and U5891 (N_5891,N_5804,N_5859);
or U5892 (N_5892,N_5755,N_5773);
and U5893 (N_5893,N_5854,N_5838);
or U5894 (N_5894,N_5780,N_5781);
xnor U5895 (N_5895,N_5787,N_5818);
xnor U5896 (N_5896,N_5797,N_5858);
nor U5897 (N_5897,N_5753,N_5815);
nor U5898 (N_5898,N_5873,N_5860);
nand U5899 (N_5899,N_5861,N_5830);
nor U5900 (N_5900,N_5868,N_5821);
nor U5901 (N_5901,N_5806,N_5794);
xnor U5902 (N_5902,N_5791,N_5789);
and U5903 (N_5903,N_5807,N_5817);
nand U5904 (N_5904,N_5844,N_5771);
nor U5905 (N_5905,N_5812,N_5855);
or U5906 (N_5906,N_5775,N_5764);
nand U5907 (N_5907,N_5819,N_5837);
nor U5908 (N_5908,N_5788,N_5802);
or U5909 (N_5909,N_5770,N_5850);
xnor U5910 (N_5910,N_5826,N_5798);
or U5911 (N_5911,N_5785,N_5800);
nand U5912 (N_5912,N_5782,N_5754);
and U5913 (N_5913,N_5765,N_5762);
nor U5914 (N_5914,N_5867,N_5799);
or U5915 (N_5915,N_5757,N_5759);
or U5916 (N_5916,N_5853,N_5835);
nor U5917 (N_5917,N_5824,N_5864);
nor U5918 (N_5918,N_5779,N_5869);
and U5919 (N_5919,N_5777,N_5849);
or U5920 (N_5920,N_5846,N_5766);
or U5921 (N_5921,N_5870,N_5857);
xnor U5922 (N_5922,N_5871,N_5842);
or U5923 (N_5923,N_5803,N_5768);
nand U5924 (N_5924,N_5862,N_5823);
and U5925 (N_5925,N_5829,N_5790);
nor U5926 (N_5926,N_5793,N_5778);
or U5927 (N_5927,N_5752,N_5872);
nor U5928 (N_5928,N_5839,N_5848);
and U5929 (N_5929,N_5774,N_5810);
xnor U5930 (N_5930,N_5820,N_5856);
nand U5931 (N_5931,N_5772,N_5776);
nor U5932 (N_5932,N_5866,N_5825);
or U5933 (N_5933,N_5756,N_5795);
nand U5934 (N_5934,N_5783,N_5751);
nand U5935 (N_5935,N_5763,N_5827);
xor U5936 (N_5936,N_5813,N_5831);
nor U5937 (N_5937,N_5750,N_5837);
nand U5938 (N_5938,N_5832,N_5837);
nor U5939 (N_5939,N_5845,N_5807);
nor U5940 (N_5940,N_5828,N_5752);
and U5941 (N_5941,N_5833,N_5772);
or U5942 (N_5942,N_5836,N_5824);
nor U5943 (N_5943,N_5777,N_5814);
xor U5944 (N_5944,N_5829,N_5775);
and U5945 (N_5945,N_5822,N_5796);
nor U5946 (N_5946,N_5807,N_5836);
nand U5947 (N_5947,N_5810,N_5817);
nor U5948 (N_5948,N_5824,N_5866);
nand U5949 (N_5949,N_5804,N_5830);
and U5950 (N_5950,N_5864,N_5870);
and U5951 (N_5951,N_5768,N_5843);
or U5952 (N_5952,N_5850,N_5792);
nand U5953 (N_5953,N_5811,N_5760);
and U5954 (N_5954,N_5858,N_5844);
nand U5955 (N_5955,N_5811,N_5856);
nor U5956 (N_5956,N_5826,N_5852);
and U5957 (N_5957,N_5754,N_5803);
or U5958 (N_5958,N_5793,N_5756);
or U5959 (N_5959,N_5788,N_5839);
or U5960 (N_5960,N_5818,N_5808);
and U5961 (N_5961,N_5811,N_5777);
xor U5962 (N_5962,N_5803,N_5789);
and U5963 (N_5963,N_5835,N_5784);
nor U5964 (N_5964,N_5786,N_5831);
xor U5965 (N_5965,N_5828,N_5866);
nand U5966 (N_5966,N_5787,N_5805);
and U5967 (N_5967,N_5781,N_5860);
or U5968 (N_5968,N_5787,N_5792);
xor U5969 (N_5969,N_5811,N_5859);
or U5970 (N_5970,N_5815,N_5775);
and U5971 (N_5971,N_5873,N_5791);
xor U5972 (N_5972,N_5787,N_5826);
nor U5973 (N_5973,N_5837,N_5828);
nand U5974 (N_5974,N_5870,N_5835);
nor U5975 (N_5975,N_5856,N_5801);
or U5976 (N_5976,N_5757,N_5750);
nor U5977 (N_5977,N_5850,N_5801);
xnor U5978 (N_5978,N_5820,N_5817);
xor U5979 (N_5979,N_5767,N_5870);
and U5980 (N_5980,N_5849,N_5863);
or U5981 (N_5981,N_5833,N_5769);
nand U5982 (N_5982,N_5817,N_5751);
nand U5983 (N_5983,N_5823,N_5819);
nor U5984 (N_5984,N_5777,N_5865);
and U5985 (N_5985,N_5771,N_5826);
or U5986 (N_5986,N_5781,N_5829);
and U5987 (N_5987,N_5805,N_5764);
nor U5988 (N_5988,N_5812,N_5845);
nand U5989 (N_5989,N_5855,N_5818);
or U5990 (N_5990,N_5853,N_5778);
nand U5991 (N_5991,N_5863,N_5814);
or U5992 (N_5992,N_5769,N_5822);
nand U5993 (N_5993,N_5780,N_5872);
and U5994 (N_5994,N_5847,N_5802);
nand U5995 (N_5995,N_5835,N_5861);
and U5996 (N_5996,N_5775,N_5841);
nand U5997 (N_5997,N_5862,N_5843);
and U5998 (N_5998,N_5760,N_5850);
nor U5999 (N_5999,N_5834,N_5782);
xnor U6000 (N_6000,N_5988,N_5991);
or U6001 (N_6001,N_5902,N_5938);
or U6002 (N_6002,N_5887,N_5973);
and U6003 (N_6003,N_5948,N_5989);
nor U6004 (N_6004,N_5882,N_5904);
nor U6005 (N_6005,N_5950,N_5924);
or U6006 (N_6006,N_5953,N_5954);
and U6007 (N_6007,N_5971,N_5998);
nor U6008 (N_6008,N_5933,N_5905);
nor U6009 (N_6009,N_5980,N_5982);
nor U6010 (N_6010,N_5936,N_5934);
or U6011 (N_6011,N_5891,N_5926);
and U6012 (N_6012,N_5955,N_5911);
nor U6013 (N_6013,N_5928,N_5910);
or U6014 (N_6014,N_5978,N_5995);
nor U6015 (N_6015,N_5990,N_5914);
and U6016 (N_6016,N_5996,N_5919);
and U6017 (N_6017,N_5906,N_5899);
xor U6018 (N_6018,N_5877,N_5916);
nand U6019 (N_6019,N_5943,N_5967);
xor U6020 (N_6020,N_5913,N_5993);
nand U6021 (N_6021,N_5875,N_5895);
nand U6022 (N_6022,N_5949,N_5927);
nor U6023 (N_6023,N_5883,N_5940);
and U6024 (N_6024,N_5884,N_5944);
nor U6025 (N_6025,N_5930,N_5897);
nor U6026 (N_6026,N_5992,N_5881);
nor U6027 (N_6027,N_5907,N_5921);
or U6028 (N_6028,N_5959,N_5970);
nand U6029 (N_6029,N_5892,N_5986);
or U6030 (N_6030,N_5908,N_5931);
or U6031 (N_6031,N_5984,N_5925);
nand U6032 (N_6032,N_5923,N_5901);
or U6033 (N_6033,N_5977,N_5947);
and U6034 (N_6034,N_5961,N_5880);
nand U6035 (N_6035,N_5885,N_5964);
and U6036 (N_6036,N_5935,N_5985);
or U6037 (N_6037,N_5975,N_5974);
nand U6038 (N_6038,N_5912,N_5965);
nor U6039 (N_6039,N_5969,N_5987);
nor U6040 (N_6040,N_5932,N_5909);
nor U6041 (N_6041,N_5879,N_5920);
nand U6042 (N_6042,N_5966,N_5886);
and U6043 (N_6043,N_5893,N_5941);
nor U6044 (N_6044,N_5979,N_5968);
or U6045 (N_6045,N_5994,N_5922);
nor U6046 (N_6046,N_5896,N_5917);
and U6047 (N_6047,N_5939,N_5937);
and U6048 (N_6048,N_5962,N_5889);
xor U6049 (N_6049,N_5956,N_5900);
nor U6050 (N_6050,N_5915,N_5999);
nor U6051 (N_6051,N_5983,N_5942);
nand U6052 (N_6052,N_5958,N_5997);
nor U6053 (N_6053,N_5952,N_5945);
nand U6054 (N_6054,N_5903,N_5894);
or U6055 (N_6055,N_5878,N_5957);
and U6056 (N_6056,N_5960,N_5976);
or U6057 (N_6057,N_5951,N_5963);
xor U6058 (N_6058,N_5946,N_5981);
nor U6059 (N_6059,N_5929,N_5876);
or U6060 (N_6060,N_5972,N_5918);
nand U6061 (N_6061,N_5898,N_5888);
nand U6062 (N_6062,N_5890,N_5905);
nor U6063 (N_6063,N_5967,N_5962);
xor U6064 (N_6064,N_5971,N_5886);
and U6065 (N_6065,N_5930,N_5943);
xor U6066 (N_6066,N_5906,N_5898);
and U6067 (N_6067,N_5978,N_5903);
nand U6068 (N_6068,N_5919,N_5928);
nor U6069 (N_6069,N_5997,N_5968);
nand U6070 (N_6070,N_5957,N_5893);
xnor U6071 (N_6071,N_5898,N_5982);
xor U6072 (N_6072,N_5900,N_5892);
nand U6073 (N_6073,N_5994,N_5897);
or U6074 (N_6074,N_5980,N_5918);
nor U6075 (N_6075,N_5938,N_5950);
and U6076 (N_6076,N_5957,N_5945);
nand U6077 (N_6077,N_5900,N_5992);
nand U6078 (N_6078,N_5998,N_5947);
nand U6079 (N_6079,N_5896,N_5990);
or U6080 (N_6080,N_5957,N_5918);
xor U6081 (N_6081,N_5926,N_5922);
nand U6082 (N_6082,N_5876,N_5972);
and U6083 (N_6083,N_5901,N_5954);
and U6084 (N_6084,N_5901,N_5922);
nand U6085 (N_6085,N_5911,N_5877);
nand U6086 (N_6086,N_5972,N_5909);
nand U6087 (N_6087,N_5914,N_5971);
nand U6088 (N_6088,N_5911,N_5992);
nand U6089 (N_6089,N_5932,N_5969);
nand U6090 (N_6090,N_5949,N_5935);
nand U6091 (N_6091,N_5968,N_5898);
nor U6092 (N_6092,N_5886,N_5926);
and U6093 (N_6093,N_5894,N_5962);
xnor U6094 (N_6094,N_5891,N_5952);
or U6095 (N_6095,N_5903,N_5919);
xor U6096 (N_6096,N_5992,N_5966);
xor U6097 (N_6097,N_5977,N_5965);
or U6098 (N_6098,N_5991,N_5973);
nand U6099 (N_6099,N_5983,N_5950);
xnor U6100 (N_6100,N_5932,N_5885);
nand U6101 (N_6101,N_5979,N_5962);
and U6102 (N_6102,N_5952,N_5977);
xor U6103 (N_6103,N_5975,N_5923);
nand U6104 (N_6104,N_5891,N_5897);
and U6105 (N_6105,N_5901,N_5936);
or U6106 (N_6106,N_5926,N_5920);
nor U6107 (N_6107,N_5970,N_5969);
or U6108 (N_6108,N_5941,N_5937);
or U6109 (N_6109,N_5940,N_5972);
nor U6110 (N_6110,N_5888,N_5970);
or U6111 (N_6111,N_5904,N_5973);
nor U6112 (N_6112,N_5980,N_5942);
nor U6113 (N_6113,N_5934,N_5982);
nand U6114 (N_6114,N_5915,N_5903);
nand U6115 (N_6115,N_5969,N_5974);
nand U6116 (N_6116,N_5883,N_5931);
xnor U6117 (N_6117,N_5995,N_5941);
and U6118 (N_6118,N_5909,N_5998);
or U6119 (N_6119,N_5955,N_5906);
nand U6120 (N_6120,N_5900,N_5969);
or U6121 (N_6121,N_5913,N_5989);
or U6122 (N_6122,N_5985,N_5930);
or U6123 (N_6123,N_5912,N_5986);
nor U6124 (N_6124,N_5949,N_5985);
nand U6125 (N_6125,N_6009,N_6027);
nand U6126 (N_6126,N_6090,N_6020);
xnor U6127 (N_6127,N_6059,N_6057);
nor U6128 (N_6128,N_6000,N_6080);
or U6129 (N_6129,N_6100,N_6033);
nor U6130 (N_6130,N_6049,N_6030);
or U6131 (N_6131,N_6052,N_6008);
or U6132 (N_6132,N_6078,N_6097);
nand U6133 (N_6133,N_6019,N_6067);
nand U6134 (N_6134,N_6086,N_6114);
nor U6135 (N_6135,N_6088,N_6031);
and U6136 (N_6136,N_6016,N_6075);
nand U6137 (N_6137,N_6021,N_6041);
xnor U6138 (N_6138,N_6110,N_6096);
nor U6139 (N_6139,N_6108,N_6112);
and U6140 (N_6140,N_6113,N_6010);
or U6141 (N_6141,N_6098,N_6048);
nor U6142 (N_6142,N_6042,N_6066);
or U6143 (N_6143,N_6087,N_6107);
or U6144 (N_6144,N_6116,N_6092);
nor U6145 (N_6145,N_6064,N_6117);
nor U6146 (N_6146,N_6068,N_6091);
nand U6147 (N_6147,N_6026,N_6013);
or U6148 (N_6148,N_6083,N_6065);
nand U6149 (N_6149,N_6085,N_6103);
or U6150 (N_6150,N_6121,N_6037);
or U6151 (N_6151,N_6109,N_6047);
nand U6152 (N_6152,N_6101,N_6040);
and U6153 (N_6153,N_6095,N_6069);
and U6154 (N_6154,N_6029,N_6028);
nor U6155 (N_6155,N_6035,N_6106);
nor U6156 (N_6156,N_6124,N_6023);
or U6157 (N_6157,N_6122,N_6012);
or U6158 (N_6158,N_6076,N_6018);
nand U6159 (N_6159,N_6062,N_6079);
and U6160 (N_6160,N_6056,N_6111);
and U6161 (N_6161,N_6054,N_6002);
nand U6162 (N_6162,N_6007,N_6017);
nand U6163 (N_6163,N_6036,N_6123);
or U6164 (N_6164,N_6077,N_6115);
or U6165 (N_6165,N_6004,N_6053);
nand U6166 (N_6166,N_6039,N_6014);
nor U6167 (N_6167,N_6038,N_6032);
nand U6168 (N_6168,N_6089,N_6072);
nor U6169 (N_6169,N_6050,N_6119);
or U6170 (N_6170,N_6055,N_6005);
xor U6171 (N_6171,N_6015,N_6043);
or U6172 (N_6172,N_6082,N_6084);
nand U6173 (N_6173,N_6003,N_6070);
nand U6174 (N_6174,N_6022,N_6081);
nor U6175 (N_6175,N_6006,N_6099);
nor U6176 (N_6176,N_6118,N_6120);
nor U6177 (N_6177,N_6044,N_6071);
nand U6178 (N_6178,N_6074,N_6024);
and U6179 (N_6179,N_6094,N_6045);
nor U6180 (N_6180,N_6061,N_6025);
nand U6181 (N_6181,N_6046,N_6105);
and U6182 (N_6182,N_6058,N_6060);
nor U6183 (N_6183,N_6001,N_6034);
and U6184 (N_6184,N_6093,N_6011);
nor U6185 (N_6185,N_6051,N_6104);
and U6186 (N_6186,N_6073,N_6102);
nor U6187 (N_6187,N_6063,N_6002);
and U6188 (N_6188,N_6019,N_6058);
xnor U6189 (N_6189,N_6035,N_6118);
and U6190 (N_6190,N_6060,N_6046);
and U6191 (N_6191,N_6118,N_6109);
or U6192 (N_6192,N_6064,N_6002);
or U6193 (N_6193,N_6066,N_6121);
xnor U6194 (N_6194,N_6039,N_6058);
nand U6195 (N_6195,N_6091,N_6107);
nor U6196 (N_6196,N_6098,N_6084);
nand U6197 (N_6197,N_6029,N_6107);
or U6198 (N_6198,N_6084,N_6075);
nor U6199 (N_6199,N_6058,N_6101);
and U6200 (N_6200,N_6102,N_6024);
and U6201 (N_6201,N_6029,N_6012);
nor U6202 (N_6202,N_6061,N_6047);
or U6203 (N_6203,N_6092,N_6108);
nor U6204 (N_6204,N_6092,N_6030);
or U6205 (N_6205,N_6112,N_6019);
nor U6206 (N_6206,N_6018,N_6093);
and U6207 (N_6207,N_6077,N_6070);
or U6208 (N_6208,N_6063,N_6003);
or U6209 (N_6209,N_6096,N_6007);
nand U6210 (N_6210,N_6048,N_6069);
or U6211 (N_6211,N_6093,N_6060);
nor U6212 (N_6212,N_6118,N_6057);
nand U6213 (N_6213,N_6023,N_6053);
and U6214 (N_6214,N_6086,N_6113);
or U6215 (N_6215,N_6034,N_6074);
or U6216 (N_6216,N_6105,N_6023);
or U6217 (N_6217,N_6037,N_6105);
and U6218 (N_6218,N_6094,N_6087);
nand U6219 (N_6219,N_6041,N_6005);
nand U6220 (N_6220,N_6014,N_6059);
xor U6221 (N_6221,N_6025,N_6031);
nand U6222 (N_6222,N_6108,N_6026);
and U6223 (N_6223,N_6023,N_6112);
xor U6224 (N_6224,N_6091,N_6089);
and U6225 (N_6225,N_6062,N_6018);
xor U6226 (N_6226,N_6081,N_6069);
nor U6227 (N_6227,N_6068,N_6115);
nor U6228 (N_6228,N_6095,N_6073);
nor U6229 (N_6229,N_6100,N_6123);
and U6230 (N_6230,N_6107,N_6079);
and U6231 (N_6231,N_6024,N_6089);
and U6232 (N_6232,N_6058,N_6029);
or U6233 (N_6233,N_6091,N_6015);
or U6234 (N_6234,N_6041,N_6109);
and U6235 (N_6235,N_6092,N_6043);
and U6236 (N_6236,N_6077,N_6028);
or U6237 (N_6237,N_6121,N_6005);
and U6238 (N_6238,N_6078,N_6053);
or U6239 (N_6239,N_6061,N_6040);
nor U6240 (N_6240,N_6025,N_6051);
or U6241 (N_6241,N_6123,N_6097);
and U6242 (N_6242,N_6085,N_6004);
nand U6243 (N_6243,N_6080,N_6005);
nor U6244 (N_6244,N_6034,N_6072);
and U6245 (N_6245,N_6033,N_6031);
and U6246 (N_6246,N_6063,N_6096);
or U6247 (N_6247,N_6108,N_6060);
and U6248 (N_6248,N_6072,N_6088);
or U6249 (N_6249,N_6019,N_6042);
nand U6250 (N_6250,N_6183,N_6193);
nand U6251 (N_6251,N_6232,N_6216);
nor U6252 (N_6252,N_6168,N_6204);
xnor U6253 (N_6253,N_6190,N_6135);
nor U6254 (N_6254,N_6208,N_6224);
nor U6255 (N_6255,N_6202,N_6182);
nand U6256 (N_6256,N_6148,N_6217);
nor U6257 (N_6257,N_6171,N_6198);
or U6258 (N_6258,N_6210,N_6241);
and U6259 (N_6259,N_6184,N_6142);
nor U6260 (N_6260,N_6235,N_6152);
nand U6261 (N_6261,N_6179,N_6128);
or U6262 (N_6262,N_6167,N_6157);
xnor U6263 (N_6263,N_6175,N_6195);
and U6264 (N_6264,N_6199,N_6219);
or U6265 (N_6265,N_6129,N_6147);
and U6266 (N_6266,N_6166,N_6130);
nor U6267 (N_6267,N_6196,N_6178);
and U6268 (N_6268,N_6159,N_6243);
or U6269 (N_6269,N_6236,N_6244);
or U6270 (N_6270,N_6212,N_6230);
nand U6271 (N_6271,N_6172,N_6247);
nor U6272 (N_6272,N_6249,N_6225);
nand U6273 (N_6273,N_6209,N_6141);
or U6274 (N_6274,N_6177,N_6211);
nand U6275 (N_6275,N_6136,N_6161);
nand U6276 (N_6276,N_6203,N_6156);
and U6277 (N_6277,N_6221,N_6189);
nor U6278 (N_6278,N_6134,N_6154);
or U6279 (N_6279,N_6197,N_6214);
nand U6280 (N_6280,N_6192,N_6242);
or U6281 (N_6281,N_6165,N_6139);
nor U6282 (N_6282,N_6133,N_6191);
nand U6283 (N_6283,N_6173,N_6215);
nor U6284 (N_6284,N_6160,N_6176);
or U6285 (N_6285,N_6213,N_6163);
nand U6286 (N_6286,N_6222,N_6145);
nor U6287 (N_6287,N_6229,N_6228);
nand U6288 (N_6288,N_6144,N_6188);
or U6289 (N_6289,N_6153,N_6180);
or U6290 (N_6290,N_6201,N_6126);
or U6291 (N_6291,N_6181,N_6187);
nor U6292 (N_6292,N_6246,N_6218);
nor U6293 (N_6293,N_6149,N_6231);
nor U6294 (N_6294,N_6169,N_6132);
and U6295 (N_6295,N_6205,N_6158);
xnor U6296 (N_6296,N_6248,N_6127);
nor U6297 (N_6297,N_6140,N_6227);
nor U6298 (N_6298,N_6137,N_6239);
nand U6299 (N_6299,N_6162,N_6245);
and U6300 (N_6300,N_6185,N_6138);
xor U6301 (N_6301,N_6226,N_6151);
nand U6302 (N_6302,N_6200,N_6237);
and U6303 (N_6303,N_6194,N_6233);
and U6304 (N_6304,N_6164,N_6146);
and U6305 (N_6305,N_6170,N_6174);
and U6306 (N_6306,N_6223,N_6206);
and U6307 (N_6307,N_6186,N_6143);
and U6308 (N_6308,N_6234,N_6131);
nand U6309 (N_6309,N_6155,N_6207);
or U6310 (N_6310,N_6150,N_6125);
and U6311 (N_6311,N_6238,N_6220);
xor U6312 (N_6312,N_6240,N_6133);
and U6313 (N_6313,N_6126,N_6164);
nor U6314 (N_6314,N_6175,N_6146);
nand U6315 (N_6315,N_6146,N_6196);
nor U6316 (N_6316,N_6154,N_6213);
nand U6317 (N_6317,N_6242,N_6178);
xor U6318 (N_6318,N_6143,N_6168);
nor U6319 (N_6319,N_6197,N_6226);
nand U6320 (N_6320,N_6245,N_6206);
and U6321 (N_6321,N_6184,N_6229);
nor U6322 (N_6322,N_6133,N_6154);
and U6323 (N_6323,N_6191,N_6137);
and U6324 (N_6324,N_6172,N_6233);
and U6325 (N_6325,N_6162,N_6170);
nand U6326 (N_6326,N_6200,N_6178);
nor U6327 (N_6327,N_6228,N_6208);
and U6328 (N_6328,N_6197,N_6223);
or U6329 (N_6329,N_6216,N_6188);
nor U6330 (N_6330,N_6242,N_6151);
or U6331 (N_6331,N_6190,N_6207);
nor U6332 (N_6332,N_6151,N_6135);
or U6333 (N_6333,N_6241,N_6146);
nor U6334 (N_6334,N_6244,N_6185);
xnor U6335 (N_6335,N_6144,N_6221);
nand U6336 (N_6336,N_6185,N_6130);
or U6337 (N_6337,N_6201,N_6137);
nand U6338 (N_6338,N_6231,N_6211);
or U6339 (N_6339,N_6188,N_6209);
nand U6340 (N_6340,N_6202,N_6139);
nor U6341 (N_6341,N_6225,N_6176);
and U6342 (N_6342,N_6197,N_6222);
nand U6343 (N_6343,N_6165,N_6191);
or U6344 (N_6344,N_6135,N_6180);
and U6345 (N_6345,N_6169,N_6205);
or U6346 (N_6346,N_6198,N_6144);
or U6347 (N_6347,N_6208,N_6222);
and U6348 (N_6348,N_6138,N_6160);
or U6349 (N_6349,N_6242,N_6146);
nor U6350 (N_6350,N_6181,N_6165);
and U6351 (N_6351,N_6200,N_6248);
nand U6352 (N_6352,N_6215,N_6245);
or U6353 (N_6353,N_6207,N_6228);
nor U6354 (N_6354,N_6211,N_6170);
nor U6355 (N_6355,N_6196,N_6169);
or U6356 (N_6356,N_6211,N_6207);
nor U6357 (N_6357,N_6216,N_6147);
xor U6358 (N_6358,N_6202,N_6189);
or U6359 (N_6359,N_6236,N_6191);
and U6360 (N_6360,N_6167,N_6204);
or U6361 (N_6361,N_6130,N_6175);
and U6362 (N_6362,N_6197,N_6163);
nand U6363 (N_6363,N_6211,N_6126);
xnor U6364 (N_6364,N_6166,N_6224);
nand U6365 (N_6365,N_6201,N_6131);
or U6366 (N_6366,N_6150,N_6142);
nand U6367 (N_6367,N_6177,N_6128);
nor U6368 (N_6368,N_6165,N_6158);
nor U6369 (N_6369,N_6143,N_6232);
xnor U6370 (N_6370,N_6184,N_6143);
nor U6371 (N_6371,N_6146,N_6208);
or U6372 (N_6372,N_6195,N_6146);
and U6373 (N_6373,N_6242,N_6126);
nand U6374 (N_6374,N_6179,N_6139);
nand U6375 (N_6375,N_6267,N_6275);
xnor U6376 (N_6376,N_6348,N_6269);
nand U6377 (N_6377,N_6273,N_6367);
or U6378 (N_6378,N_6317,N_6305);
nor U6379 (N_6379,N_6351,N_6300);
nor U6380 (N_6380,N_6293,N_6349);
or U6381 (N_6381,N_6330,N_6289);
nor U6382 (N_6382,N_6355,N_6327);
or U6383 (N_6383,N_6320,N_6254);
nand U6384 (N_6384,N_6308,N_6279);
nand U6385 (N_6385,N_6360,N_6363);
nand U6386 (N_6386,N_6372,N_6331);
or U6387 (N_6387,N_6288,N_6298);
nand U6388 (N_6388,N_6371,N_6303);
and U6389 (N_6389,N_6359,N_6272);
nand U6390 (N_6390,N_6294,N_6335);
xor U6391 (N_6391,N_6336,N_6256);
xor U6392 (N_6392,N_6265,N_6270);
nor U6393 (N_6393,N_6292,N_6324);
xor U6394 (N_6394,N_6304,N_6326);
and U6395 (N_6395,N_6319,N_6295);
or U6396 (N_6396,N_6352,N_6358);
and U6397 (N_6397,N_6350,N_6291);
nor U6398 (N_6398,N_6338,N_6345);
nand U6399 (N_6399,N_6339,N_6285);
nand U6400 (N_6400,N_6318,N_6301);
and U6401 (N_6401,N_6356,N_6344);
nor U6402 (N_6402,N_6364,N_6365);
xnor U6403 (N_6403,N_6252,N_6260);
nand U6404 (N_6404,N_6347,N_6284);
nor U6405 (N_6405,N_6354,N_6334);
or U6406 (N_6406,N_6374,N_6313);
nand U6407 (N_6407,N_6307,N_6309);
and U6408 (N_6408,N_6258,N_6312);
nor U6409 (N_6409,N_6268,N_6302);
xnor U6410 (N_6410,N_6253,N_6266);
or U6411 (N_6411,N_6286,N_6337);
xnor U6412 (N_6412,N_6251,N_6287);
or U6413 (N_6413,N_6353,N_6373);
nor U6414 (N_6414,N_6263,N_6277);
xnor U6415 (N_6415,N_6362,N_6370);
and U6416 (N_6416,N_6264,N_6257);
nor U6417 (N_6417,N_6280,N_6290);
and U6418 (N_6418,N_6278,N_6341);
nor U6419 (N_6419,N_6321,N_6281);
nor U6420 (N_6420,N_6296,N_6297);
or U6421 (N_6421,N_6274,N_6306);
and U6422 (N_6422,N_6333,N_6342);
or U6423 (N_6423,N_6361,N_6314);
or U6424 (N_6424,N_6271,N_6316);
nor U6425 (N_6425,N_6332,N_6283);
nor U6426 (N_6426,N_6346,N_6322);
or U6427 (N_6427,N_6343,N_6328);
and U6428 (N_6428,N_6299,N_6357);
nor U6429 (N_6429,N_6329,N_6366);
nand U6430 (N_6430,N_6340,N_6315);
and U6431 (N_6431,N_6368,N_6259);
nand U6432 (N_6432,N_6282,N_6262);
xor U6433 (N_6433,N_6255,N_6311);
and U6434 (N_6434,N_6323,N_6310);
nor U6435 (N_6435,N_6276,N_6261);
or U6436 (N_6436,N_6369,N_6325);
or U6437 (N_6437,N_6250,N_6265);
or U6438 (N_6438,N_6294,N_6350);
nand U6439 (N_6439,N_6371,N_6276);
nor U6440 (N_6440,N_6345,N_6370);
or U6441 (N_6441,N_6364,N_6366);
or U6442 (N_6442,N_6368,N_6318);
or U6443 (N_6443,N_6295,N_6310);
and U6444 (N_6444,N_6345,N_6364);
xor U6445 (N_6445,N_6304,N_6275);
nand U6446 (N_6446,N_6313,N_6295);
xnor U6447 (N_6447,N_6350,N_6284);
nand U6448 (N_6448,N_6321,N_6255);
xnor U6449 (N_6449,N_6270,N_6296);
and U6450 (N_6450,N_6361,N_6255);
nand U6451 (N_6451,N_6343,N_6278);
nor U6452 (N_6452,N_6306,N_6323);
nand U6453 (N_6453,N_6259,N_6357);
or U6454 (N_6454,N_6266,N_6325);
nand U6455 (N_6455,N_6373,N_6251);
and U6456 (N_6456,N_6324,N_6286);
or U6457 (N_6457,N_6289,N_6358);
and U6458 (N_6458,N_6355,N_6330);
xor U6459 (N_6459,N_6314,N_6318);
and U6460 (N_6460,N_6369,N_6311);
nand U6461 (N_6461,N_6370,N_6368);
nor U6462 (N_6462,N_6279,N_6250);
xor U6463 (N_6463,N_6292,N_6260);
or U6464 (N_6464,N_6322,N_6251);
and U6465 (N_6465,N_6340,N_6305);
or U6466 (N_6466,N_6317,N_6360);
or U6467 (N_6467,N_6321,N_6347);
nor U6468 (N_6468,N_6272,N_6314);
or U6469 (N_6469,N_6364,N_6372);
and U6470 (N_6470,N_6255,N_6337);
and U6471 (N_6471,N_6359,N_6349);
or U6472 (N_6472,N_6332,N_6267);
nand U6473 (N_6473,N_6341,N_6347);
or U6474 (N_6474,N_6276,N_6289);
nand U6475 (N_6475,N_6352,N_6343);
xnor U6476 (N_6476,N_6309,N_6327);
nand U6477 (N_6477,N_6349,N_6280);
nand U6478 (N_6478,N_6289,N_6309);
nand U6479 (N_6479,N_6250,N_6303);
xnor U6480 (N_6480,N_6297,N_6331);
nand U6481 (N_6481,N_6333,N_6264);
and U6482 (N_6482,N_6341,N_6366);
xnor U6483 (N_6483,N_6314,N_6277);
nand U6484 (N_6484,N_6350,N_6311);
and U6485 (N_6485,N_6325,N_6367);
xor U6486 (N_6486,N_6266,N_6292);
and U6487 (N_6487,N_6354,N_6310);
nor U6488 (N_6488,N_6296,N_6288);
nand U6489 (N_6489,N_6328,N_6292);
or U6490 (N_6490,N_6282,N_6297);
and U6491 (N_6491,N_6292,N_6335);
or U6492 (N_6492,N_6298,N_6369);
nand U6493 (N_6493,N_6364,N_6339);
nand U6494 (N_6494,N_6321,N_6361);
nor U6495 (N_6495,N_6341,N_6355);
and U6496 (N_6496,N_6267,N_6256);
or U6497 (N_6497,N_6265,N_6311);
nand U6498 (N_6498,N_6309,N_6274);
and U6499 (N_6499,N_6341,N_6311);
or U6500 (N_6500,N_6436,N_6483);
and U6501 (N_6501,N_6450,N_6409);
nor U6502 (N_6502,N_6490,N_6402);
or U6503 (N_6503,N_6401,N_6378);
nor U6504 (N_6504,N_6481,N_6474);
and U6505 (N_6505,N_6434,N_6375);
nand U6506 (N_6506,N_6385,N_6485);
and U6507 (N_6507,N_6384,N_6423);
nor U6508 (N_6508,N_6477,N_6388);
nand U6509 (N_6509,N_6480,N_6496);
and U6510 (N_6510,N_6499,N_6445);
nor U6511 (N_6511,N_6426,N_6397);
nand U6512 (N_6512,N_6387,N_6458);
or U6513 (N_6513,N_6430,N_6392);
and U6514 (N_6514,N_6396,N_6449);
or U6515 (N_6515,N_6439,N_6417);
nor U6516 (N_6516,N_6443,N_6420);
nand U6517 (N_6517,N_6455,N_6461);
and U6518 (N_6518,N_6414,N_6473);
or U6519 (N_6519,N_6383,N_6429);
nand U6520 (N_6520,N_6408,N_6379);
or U6521 (N_6521,N_6448,N_6482);
and U6522 (N_6522,N_6451,N_6465);
and U6523 (N_6523,N_6433,N_6484);
nand U6524 (N_6524,N_6390,N_6425);
and U6525 (N_6525,N_6400,N_6488);
nor U6526 (N_6526,N_6467,N_6459);
nor U6527 (N_6527,N_6492,N_6469);
and U6528 (N_6528,N_6386,N_6494);
and U6529 (N_6529,N_6447,N_6438);
xnor U6530 (N_6530,N_6446,N_6435);
and U6531 (N_6531,N_6395,N_6454);
and U6532 (N_6532,N_6464,N_6486);
nor U6533 (N_6533,N_6413,N_6498);
nand U6534 (N_6534,N_6380,N_6478);
nand U6535 (N_6535,N_6419,N_6431);
and U6536 (N_6536,N_6416,N_6406);
and U6537 (N_6537,N_6381,N_6410);
and U6538 (N_6538,N_6489,N_6412);
nor U6539 (N_6539,N_6432,N_6428);
xnor U6540 (N_6540,N_6457,N_6391);
or U6541 (N_6541,N_6415,N_6437);
nor U6542 (N_6542,N_6422,N_6495);
or U6543 (N_6543,N_6475,N_6441);
xor U6544 (N_6544,N_6398,N_6377);
and U6545 (N_6545,N_6479,N_6407);
or U6546 (N_6546,N_6487,N_6421);
and U6547 (N_6547,N_6382,N_6453);
and U6548 (N_6548,N_6404,N_6440);
and U6549 (N_6549,N_6393,N_6442);
and U6550 (N_6550,N_6405,N_6468);
or U6551 (N_6551,N_6476,N_6394);
or U6552 (N_6552,N_6491,N_6497);
and U6553 (N_6553,N_6403,N_6389);
nand U6554 (N_6554,N_6418,N_6399);
or U6555 (N_6555,N_6427,N_6376);
nand U6556 (N_6556,N_6424,N_6472);
or U6557 (N_6557,N_6466,N_6471);
or U6558 (N_6558,N_6493,N_6411);
nor U6559 (N_6559,N_6460,N_6463);
nand U6560 (N_6560,N_6444,N_6462);
nand U6561 (N_6561,N_6452,N_6456);
xnor U6562 (N_6562,N_6470,N_6439);
nand U6563 (N_6563,N_6483,N_6382);
and U6564 (N_6564,N_6421,N_6404);
nor U6565 (N_6565,N_6448,N_6437);
and U6566 (N_6566,N_6386,N_6488);
nand U6567 (N_6567,N_6381,N_6478);
or U6568 (N_6568,N_6443,N_6422);
nand U6569 (N_6569,N_6482,N_6412);
nand U6570 (N_6570,N_6474,N_6467);
xnor U6571 (N_6571,N_6390,N_6454);
nor U6572 (N_6572,N_6408,N_6494);
nor U6573 (N_6573,N_6447,N_6423);
nor U6574 (N_6574,N_6442,N_6417);
or U6575 (N_6575,N_6472,N_6431);
xor U6576 (N_6576,N_6445,N_6386);
nand U6577 (N_6577,N_6443,N_6415);
and U6578 (N_6578,N_6468,N_6459);
and U6579 (N_6579,N_6492,N_6399);
xnor U6580 (N_6580,N_6448,N_6447);
nand U6581 (N_6581,N_6470,N_6384);
or U6582 (N_6582,N_6457,N_6460);
or U6583 (N_6583,N_6401,N_6490);
nand U6584 (N_6584,N_6488,N_6443);
and U6585 (N_6585,N_6431,N_6478);
or U6586 (N_6586,N_6445,N_6424);
nand U6587 (N_6587,N_6442,N_6482);
or U6588 (N_6588,N_6416,N_6418);
nand U6589 (N_6589,N_6497,N_6484);
or U6590 (N_6590,N_6463,N_6414);
and U6591 (N_6591,N_6453,N_6485);
nor U6592 (N_6592,N_6402,N_6408);
and U6593 (N_6593,N_6428,N_6486);
xnor U6594 (N_6594,N_6462,N_6441);
and U6595 (N_6595,N_6406,N_6427);
and U6596 (N_6596,N_6375,N_6451);
nor U6597 (N_6597,N_6426,N_6377);
or U6598 (N_6598,N_6499,N_6456);
xnor U6599 (N_6599,N_6477,N_6495);
nor U6600 (N_6600,N_6420,N_6421);
or U6601 (N_6601,N_6397,N_6420);
and U6602 (N_6602,N_6439,N_6445);
and U6603 (N_6603,N_6491,N_6435);
and U6604 (N_6604,N_6496,N_6459);
and U6605 (N_6605,N_6451,N_6478);
or U6606 (N_6606,N_6420,N_6449);
or U6607 (N_6607,N_6485,N_6436);
or U6608 (N_6608,N_6411,N_6491);
nor U6609 (N_6609,N_6421,N_6446);
xor U6610 (N_6610,N_6479,N_6485);
and U6611 (N_6611,N_6390,N_6401);
nand U6612 (N_6612,N_6407,N_6413);
xnor U6613 (N_6613,N_6478,N_6387);
nand U6614 (N_6614,N_6395,N_6493);
nand U6615 (N_6615,N_6454,N_6409);
xor U6616 (N_6616,N_6384,N_6426);
nor U6617 (N_6617,N_6457,N_6465);
xnor U6618 (N_6618,N_6436,N_6413);
or U6619 (N_6619,N_6421,N_6408);
nor U6620 (N_6620,N_6448,N_6391);
nor U6621 (N_6621,N_6495,N_6418);
nand U6622 (N_6622,N_6472,N_6465);
and U6623 (N_6623,N_6484,N_6421);
nor U6624 (N_6624,N_6386,N_6427);
nand U6625 (N_6625,N_6547,N_6553);
nor U6626 (N_6626,N_6533,N_6516);
or U6627 (N_6627,N_6562,N_6605);
or U6628 (N_6628,N_6524,N_6592);
and U6629 (N_6629,N_6612,N_6613);
nor U6630 (N_6630,N_6567,N_6578);
or U6631 (N_6631,N_6510,N_6502);
or U6632 (N_6632,N_6585,N_6616);
nand U6633 (N_6633,N_6604,N_6596);
or U6634 (N_6634,N_6588,N_6581);
nor U6635 (N_6635,N_6580,N_6610);
or U6636 (N_6636,N_6545,N_6526);
and U6637 (N_6637,N_6563,N_6621);
nand U6638 (N_6638,N_6505,N_6539);
and U6639 (N_6639,N_6538,N_6556);
nand U6640 (N_6640,N_6515,N_6517);
nand U6641 (N_6641,N_6622,N_6614);
or U6642 (N_6642,N_6531,N_6608);
nand U6643 (N_6643,N_6541,N_6529);
nor U6644 (N_6644,N_6518,N_6606);
nand U6645 (N_6645,N_6551,N_6532);
nand U6646 (N_6646,N_6591,N_6575);
nand U6647 (N_6647,N_6561,N_6600);
nand U6648 (N_6648,N_6564,N_6570);
and U6649 (N_6649,N_6530,N_6560);
nor U6650 (N_6650,N_6589,N_6597);
nand U6651 (N_6651,N_6595,N_6572);
or U6652 (N_6652,N_6542,N_6579);
nand U6653 (N_6653,N_6619,N_6593);
nor U6654 (N_6654,N_6500,N_6558);
nor U6655 (N_6655,N_6624,N_6513);
nand U6656 (N_6656,N_6590,N_6543);
or U6657 (N_6657,N_6512,N_6501);
and U6658 (N_6658,N_6576,N_6523);
nor U6659 (N_6659,N_6611,N_6536);
or U6660 (N_6660,N_6594,N_6603);
and U6661 (N_6661,N_6520,N_6617);
nand U6662 (N_6662,N_6537,N_6557);
nor U6663 (N_6663,N_6514,N_6615);
or U6664 (N_6664,N_6574,N_6527);
and U6665 (N_6665,N_6544,N_6620);
and U6666 (N_6666,N_6528,N_6507);
or U6667 (N_6667,N_6586,N_6555);
nor U6668 (N_6668,N_6511,N_6522);
nand U6669 (N_6669,N_6552,N_6508);
and U6670 (N_6670,N_6569,N_6550);
xnor U6671 (N_6671,N_6546,N_6568);
nand U6672 (N_6672,N_6503,N_6577);
and U6673 (N_6673,N_6583,N_6548);
nand U6674 (N_6674,N_6504,N_6582);
and U6675 (N_6675,N_6559,N_6598);
nor U6676 (N_6676,N_6540,N_6554);
nor U6677 (N_6677,N_6525,N_6609);
or U6678 (N_6678,N_6599,N_6623);
nor U6679 (N_6679,N_6519,N_6534);
or U6680 (N_6680,N_6587,N_6565);
xnor U6681 (N_6681,N_6566,N_6618);
or U6682 (N_6682,N_6607,N_6521);
nand U6683 (N_6683,N_6549,N_6584);
xnor U6684 (N_6684,N_6573,N_6509);
nor U6685 (N_6685,N_6506,N_6571);
or U6686 (N_6686,N_6535,N_6602);
and U6687 (N_6687,N_6601,N_6603);
or U6688 (N_6688,N_6504,N_6528);
nor U6689 (N_6689,N_6547,N_6568);
and U6690 (N_6690,N_6546,N_6622);
nor U6691 (N_6691,N_6534,N_6547);
xor U6692 (N_6692,N_6582,N_6598);
nand U6693 (N_6693,N_6600,N_6605);
nor U6694 (N_6694,N_6592,N_6591);
nor U6695 (N_6695,N_6573,N_6566);
nand U6696 (N_6696,N_6531,N_6533);
or U6697 (N_6697,N_6544,N_6568);
nand U6698 (N_6698,N_6558,N_6597);
nand U6699 (N_6699,N_6539,N_6524);
or U6700 (N_6700,N_6617,N_6623);
or U6701 (N_6701,N_6623,N_6506);
nand U6702 (N_6702,N_6556,N_6560);
and U6703 (N_6703,N_6612,N_6588);
nand U6704 (N_6704,N_6592,N_6560);
and U6705 (N_6705,N_6585,N_6571);
or U6706 (N_6706,N_6524,N_6603);
nor U6707 (N_6707,N_6551,N_6624);
and U6708 (N_6708,N_6536,N_6592);
or U6709 (N_6709,N_6587,N_6563);
nor U6710 (N_6710,N_6538,N_6521);
and U6711 (N_6711,N_6516,N_6576);
or U6712 (N_6712,N_6533,N_6549);
nand U6713 (N_6713,N_6524,N_6506);
nand U6714 (N_6714,N_6514,N_6565);
and U6715 (N_6715,N_6579,N_6621);
nand U6716 (N_6716,N_6525,N_6511);
nor U6717 (N_6717,N_6572,N_6618);
nor U6718 (N_6718,N_6542,N_6590);
nor U6719 (N_6719,N_6582,N_6624);
nand U6720 (N_6720,N_6611,N_6618);
nor U6721 (N_6721,N_6595,N_6507);
or U6722 (N_6722,N_6563,N_6546);
nand U6723 (N_6723,N_6592,N_6594);
nand U6724 (N_6724,N_6554,N_6568);
or U6725 (N_6725,N_6612,N_6502);
nand U6726 (N_6726,N_6574,N_6559);
nor U6727 (N_6727,N_6561,N_6595);
or U6728 (N_6728,N_6512,N_6616);
or U6729 (N_6729,N_6601,N_6616);
nor U6730 (N_6730,N_6602,N_6568);
and U6731 (N_6731,N_6602,N_6596);
or U6732 (N_6732,N_6571,N_6521);
xor U6733 (N_6733,N_6540,N_6552);
nor U6734 (N_6734,N_6526,N_6596);
or U6735 (N_6735,N_6535,N_6538);
or U6736 (N_6736,N_6569,N_6558);
and U6737 (N_6737,N_6546,N_6623);
or U6738 (N_6738,N_6581,N_6526);
nor U6739 (N_6739,N_6610,N_6591);
nor U6740 (N_6740,N_6558,N_6549);
or U6741 (N_6741,N_6532,N_6510);
and U6742 (N_6742,N_6579,N_6546);
nor U6743 (N_6743,N_6586,N_6522);
or U6744 (N_6744,N_6534,N_6557);
nor U6745 (N_6745,N_6592,N_6537);
and U6746 (N_6746,N_6578,N_6536);
nand U6747 (N_6747,N_6572,N_6527);
and U6748 (N_6748,N_6537,N_6532);
or U6749 (N_6749,N_6555,N_6614);
and U6750 (N_6750,N_6653,N_6704);
and U6751 (N_6751,N_6724,N_6721);
or U6752 (N_6752,N_6627,N_6714);
xnor U6753 (N_6753,N_6715,N_6700);
and U6754 (N_6754,N_6668,N_6719);
nor U6755 (N_6755,N_6744,N_6691);
nand U6756 (N_6756,N_6686,N_6655);
nand U6757 (N_6757,N_6687,N_6651);
and U6758 (N_6758,N_6736,N_6711);
xnor U6759 (N_6759,N_6663,N_6664);
nand U6760 (N_6760,N_6732,N_6746);
nand U6761 (N_6761,N_6693,N_6670);
nor U6762 (N_6762,N_6669,N_6625);
nor U6763 (N_6763,N_6696,N_6679);
nor U6764 (N_6764,N_6705,N_6713);
nor U6765 (N_6765,N_6685,N_6649);
or U6766 (N_6766,N_6688,N_6676);
or U6767 (N_6767,N_6647,N_6709);
or U6768 (N_6768,N_6675,N_6698);
nor U6769 (N_6769,N_6712,N_6660);
nor U6770 (N_6770,N_6629,N_6661);
nor U6771 (N_6771,N_6692,N_6654);
nand U6772 (N_6772,N_6718,N_6717);
nand U6773 (N_6773,N_6730,N_6729);
nand U6774 (N_6774,N_6684,N_6652);
and U6775 (N_6775,N_6681,N_6722);
and U6776 (N_6776,N_6690,N_6701);
nor U6777 (N_6777,N_6699,N_6633);
or U6778 (N_6778,N_6674,N_6638);
nand U6779 (N_6779,N_6642,N_6644);
or U6780 (N_6780,N_6657,N_6737);
or U6781 (N_6781,N_6659,N_6689);
xnor U6782 (N_6782,N_6749,N_6645);
or U6783 (N_6783,N_6726,N_6695);
xnor U6784 (N_6784,N_6636,N_6665);
and U6785 (N_6785,N_6703,N_6725);
nor U6786 (N_6786,N_6667,N_6694);
nand U6787 (N_6787,N_6648,N_6742);
nand U6788 (N_6788,N_6716,N_6631);
xor U6789 (N_6789,N_6702,N_6632);
nand U6790 (N_6790,N_6735,N_6743);
nor U6791 (N_6791,N_6662,N_6628);
nand U6792 (N_6792,N_6723,N_6682);
nor U6793 (N_6793,N_6643,N_6677);
xor U6794 (N_6794,N_6683,N_6671);
and U6795 (N_6795,N_6658,N_6640);
nand U6796 (N_6796,N_6678,N_6728);
nor U6797 (N_6797,N_6708,N_6740);
nor U6798 (N_6798,N_6641,N_6666);
nor U6799 (N_6799,N_6748,N_6706);
and U6800 (N_6800,N_6639,N_6739);
and U6801 (N_6801,N_6635,N_6680);
or U6802 (N_6802,N_6646,N_6710);
xor U6803 (N_6803,N_6637,N_6747);
and U6804 (N_6804,N_6626,N_6656);
nor U6805 (N_6805,N_6733,N_6727);
nand U6806 (N_6806,N_6741,N_6650);
nor U6807 (N_6807,N_6707,N_6731);
or U6808 (N_6808,N_6720,N_6738);
nor U6809 (N_6809,N_6673,N_6745);
nor U6810 (N_6810,N_6630,N_6734);
or U6811 (N_6811,N_6672,N_6634);
nor U6812 (N_6812,N_6697,N_6693);
nand U6813 (N_6813,N_6701,N_6646);
nand U6814 (N_6814,N_6736,N_6634);
and U6815 (N_6815,N_6685,N_6666);
xnor U6816 (N_6816,N_6643,N_6707);
or U6817 (N_6817,N_6639,N_6745);
or U6818 (N_6818,N_6715,N_6710);
and U6819 (N_6819,N_6628,N_6642);
nor U6820 (N_6820,N_6663,N_6649);
nor U6821 (N_6821,N_6654,N_6667);
nand U6822 (N_6822,N_6642,N_6716);
or U6823 (N_6823,N_6671,N_6641);
and U6824 (N_6824,N_6625,N_6644);
nor U6825 (N_6825,N_6642,N_6717);
or U6826 (N_6826,N_6640,N_6726);
or U6827 (N_6827,N_6639,N_6703);
nor U6828 (N_6828,N_6693,N_6681);
or U6829 (N_6829,N_6649,N_6700);
nor U6830 (N_6830,N_6668,N_6683);
and U6831 (N_6831,N_6697,N_6736);
nor U6832 (N_6832,N_6642,N_6701);
or U6833 (N_6833,N_6682,N_6741);
or U6834 (N_6834,N_6650,N_6732);
and U6835 (N_6835,N_6715,N_6640);
or U6836 (N_6836,N_6667,N_6628);
or U6837 (N_6837,N_6691,N_6702);
xnor U6838 (N_6838,N_6735,N_6640);
nand U6839 (N_6839,N_6729,N_6653);
or U6840 (N_6840,N_6717,N_6667);
and U6841 (N_6841,N_6643,N_6701);
or U6842 (N_6842,N_6696,N_6723);
nor U6843 (N_6843,N_6705,N_6668);
nand U6844 (N_6844,N_6632,N_6657);
nand U6845 (N_6845,N_6680,N_6637);
nand U6846 (N_6846,N_6720,N_6694);
nand U6847 (N_6847,N_6653,N_6644);
or U6848 (N_6848,N_6658,N_6724);
nor U6849 (N_6849,N_6675,N_6649);
or U6850 (N_6850,N_6708,N_6714);
or U6851 (N_6851,N_6722,N_6710);
or U6852 (N_6852,N_6629,N_6679);
and U6853 (N_6853,N_6719,N_6656);
and U6854 (N_6854,N_6729,N_6742);
nor U6855 (N_6855,N_6638,N_6706);
or U6856 (N_6856,N_6694,N_6703);
nand U6857 (N_6857,N_6666,N_6654);
xor U6858 (N_6858,N_6701,N_6705);
and U6859 (N_6859,N_6626,N_6711);
nand U6860 (N_6860,N_6695,N_6642);
xor U6861 (N_6861,N_6701,N_6722);
nor U6862 (N_6862,N_6661,N_6734);
and U6863 (N_6863,N_6730,N_6654);
or U6864 (N_6864,N_6745,N_6729);
nor U6865 (N_6865,N_6748,N_6737);
nand U6866 (N_6866,N_6721,N_6729);
or U6867 (N_6867,N_6664,N_6639);
or U6868 (N_6868,N_6702,N_6706);
nand U6869 (N_6869,N_6656,N_6744);
nor U6870 (N_6870,N_6722,N_6674);
nand U6871 (N_6871,N_6680,N_6699);
or U6872 (N_6872,N_6660,N_6672);
nor U6873 (N_6873,N_6627,N_6740);
nor U6874 (N_6874,N_6640,N_6718);
nor U6875 (N_6875,N_6771,N_6853);
nor U6876 (N_6876,N_6756,N_6812);
nand U6877 (N_6877,N_6810,N_6807);
xor U6878 (N_6878,N_6844,N_6786);
nand U6879 (N_6879,N_6798,N_6848);
nand U6880 (N_6880,N_6790,N_6849);
or U6881 (N_6881,N_6872,N_6856);
and U6882 (N_6882,N_6871,N_6837);
nand U6883 (N_6883,N_6847,N_6860);
and U6884 (N_6884,N_6787,N_6760);
nand U6885 (N_6885,N_6797,N_6809);
and U6886 (N_6886,N_6846,N_6829);
nor U6887 (N_6887,N_6818,N_6781);
xor U6888 (N_6888,N_6795,N_6811);
or U6889 (N_6889,N_6834,N_6855);
nor U6890 (N_6890,N_6841,N_6751);
nor U6891 (N_6891,N_6789,N_6803);
nor U6892 (N_6892,N_6769,N_6838);
nor U6893 (N_6893,N_6788,N_6765);
nor U6894 (N_6894,N_6822,N_6801);
nor U6895 (N_6895,N_6868,N_6861);
nor U6896 (N_6896,N_6782,N_6842);
or U6897 (N_6897,N_6815,N_6859);
and U6898 (N_6898,N_6796,N_6831);
nand U6899 (N_6899,N_6773,N_6770);
nor U6900 (N_6900,N_6759,N_6823);
and U6901 (N_6901,N_6791,N_6852);
nor U6902 (N_6902,N_6779,N_6830);
or U6903 (N_6903,N_6850,N_6863);
and U6904 (N_6904,N_6775,N_6780);
nor U6905 (N_6905,N_6862,N_6778);
and U6906 (N_6906,N_6828,N_6814);
nor U6907 (N_6907,N_6794,N_6776);
nor U6908 (N_6908,N_6833,N_6858);
and U6909 (N_6909,N_6799,N_6820);
nor U6910 (N_6910,N_6864,N_6819);
or U6911 (N_6911,N_6845,N_6869);
nand U6912 (N_6912,N_6826,N_6774);
nand U6913 (N_6913,N_6761,N_6866);
nor U6914 (N_6914,N_6808,N_6806);
and U6915 (N_6915,N_6825,N_6817);
nand U6916 (N_6916,N_6758,N_6804);
or U6917 (N_6917,N_6865,N_6750);
and U6918 (N_6918,N_6827,N_6802);
and U6919 (N_6919,N_6763,N_6873);
nand U6920 (N_6920,N_6854,N_6768);
and U6921 (N_6921,N_6755,N_6870);
nand U6922 (N_6922,N_6764,N_6793);
nand U6923 (N_6923,N_6805,N_6783);
nand U6924 (N_6924,N_6836,N_6785);
nand U6925 (N_6925,N_6874,N_6816);
nand U6926 (N_6926,N_6752,N_6821);
or U6927 (N_6927,N_6824,N_6857);
and U6928 (N_6928,N_6767,N_6800);
xor U6929 (N_6929,N_6757,N_6777);
or U6930 (N_6930,N_6784,N_6867);
nand U6931 (N_6931,N_6772,N_6792);
xnor U6932 (N_6932,N_6762,N_6839);
nand U6933 (N_6933,N_6840,N_6843);
nor U6934 (N_6934,N_6851,N_6754);
and U6935 (N_6935,N_6832,N_6753);
and U6936 (N_6936,N_6766,N_6813);
or U6937 (N_6937,N_6835,N_6829);
or U6938 (N_6938,N_6855,N_6810);
nor U6939 (N_6939,N_6859,N_6852);
and U6940 (N_6940,N_6804,N_6855);
or U6941 (N_6941,N_6838,N_6785);
nand U6942 (N_6942,N_6859,N_6866);
nand U6943 (N_6943,N_6837,N_6753);
and U6944 (N_6944,N_6865,N_6814);
or U6945 (N_6945,N_6841,N_6873);
xnor U6946 (N_6946,N_6764,N_6760);
nor U6947 (N_6947,N_6844,N_6801);
xnor U6948 (N_6948,N_6755,N_6862);
nand U6949 (N_6949,N_6816,N_6830);
nor U6950 (N_6950,N_6826,N_6850);
or U6951 (N_6951,N_6842,N_6797);
or U6952 (N_6952,N_6814,N_6872);
and U6953 (N_6953,N_6869,N_6822);
or U6954 (N_6954,N_6794,N_6805);
nor U6955 (N_6955,N_6813,N_6839);
nor U6956 (N_6956,N_6805,N_6837);
or U6957 (N_6957,N_6793,N_6751);
nor U6958 (N_6958,N_6750,N_6810);
and U6959 (N_6959,N_6856,N_6821);
and U6960 (N_6960,N_6755,N_6770);
nor U6961 (N_6961,N_6813,N_6810);
or U6962 (N_6962,N_6837,N_6844);
or U6963 (N_6963,N_6763,N_6818);
or U6964 (N_6964,N_6851,N_6856);
or U6965 (N_6965,N_6751,N_6840);
and U6966 (N_6966,N_6756,N_6841);
nor U6967 (N_6967,N_6814,N_6822);
or U6968 (N_6968,N_6834,N_6810);
xnor U6969 (N_6969,N_6777,N_6828);
nand U6970 (N_6970,N_6826,N_6786);
nand U6971 (N_6971,N_6844,N_6873);
nand U6972 (N_6972,N_6782,N_6807);
and U6973 (N_6973,N_6752,N_6766);
and U6974 (N_6974,N_6854,N_6800);
nor U6975 (N_6975,N_6858,N_6764);
and U6976 (N_6976,N_6751,N_6847);
and U6977 (N_6977,N_6765,N_6799);
nand U6978 (N_6978,N_6750,N_6874);
or U6979 (N_6979,N_6827,N_6782);
xnor U6980 (N_6980,N_6772,N_6819);
or U6981 (N_6981,N_6872,N_6808);
nor U6982 (N_6982,N_6820,N_6830);
nand U6983 (N_6983,N_6851,N_6874);
and U6984 (N_6984,N_6829,N_6798);
or U6985 (N_6985,N_6808,N_6823);
xor U6986 (N_6986,N_6775,N_6823);
nand U6987 (N_6987,N_6841,N_6816);
and U6988 (N_6988,N_6816,N_6814);
nand U6989 (N_6989,N_6849,N_6823);
and U6990 (N_6990,N_6802,N_6821);
nor U6991 (N_6991,N_6852,N_6772);
or U6992 (N_6992,N_6874,N_6868);
nand U6993 (N_6993,N_6754,N_6841);
nand U6994 (N_6994,N_6754,N_6815);
and U6995 (N_6995,N_6818,N_6854);
nand U6996 (N_6996,N_6859,N_6809);
nand U6997 (N_6997,N_6868,N_6823);
and U6998 (N_6998,N_6855,N_6854);
or U6999 (N_6999,N_6752,N_6794);
nor U7000 (N_7000,N_6953,N_6932);
nand U7001 (N_7001,N_6876,N_6975);
or U7002 (N_7002,N_6985,N_6963);
nand U7003 (N_7003,N_6915,N_6998);
or U7004 (N_7004,N_6983,N_6904);
nand U7005 (N_7005,N_6965,N_6935);
and U7006 (N_7006,N_6942,N_6883);
nand U7007 (N_7007,N_6956,N_6955);
or U7008 (N_7008,N_6991,N_6971);
xor U7009 (N_7009,N_6972,N_6996);
nand U7010 (N_7010,N_6959,N_6990);
and U7011 (N_7011,N_6978,N_6969);
and U7012 (N_7012,N_6882,N_6879);
nor U7013 (N_7013,N_6892,N_6887);
nor U7014 (N_7014,N_6910,N_6896);
nor U7015 (N_7015,N_6938,N_6957);
nand U7016 (N_7016,N_6878,N_6908);
or U7017 (N_7017,N_6886,N_6954);
xnor U7018 (N_7018,N_6970,N_6977);
nand U7019 (N_7019,N_6937,N_6961);
nor U7020 (N_7020,N_6951,N_6987);
nand U7021 (N_7021,N_6894,N_6888);
or U7022 (N_7022,N_6907,N_6993);
xnor U7023 (N_7023,N_6921,N_6960);
or U7024 (N_7024,N_6901,N_6931);
nand U7025 (N_7025,N_6939,N_6919);
or U7026 (N_7026,N_6881,N_6974);
or U7027 (N_7027,N_6999,N_6893);
and U7028 (N_7028,N_6944,N_6925);
nand U7029 (N_7029,N_6988,N_6913);
or U7030 (N_7030,N_6895,N_6890);
nand U7031 (N_7031,N_6958,N_6980);
xor U7032 (N_7032,N_6967,N_6885);
or U7033 (N_7033,N_6926,N_6945);
nor U7034 (N_7034,N_6900,N_6943);
or U7035 (N_7035,N_6941,N_6929);
or U7036 (N_7036,N_6947,N_6995);
nand U7037 (N_7037,N_6949,N_6986);
and U7038 (N_7038,N_6916,N_6880);
and U7039 (N_7039,N_6903,N_6934);
or U7040 (N_7040,N_6912,N_6898);
or U7041 (N_7041,N_6906,N_6973);
and U7042 (N_7042,N_6884,N_6936);
or U7043 (N_7043,N_6889,N_6984);
nor U7044 (N_7044,N_6920,N_6902);
nor U7045 (N_7045,N_6930,N_6875);
and U7046 (N_7046,N_6952,N_6918);
or U7047 (N_7047,N_6927,N_6994);
and U7048 (N_7048,N_6992,N_6923);
and U7049 (N_7049,N_6924,N_6976);
xor U7050 (N_7050,N_6940,N_6946);
and U7051 (N_7051,N_6968,N_6989);
nor U7052 (N_7052,N_6891,N_6982);
or U7053 (N_7053,N_6928,N_6914);
nand U7054 (N_7054,N_6950,N_6917);
nand U7055 (N_7055,N_6997,N_6911);
or U7056 (N_7056,N_6979,N_6964);
nand U7057 (N_7057,N_6877,N_6905);
and U7058 (N_7058,N_6962,N_6981);
and U7059 (N_7059,N_6909,N_6933);
or U7060 (N_7060,N_6966,N_6897);
nand U7061 (N_7061,N_6922,N_6948);
or U7062 (N_7062,N_6899,N_6986);
and U7063 (N_7063,N_6951,N_6903);
xor U7064 (N_7064,N_6881,N_6982);
or U7065 (N_7065,N_6944,N_6911);
nor U7066 (N_7066,N_6901,N_6894);
and U7067 (N_7067,N_6893,N_6875);
and U7068 (N_7068,N_6906,N_6942);
xor U7069 (N_7069,N_6946,N_6922);
or U7070 (N_7070,N_6888,N_6887);
or U7071 (N_7071,N_6980,N_6984);
and U7072 (N_7072,N_6907,N_6908);
nor U7073 (N_7073,N_6968,N_6916);
and U7074 (N_7074,N_6927,N_6896);
nand U7075 (N_7075,N_6978,N_6886);
and U7076 (N_7076,N_6983,N_6985);
or U7077 (N_7077,N_6900,N_6904);
nand U7078 (N_7078,N_6879,N_6993);
nor U7079 (N_7079,N_6916,N_6903);
nand U7080 (N_7080,N_6912,N_6972);
and U7081 (N_7081,N_6894,N_6877);
nor U7082 (N_7082,N_6978,N_6972);
nor U7083 (N_7083,N_6956,N_6957);
nor U7084 (N_7084,N_6909,N_6961);
nor U7085 (N_7085,N_6883,N_6956);
nor U7086 (N_7086,N_6902,N_6952);
nand U7087 (N_7087,N_6890,N_6915);
or U7088 (N_7088,N_6989,N_6985);
and U7089 (N_7089,N_6986,N_6944);
nor U7090 (N_7090,N_6905,N_6975);
or U7091 (N_7091,N_6960,N_6894);
nor U7092 (N_7092,N_6954,N_6970);
or U7093 (N_7093,N_6954,N_6878);
nand U7094 (N_7094,N_6999,N_6883);
nand U7095 (N_7095,N_6955,N_6925);
nand U7096 (N_7096,N_6976,N_6889);
nand U7097 (N_7097,N_6962,N_6918);
nand U7098 (N_7098,N_6879,N_6939);
and U7099 (N_7099,N_6955,N_6946);
or U7100 (N_7100,N_6928,N_6887);
xor U7101 (N_7101,N_6952,N_6898);
and U7102 (N_7102,N_6899,N_6879);
and U7103 (N_7103,N_6999,N_6971);
nor U7104 (N_7104,N_6982,N_6971);
nand U7105 (N_7105,N_6915,N_6880);
and U7106 (N_7106,N_6926,N_6877);
or U7107 (N_7107,N_6958,N_6903);
or U7108 (N_7108,N_6898,N_6966);
and U7109 (N_7109,N_6945,N_6909);
xor U7110 (N_7110,N_6896,N_6983);
or U7111 (N_7111,N_6947,N_6969);
nand U7112 (N_7112,N_6945,N_6959);
or U7113 (N_7113,N_6979,N_6930);
xor U7114 (N_7114,N_6904,N_6997);
xor U7115 (N_7115,N_6990,N_6945);
nor U7116 (N_7116,N_6985,N_6957);
nand U7117 (N_7117,N_6997,N_6890);
nand U7118 (N_7118,N_6961,N_6974);
nor U7119 (N_7119,N_6953,N_6982);
nand U7120 (N_7120,N_6896,N_6999);
nand U7121 (N_7121,N_6924,N_6968);
and U7122 (N_7122,N_6970,N_6926);
nand U7123 (N_7123,N_6916,N_6998);
nand U7124 (N_7124,N_6896,N_6987);
nand U7125 (N_7125,N_7042,N_7003);
or U7126 (N_7126,N_7087,N_7033);
xnor U7127 (N_7127,N_7001,N_7059);
or U7128 (N_7128,N_7072,N_7050);
nand U7129 (N_7129,N_7104,N_7077);
and U7130 (N_7130,N_7119,N_7100);
and U7131 (N_7131,N_7036,N_7099);
and U7132 (N_7132,N_7081,N_7020);
and U7133 (N_7133,N_7017,N_7067);
nand U7134 (N_7134,N_7041,N_7015);
nand U7135 (N_7135,N_7097,N_7117);
or U7136 (N_7136,N_7108,N_7115);
nor U7137 (N_7137,N_7037,N_7044);
or U7138 (N_7138,N_7110,N_7027);
nand U7139 (N_7139,N_7019,N_7073);
and U7140 (N_7140,N_7066,N_7094);
nor U7141 (N_7141,N_7076,N_7064);
nand U7142 (N_7142,N_7048,N_7032);
nor U7143 (N_7143,N_7011,N_7046);
and U7144 (N_7144,N_7079,N_7025);
and U7145 (N_7145,N_7089,N_7085);
and U7146 (N_7146,N_7047,N_7012);
nor U7147 (N_7147,N_7088,N_7004);
and U7148 (N_7148,N_7091,N_7061);
nor U7149 (N_7149,N_7121,N_7038);
and U7150 (N_7150,N_7086,N_7028);
nand U7151 (N_7151,N_7009,N_7008);
and U7152 (N_7152,N_7060,N_7093);
and U7153 (N_7153,N_7056,N_7051);
or U7154 (N_7154,N_7123,N_7084);
or U7155 (N_7155,N_7018,N_7049);
nand U7156 (N_7156,N_7103,N_7071);
nand U7157 (N_7157,N_7078,N_7029);
nor U7158 (N_7158,N_7000,N_7023);
and U7159 (N_7159,N_7070,N_7114);
nand U7160 (N_7160,N_7010,N_7022);
and U7161 (N_7161,N_7069,N_7040);
nand U7162 (N_7162,N_7106,N_7120);
xor U7163 (N_7163,N_7095,N_7052);
nand U7164 (N_7164,N_7007,N_7102);
or U7165 (N_7165,N_7080,N_7035);
xnor U7166 (N_7166,N_7045,N_7043);
nand U7167 (N_7167,N_7068,N_7075);
or U7168 (N_7168,N_7057,N_7024);
xnor U7169 (N_7169,N_7101,N_7014);
nand U7170 (N_7170,N_7098,N_7113);
or U7171 (N_7171,N_7062,N_7058);
or U7172 (N_7172,N_7031,N_7124);
and U7173 (N_7173,N_7116,N_7107);
nand U7174 (N_7174,N_7013,N_7109);
or U7175 (N_7175,N_7054,N_7090);
and U7176 (N_7176,N_7026,N_7082);
and U7177 (N_7177,N_7006,N_7065);
nand U7178 (N_7178,N_7039,N_7016);
and U7179 (N_7179,N_7002,N_7118);
nand U7180 (N_7180,N_7030,N_7122);
or U7181 (N_7181,N_7055,N_7034);
nor U7182 (N_7182,N_7074,N_7021);
or U7183 (N_7183,N_7005,N_7112);
nand U7184 (N_7184,N_7092,N_7111);
or U7185 (N_7185,N_7063,N_7105);
and U7186 (N_7186,N_7096,N_7083);
and U7187 (N_7187,N_7053,N_7049);
nand U7188 (N_7188,N_7055,N_7079);
and U7189 (N_7189,N_7064,N_7008);
nand U7190 (N_7190,N_7052,N_7077);
or U7191 (N_7191,N_7020,N_7070);
and U7192 (N_7192,N_7002,N_7051);
nand U7193 (N_7193,N_7025,N_7097);
or U7194 (N_7194,N_7061,N_7013);
nor U7195 (N_7195,N_7121,N_7064);
xor U7196 (N_7196,N_7106,N_7032);
nand U7197 (N_7197,N_7054,N_7085);
and U7198 (N_7198,N_7013,N_7113);
nor U7199 (N_7199,N_7008,N_7085);
nand U7200 (N_7200,N_7019,N_7098);
nand U7201 (N_7201,N_7038,N_7087);
or U7202 (N_7202,N_7095,N_7104);
nand U7203 (N_7203,N_7088,N_7084);
xnor U7204 (N_7204,N_7019,N_7030);
nor U7205 (N_7205,N_7122,N_7051);
xnor U7206 (N_7206,N_7069,N_7014);
or U7207 (N_7207,N_7121,N_7102);
and U7208 (N_7208,N_7092,N_7089);
nand U7209 (N_7209,N_7025,N_7109);
or U7210 (N_7210,N_7031,N_7022);
and U7211 (N_7211,N_7098,N_7003);
xor U7212 (N_7212,N_7094,N_7045);
nor U7213 (N_7213,N_7120,N_7043);
nor U7214 (N_7214,N_7097,N_7050);
nand U7215 (N_7215,N_7007,N_7001);
and U7216 (N_7216,N_7108,N_7041);
nand U7217 (N_7217,N_7121,N_7058);
nand U7218 (N_7218,N_7061,N_7080);
and U7219 (N_7219,N_7109,N_7028);
nand U7220 (N_7220,N_7078,N_7018);
or U7221 (N_7221,N_7040,N_7060);
or U7222 (N_7222,N_7074,N_7116);
and U7223 (N_7223,N_7013,N_7027);
and U7224 (N_7224,N_7007,N_7098);
nand U7225 (N_7225,N_7117,N_7057);
nor U7226 (N_7226,N_7028,N_7115);
nand U7227 (N_7227,N_7014,N_7120);
xnor U7228 (N_7228,N_7036,N_7063);
nor U7229 (N_7229,N_7088,N_7058);
xor U7230 (N_7230,N_7119,N_7038);
xor U7231 (N_7231,N_7078,N_7071);
or U7232 (N_7232,N_7094,N_7100);
nor U7233 (N_7233,N_7003,N_7104);
and U7234 (N_7234,N_7045,N_7121);
nand U7235 (N_7235,N_7084,N_7005);
nor U7236 (N_7236,N_7044,N_7045);
and U7237 (N_7237,N_7029,N_7006);
nor U7238 (N_7238,N_7024,N_7111);
or U7239 (N_7239,N_7073,N_7014);
and U7240 (N_7240,N_7004,N_7109);
and U7241 (N_7241,N_7084,N_7074);
or U7242 (N_7242,N_7104,N_7103);
nand U7243 (N_7243,N_7120,N_7013);
or U7244 (N_7244,N_7106,N_7117);
nand U7245 (N_7245,N_7019,N_7097);
or U7246 (N_7246,N_7049,N_7031);
nor U7247 (N_7247,N_7043,N_7020);
and U7248 (N_7248,N_7074,N_7079);
nand U7249 (N_7249,N_7109,N_7107);
and U7250 (N_7250,N_7169,N_7135);
and U7251 (N_7251,N_7246,N_7243);
nand U7252 (N_7252,N_7154,N_7183);
xor U7253 (N_7253,N_7210,N_7225);
and U7254 (N_7254,N_7245,N_7140);
and U7255 (N_7255,N_7167,N_7227);
and U7256 (N_7256,N_7223,N_7239);
or U7257 (N_7257,N_7238,N_7205);
nor U7258 (N_7258,N_7193,N_7229);
nand U7259 (N_7259,N_7248,N_7161);
nor U7260 (N_7260,N_7217,N_7208);
or U7261 (N_7261,N_7247,N_7165);
nand U7262 (N_7262,N_7130,N_7236);
nor U7263 (N_7263,N_7241,N_7178);
xnor U7264 (N_7264,N_7197,N_7182);
xor U7265 (N_7265,N_7163,N_7147);
or U7266 (N_7266,N_7173,N_7166);
nand U7267 (N_7267,N_7237,N_7222);
or U7268 (N_7268,N_7171,N_7230);
xnor U7269 (N_7269,N_7196,N_7153);
nand U7270 (N_7270,N_7145,N_7242);
nor U7271 (N_7271,N_7207,N_7187);
and U7272 (N_7272,N_7213,N_7233);
xnor U7273 (N_7273,N_7191,N_7200);
xor U7274 (N_7274,N_7172,N_7249);
or U7275 (N_7275,N_7141,N_7198);
nand U7276 (N_7276,N_7244,N_7221);
and U7277 (N_7277,N_7206,N_7219);
nor U7278 (N_7278,N_7152,N_7159);
or U7279 (N_7279,N_7194,N_7127);
xor U7280 (N_7280,N_7150,N_7190);
xnor U7281 (N_7281,N_7125,N_7204);
and U7282 (N_7282,N_7211,N_7228);
xor U7283 (N_7283,N_7192,N_7136);
or U7284 (N_7284,N_7179,N_7231);
or U7285 (N_7285,N_7160,N_7181);
and U7286 (N_7286,N_7128,N_7224);
or U7287 (N_7287,N_7133,N_7132);
or U7288 (N_7288,N_7201,N_7155);
nand U7289 (N_7289,N_7144,N_7162);
nand U7290 (N_7290,N_7186,N_7203);
or U7291 (N_7291,N_7202,N_7142);
and U7292 (N_7292,N_7134,N_7184);
nand U7293 (N_7293,N_7174,N_7199);
nand U7294 (N_7294,N_7176,N_7180);
nand U7295 (N_7295,N_7148,N_7212);
and U7296 (N_7296,N_7215,N_7177);
and U7297 (N_7297,N_7175,N_7156);
nand U7298 (N_7298,N_7195,N_7226);
nor U7299 (N_7299,N_7209,N_7139);
nor U7300 (N_7300,N_7170,N_7234);
nor U7301 (N_7301,N_7157,N_7240);
or U7302 (N_7302,N_7158,N_7151);
nor U7303 (N_7303,N_7220,N_7143);
nor U7304 (N_7304,N_7235,N_7214);
nor U7305 (N_7305,N_7129,N_7232);
nor U7306 (N_7306,N_7126,N_7216);
and U7307 (N_7307,N_7218,N_7146);
and U7308 (N_7308,N_7137,N_7138);
nand U7309 (N_7309,N_7164,N_7131);
and U7310 (N_7310,N_7185,N_7189);
nand U7311 (N_7311,N_7188,N_7149);
xnor U7312 (N_7312,N_7168,N_7127);
nand U7313 (N_7313,N_7199,N_7233);
nor U7314 (N_7314,N_7196,N_7237);
nand U7315 (N_7315,N_7132,N_7204);
or U7316 (N_7316,N_7164,N_7183);
or U7317 (N_7317,N_7132,N_7207);
nand U7318 (N_7318,N_7190,N_7185);
nor U7319 (N_7319,N_7204,N_7170);
or U7320 (N_7320,N_7181,N_7174);
or U7321 (N_7321,N_7152,N_7157);
xnor U7322 (N_7322,N_7174,N_7222);
nor U7323 (N_7323,N_7193,N_7225);
or U7324 (N_7324,N_7188,N_7183);
or U7325 (N_7325,N_7175,N_7214);
and U7326 (N_7326,N_7233,N_7236);
or U7327 (N_7327,N_7128,N_7148);
nand U7328 (N_7328,N_7158,N_7187);
or U7329 (N_7329,N_7189,N_7146);
nand U7330 (N_7330,N_7245,N_7129);
and U7331 (N_7331,N_7158,N_7204);
and U7332 (N_7332,N_7170,N_7228);
nand U7333 (N_7333,N_7201,N_7203);
xnor U7334 (N_7334,N_7214,N_7188);
nor U7335 (N_7335,N_7164,N_7193);
nand U7336 (N_7336,N_7166,N_7224);
xor U7337 (N_7337,N_7191,N_7153);
nand U7338 (N_7338,N_7184,N_7202);
or U7339 (N_7339,N_7172,N_7163);
nor U7340 (N_7340,N_7186,N_7187);
xnor U7341 (N_7341,N_7144,N_7219);
xnor U7342 (N_7342,N_7235,N_7161);
nor U7343 (N_7343,N_7183,N_7142);
nand U7344 (N_7344,N_7171,N_7128);
or U7345 (N_7345,N_7130,N_7129);
nor U7346 (N_7346,N_7139,N_7181);
or U7347 (N_7347,N_7227,N_7163);
and U7348 (N_7348,N_7174,N_7130);
or U7349 (N_7349,N_7214,N_7156);
nor U7350 (N_7350,N_7192,N_7166);
or U7351 (N_7351,N_7230,N_7184);
or U7352 (N_7352,N_7167,N_7131);
nand U7353 (N_7353,N_7226,N_7154);
nand U7354 (N_7354,N_7187,N_7240);
or U7355 (N_7355,N_7144,N_7185);
nand U7356 (N_7356,N_7240,N_7163);
nand U7357 (N_7357,N_7215,N_7196);
and U7358 (N_7358,N_7175,N_7226);
and U7359 (N_7359,N_7176,N_7239);
nand U7360 (N_7360,N_7199,N_7223);
nor U7361 (N_7361,N_7133,N_7232);
and U7362 (N_7362,N_7182,N_7136);
or U7363 (N_7363,N_7137,N_7220);
nor U7364 (N_7364,N_7221,N_7207);
nor U7365 (N_7365,N_7240,N_7170);
or U7366 (N_7366,N_7169,N_7142);
nor U7367 (N_7367,N_7154,N_7203);
nand U7368 (N_7368,N_7237,N_7161);
nand U7369 (N_7369,N_7135,N_7247);
nand U7370 (N_7370,N_7248,N_7174);
and U7371 (N_7371,N_7180,N_7135);
and U7372 (N_7372,N_7220,N_7201);
and U7373 (N_7373,N_7248,N_7203);
nand U7374 (N_7374,N_7146,N_7170);
or U7375 (N_7375,N_7313,N_7339);
xnor U7376 (N_7376,N_7276,N_7266);
nand U7377 (N_7377,N_7336,N_7306);
or U7378 (N_7378,N_7263,N_7372);
nor U7379 (N_7379,N_7329,N_7291);
and U7380 (N_7380,N_7275,N_7290);
nor U7381 (N_7381,N_7271,N_7315);
or U7382 (N_7382,N_7337,N_7273);
or U7383 (N_7383,N_7333,N_7331);
and U7384 (N_7384,N_7345,N_7314);
or U7385 (N_7385,N_7277,N_7294);
and U7386 (N_7386,N_7360,N_7289);
nand U7387 (N_7387,N_7278,N_7367);
xor U7388 (N_7388,N_7309,N_7264);
or U7389 (N_7389,N_7252,N_7260);
nor U7390 (N_7390,N_7369,N_7303);
nor U7391 (N_7391,N_7304,N_7327);
and U7392 (N_7392,N_7352,N_7310);
nor U7393 (N_7393,N_7284,N_7356);
nand U7394 (N_7394,N_7362,N_7318);
nor U7395 (N_7395,N_7346,N_7351);
nand U7396 (N_7396,N_7259,N_7302);
and U7397 (N_7397,N_7297,N_7355);
nor U7398 (N_7398,N_7341,N_7374);
nand U7399 (N_7399,N_7349,N_7370);
and U7400 (N_7400,N_7300,N_7324);
and U7401 (N_7401,N_7262,N_7296);
nor U7402 (N_7402,N_7272,N_7348);
nor U7403 (N_7403,N_7335,N_7361);
or U7404 (N_7404,N_7330,N_7261);
nand U7405 (N_7405,N_7373,N_7353);
nor U7406 (N_7406,N_7251,N_7254);
nor U7407 (N_7407,N_7342,N_7364);
nand U7408 (N_7408,N_7366,N_7326);
or U7409 (N_7409,N_7256,N_7286);
nor U7410 (N_7410,N_7268,N_7283);
or U7411 (N_7411,N_7267,N_7307);
and U7412 (N_7412,N_7293,N_7371);
nand U7413 (N_7413,N_7354,N_7332);
and U7414 (N_7414,N_7319,N_7298);
and U7415 (N_7415,N_7257,N_7316);
and U7416 (N_7416,N_7350,N_7347);
nor U7417 (N_7417,N_7368,N_7325);
nor U7418 (N_7418,N_7320,N_7321);
and U7419 (N_7419,N_7322,N_7282);
nand U7420 (N_7420,N_7288,N_7281);
nor U7421 (N_7421,N_7308,N_7312);
or U7422 (N_7422,N_7340,N_7280);
or U7423 (N_7423,N_7334,N_7295);
or U7424 (N_7424,N_7328,N_7285);
or U7425 (N_7425,N_7358,N_7323);
nand U7426 (N_7426,N_7270,N_7269);
or U7427 (N_7427,N_7359,N_7338);
or U7428 (N_7428,N_7287,N_7292);
and U7429 (N_7429,N_7301,N_7250);
nand U7430 (N_7430,N_7258,N_7311);
nand U7431 (N_7431,N_7363,N_7265);
nand U7432 (N_7432,N_7299,N_7305);
or U7433 (N_7433,N_7365,N_7344);
nand U7434 (N_7434,N_7253,N_7317);
and U7435 (N_7435,N_7279,N_7357);
or U7436 (N_7436,N_7343,N_7274);
nor U7437 (N_7437,N_7255,N_7276);
or U7438 (N_7438,N_7353,N_7356);
and U7439 (N_7439,N_7339,N_7252);
or U7440 (N_7440,N_7290,N_7291);
nand U7441 (N_7441,N_7252,N_7359);
nor U7442 (N_7442,N_7352,N_7357);
and U7443 (N_7443,N_7328,N_7354);
nand U7444 (N_7444,N_7270,N_7258);
or U7445 (N_7445,N_7292,N_7353);
nor U7446 (N_7446,N_7310,N_7331);
and U7447 (N_7447,N_7286,N_7275);
or U7448 (N_7448,N_7329,N_7268);
nor U7449 (N_7449,N_7348,N_7300);
nor U7450 (N_7450,N_7346,N_7305);
or U7451 (N_7451,N_7273,N_7327);
xor U7452 (N_7452,N_7296,N_7290);
and U7453 (N_7453,N_7259,N_7370);
nand U7454 (N_7454,N_7306,N_7366);
and U7455 (N_7455,N_7284,N_7311);
or U7456 (N_7456,N_7370,N_7301);
nor U7457 (N_7457,N_7252,N_7368);
or U7458 (N_7458,N_7340,N_7358);
nor U7459 (N_7459,N_7349,N_7259);
nand U7460 (N_7460,N_7352,N_7318);
nand U7461 (N_7461,N_7309,N_7315);
nand U7462 (N_7462,N_7285,N_7335);
or U7463 (N_7463,N_7367,N_7368);
nand U7464 (N_7464,N_7254,N_7298);
or U7465 (N_7465,N_7296,N_7322);
nor U7466 (N_7466,N_7306,N_7329);
and U7467 (N_7467,N_7315,N_7286);
or U7468 (N_7468,N_7344,N_7282);
xor U7469 (N_7469,N_7265,N_7257);
or U7470 (N_7470,N_7298,N_7327);
or U7471 (N_7471,N_7334,N_7336);
or U7472 (N_7472,N_7254,N_7278);
or U7473 (N_7473,N_7267,N_7342);
or U7474 (N_7474,N_7263,N_7307);
nand U7475 (N_7475,N_7302,N_7279);
and U7476 (N_7476,N_7354,N_7303);
and U7477 (N_7477,N_7372,N_7341);
nor U7478 (N_7478,N_7315,N_7250);
nand U7479 (N_7479,N_7360,N_7254);
nor U7480 (N_7480,N_7314,N_7272);
nand U7481 (N_7481,N_7312,N_7326);
and U7482 (N_7482,N_7280,N_7361);
nand U7483 (N_7483,N_7331,N_7365);
and U7484 (N_7484,N_7277,N_7342);
and U7485 (N_7485,N_7285,N_7372);
nand U7486 (N_7486,N_7314,N_7324);
xnor U7487 (N_7487,N_7271,N_7334);
and U7488 (N_7488,N_7259,N_7330);
nand U7489 (N_7489,N_7359,N_7315);
and U7490 (N_7490,N_7290,N_7341);
and U7491 (N_7491,N_7325,N_7341);
nand U7492 (N_7492,N_7300,N_7362);
nand U7493 (N_7493,N_7350,N_7366);
or U7494 (N_7494,N_7290,N_7372);
nor U7495 (N_7495,N_7357,N_7268);
or U7496 (N_7496,N_7276,N_7358);
nand U7497 (N_7497,N_7361,N_7263);
nand U7498 (N_7498,N_7273,N_7323);
nor U7499 (N_7499,N_7273,N_7271);
nand U7500 (N_7500,N_7497,N_7444);
nor U7501 (N_7501,N_7433,N_7447);
or U7502 (N_7502,N_7394,N_7415);
xnor U7503 (N_7503,N_7471,N_7428);
or U7504 (N_7504,N_7409,N_7465);
nand U7505 (N_7505,N_7486,N_7376);
or U7506 (N_7506,N_7387,N_7420);
nand U7507 (N_7507,N_7457,N_7439);
nand U7508 (N_7508,N_7395,N_7449);
or U7509 (N_7509,N_7386,N_7375);
or U7510 (N_7510,N_7410,N_7424);
nor U7511 (N_7511,N_7499,N_7495);
nand U7512 (N_7512,N_7381,N_7430);
and U7513 (N_7513,N_7451,N_7392);
nand U7514 (N_7514,N_7453,N_7464);
nand U7515 (N_7515,N_7480,N_7458);
or U7516 (N_7516,N_7399,N_7483);
or U7517 (N_7517,N_7432,N_7389);
or U7518 (N_7518,N_7377,N_7418);
nand U7519 (N_7519,N_7490,N_7456);
or U7520 (N_7520,N_7467,N_7398);
nand U7521 (N_7521,N_7385,N_7446);
nor U7522 (N_7522,N_7494,N_7474);
and U7523 (N_7523,N_7379,N_7462);
nand U7524 (N_7524,N_7404,N_7393);
or U7525 (N_7525,N_7472,N_7431);
or U7526 (N_7526,N_7476,N_7461);
nand U7527 (N_7527,N_7419,N_7481);
and U7528 (N_7528,N_7441,N_7440);
nor U7529 (N_7529,N_7382,N_7459);
xor U7530 (N_7530,N_7498,N_7455);
and U7531 (N_7531,N_7436,N_7487);
or U7532 (N_7532,N_7427,N_7442);
or U7533 (N_7533,N_7496,N_7470);
and U7534 (N_7534,N_7400,N_7489);
and U7535 (N_7535,N_7493,N_7488);
or U7536 (N_7536,N_7407,N_7469);
nor U7537 (N_7537,N_7391,N_7448);
nand U7538 (N_7538,N_7417,N_7423);
or U7539 (N_7539,N_7388,N_7443);
or U7540 (N_7540,N_7482,N_7484);
and U7541 (N_7541,N_7406,N_7408);
nor U7542 (N_7542,N_7466,N_7445);
nor U7543 (N_7543,N_7401,N_7478);
nor U7544 (N_7544,N_7426,N_7485);
and U7545 (N_7545,N_7437,N_7435);
and U7546 (N_7546,N_7460,N_7403);
nand U7547 (N_7547,N_7454,N_7396);
and U7548 (N_7548,N_7416,N_7397);
nand U7549 (N_7549,N_7434,N_7384);
and U7550 (N_7550,N_7413,N_7412);
or U7551 (N_7551,N_7380,N_7492);
nand U7552 (N_7552,N_7473,N_7414);
xor U7553 (N_7553,N_7491,N_7402);
nor U7554 (N_7554,N_7468,N_7463);
nor U7555 (N_7555,N_7450,N_7421);
and U7556 (N_7556,N_7438,N_7383);
or U7557 (N_7557,N_7479,N_7378);
or U7558 (N_7558,N_7452,N_7405);
and U7559 (N_7559,N_7429,N_7422);
or U7560 (N_7560,N_7390,N_7411);
nand U7561 (N_7561,N_7475,N_7425);
xnor U7562 (N_7562,N_7477,N_7411);
or U7563 (N_7563,N_7408,N_7444);
nand U7564 (N_7564,N_7443,N_7449);
xnor U7565 (N_7565,N_7422,N_7457);
xnor U7566 (N_7566,N_7415,N_7485);
or U7567 (N_7567,N_7465,N_7478);
and U7568 (N_7568,N_7477,N_7465);
nand U7569 (N_7569,N_7381,N_7404);
and U7570 (N_7570,N_7387,N_7489);
nand U7571 (N_7571,N_7396,N_7485);
and U7572 (N_7572,N_7424,N_7419);
nand U7573 (N_7573,N_7471,N_7392);
nor U7574 (N_7574,N_7417,N_7472);
and U7575 (N_7575,N_7391,N_7426);
nand U7576 (N_7576,N_7491,N_7435);
or U7577 (N_7577,N_7397,N_7403);
nor U7578 (N_7578,N_7457,N_7469);
nor U7579 (N_7579,N_7384,N_7433);
and U7580 (N_7580,N_7395,N_7401);
nor U7581 (N_7581,N_7497,N_7434);
xor U7582 (N_7582,N_7375,N_7498);
nand U7583 (N_7583,N_7392,N_7432);
or U7584 (N_7584,N_7383,N_7444);
nand U7585 (N_7585,N_7466,N_7406);
or U7586 (N_7586,N_7450,N_7420);
nor U7587 (N_7587,N_7482,N_7378);
and U7588 (N_7588,N_7494,N_7408);
and U7589 (N_7589,N_7438,N_7429);
and U7590 (N_7590,N_7463,N_7449);
or U7591 (N_7591,N_7381,N_7422);
nor U7592 (N_7592,N_7453,N_7475);
or U7593 (N_7593,N_7379,N_7457);
or U7594 (N_7594,N_7476,N_7449);
nor U7595 (N_7595,N_7432,N_7388);
nor U7596 (N_7596,N_7495,N_7485);
xor U7597 (N_7597,N_7392,N_7462);
nand U7598 (N_7598,N_7462,N_7477);
nor U7599 (N_7599,N_7386,N_7403);
and U7600 (N_7600,N_7394,N_7437);
and U7601 (N_7601,N_7445,N_7481);
or U7602 (N_7602,N_7476,N_7390);
or U7603 (N_7603,N_7423,N_7481);
nor U7604 (N_7604,N_7472,N_7483);
nor U7605 (N_7605,N_7397,N_7464);
nor U7606 (N_7606,N_7410,N_7494);
and U7607 (N_7607,N_7485,N_7466);
nor U7608 (N_7608,N_7388,N_7467);
nor U7609 (N_7609,N_7464,N_7378);
nand U7610 (N_7610,N_7443,N_7429);
nor U7611 (N_7611,N_7394,N_7490);
and U7612 (N_7612,N_7465,N_7419);
nor U7613 (N_7613,N_7396,N_7448);
nor U7614 (N_7614,N_7424,N_7470);
nand U7615 (N_7615,N_7418,N_7447);
and U7616 (N_7616,N_7483,N_7453);
nor U7617 (N_7617,N_7416,N_7456);
xor U7618 (N_7618,N_7464,N_7486);
and U7619 (N_7619,N_7402,N_7385);
nand U7620 (N_7620,N_7436,N_7425);
nand U7621 (N_7621,N_7394,N_7378);
or U7622 (N_7622,N_7410,N_7495);
xnor U7623 (N_7623,N_7400,N_7491);
nor U7624 (N_7624,N_7463,N_7489);
xnor U7625 (N_7625,N_7522,N_7540);
nor U7626 (N_7626,N_7586,N_7559);
and U7627 (N_7627,N_7569,N_7581);
and U7628 (N_7628,N_7538,N_7536);
nand U7629 (N_7629,N_7619,N_7552);
or U7630 (N_7630,N_7604,N_7623);
nor U7631 (N_7631,N_7537,N_7579);
nor U7632 (N_7632,N_7547,N_7595);
or U7633 (N_7633,N_7613,N_7525);
nor U7634 (N_7634,N_7592,N_7611);
nand U7635 (N_7635,N_7521,N_7618);
nor U7636 (N_7636,N_7503,N_7609);
nand U7637 (N_7637,N_7517,N_7535);
and U7638 (N_7638,N_7549,N_7597);
and U7639 (N_7639,N_7583,N_7582);
nand U7640 (N_7640,N_7594,N_7548);
or U7641 (N_7641,N_7501,N_7590);
xnor U7642 (N_7642,N_7577,N_7515);
nor U7643 (N_7643,N_7512,N_7511);
or U7644 (N_7644,N_7578,N_7530);
nand U7645 (N_7645,N_7572,N_7617);
nor U7646 (N_7646,N_7607,N_7622);
nand U7647 (N_7647,N_7542,N_7561);
xnor U7648 (N_7648,N_7614,N_7504);
nand U7649 (N_7649,N_7556,N_7516);
or U7650 (N_7650,N_7566,N_7585);
nor U7651 (N_7651,N_7544,N_7624);
and U7652 (N_7652,N_7505,N_7555);
nor U7653 (N_7653,N_7576,N_7508);
and U7654 (N_7654,N_7514,N_7509);
nand U7655 (N_7655,N_7528,N_7502);
nor U7656 (N_7656,N_7567,N_7520);
and U7657 (N_7657,N_7571,N_7531);
or U7658 (N_7658,N_7558,N_7527);
nor U7659 (N_7659,N_7534,N_7621);
nand U7660 (N_7660,N_7518,N_7612);
nor U7661 (N_7661,N_7600,N_7539);
nand U7662 (N_7662,N_7620,N_7573);
or U7663 (N_7663,N_7543,N_7564);
nand U7664 (N_7664,N_7575,N_7598);
or U7665 (N_7665,N_7519,N_7599);
xor U7666 (N_7666,N_7580,N_7587);
or U7667 (N_7667,N_7591,N_7523);
and U7668 (N_7668,N_7526,N_7602);
nand U7669 (N_7669,N_7589,N_7500);
nor U7670 (N_7670,N_7524,N_7601);
nor U7671 (N_7671,N_7603,N_7574);
nor U7672 (N_7672,N_7541,N_7605);
and U7673 (N_7673,N_7606,N_7545);
nor U7674 (N_7674,N_7513,N_7588);
or U7675 (N_7675,N_7546,N_7529);
and U7676 (N_7676,N_7562,N_7570);
xor U7677 (N_7677,N_7615,N_7551);
and U7678 (N_7678,N_7550,N_7563);
or U7679 (N_7679,N_7553,N_7584);
or U7680 (N_7680,N_7510,N_7533);
and U7681 (N_7681,N_7560,N_7554);
and U7682 (N_7682,N_7608,N_7568);
or U7683 (N_7683,N_7506,N_7557);
and U7684 (N_7684,N_7616,N_7565);
nand U7685 (N_7685,N_7596,N_7507);
and U7686 (N_7686,N_7532,N_7610);
and U7687 (N_7687,N_7593,N_7520);
or U7688 (N_7688,N_7568,N_7616);
nand U7689 (N_7689,N_7553,N_7562);
nor U7690 (N_7690,N_7541,N_7554);
and U7691 (N_7691,N_7576,N_7502);
nand U7692 (N_7692,N_7581,N_7554);
or U7693 (N_7693,N_7573,N_7594);
nor U7694 (N_7694,N_7621,N_7541);
nand U7695 (N_7695,N_7538,N_7610);
and U7696 (N_7696,N_7525,N_7585);
nor U7697 (N_7697,N_7575,N_7617);
and U7698 (N_7698,N_7606,N_7557);
and U7699 (N_7699,N_7536,N_7598);
nand U7700 (N_7700,N_7519,N_7604);
nand U7701 (N_7701,N_7608,N_7530);
nor U7702 (N_7702,N_7601,N_7516);
and U7703 (N_7703,N_7567,N_7623);
nand U7704 (N_7704,N_7597,N_7505);
and U7705 (N_7705,N_7595,N_7616);
xnor U7706 (N_7706,N_7597,N_7535);
nor U7707 (N_7707,N_7624,N_7536);
or U7708 (N_7708,N_7521,N_7515);
and U7709 (N_7709,N_7516,N_7537);
and U7710 (N_7710,N_7583,N_7588);
nand U7711 (N_7711,N_7618,N_7606);
nor U7712 (N_7712,N_7502,N_7520);
and U7713 (N_7713,N_7529,N_7545);
or U7714 (N_7714,N_7566,N_7530);
and U7715 (N_7715,N_7558,N_7518);
nor U7716 (N_7716,N_7502,N_7538);
xor U7717 (N_7717,N_7554,N_7579);
nand U7718 (N_7718,N_7587,N_7567);
xnor U7719 (N_7719,N_7602,N_7605);
nand U7720 (N_7720,N_7599,N_7594);
nor U7721 (N_7721,N_7557,N_7554);
or U7722 (N_7722,N_7601,N_7534);
nand U7723 (N_7723,N_7588,N_7608);
xnor U7724 (N_7724,N_7552,N_7584);
or U7725 (N_7725,N_7513,N_7618);
xnor U7726 (N_7726,N_7564,N_7579);
or U7727 (N_7727,N_7523,N_7515);
and U7728 (N_7728,N_7618,N_7552);
nand U7729 (N_7729,N_7596,N_7624);
nand U7730 (N_7730,N_7541,N_7547);
and U7731 (N_7731,N_7508,N_7563);
or U7732 (N_7732,N_7604,N_7545);
or U7733 (N_7733,N_7520,N_7586);
nand U7734 (N_7734,N_7599,N_7624);
nor U7735 (N_7735,N_7572,N_7598);
nand U7736 (N_7736,N_7591,N_7501);
or U7737 (N_7737,N_7565,N_7569);
nand U7738 (N_7738,N_7587,N_7608);
nand U7739 (N_7739,N_7517,N_7527);
nor U7740 (N_7740,N_7511,N_7569);
nand U7741 (N_7741,N_7595,N_7582);
nand U7742 (N_7742,N_7613,N_7564);
and U7743 (N_7743,N_7613,N_7549);
nand U7744 (N_7744,N_7573,N_7611);
nand U7745 (N_7745,N_7575,N_7587);
nor U7746 (N_7746,N_7549,N_7622);
nor U7747 (N_7747,N_7530,N_7518);
nand U7748 (N_7748,N_7538,N_7545);
nand U7749 (N_7749,N_7535,N_7557);
and U7750 (N_7750,N_7639,N_7719);
xnor U7751 (N_7751,N_7652,N_7696);
or U7752 (N_7752,N_7736,N_7698);
xnor U7753 (N_7753,N_7735,N_7745);
and U7754 (N_7754,N_7733,N_7635);
nand U7755 (N_7755,N_7728,N_7711);
or U7756 (N_7756,N_7723,N_7742);
and U7757 (N_7757,N_7706,N_7722);
or U7758 (N_7758,N_7665,N_7682);
xor U7759 (N_7759,N_7681,N_7721);
or U7760 (N_7760,N_7744,N_7734);
xor U7761 (N_7761,N_7661,N_7641);
nor U7762 (N_7762,N_7725,N_7631);
nor U7763 (N_7763,N_7697,N_7694);
or U7764 (N_7764,N_7701,N_7731);
nand U7765 (N_7765,N_7668,N_7678);
and U7766 (N_7766,N_7656,N_7692);
and U7767 (N_7767,N_7677,N_7645);
nand U7768 (N_7768,N_7649,N_7704);
and U7769 (N_7769,N_7655,N_7640);
and U7770 (N_7770,N_7663,N_7638);
nand U7771 (N_7771,N_7673,N_7651);
nor U7772 (N_7772,N_7710,N_7659);
and U7773 (N_7773,N_7695,N_7708);
nor U7774 (N_7774,N_7674,N_7690);
nor U7775 (N_7775,N_7627,N_7684);
nor U7776 (N_7776,N_7644,N_7630);
or U7777 (N_7777,N_7703,N_7626);
nor U7778 (N_7778,N_7686,N_7737);
nor U7779 (N_7779,N_7743,N_7625);
or U7780 (N_7780,N_7741,N_7648);
and U7781 (N_7781,N_7693,N_7748);
and U7782 (N_7782,N_7680,N_7702);
and U7783 (N_7783,N_7628,N_7747);
or U7784 (N_7784,N_7636,N_7730);
xnor U7785 (N_7785,N_7650,N_7664);
nand U7786 (N_7786,N_7646,N_7671);
and U7787 (N_7787,N_7670,N_7700);
nor U7788 (N_7788,N_7718,N_7662);
nand U7789 (N_7789,N_7634,N_7666);
nor U7790 (N_7790,N_7647,N_7629);
or U7791 (N_7791,N_7739,N_7713);
nor U7792 (N_7792,N_7683,N_7633);
nand U7793 (N_7793,N_7654,N_7672);
nand U7794 (N_7794,N_7643,N_7679);
or U7795 (N_7795,N_7749,N_7688);
nor U7796 (N_7796,N_7669,N_7676);
and U7797 (N_7797,N_7712,N_7720);
or U7798 (N_7798,N_7642,N_7707);
and U7799 (N_7799,N_7740,N_7675);
and U7800 (N_7800,N_7724,N_7746);
nand U7801 (N_7801,N_7660,N_7717);
nor U7802 (N_7802,N_7653,N_7637);
and U7803 (N_7803,N_7689,N_7685);
and U7804 (N_7804,N_7727,N_7687);
or U7805 (N_7805,N_7667,N_7714);
xor U7806 (N_7806,N_7658,N_7726);
and U7807 (N_7807,N_7738,N_7709);
or U7808 (N_7808,N_7632,N_7729);
nor U7809 (N_7809,N_7705,N_7716);
nand U7810 (N_7810,N_7657,N_7699);
nand U7811 (N_7811,N_7715,N_7691);
and U7812 (N_7812,N_7732,N_7712);
xnor U7813 (N_7813,N_7706,N_7743);
nor U7814 (N_7814,N_7718,N_7638);
or U7815 (N_7815,N_7686,N_7625);
nand U7816 (N_7816,N_7712,N_7746);
and U7817 (N_7817,N_7706,N_7724);
or U7818 (N_7818,N_7712,N_7716);
xnor U7819 (N_7819,N_7676,N_7697);
and U7820 (N_7820,N_7747,N_7696);
nor U7821 (N_7821,N_7672,N_7699);
or U7822 (N_7822,N_7740,N_7700);
or U7823 (N_7823,N_7717,N_7732);
xor U7824 (N_7824,N_7628,N_7663);
and U7825 (N_7825,N_7748,N_7652);
or U7826 (N_7826,N_7632,N_7662);
nand U7827 (N_7827,N_7676,N_7721);
nor U7828 (N_7828,N_7673,N_7741);
nor U7829 (N_7829,N_7657,N_7648);
xnor U7830 (N_7830,N_7720,N_7634);
nor U7831 (N_7831,N_7648,N_7739);
xor U7832 (N_7832,N_7628,N_7688);
nor U7833 (N_7833,N_7626,N_7714);
and U7834 (N_7834,N_7703,N_7685);
xor U7835 (N_7835,N_7701,N_7691);
nor U7836 (N_7836,N_7697,N_7678);
or U7837 (N_7837,N_7703,N_7718);
nor U7838 (N_7838,N_7687,N_7631);
or U7839 (N_7839,N_7710,N_7670);
and U7840 (N_7840,N_7698,N_7649);
nand U7841 (N_7841,N_7733,N_7740);
nor U7842 (N_7842,N_7626,N_7683);
xnor U7843 (N_7843,N_7721,N_7663);
or U7844 (N_7844,N_7669,N_7721);
and U7845 (N_7845,N_7720,N_7737);
nand U7846 (N_7846,N_7636,N_7725);
nor U7847 (N_7847,N_7692,N_7675);
nand U7848 (N_7848,N_7695,N_7636);
and U7849 (N_7849,N_7691,N_7739);
and U7850 (N_7850,N_7705,N_7728);
xnor U7851 (N_7851,N_7676,N_7630);
and U7852 (N_7852,N_7732,N_7647);
nand U7853 (N_7853,N_7746,N_7690);
or U7854 (N_7854,N_7702,N_7662);
and U7855 (N_7855,N_7744,N_7716);
nor U7856 (N_7856,N_7684,N_7687);
or U7857 (N_7857,N_7658,N_7650);
nor U7858 (N_7858,N_7723,N_7664);
or U7859 (N_7859,N_7704,N_7694);
and U7860 (N_7860,N_7685,N_7720);
nor U7861 (N_7861,N_7734,N_7721);
and U7862 (N_7862,N_7641,N_7696);
or U7863 (N_7863,N_7696,N_7684);
or U7864 (N_7864,N_7690,N_7712);
nor U7865 (N_7865,N_7704,N_7731);
and U7866 (N_7866,N_7625,N_7652);
xor U7867 (N_7867,N_7684,N_7719);
nand U7868 (N_7868,N_7669,N_7686);
nand U7869 (N_7869,N_7639,N_7685);
xor U7870 (N_7870,N_7667,N_7719);
xnor U7871 (N_7871,N_7693,N_7712);
or U7872 (N_7872,N_7634,N_7654);
or U7873 (N_7873,N_7714,N_7631);
xor U7874 (N_7874,N_7709,N_7706);
and U7875 (N_7875,N_7755,N_7848);
or U7876 (N_7876,N_7781,N_7845);
nor U7877 (N_7877,N_7806,N_7833);
and U7878 (N_7878,N_7772,N_7842);
xnor U7879 (N_7879,N_7849,N_7817);
or U7880 (N_7880,N_7836,N_7767);
and U7881 (N_7881,N_7778,N_7759);
nand U7882 (N_7882,N_7840,N_7805);
or U7883 (N_7883,N_7799,N_7780);
and U7884 (N_7884,N_7761,N_7847);
or U7885 (N_7885,N_7754,N_7791);
nand U7886 (N_7886,N_7820,N_7771);
or U7887 (N_7887,N_7752,N_7773);
nor U7888 (N_7888,N_7852,N_7867);
nand U7889 (N_7889,N_7783,N_7834);
or U7890 (N_7890,N_7819,N_7800);
nand U7891 (N_7891,N_7774,N_7818);
or U7892 (N_7892,N_7786,N_7868);
nor U7893 (N_7893,N_7787,N_7830);
nor U7894 (N_7894,N_7853,N_7821);
or U7895 (N_7895,N_7766,N_7782);
nor U7896 (N_7896,N_7813,N_7779);
and U7897 (N_7897,N_7765,N_7757);
nand U7898 (N_7898,N_7860,N_7784);
xnor U7899 (N_7899,N_7871,N_7844);
and U7900 (N_7900,N_7753,N_7762);
or U7901 (N_7901,N_7810,N_7763);
nor U7902 (N_7902,N_7866,N_7797);
xor U7903 (N_7903,N_7768,N_7851);
and U7904 (N_7904,N_7812,N_7815);
and U7905 (N_7905,N_7794,N_7764);
and U7906 (N_7906,N_7822,N_7756);
and U7907 (N_7907,N_7859,N_7827);
nor U7908 (N_7908,N_7795,N_7856);
nand U7909 (N_7909,N_7850,N_7828);
xnor U7910 (N_7910,N_7770,N_7808);
nor U7911 (N_7911,N_7832,N_7872);
nand U7912 (N_7912,N_7793,N_7758);
nor U7913 (N_7913,N_7838,N_7809);
nor U7914 (N_7914,N_7826,N_7874);
or U7915 (N_7915,N_7798,N_7796);
or U7916 (N_7916,N_7750,N_7789);
nand U7917 (N_7917,N_7843,N_7825);
or U7918 (N_7918,N_7814,N_7777);
xor U7919 (N_7919,N_7769,N_7816);
or U7920 (N_7920,N_7864,N_7855);
or U7921 (N_7921,N_7776,N_7792);
or U7922 (N_7922,N_7837,N_7869);
or U7923 (N_7923,N_7854,N_7865);
nand U7924 (N_7924,N_7807,N_7829);
nor U7925 (N_7925,N_7790,N_7831);
nor U7926 (N_7926,N_7811,N_7823);
nand U7927 (N_7927,N_7858,N_7841);
nand U7928 (N_7928,N_7788,N_7785);
xor U7929 (N_7929,N_7839,N_7863);
or U7930 (N_7930,N_7846,N_7824);
nand U7931 (N_7931,N_7870,N_7862);
nor U7932 (N_7932,N_7873,N_7802);
or U7933 (N_7933,N_7801,N_7760);
nor U7934 (N_7934,N_7857,N_7751);
and U7935 (N_7935,N_7775,N_7861);
and U7936 (N_7936,N_7835,N_7803);
nor U7937 (N_7937,N_7804,N_7834);
nor U7938 (N_7938,N_7765,N_7848);
and U7939 (N_7939,N_7777,N_7753);
nor U7940 (N_7940,N_7855,N_7777);
nand U7941 (N_7941,N_7847,N_7784);
nor U7942 (N_7942,N_7871,N_7798);
nor U7943 (N_7943,N_7790,N_7765);
or U7944 (N_7944,N_7813,N_7810);
nand U7945 (N_7945,N_7872,N_7800);
nand U7946 (N_7946,N_7755,N_7831);
xor U7947 (N_7947,N_7767,N_7757);
xnor U7948 (N_7948,N_7806,N_7793);
xor U7949 (N_7949,N_7813,N_7832);
or U7950 (N_7950,N_7769,N_7865);
nor U7951 (N_7951,N_7810,N_7753);
and U7952 (N_7952,N_7804,N_7771);
nor U7953 (N_7953,N_7818,N_7874);
and U7954 (N_7954,N_7843,N_7835);
nor U7955 (N_7955,N_7793,N_7805);
nor U7956 (N_7956,N_7785,N_7867);
nand U7957 (N_7957,N_7795,N_7823);
nor U7958 (N_7958,N_7778,N_7854);
nand U7959 (N_7959,N_7852,N_7796);
and U7960 (N_7960,N_7800,N_7781);
and U7961 (N_7961,N_7803,N_7753);
nor U7962 (N_7962,N_7807,N_7788);
or U7963 (N_7963,N_7789,N_7866);
or U7964 (N_7964,N_7758,N_7862);
and U7965 (N_7965,N_7777,N_7835);
xnor U7966 (N_7966,N_7858,N_7814);
and U7967 (N_7967,N_7819,N_7766);
xnor U7968 (N_7968,N_7771,N_7867);
or U7969 (N_7969,N_7761,N_7872);
or U7970 (N_7970,N_7759,N_7763);
nor U7971 (N_7971,N_7870,N_7832);
or U7972 (N_7972,N_7753,N_7820);
nand U7973 (N_7973,N_7794,N_7855);
or U7974 (N_7974,N_7812,N_7779);
nor U7975 (N_7975,N_7798,N_7829);
nand U7976 (N_7976,N_7774,N_7827);
nor U7977 (N_7977,N_7813,N_7806);
nor U7978 (N_7978,N_7753,N_7824);
nand U7979 (N_7979,N_7799,N_7778);
or U7980 (N_7980,N_7829,N_7762);
or U7981 (N_7981,N_7859,N_7769);
and U7982 (N_7982,N_7848,N_7824);
or U7983 (N_7983,N_7865,N_7862);
and U7984 (N_7984,N_7762,N_7782);
or U7985 (N_7985,N_7842,N_7874);
nand U7986 (N_7986,N_7763,N_7869);
and U7987 (N_7987,N_7771,N_7751);
nor U7988 (N_7988,N_7862,N_7826);
xnor U7989 (N_7989,N_7846,N_7778);
nand U7990 (N_7990,N_7795,N_7787);
nand U7991 (N_7991,N_7781,N_7757);
or U7992 (N_7992,N_7824,N_7874);
and U7993 (N_7993,N_7795,N_7814);
or U7994 (N_7994,N_7817,N_7834);
nand U7995 (N_7995,N_7810,N_7779);
or U7996 (N_7996,N_7788,N_7871);
nor U7997 (N_7997,N_7809,N_7839);
xor U7998 (N_7998,N_7825,N_7832);
nor U7999 (N_7999,N_7758,N_7860);
nand U8000 (N_8000,N_7895,N_7977);
nand U8001 (N_8001,N_7887,N_7879);
nor U8002 (N_8002,N_7991,N_7985);
nor U8003 (N_8003,N_7963,N_7877);
or U8004 (N_8004,N_7936,N_7982);
xnor U8005 (N_8005,N_7989,N_7968);
and U8006 (N_8006,N_7929,N_7987);
or U8007 (N_8007,N_7939,N_7994);
or U8008 (N_8008,N_7918,N_7955);
nor U8009 (N_8009,N_7917,N_7978);
nor U8010 (N_8010,N_7992,N_7941);
nand U8011 (N_8011,N_7942,N_7973);
nor U8012 (N_8012,N_7935,N_7954);
or U8013 (N_8013,N_7974,N_7947);
xor U8014 (N_8014,N_7892,N_7884);
or U8015 (N_8015,N_7898,N_7916);
or U8016 (N_8016,N_7949,N_7904);
or U8017 (N_8017,N_7880,N_7931);
nand U8018 (N_8018,N_7927,N_7890);
nand U8019 (N_8019,N_7970,N_7993);
nor U8020 (N_8020,N_7938,N_7934);
xnor U8021 (N_8021,N_7889,N_7988);
nor U8022 (N_8022,N_7975,N_7925);
and U8023 (N_8023,N_7893,N_7894);
nand U8024 (N_8024,N_7946,N_7971);
and U8025 (N_8025,N_7932,N_7961);
or U8026 (N_8026,N_7897,N_7979);
xnor U8027 (N_8027,N_7958,N_7986);
and U8028 (N_8028,N_7933,N_7906);
nor U8029 (N_8029,N_7937,N_7909);
nand U8030 (N_8030,N_7959,N_7996);
nand U8031 (N_8031,N_7984,N_7998);
or U8032 (N_8032,N_7923,N_7957);
nand U8033 (N_8033,N_7976,N_7969);
nand U8034 (N_8034,N_7891,N_7997);
and U8035 (N_8035,N_7883,N_7930);
nand U8036 (N_8036,N_7912,N_7915);
or U8037 (N_8037,N_7911,N_7896);
nor U8038 (N_8038,N_7899,N_7951);
or U8039 (N_8039,N_7999,N_7924);
or U8040 (N_8040,N_7920,N_7960);
nand U8041 (N_8041,N_7950,N_7907);
nand U8042 (N_8042,N_7888,N_7943);
xnor U8043 (N_8043,N_7882,N_7983);
and U8044 (N_8044,N_7972,N_7944);
or U8045 (N_8045,N_7953,N_7913);
nor U8046 (N_8046,N_7962,N_7980);
nand U8047 (N_8047,N_7900,N_7926);
or U8048 (N_8048,N_7965,N_7901);
and U8049 (N_8049,N_7922,N_7881);
nor U8050 (N_8050,N_7875,N_7886);
nand U8051 (N_8051,N_7956,N_7995);
and U8052 (N_8052,N_7948,N_7921);
xor U8053 (N_8053,N_7966,N_7903);
and U8054 (N_8054,N_7964,N_7945);
or U8055 (N_8055,N_7910,N_7876);
nand U8056 (N_8056,N_7967,N_7919);
nor U8057 (N_8057,N_7940,N_7902);
nor U8058 (N_8058,N_7908,N_7990);
or U8059 (N_8059,N_7981,N_7952);
nand U8060 (N_8060,N_7885,N_7905);
nand U8061 (N_8061,N_7928,N_7878);
nor U8062 (N_8062,N_7914,N_7889);
nor U8063 (N_8063,N_7913,N_7990);
or U8064 (N_8064,N_7987,N_7994);
and U8065 (N_8065,N_7955,N_7912);
xnor U8066 (N_8066,N_7944,N_7900);
nand U8067 (N_8067,N_7937,N_7936);
nor U8068 (N_8068,N_7962,N_7910);
or U8069 (N_8069,N_7988,N_7983);
nor U8070 (N_8070,N_7971,N_7964);
or U8071 (N_8071,N_7959,N_7916);
or U8072 (N_8072,N_7938,N_7883);
nand U8073 (N_8073,N_7980,N_7952);
xnor U8074 (N_8074,N_7887,N_7914);
nor U8075 (N_8075,N_7974,N_7988);
and U8076 (N_8076,N_7984,N_7936);
and U8077 (N_8077,N_7938,N_7900);
and U8078 (N_8078,N_7947,N_7882);
and U8079 (N_8079,N_7903,N_7992);
and U8080 (N_8080,N_7878,N_7923);
nor U8081 (N_8081,N_7928,N_7932);
or U8082 (N_8082,N_7997,N_7885);
nor U8083 (N_8083,N_7919,N_7970);
or U8084 (N_8084,N_7894,N_7973);
or U8085 (N_8085,N_7881,N_7924);
nor U8086 (N_8086,N_7909,N_7878);
or U8087 (N_8087,N_7960,N_7897);
and U8088 (N_8088,N_7957,N_7975);
or U8089 (N_8089,N_7876,N_7905);
and U8090 (N_8090,N_7922,N_7907);
nand U8091 (N_8091,N_7930,N_7974);
nor U8092 (N_8092,N_7888,N_7905);
or U8093 (N_8093,N_7995,N_7886);
or U8094 (N_8094,N_7916,N_7922);
nand U8095 (N_8095,N_7981,N_7925);
or U8096 (N_8096,N_7933,N_7997);
nand U8097 (N_8097,N_7898,N_7986);
nor U8098 (N_8098,N_7932,N_7911);
xnor U8099 (N_8099,N_7891,N_7921);
nor U8100 (N_8100,N_7953,N_7918);
nand U8101 (N_8101,N_7875,N_7937);
nand U8102 (N_8102,N_7900,N_7915);
or U8103 (N_8103,N_7923,N_7920);
xnor U8104 (N_8104,N_7911,N_7954);
nor U8105 (N_8105,N_7879,N_7876);
xor U8106 (N_8106,N_7911,N_7930);
xor U8107 (N_8107,N_7913,N_7951);
or U8108 (N_8108,N_7907,N_7972);
or U8109 (N_8109,N_7951,N_7941);
and U8110 (N_8110,N_7973,N_7939);
and U8111 (N_8111,N_7916,N_7936);
or U8112 (N_8112,N_7989,N_7919);
nor U8113 (N_8113,N_7958,N_7899);
nand U8114 (N_8114,N_7922,N_7917);
and U8115 (N_8115,N_7947,N_7990);
nand U8116 (N_8116,N_7971,N_7934);
nand U8117 (N_8117,N_7923,N_7917);
xor U8118 (N_8118,N_7926,N_7882);
nor U8119 (N_8119,N_7885,N_7883);
nand U8120 (N_8120,N_7918,N_7888);
nor U8121 (N_8121,N_7891,N_7931);
nor U8122 (N_8122,N_7932,N_7990);
or U8123 (N_8123,N_7913,N_7962);
or U8124 (N_8124,N_7980,N_7876);
nor U8125 (N_8125,N_8106,N_8083);
xnor U8126 (N_8126,N_8028,N_8107);
and U8127 (N_8127,N_8097,N_8091);
nor U8128 (N_8128,N_8010,N_8058);
and U8129 (N_8129,N_8071,N_8085);
or U8130 (N_8130,N_8101,N_8076);
nand U8131 (N_8131,N_8017,N_8096);
nor U8132 (N_8132,N_8030,N_8117);
and U8133 (N_8133,N_8059,N_8092);
nand U8134 (N_8134,N_8122,N_8088);
or U8135 (N_8135,N_8015,N_8000);
and U8136 (N_8136,N_8074,N_8124);
and U8137 (N_8137,N_8061,N_8026);
or U8138 (N_8138,N_8042,N_8093);
xnor U8139 (N_8139,N_8020,N_8084);
nor U8140 (N_8140,N_8113,N_8048);
and U8141 (N_8141,N_8032,N_8060);
nand U8142 (N_8142,N_8082,N_8039);
nand U8143 (N_8143,N_8123,N_8105);
or U8144 (N_8144,N_8027,N_8014);
and U8145 (N_8145,N_8099,N_8034);
nor U8146 (N_8146,N_8072,N_8004);
xor U8147 (N_8147,N_8067,N_8005);
and U8148 (N_8148,N_8073,N_8043);
and U8149 (N_8149,N_8049,N_8018);
and U8150 (N_8150,N_8013,N_8033);
xnor U8151 (N_8151,N_8053,N_8104);
xor U8152 (N_8152,N_8006,N_8008);
or U8153 (N_8153,N_8029,N_8080);
xnor U8154 (N_8154,N_8098,N_8016);
xor U8155 (N_8155,N_8055,N_8051);
or U8156 (N_8156,N_8041,N_8095);
nand U8157 (N_8157,N_8109,N_8050);
nand U8158 (N_8158,N_8023,N_8116);
nand U8159 (N_8159,N_8040,N_8002);
xor U8160 (N_8160,N_8115,N_8100);
and U8161 (N_8161,N_8038,N_8035);
and U8162 (N_8162,N_8022,N_8025);
nor U8163 (N_8163,N_8112,N_8031);
nor U8164 (N_8164,N_8057,N_8064);
nand U8165 (N_8165,N_8079,N_8068);
xor U8166 (N_8166,N_8111,N_8052);
nor U8167 (N_8167,N_8081,N_8078);
nand U8168 (N_8168,N_8077,N_8044);
xnor U8169 (N_8169,N_8003,N_8119);
xnor U8170 (N_8170,N_8037,N_8054);
nor U8171 (N_8171,N_8090,N_8066);
nor U8172 (N_8172,N_8094,N_8086);
nor U8173 (N_8173,N_8110,N_8011);
or U8174 (N_8174,N_8102,N_8075);
nor U8175 (N_8175,N_8062,N_8063);
and U8176 (N_8176,N_8046,N_8001);
nor U8177 (N_8177,N_8087,N_8121);
or U8178 (N_8178,N_8065,N_8120);
nand U8179 (N_8179,N_8045,N_8103);
nor U8180 (N_8180,N_8019,N_8024);
or U8181 (N_8181,N_8007,N_8089);
nand U8182 (N_8182,N_8012,N_8114);
nand U8183 (N_8183,N_8070,N_8047);
or U8184 (N_8184,N_8036,N_8021);
nand U8185 (N_8185,N_8056,N_8118);
nand U8186 (N_8186,N_8108,N_8069);
or U8187 (N_8187,N_8009,N_8048);
or U8188 (N_8188,N_8066,N_8059);
nor U8189 (N_8189,N_8029,N_8039);
nand U8190 (N_8190,N_8095,N_8040);
and U8191 (N_8191,N_8015,N_8088);
xnor U8192 (N_8192,N_8023,N_8079);
or U8193 (N_8193,N_8011,N_8120);
xnor U8194 (N_8194,N_8121,N_8011);
nor U8195 (N_8195,N_8054,N_8066);
and U8196 (N_8196,N_8032,N_8111);
or U8197 (N_8197,N_8051,N_8008);
nor U8198 (N_8198,N_8088,N_8037);
and U8199 (N_8199,N_8111,N_8018);
xnor U8200 (N_8200,N_8058,N_8080);
nor U8201 (N_8201,N_8003,N_8025);
nor U8202 (N_8202,N_8073,N_8053);
nor U8203 (N_8203,N_8030,N_8060);
nand U8204 (N_8204,N_8124,N_8030);
nor U8205 (N_8205,N_8053,N_8043);
nor U8206 (N_8206,N_8047,N_8017);
nand U8207 (N_8207,N_8055,N_8081);
nor U8208 (N_8208,N_8054,N_8095);
nand U8209 (N_8209,N_8118,N_8046);
nor U8210 (N_8210,N_8065,N_8030);
and U8211 (N_8211,N_8099,N_8082);
nand U8212 (N_8212,N_8003,N_8020);
or U8213 (N_8213,N_8122,N_8019);
and U8214 (N_8214,N_8001,N_8000);
and U8215 (N_8215,N_8068,N_8087);
and U8216 (N_8216,N_8055,N_8082);
and U8217 (N_8217,N_8094,N_8002);
or U8218 (N_8218,N_8003,N_8093);
or U8219 (N_8219,N_8041,N_8061);
or U8220 (N_8220,N_8106,N_8110);
and U8221 (N_8221,N_8108,N_8015);
nand U8222 (N_8222,N_8002,N_8086);
and U8223 (N_8223,N_8066,N_8085);
nor U8224 (N_8224,N_8076,N_8033);
nor U8225 (N_8225,N_8120,N_8068);
nand U8226 (N_8226,N_8045,N_8082);
nor U8227 (N_8227,N_8032,N_8029);
or U8228 (N_8228,N_8007,N_8083);
nor U8229 (N_8229,N_8039,N_8092);
and U8230 (N_8230,N_8083,N_8060);
and U8231 (N_8231,N_8092,N_8098);
nand U8232 (N_8232,N_8039,N_8020);
nand U8233 (N_8233,N_8024,N_8039);
xnor U8234 (N_8234,N_8110,N_8045);
nand U8235 (N_8235,N_8034,N_8049);
and U8236 (N_8236,N_8001,N_8040);
nand U8237 (N_8237,N_8075,N_8096);
and U8238 (N_8238,N_8088,N_8110);
or U8239 (N_8239,N_8047,N_8100);
nor U8240 (N_8240,N_8077,N_8020);
nor U8241 (N_8241,N_8046,N_8120);
and U8242 (N_8242,N_8055,N_8094);
and U8243 (N_8243,N_8020,N_8081);
xor U8244 (N_8244,N_8066,N_8041);
nand U8245 (N_8245,N_8041,N_8115);
nor U8246 (N_8246,N_8048,N_8109);
or U8247 (N_8247,N_8085,N_8106);
or U8248 (N_8248,N_8103,N_8007);
xnor U8249 (N_8249,N_8075,N_8047);
and U8250 (N_8250,N_8245,N_8208);
and U8251 (N_8251,N_8178,N_8154);
xnor U8252 (N_8252,N_8236,N_8218);
nand U8253 (N_8253,N_8186,N_8222);
or U8254 (N_8254,N_8189,N_8162);
and U8255 (N_8255,N_8157,N_8177);
and U8256 (N_8256,N_8207,N_8130);
and U8257 (N_8257,N_8200,N_8224);
or U8258 (N_8258,N_8247,N_8143);
xnor U8259 (N_8259,N_8175,N_8174);
and U8260 (N_8260,N_8201,N_8197);
nor U8261 (N_8261,N_8226,N_8182);
and U8262 (N_8262,N_8138,N_8128);
nor U8263 (N_8263,N_8223,N_8241);
nand U8264 (N_8264,N_8229,N_8131);
or U8265 (N_8265,N_8134,N_8126);
and U8266 (N_8266,N_8146,N_8181);
nor U8267 (N_8267,N_8161,N_8129);
nor U8268 (N_8268,N_8139,N_8219);
nand U8269 (N_8269,N_8176,N_8204);
or U8270 (N_8270,N_8145,N_8155);
or U8271 (N_8271,N_8215,N_8240);
xnor U8272 (N_8272,N_8137,N_8170);
and U8273 (N_8273,N_8212,N_8239);
nor U8274 (N_8274,N_8172,N_8190);
or U8275 (N_8275,N_8193,N_8135);
nand U8276 (N_8276,N_8237,N_8214);
nor U8277 (N_8277,N_8202,N_8141);
nor U8278 (N_8278,N_8169,N_8230);
or U8279 (N_8279,N_8185,N_8152);
nand U8280 (N_8280,N_8149,N_8248);
and U8281 (N_8281,N_8133,N_8184);
and U8282 (N_8282,N_8159,N_8140);
nand U8283 (N_8283,N_8166,N_8188);
nor U8284 (N_8284,N_8187,N_8179);
nor U8285 (N_8285,N_8125,N_8173);
or U8286 (N_8286,N_8191,N_8249);
xor U8287 (N_8287,N_8216,N_8232);
nor U8288 (N_8288,N_8167,N_8151);
or U8289 (N_8289,N_8220,N_8156);
and U8290 (N_8290,N_8244,N_8210);
nand U8291 (N_8291,N_8153,N_8233);
or U8292 (N_8292,N_8235,N_8228);
nor U8293 (N_8293,N_8238,N_8192);
and U8294 (N_8294,N_8234,N_8221);
or U8295 (N_8295,N_8195,N_8158);
nor U8296 (N_8296,N_8198,N_8163);
or U8297 (N_8297,N_8132,N_8199);
and U8298 (N_8298,N_8127,N_8150);
and U8299 (N_8299,N_8194,N_8231);
nand U8300 (N_8300,N_8164,N_8144);
and U8301 (N_8301,N_8136,N_8242);
and U8302 (N_8302,N_8147,N_8203);
nor U8303 (N_8303,N_8211,N_8217);
nor U8304 (N_8304,N_8209,N_8243);
or U8305 (N_8305,N_8160,N_8246);
and U8306 (N_8306,N_8183,N_8148);
or U8307 (N_8307,N_8165,N_8180);
or U8308 (N_8308,N_8168,N_8196);
and U8309 (N_8309,N_8225,N_8213);
or U8310 (N_8310,N_8206,N_8227);
nor U8311 (N_8311,N_8171,N_8205);
and U8312 (N_8312,N_8142,N_8199);
nor U8313 (N_8313,N_8226,N_8221);
xnor U8314 (N_8314,N_8181,N_8166);
nand U8315 (N_8315,N_8158,N_8241);
nand U8316 (N_8316,N_8198,N_8239);
or U8317 (N_8317,N_8202,N_8207);
nor U8318 (N_8318,N_8145,N_8232);
nand U8319 (N_8319,N_8135,N_8200);
nand U8320 (N_8320,N_8185,N_8199);
and U8321 (N_8321,N_8193,N_8208);
and U8322 (N_8322,N_8161,N_8178);
nand U8323 (N_8323,N_8214,N_8134);
nor U8324 (N_8324,N_8166,N_8194);
nand U8325 (N_8325,N_8222,N_8174);
nand U8326 (N_8326,N_8205,N_8148);
and U8327 (N_8327,N_8247,N_8148);
nand U8328 (N_8328,N_8202,N_8163);
or U8329 (N_8329,N_8218,N_8174);
and U8330 (N_8330,N_8159,N_8180);
or U8331 (N_8331,N_8149,N_8201);
or U8332 (N_8332,N_8167,N_8247);
nor U8333 (N_8333,N_8239,N_8133);
xnor U8334 (N_8334,N_8235,N_8180);
nand U8335 (N_8335,N_8218,N_8194);
and U8336 (N_8336,N_8155,N_8144);
or U8337 (N_8337,N_8197,N_8237);
xor U8338 (N_8338,N_8147,N_8192);
and U8339 (N_8339,N_8237,N_8209);
or U8340 (N_8340,N_8224,N_8216);
nand U8341 (N_8341,N_8194,N_8217);
or U8342 (N_8342,N_8132,N_8247);
nand U8343 (N_8343,N_8143,N_8216);
or U8344 (N_8344,N_8194,N_8191);
or U8345 (N_8345,N_8229,N_8190);
and U8346 (N_8346,N_8200,N_8219);
nor U8347 (N_8347,N_8210,N_8127);
and U8348 (N_8348,N_8223,N_8172);
xnor U8349 (N_8349,N_8129,N_8247);
or U8350 (N_8350,N_8226,N_8200);
nor U8351 (N_8351,N_8129,N_8242);
and U8352 (N_8352,N_8139,N_8209);
nand U8353 (N_8353,N_8191,N_8161);
or U8354 (N_8354,N_8163,N_8214);
or U8355 (N_8355,N_8174,N_8249);
nand U8356 (N_8356,N_8157,N_8179);
xnor U8357 (N_8357,N_8193,N_8130);
xor U8358 (N_8358,N_8183,N_8208);
or U8359 (N_8359,N_8226,N_8175);
and U8360 (N_8360,N_8155,N_8175);
and U8361 (N_8361,N_8138,N_8234);
xnor U8362 (N_8362,N_8180,N_8170);
or U8363 (N_8363,N_8148,N_8143);
nand U8364 (N_8364,N_8133,N_8129);
nor U8365 (N_8365,N_8136,N_8206);
and U8366 (N_8366,N_8161,N_8195);
xor U8367 (N_8367,N_8161,N_8151);
nor U8368 (N_8368,N_8161,N_8139);
nor U8369 (N_8369,N_8171,N_8167);
and U8370 (N_8370,N_8132,N_8228);
nand U8371 (N_8371,N_8157,N_8194);
or U8372 (N_8372,N_8160,N_8219);
xor U8373 (N_8373,N_8162,N_8217);
and U8374 (N_8374,N_8132,N_8191);
xor U8375 (N_8375,N_8271,N_8327);
nor U8376 (N_8376,N_8251,N_8335);
nand U8377 (N_8377,N_8363,N_8337);
nor U8378 (N_8378,N_8319,N_8302);
or U8379 (N_8379,N_8310,N_8318);
or U8380 (N_8380,N_8270,N_8275);
and U8381 (N_8381,N_8358,N_8258);
nor U8382 (N_8382,N_8315,N_8280);
or U8383 (N_8383,N_8344,N_8353);
and U8384 (N_8384,N_8326,N_8305);
and U8385 (N_8385,N_8341,N_8295);
xnor U8386 (N_8386,N_8265,N_8329);
xor U8387 (N_8387,N_8346,N_8303);
nor U8388 (N_8388,N_8347,N_8334);
nor U8389 (N_8389,N_8304,N_8355);
nor U8390 (N_8390,N_8373,N_8264);
nand U8391 (N_8391,N_8250,N_8374);
nor U8392 (N_8392,N_8311,N_8306);
nand U8393 (N_8393,N_8356,N_8364);
or U8394 (N_8394,N_8368,N_8320);
and U8395 (N_8395,N_8279,N_8338);
and U8396 (N_8396,N_8345,N_8299);
nand U8397 (N_8397,N_8289,N_8253);
nand U8398 (N_8398,N_8312,N_8357);
and U8399 (N_8399,N_8331,N_8263);
nor U8400 (N_8400,N_8294,N_8301);
nor U8401 (N_8401,N_8369,N_8309);
and U8402 (N_8402,N_8323,N_8261);
xnor U8403 (N_8403,N_8325,N_8367);
nand U8404 (N_8404,N_8308,N_8350);
nor U8405 (N_8405,N_8296,N_8360);
or U8406 (N_8406,N_8361,N_8307);
xnor U8407 (N_8407,N_8278,N_8370);
nor U8408 (N_8408,N_8257,N_8314);
nor U8409 (N_8409,N_8297,N_8267);
nor U8410 (N_8410,N_8313,N_8333);
and U8411 (N_8411,N_8277,N_8252);
nor U8412 (N_8412,N_8365,N_8290);
nor U8413 (N_8413,N_8272,N_8371);
or U8414 (N_8414,N_8291,N_8288);
nor U8415 (N_8415,N_8362,N_8339);
or U8416 (N_8416,N_8322,N_8255);
or U8417 (N_8417,N_8330,N_8343);
and U8418 (N_8418,N_8298,N_8281);
nor U8419 (N_8419,N_8260,N_8254);
xnor U8420 (N_8420,N_8284,N_8352);
or U8421 (N_8421,N_8332,N_8282);
or U8422 (N_8422,N_8336,N_8293);
nor U8423 (N_8423,N_8276,N_8321);
and U8424 (N_8424,N_8359,N_8268);
or U8425 (N_8425,N_8285,N_8328);
xor U8426 (N_8426,N_8349,N_8259);
nor U8427 (N_8427,N_8354,N_8283);
and U8428 (N_8428,N_8273,N_8342);
and U8429 (N_8429,N_8372,N_8348);
nand U8430 (N_8430,N_8317,N_8287);
or U8431 (N_8431,N_8269,N_8286);
or U8432 (N_8432,N_8340,N_8300);
nand U8433 (N_8433,N_8316,N_8351);
nor U8434 (N_8434,N_8366,N_8256);
nand U8435 (N_8435,N_8266,N_8292);
nand U8436 (N_8436,N_8262,N_8324);
and U8437 (N_8437,N_8274,N_8346);
and U8438 (N_8438,N_8279,N_8291);
xnor U8439 (N_8439,N_8338,N_8356);
or U8440 (N_8440,N_8259,N_8305);
and U8441 (N_8441,N_8368,N_8343);
or U8442 (N_8442,N_8266,N_8288);
xor U8443 (N_8443,N_8347,N_8265);
nor U8444 (N_8444,N_8361,N_8336);
xor U8445 (N_8445,N_8312,N_8372);
nor U8446 (N_8446,N_8367,N_8266);
xor U8447 (N_8447,N_8289,N_8309);
nand U8448 (N_8448,N_8257,N_8261);
and U8449 (N_8449,N_8270,N_8352);
nand U8450 (N_8450,N_8293,N_8268);
or U8451 (N_8451,N_8365,N_8318);
nor U8452 (N_8452,N_8284,N_8364);
nand U8453 (N_8453,N_8330,N_8262);
xor U8454 (N_8454,N_8302,N_8355);
nand U8455 (N_8455,N_8266,N_8282);
and U8456 (N_8456,N_8341,N_8280);
and U8457 (N_8457,N_8325,N_8337);
nor U8458 (N_8458,N_8372,N_8371);
or U8459 (N_8459,N_8276,N_8293);
nor U8460 (N_8460,N_8374,N_8319);
or U8461 (N_8461,N_8266,N_8284);
and U8462 (N_8462,N_8259,N_8346);
nor U8463 (N_8463,N_8286,N_8309);
nand U8464 (N_8464,N_8343,N_8324);
nand U8465 (N_8465,N_8358,N_8360);
nor U8466 (N_8466,N_8363,N_8274);
xnor U8467 (N_8467,N_8295,N_8281);
or U8468 (N_8468,N_8340,N_8315);
or U8469 (N_8469,N_8322,N_8344);
or U8470 (N_8470,N_8349,N_8316);
and U8471 (N_8471,N_8300,N_8282);
or U8472 (N_8472,N_8274,N_8288);
nor U8473 (N_8473,N_8370,N_8374);
or U8474 (N_8474,N_8259,N_8263);
nand U8475 (N_8475,N_8372,N_8283);
nand U8476 (N_8476,N_8333,N_8356);
or U8477 (N_8477,N_8313,N_8331);
nand U8478 (N_8478,N_8274,N_8339);
nor U8479 (N_8479,N_8370,N_8264);
nor U8480 (N_8480,N_8258,N_8272);
and U8481 (N_8481,N_8359,N_8307);
and U8482 (N_8482,N_8352,N_8372);
nor U8483 (N_8483,N_8362,N_8332);
nand U8484 (N_8484,N_8369,N_8344);
nand U8485 (N_8485,N_8258,N_8347);
and U8486 (N_8486,N_8309,N_8284);
nor U8487 (N_8487,N_8261,N_8300);
and U8488 (N_8488,N_8308,N_8274);
xnor U8489 (N_8489,N_8320,N_8351);
nor U8490 (N_8490,N_8325,N_8269);
and U8491 (N_8491,N_8304,N_8299);
nor U8492 (N_8492,N_8339,N_8283);
or U8493 (N_8493,N_8367,N_8329);
or U8494 (N_8494,N_8366,N_8339);
nor U8495 (N_8495,N_8357,N_8250);
xor U8496 (N_8496,N_8293,N_8326);
and U8497 (N_8497,N_8358,N_8369);
nand U8498 (N_8498,N_8366,N_8353);
and U8499 (N_8499,N_8290,N_8307);
and U8500 (N_8500,N_8474,N_8472);
nor U8501 (N_8501,N_8427,N_8492);
nor U8502 (N_8502,N_8449,N_8450);
nand U8503 (N_8503,N_8393,N_8421);
or U8504 (N_8504,N_8414,N_8455);
and U8505 (N_8505,N_8392,N_8398);
xnor U8506 (N_8506,N_8426,N_8476);
nand U8507 (N_8507,N_8378,N_8382);
and U8508 (N_8508,N_8428,N_8403);
nand U8509 (N_8509,N_8446,N_8442);
and U8510 (N_8510,N_8473,N_8420);
nor U8511 (N_8511,N_8431,N_8443);
xnor U8512 (N_8512,N_8439,N_8425);
or U8513 (N_8513,N_8485,N_8497);
and U8514 (N_8514,N_8409,N_8397);
xnor U8515 (N_8515,N_8433,N_8438);
nor U8516 (N_8516,N_8459,N_8386);
or U8517 (N_8517,N_8495,N_8417);
nand U8518 (N_8518,N_8379,N_8434);
and U8519 (N_8519,N_8375,N_8405);
nor U8520 (N_8520,N_8482,N_8488);
xnor U8521 (N_8521,N_8467,N_8387);
xor U8522 (N_8522,N_8452,N_8479);
or U8523 (N_8523,N_8404,N_8401);
and U8524 (N_8524,N_8462,N_8481);
nand U8525 (N_8525,N_8410,N_8498);
and U8526 (N_8526,N_8463,N_8395);
nand U8527 (N_8527,N_8470,N_8406);
nand U8528 (N_8528,N_8388,N_8454);
nor U8529 (N_8529,N_8453,N_8419);
or U8530 (N_8530,N_8432,N_8456);
or U8531 (N_8531,N_8412,N_8391);
nand U8532 (N_8532,N_8437,N_8486);
or U8533 (N_8533,N_8487,N_8468);
nand U8534 (N_8534,N_8376,N_8411);
xor U8535 (N_8535,N_8471,N_8491);
nand U8536 (N_8536,N_8494,N_8384);
nand U8537 (N_8537,N_8493,N_8483);
and U8538 (N_8538,N_8415,N_8416);
or U8539 (N_8539,N_8445,N_8390);
nand U8540 (N_8540,N_8385,N_8381);
nor U8541 (N_8541,N_8480,N_8413);
nor U8542 (N_8542,N_8461,N_8477);
nand U8543 (N_8543,N_8407,N_8464);
nor U8544 (N_8544,N_8469,N_8465);
xnor U8545 (N_8545,N_8475,N_8496);
and U8546 (N_8546,N_8389,N_8430);
or U8547 (N_8547,N_8441,N_8418);
nand U8548 (N_8548,N_8377,N_8478);
and U8549 (N_8549,N_8460,N_8444);
nand U8550 (N_8550,N_8394,N_8422);
nor U8551 (N_8551,N_8440,N_8424);
nand U8552 (N_8552,N_8396,N_8402);
and U8553 (N_8553,N_8490,N_8383);
nor U8554 (N_8554,N_8457,N_8399);
xor U8555 (N_8555,N_8408,N_8484);
and U8556 (N_8556,N_8458,N_8380);
nor U8557 (N_8557,N_8400,N_8499);
nand U8558 (N_8558,N_8423,N_8451);
and U8559 (N_8559,N_8447,N_8429);
and U8560 (N_8560,N_8466,N_8436);
nand U8561 (N_8561,N_8489,N_8435);
nor U8562 (N_8562,N_8448,N_8437);
nor U8563 (N_8563,N_8429,N_8438);
nor U8564 (N_8564,N_8474,N_8470);
and U8565 (N_8565,N_8463,N_8430);
nand U8566 (N_8566,N_8442,N_8428);
nor U8567 (N_8567,N_8377,N_8423);
and U8568 (N_8568,N_8452,N_8428);
and U8569 (N_8569,N_8440,N_8485);
and U8570 (N_8570,N_8406,N_8387);
or U8571 (N_8571,N_8456,N_8453);
or U8572 (N_8572,N_8423,N_8399);
nor U8573 (N_8573,N_8435,N_8466);
and U8574 (N_8574,N_8400,N_8462);
and U8575 (N_8575,N_8422,N_8387);
or U8576 (N_8576,N_8499,N_8489);
and U8577 (N_8577,N_8486,N_8457);
and U8578 (N_8578,N_8499,N_8376);
or U8579 (N_8579,N_8377,N_8433);
and U8580 (N_8580,N_8441,N_8491);
nand U8581 (N_8581,N_8454,N_8384);
or U8582 (N_8582,N_8414,N_8423);
nor U8583 (N_8583,N_8414,N_8463);
or U8584 (N_8584,N_8476,N_8439);
and U8585 (N_8585,N_8417,N_8432);
or U8586 (N_8586,N_8473,N_8459);
nand U8587 (N_8587,N_8445,N_8382);
nor U8588 (N_8588,N_8388,N_8434);
xnor U8589 (N_8589,N_8405,N_8430);
nor U8590 (N_8590,N_8464,N_8380);
or U8591 (N_8591,N_8424,N_8387);
nor U8592 (N_8592,N_8376,N_8475);
nor U8593 (N_8593,N_8470,N_8383);
nor U8594 (N_8594,N_8380,N_8432);
nor U8595 (N_8595,N_8484,N_8491);
and U8596 (N_8596,N_8480,N_8414);
nor U8597 (N_8597,N_8432,N_8490);
or U8598 (N_8598,N_8424,N_8389);
and U8599 (N_8599,N_8441,N_8498);
or U8600 (N_8600,N_8482,N_8377);
or U8601 (N_8601,N_8449,N_8377);
or U8602 (N_8602,N_8398,N_8469);
and U8603 (N_8603,N_8405,N_8479);
xor U8604 (N_8604,N_8414,N_8401);
nand U8605 (N_8605,N_8476,N_8414);
nor U8606 (N_8606,N_8455,N_8420);
xor U8607 (N_8607,N_8481,N_8450);
nor U8608 (N_8608,N_8481,N_8437);
and U8609 (N_8609,N_8430,N_8436);
and U8610 (N_8610,N_8394,N_8388);
nand U8611 (N_8611,N_8399,N_8475);
nor U8612 (N_8612,N_8405,N_8496);
or U8613 (N_8613,N_8489,N_8425);
or U8614 (N_8614,N_8444,N_8397);
nor U8615 (N_8615,N_8376,N_8391);
nor U8616 (N_8616,N_8391,N_8440);
or U8617 (N_8617,N_8463,N_8392);
and U8618 (N_8618,N_8437,N_8465);
nand U8619 (N_8619,N_8444,N_8492);
or U8620 (N_8620,N_8419,N_8474);
or U8621 (N_8621,N_8459,N_8393);
and U8622 (N_8622,N_8425,N_8453);
and U8623 (N_8623,N_8425,N_8496);
or U8624 (N_8624,N_8499,N_8408);
and U8625 (N_8625,N_8526,N_8522);
or U8626 (N_8626,N_8502,N_8572);
or U8627 (N_8627,N_8614,N_8509);
xnor U8628 (N_8628,N_8547,N_8503);
nand U8629 (N_8629,N_8543,N_8604);
and U8630 (N_8630,N_8546,N_8542);
or U8631 (N_8631,N_8573,N_8527);
nor U8632 (N_8632,N_8560,N_8515);
and U8633 (N_8633,N_8574,N_8562);
or U8634 (N_8634,N_8514,N_8592);
nand U8635 (N_8635,N_8508,N_8584);
and U8636 (N_8636,N_8511,N_8611);
nand U8637 (N_8637,N_8599,N_8519);
nor U8638 (N_8638,N_8556,N_8510);
and U8639 (N_8639,N_8536,N_8620);
nand U8640 (N_8640,N_8597,N_8593);
and U8641 (N_8641,N_8587,N_8533);
and U8642 (N_8642,N_8512,N_8610);
or U8643 (N_8643,N_8532,N_8529);
xnor U8644 (N_8644,N_8571,N_8605);
nor U8645 (N_8645,N_8557,N_8570);
or U8646 (N_8646,N_8606,N_8538);
nor U8647 (N_8647,N_8521,N_8615);
nand U8648 (N_8648,N_8520,N_8530);
or U8649 (N_8649,N_8551,N_8579);
nand U8650 (N_8650,N_8565,N_8517);
and U8651 (N_8651,N_8505,N_8552);
nand U8652 (N_8652,N_8545,N_8567);
nor U8653 (N_8653,N_8554,N_8589);
and U8654 (N_8654,N_8504,N_8612);
or U8655 (N_8655,N_8535,N_8506);
nor U8656 (N_8656,N_8590,N_8525);
and U8657 (N_8657,N_8564,N_8539);
or U8658 (N_8658,N_8617,N_8588);
or U8659 (N_8659,N_8623,N_8534);
nand U8660 (N_8660,N_8583,N_8576);
nand U8661 (N_8661,N_8524,N_8523);
xnor U8662 (N_8662,N_8501,N_8598);
nor U8663 (N_8663,N_8553,N_8548);
nand U8664 (N_8664,N_8603,N_8544);
nand U8665 (N_8665,N_8582,N_8600);
and U8666 (N_8666,N_8607,N_8578);
nand U8667 (N_8667,N_8500,N_8550);
nand U8668 (N_8668,N_8537,N_8566);
nor U8669 (N_8669,N_8575,N_8531);
and U8670 (N_8670,N_8595,N_8540);
or U8671 (N_8671,N_8549,N_8561);
nor U8672 (N_8672,N_8594,N_8580);
and U8673 (N_8673,N_8541,N_8601);
nor U8674 (N_8674,N_8609,N_8507);
or U8675 (N_8675,N_8621,N_8563);
nand U8676 (N_8676,N_8581,N_8585);
or U8677 (N_8677,N_8596,N_8516);
and U8678 (N_8678,N_8619,N_8602);
nand U8679 (N_8679,N_8528,N_8569);
and U8680 (N_8680,N_8616,N_8622);
and U8681 (N_8681,N_8613,N_8591);
xor U8682 (N_8682,N_8558,N_8577);
and U8683 (N_8683,N_8518,N_8586);
nand U8684 (N_8684,N_8608,N_8555);
nor U8685 (N_8685,N_8513,N_8624);
or U8686 (N_8686,N_8568,N_8559);
and U8687 (N_8687,N_8618,N_8580);
or U8688 (N_8688,N_8586,N_8561);
nor U8689 (N_8689,N_8523,N_8600);
nor U8690 (N_8690,N_8606,N_8590);
and U8691 (N_8691,N_8592,N_8545);
nand U8692 (N_8692,N_8574,N_8618);
and U8693 (N_8693,N_8517,N_8562);
nor U8694 (N_8694,N_8584,N_8553);
or U8695 (N_8695,N_8610,N_8534);
or U8696 (N_8696,N_8503,N_8535);
nor U8697 (N_8697,N_8565,N_8581);
xor U8698 (N_8698,N_8516,N_8524);
and U8699 (N_8699,N_8599,N_8503);
and U8700 (N_8700,N_8603,N_8613);
and U8701 (N_8701,N_8528,N_8577);
and U8702 (N_8702,N_8601,N_8591);
or U8703 (N_8703,N_8516,N_8620);
nand U8704 (N_8704,N_8555,N_8621);
nand U8705 (N_8705,N_8545,N_8591);
or U8706 (N_8706,N_8595,N_8624);
and U8707 (N_8707,N_8581,N_8505);
and U8708 (N_8708,N_8569,N_8502);
nand U8709 (N_8709,N_8556,N_8554);
nor U8710 (N_8710,N_8603,N_8561);
or U8711 (N_8711,N_8609,N_8549);
nor U8712 (N_8712,N_8556,N_8583);
and U8713 (N_8713,N_8590,N_8597);
or U8714 (N_8714,N_8578,N_8603);
or U8715 (N_8715,N_8599,N_8536);
and U8716 (N_8716,N_8605,N_8559);
and U8717 (N_8717,N_8586,N_8567);
nand U8718 (N_8718,N_8555,N_8612);
nand U8719 (N_8719,N_8567,N_8522);
nor U8720 (N_8720,N_8501,N_8581);
nand U8721 (N_8721,N_8515,N_8618);
or U8722 (N_8722,N_8561,N_8621);
nand U8723 (N_8723,N_8506,N_8582);
nor U8724 (N_8724,N_8605,N_8555);
or U8725 (N_8725,N_8528,N_8504);
nand U8726 (N_8726,N_8609,N_8558);
and U8727 (N_8727,N_8538,N_8598);
nand U8728 (N_8728,N_8612,N_8597);
and U8729 (N_8729,N_8539,N_8583);
nand U8730 (N_8730,N_8610,N_8578);
and U8731 (N_8731,N_8590,N_8624);
nor U8732 (N_8732,N_8570,N_8555);
or U8733 (N_8733,N_8519,N_8598);
nor U8734 (N_8734,N_8599,N_8540);
or U8735 (N_8735,N_8504,N_8542);
nor U8736 (N_8736,N_8558,N_8567);
nand U8737 (N_8737,N_8593,N_8512);
or U8738 (N_8738,N_8549,N_8611);
and U8739 (N_8739,N_8507,N_8571);
or U8740 (N_8740,N_8584,N_8506);
xor U8741 (N_8741,N_8591,N_8544);
nand U8742 (N_8742,N_8509,N_8525);
and U8743 (N_8743,N_8525,N_8502);
nor U8744 (N_8744,N_8599,N_8614);
nand U8745 (N_8745,N_8511,N_8537);
or U8746 (N_8746,N_8580,N_8615);
xnor U8747 (N_8747,N_8608,N_8566);
nand U8748 (N_8748,N_8523,N_8585);
or U8749 (N_8749,N_8512,N_8502);
and U8750 (N_8750,N_8715,N_8655);
nand U8751 (N_8751,N_8685,N_8739);
nand U8752 (N_8752,N_8703,N_8707);
nand U8753 (N_8753,N_8690,N_8675);
xnor U8754 (N_8754,N_8664,N_8700);
and U8755 (N_8755,N_8629,N_8696);
or U8756 (N_8756,N_8633,N_8747);
nand U8757 (N_8757,N_8738,N_8639);
xor U8758 (N_8758,N_8745,N_8632);
nand U8759 (N_8759,N_8638,N_8673);
nand U8760 (N_8760,N_8714,N_8677);
and U8761 (N_8761,N_8669,N_8720);
xor U8762 (N_8762,N_8708,N_8680);
and U8763 (N_8763,N_8697,N_8736);
and U8764 (N_8764,N_8647,N_8705);
nor U8765 (N_8765,N_8702,N_8635);
and U8766 (N_8766,N_8695,N_8671);
nor U8767 (N_8767,N_8627,N_8746);
or U8768 (N_8768,N_8744,N_8688);
nor U8769 (N_8769,N_8676,N_8704);
or U8770 (N_8770,N_8734,N_8656);
xnor U8771 (N_8771,N_8661,N_8733);
or U8772 (N_8772,N_8686,N_8725);
nand U8773 (N_8773,N_8645,N_8640);
and U8774 (N_8774,N_8653,N_8679);
nor U8775 (N_8775,N_8728,N_8730);
or U8776 (N_8776,N_8654,N_8735);
or U8777 (N_8777,N_8668,N_8648);
nand U8778 (N_8778,N_8709,N_8699);
xnor U8779 (N_8779,N_8643,N_8634);
and U8780 (N_8780,N_8716,N_8749);
nand U8781 (N_8781,N_8641,N_8748);
nor U8782 (N_8782,N_8722,N_8742);
nand U8783 (N_8783,N_8717,N_8663);
or U8784 (N_8784,N_8689,N_8678);
or U8785 (N_8785,N_8682,N_8710);
or U8786 (N_8786,N_8642,N_8659);
xor U8787 (N_8787,N_8683,N_8681);
nor U8788 (N_8788,N_8652,N_8692);
and U8789 (N_8789,N_8672,N_8646);
nand U8790 (N_8790,N_8724,N_8694);
nor U8791 (N_8791,N_8729,N_8674);
or U8792 (N_8792,N_8666,N_8636);
xnor U8793 (N_8793,N_8665,N_8660);
and U8794 (N_8794,N_8732,N_8684);
or U8795 (N_8795,N_8651,N_8718);
nor U8796 (N_8796,N_8737,N_8698);
nor U8797 (N_8797,N_8691,N_8670);
xor U8798 (N_8798,N_8626,N_8726);
and U8799 (N_8799,N_8657,N_8667);
nor U8800 (N_8800,N_8723,N_8658);
or U8801 (N_8801,N_8662,N_8628);
or U8802 (N_8802,N_8711,N_8706);
nor U8803 (N_8803,N_8687,N_8740);
and U8804 (N_8804,N_8701,N_8741);
nor U8805 (N_8805,N_8721,N_8731);
xor U8806 (N_8806,N_8644,N_8630);
and U8807 (N_8807,N_8743,N_8693);
nor U8808 (N_8808,N_8631,N_8727);
or U8809 (N_8809,N_8625,N_8650);
and U8810 (N_8810,N_8719,N_8649);
and U8811 (N_8811,N_8713,N_8637);
and U8812 (N_8812,N_8712,N_8714);
nor U8813 (N_8813,N_8698,N_8693);
or U8814 (N_8814,N_8719,N_8723);
nor U8815 (N_8815,N_8673,N_8683);
and U8816 (N_8816,N_8648,N_8729);
or U8817 (N_8817,N_8682,N_8677);
nand U8818 (N_8818,N_8733,N_8654);
nand U8819 (N_8819,N_8664,N_8657);
xnor U8820 (N_8820,N_8638,N_8745);
or U8821 (N_8821,N_8747,N_8636);
nand U8822 (N_8822,N_8735,N_8725);
or U8823 (N_8823,N_8631,N_8710);
or U8824 (N_8824,N_8688,N_8663);
nand U8825 (N_8825,N_8657,N_8627);
nor U8826 (N_8826,N_8707,N_8666);
and U8827 (N_8827,N_8675,N_8631);
and U8828 (N_8828,N_8661,N_8702);
nor U8829 (N_8829,N_8683,N_8730);
xor U8830 (N_8830,N_8719,N_8736);
and U8831 (N_8831,N_8703,N_8705);
nand U8832 (N_8832,N_8656,N_8720);
or U8833 (N_8833,N_8714,N_8682);
nor U8834 (N_8834,N_8710,N_8660);
xnor U8835 (N_8835,N_8711,N_8690);
nand U8836 (N_8836,N_8739,N_8724);
or U8837 (N_8837,N_8724,N_8700);
and U8838 (N_8838,N_8715,N_8673);
xnor U8839 (N_8839,N_8727,N_8646);
and U8840 (N_8840,N_8641,N_8742);
and U8841 (N_8841,N_8707,N_8745);
and U8842 (N_8842,N_8669,N_8633);
nor U8843 (N_8843,N_8709,N_8729);
nand U8844 (N_8844,N_8735,N_8687);
xnor U8845 (N_8845,N_8707,N_8702);
nand U8846 (N_8846,N_8693,N_8625);
nand U8847 (N_8847,N_8656,N_8652);
and U8848 (N_8848,N_8718,N_8695);
nor U8849 (N_8849,N_8648,N_8670);
or U8850 (N_8850,N_8686,N_8649);
nand U8851 (N_8851,N_8704,N_8721);
nand U8852 (N_8852,N_8677,N_8727);
nand U8853 (N_8853,N_8642,N_8675);
nand U8854 (N_8854,N_8651,N_8668);
nor U8855 (N_8855,N_8727,N_8732);
and U8856 (N_8856,N_8665,N_8698);
nand U8857 (N_8857,N_8713,N_8729);
nand U8858 (N_8858,N_8718,N_8700);
xor U8859 (N_8859,N_8651,N_8653);
or U8860 (N_8860,N_8733,N_8722);
or U8861 (N_8861,N_8699,N_8691);
nand U8862 (N_8862,N_8684,N_8631);
nor U8863 (N_8863,N_8683,N_8670);
and U8864 (N_8864,N_8630,N_8707);
nand U8865 (N_8865,N_8650,N_8720);
nor U8866 (N_8866,N_8683,N_8734);
nand U8867 (N_8867,N_8692,N_8686);
nand U8868 (N_8868,N_8715,N_8686);
nor U8869 (N_8869,N_8644,N_8696);
nand U8870 (N_8870,N_8661,N_8675);
nor U8871 (N_8871,N_8697,N_8671);
nand U8872 (N_8872,N_8748,N_8706);
and U8873 (N_8873,N_8659,N_8626);
nand U8874 (N_8874,N_8629,N_8746);
and U8875 (N_8875,N_8854,N_8814);
and U8876 (N_8876,N_8873,N_8813);
nor U8877 (N_8877,N_8797,N_8829);
xor U8878 (N_8878,N_8780,N_8790);
nor U8879 (N_8879,N_8799,N_8754);
and U8880 (N_8880,N_8807,N_8871);
nor U8881 (N_8881,N_8779,N_8784);
and U8882 (N_8882,N_8770,N_8847);
or U8883 (N_8883,N_8806,N_8768);
and U8884 (N_8884,N_8809,N_8793);
xnor U8885 (N_8885,N_8822,N_8868);
nor U8886 (N_8886,N_8838,N_8850);
or U8887 (N_8887,N_8858,N_8802);
and U8888 (N_8888,N_8837,N_8774);
nand U8889 (N_8889,N_8843,N_8817);
nor U8890 (N_8890,N_8821,N_8798);
nor U8891 (N_8891,N_8846,N_8786);
xor U8892 (N_8892,N_8766,N_8763);
nor U8893 (N_8893,N_8787,N_8783);
xnor U8894 (N_8894,N_8866,N_8857);
nor U8895 (N_8895,N_8864,N_8848);
nand U8896 (N_8896,N_8757,N_8870);
and U8897 (N_8897,N_8835,N_8861);
and U8898 (N_8898,N_8859,N_8800);
nor U8899 (N_8899,N_8855,N_8791);
nand U8900 (N_8900,N_8831,N_8825);
or U8901 (N_8901,N_8771,N_8767);
nand U8902 (N_8902,N_8853,N_8820);
and U8903 (N_8903,N_8795,N_8867);
and U8904 (N_8904,N_8863,N_8874);
xnor U8905 (N_8905,N_8789,N_8862);
and U8906 (N_8906,N_8788,N_8801);
xnor U8907 (N_8907,N_8851,N_8823);
nor U8908 (N_8908,N_8852,N_8812);
nor U8909 (N_8909,N_8815,N_8844);
nor U8910 (N_8910,N_8777,N_8839);
nor U8911 (N_8911,N_8775,N_8808);
nand U8912 (N_8912,N_8830,N_8832);
and U8913 (N_8913,N_8872,N_8794);
xnor U8914 (N_8914,N_8764,N_8824);
nand U8915 (N_8915,N_8842,N_8841);
nor U8916 (N_8916,N_8833,N_8865);
nor U8917 (N_8917,N_8772,N_8758);
and U8918 (N_8918,N_8828,N_8869);
nand U8919 (N_8919,N_8755,N_8804);
or U8920 (N_8920,N_8826,N_8785);
or U8921 (N_8921,N_8781,N_8827);
nand U8922 (N_8922,N_8849,N_8818);
or U8923 (N_8923,N_8845,N_8792);
and U8924 (N_8924,N_8753,N_8759);
xor U8925 (N_8925,N_8760,N_8836);
or U8926 (N_8926,N_8778,N_8776);
nand U8927 (N_8927,N_8752,N_8782);
and U8928 (N_8928,N_8840,N_8751);
xnor U8929 (N_8929,N_8860,N_8769);
or U8930 (N_8930,N_8816,N_8819);
and U8931 (N_8931,N_8765,N_8803);
xnor U8932 (N_8932,N_8805,N_8856);
nand U8933 (N_8933,N_8773,N_8761);
nor U8934 (N_8934,N_8810,N_8762);
and U8935 (N_8935,N_8756,N_8811);
nand U8936 (N_8936,N_8750,N_8834);
nor U8937 (N_8937,N_8796,N_8857);
xor U8938 (N_8938,N_8814,N_8793);
and U8939 (N_8939,N_8784,N_8865);
or U8940 (N_8940,N_8819,N_8809);
xnor U8941 (N_8941,N_8860,N_8812);
nor U8942 (N_8942,N_8867,N_8804);
nor U8943 (N_8943,N_8805,N_8769);
or U8944 (N_8944,N_8826,N_8792);
nand U8945 (N_8945,N_8778,N_8762);
and U8946 (N_8946,N_8854,N_8770);
or U8947 (N_8947,N_8812,N_8801);
and U8948 (N_8948,N_8750,N_8849);
and U8949 (N_8949,N_8856,N_8767);
nand U8950 (N_8950,N_8768,N_8805);
or U8951 (N_8951,N_8866,N_8761);
or U8952 (N_8952,N_8780,N_8756);
nor U8953 (N_8953,N_8759,N_8783);
nand U8954 (N_8954,N_8868,N_8837);
and U8955 (N_8955,N_8840,N_8843);
and U8956 (N_8956,N_8845,N_8867);
nand U8957 (N_8957,N_8807,N_8822);
and U8958 (N_8958,N_8863,N_8792);
xnor U8959 (N_8959,N_8759,N_8790);
nand U8960 (N_8960,N_8779,N_8781);
nand U8961 (N_8961,N_8864,N_8866);
and U8962 (N_8962,N_8784,N_8845);
nor U8963 (N_8963,N_8758,N_8770);
nor U8964 (N_8964,N_8835,N_8859);
and U8965 (N_8965,N_8819,N_8821);
nand U8966 (N_8966,N_8861,N_8756);
nand U8967 (N_8967,N_8866,N_8770);
and U8968 (N_8968,N_8774,N_8867);
or U8969 (N_8969,N_8810,N_8852);
nand U8970 (N_8970,N_8765,N_8872);
nand U8971 (N_8971,N_8839,N_8766);
or U8972 (N_8972,N_8815,N_8841);
or U8973 (N_8973,N_8813,N_8762);
nor U8974 (N_8974,N_8873,N_8756);
nor U8975 (N_8975,N_8785,N_8755);
or U8976 (N_8976,N_8865,N_8829);
or U8977 (N_8977,N_8824,N_8750);
or U8978 (N_8978,N_8814,N_8754);
xnor U8979 (N_8979,N_8843,N_8865);
or U8980 (N_8980,N_8824,N_8857);
nand U8981 (N_8981,N_8761,N_8840);
nor U8982 (N_8982,N_8797,N_8858);
xnor U8983 (N_8983,N_8843,N_8805);
nand U8984 (N_8984,N_8857,N_8773);
and U8985 (N_8985,N_8871,N_8772);
and U8986 (N_8986,N_8861,N_8803);
nor U8987 (N_8987,N_8808,N_8816);
or U8988 (N_8988,N_8807,N_8866);
nor U8989 (N_8989,N_8856,N_8784);
nand U8990 (N_8990,N_8761,N_8865);
and U8991 (N_8991,N_8866,N_8833);
or U8992 (N_8992,N_8821,N_8843);
nor U8993 (N_8993,N_8785,N_8820);
nand U8994 (N_8994,N_8767,N_8807);
and U8995 (N_8995,N_8858,N_8833);
nor U8996 (N_8996,N_8758,N_8805);
xor U8997 (N_8997,N_8838,N_8767);
nor U8998 (N_8998,N_8873,N_8751);
nand U8999 (N_8999,N_8870,N_8866);
xor U9000 (N_9000,N_8945,N_8996);
and U9001 (N_9001,N_8989,N_8986);
nand U9002 (N_9002,N_8944,N_8993);
or U9003 (N_9003,N_8902,N_8886);
nand U9004 (N_9004,N_8966,N_8925);
nor U9005 (N_9005,N_8958,N_8878);
nor U9006 (N_9006,N_8926,N_8938);
and U9007 (N_9007,N_8943,N_8909);
nand U9008 (N_9008,N_8931,N_8968);
nand U9009 (N_9009,N_8877,N_8954);
nand U9010 (N_9010,N_8880,N_8948);
and U9011 (N_9011,N_8881,N_8899);
nand U9012 (N_9012,N_8999,N_8947);
xnor U9013 (N_9013,N_8949,N_8906);
nand U9014 (N_9014,N_8898,N_8932);
nand U9015 (N_9015,N_8981,N_8942);
or U9016 (N_9016,N_8893,N_8919);
nand U9017 (N_9017,N_8978,N_8963);
nor U9018 (N_9018,N_8875,N_8888);
xnor U9019 (N_9019,N_8983,N_8971);
or U9020 (N_9020,N_8998,N_8951);
nor U9021 (N_9021,N_8905,N_8959);
and U9022 (N_9022,N_8937,N_8972);
nor U9023 (N_9023,N_8992,N_8997);
nand U9024 (N_9024,N_8914,N_8930);
and U9025 (N_9025,N_8918,N_8962);
nor U9026 (N_9026,N_8911,N_8979);
nor U9027 (N_9027,N_8900,N_8913);
nor U9028 (N_9028,N_8923,N_8892);
and U9029 (N_9029,N_8967,N_8916);
or U9030 (N_9030,N_8912,N_8922);
and U9031 (N_9031,N_8969,N_8936);
and U9032 (N_9032,N_8953,N_8955);
nor U9033 (N_9033,N_8946,N_8987);
nor U9034 (N_9034,N_8928,N_8897);
and U9035 (N_9035,N_8940,N_8920);
nor U9036 (N_9036,N_8974,N_8934);
nand U9037 (N_9037,N_8984,N_8910);
nor U9038 (N_9038,N_8884,N_8895);
or U9039 (N_9039,N_8917,N_8883);
nor U9040 (N_9040,N_8935,N_8896);
and U9041 (N_9041,N_8973,N_8879);
xnor U9042 (N_9042,N_8939,N_8876);
nand U9043 (N_9043,N_8929,N_8995);
nor U9044 (N_9044,N_8921,N_8982);
and U9045 (N_9045,N_8891,N_8915);
or U9046 (N_9046,N_8994,N_8950);
nor U9047 (N_9047,N_8887,N_8890);
nand U9048 (N_9048,N_8964,N_8960);
or U9049 (N_9049,N_8907,N_8961);
xnor U9050 (N_9050,N_8991,N_8933);
or U9051 (N_9051,N_8924,N_8894);
and U9052 (N_9052,N_8903,N_8957);
nor U9053 (N_9053,N_8882,N_8952);
nor U9054 (N_9054,N_8980,N_8885);
nand U9055 (N_9055,N_8956,N_8904);
nor U9056 (N_9056,N_8976,N_8985);
nor U9057 (N_9057,N_8990,N_8988);
and U9058 (N_9058,N_8889,N_8901);
nand U9059 (N_9059,N_8975,N_8908);
nor U9060 (N_9060,N_8927,N_8977);
and U9061 (N_9061,N_8965,N_8941);
or U9062 (N_9062,N_8970,N_8996);
and U9063 (N_9063,N_8895,N_8878);
or U9064 (N_9064,N_8907,N_8994);
and U9065 (N_9065,N_8886,N_8889);
nor U9066 (N_9066,N_8936,N_8950);
and U9067 (N_9067,N_8939,N_8942);
or U9068 (N_9068,N_8927,N_8926);
or U9069 (N_9069,N_8984,N_8945);
nand U9070 (N_9070,N_8888,N_8986);
and U9071 (N_9071,N_8998,N_8993);
nor U9072 (N_9072,N_8976,N_8887);
or U9073 (N_9073,N_8930,N_8986);
and U9074 (N_9074,N_8887,N_8939);
or U9075 (N_9075,N_8918,N_8998);
xor U9076 (N_9076,N_8905,N_8900);
and U9077 (N_9077,N_8941,N_8903);
nor U9078 (N_9078,N_8897,N_8985);
nand U9079 (N_9079,N_8970,N_8971);
xor U9080 (N_9080,N_8926,N_8878);
nor U9081 (N_9081,N_8999,N_8983);
nor U9082 (N_9082,N_8946,N_8977);
nand U9083 (N_9083,N_8958,N_8923);
and U9084 (N_9084,N_8944,N_8997);
nor U9085 (N_9085,N_8910,N_8912);
or U9086 (N_9086,N_8876,N_8981);
xnor U9087 (N_9087,N_8897,N_8982);
nand U9088 (N_9088,N_8899,N_8976);
or U9089 (N_9089,N_8905,N_8890);
and U9090 (N_9090,N_8989,N_8898);
xnor U9091 (N_9091,N_8900,N_8908);
and U9092 (N_9092,N_8931,N_8973);
and U9093 (N_9093,N_8988,N_8890);
nor U9094 (N_9094,N_8974,N_8880);
nand U9095 (N_9095,N_8985,N_8990);
nand U9096 (N_9096,N_8986,N_8942);
nand U9097 (N_9097,N_8973,N_8933);
and U9098 (N_9098,N_8884,N_8957);
xnor U9099 (N_9099,N_8910,N_8976);
nor U9100 (N_9100,N_8963,N_8994);
or U9101 (N_9101,N_8928,N_8908);
nor U9102 (N_9102,N_8999,N_8992);
and U9103 (N_9103,N_8931,N_8994);
nor U9104 (N_9104,N_8875,N_8878);
xor U9105 (N_9105,N_8981,N_8940);
nand U9106 (N_9106,N_8950,N_8995);
nor U9107 (N_9107,N_8976,N_8919);
or U9108 (N_9108,N_8891,N_8884);
or U9109 (N_9109,N_8896,N_8964);
nor U9110 (N_9110,N_8924,N_8937);
or U9111 (N_9111,N_8906,N_8931);
or U9112 (N_9112,N_8949,N_8952);
nand U9113 (N_9113,N_8991,N_8974);
or U9114 (N_9114,N_8903,N_8925);
or U9115 (N_9115,N_8896,N_8978);
nor U9116 (N_9116,N_8879,N_8877);
nand U9117 (N_9117,N_8899,N_8883);
and U9118 (N_9118,N_8985,N_8943);
nor U9119 (N_9119,N_8934,N_8963);
nand U9120 (N_9120,N_8881,N_8924);
nand U9121 (N_9121,N_8920,N_8897);
or U9122 (N_9122,N_8932,N_8901);
nor U9123 (N_9123,N_8909,N_8955);
and U9124 (N_9124,N_8957,N_8917);
nor U9125 (N_9125,N_9029,N_9117);
or U9126 (N_9126,N_9017,N_9062);
xor U9127 (N_9127,N_9119,N_9058);
nand U9128 (N_9128,N_9065,N_9122);
or U9129 (N_9129,N_9104,N_9099);
nand U9130 (N_9130,N_9024,N_9032);
nand U9131 (N_9131,N_9098,N_9023);
and U9132 (N_9132,N_9038,N_9041);
nand U9133 (N_9133,N_9031,N_9107);
nand U9134 (N_9134,N_9069,N_9025);
or U9135 (N_9135,N_9063,N_9040);
and U9136 (N_9136,N_9015,N_9042);
or U9137 (N_9137,N_9039,N_9090);
nor U9138 (N_9138,N_9060,N_9114);
or U9139 (N_9139,N_9046,N_9050);
nor U9140 (N_9140,N_9115,N_9066);
and U9141 (N_9141,N_9001,N_9006);
and U9142 (N_9142,N_9085,N_9079);
xor U9143 (N_9143,N_9100,N_9056);
nor U9144 (N_9144,N_9088,N_9086);
and U9145 (N_9145,N_9000,N_9070);
xnor U9146 (N_9146,N_9103,N_9078);
nand U9147 (N_9147,N_9097,N_9013);
and U9148 (N_9148,N_9022,N_9089);
and U9149 (N_9149,N_9077,N_9095);
or U9150 (N_9150,N_9035,N_9048);
xor U9151 (N_9151,N_9003,N_9053);
nand U9152 (N_9152,N_9082,N_9118);
and U9153 (N_9153,N_9034,N_9037);
or U9154 (N_9154,N_9123,N_9054);
or U9155 (N_9155,N_9061,N_9110);
and U9156 (N_9156,N_9074,N_9047);
or U9157 (N_9157,N_9021,N_9018);
or U9158 (N_9158,N_9111,N_9059);
nor U9159 (N_9159,N_9009,N_9076);
xor U9160 (N_9160,N_9092,N_9067);
and U9161 (N_9161,N_9108,N_9084);
xnor U9162 (N_9162,N_9087,N_9036);
nand U9163 (N_9163,N_9030,N_9045);
nand U9164 (N_9164,N_9071,N_9094);
nor U9165 (N_9165,N_9051,N_9052);
or U9166 (N_9166,N_9105,N_9120);
nand U9167 (N_9167,N_9101,N_9102);
and U9168 (N_9168,N_9055,N_9007);
nor U9169 (N_9169,N_9106,N_9116);
nand U9170 (N_9170,N_9008,N_9020);
or U9171 (N_9171,N_9010,N_9049);
nand U9172 (N_9172,N_9083,N_9112);
nor U9173 (N_9173,N_9109,N_9080);
nand U9174 (N_9174,N_9091,N_9124);
xor U9175 (N_9175,N_9004,N_9028);
nand U9176 (N_9176,N_9026,N_9005);
xnor U9177 (N_9177,N_9081,N_9012);
nor U9178 (N_9178,N_9019,N_9113);
nand U9179 (N_9179,N_9068,N_9093);
nand U9180 (N_9180,N_9044,N_9064);
xnor U9181 (N_9181,N_9043,N_9027);
xor U9182 (N_9182,N_9033,N_9075);
and U9183 (N_9183,N_9073,N_9016);
nand U9184 (N_9184,N_9002,N_9121);
or U9185 (N_9185,N_9072,N_9096);
nor U9186 (N_9186,N_9057,N_9011);
or U9187 (N_9187,N_9014,N_9021);
nor U9188 (N_9188,N_9094,N_9003);
xnor U9189 (N_9189,N_9031,N_9109);
nand U9190 (N_9190,N_9027,N_9023);
and U9191 (N_9191,N_9115,N_9036);
nand U9192 (N_9192,N_9108,N_9072);
or U9193 (N_9193,N_9052,N_9015);
nand U9194 (N_9194,N_9050,N_9058);
nand U9195 (N_9195,N_9032,N_9059);
and U9196 (N_9196,N_9037,N_9033);
nor U9197 (N_9197,N_9060,N_9020);
or U9198 (N_9198,N_9123,N_9104);
nor U9199 (N_9199,N_9001,N_9088);
or U9200 (N_9200,N_9120,N_9027);
nand U9201 (N_9201,N_9039,N_9010);
and U9202 (N_9202,N_9027,N_9049);
or U9203 (N_9203,N_9058,N_9016);
nor U9204 (N_9204,N_9104,N_9033);
nor U9205 (N_9205,N_9095,N_9083);
nor U9206 (N_9206,N_9013,N_9071);
nand U9207 (N_9207,N_9079,N_9077);
nor U9208 (N_9208,N_9030,N_9037);
xnor U9209 (N_9209,N_9005,N_9035);
nor U9210 (N_9210,N_9093,N_9057);
nand U9211 (N_9211,N_9020,N_9021);
and U9212 (N_9212,N_9030,N_9049);
nand U9213 (N_9213,N_9029,N_9027);
or U9214 (N_9214,N_9054,N_9069);
nand U9215 (N_9215,N_9085,N_9078);
nor U9216 (N_9216,N_9019,N_9010);
nand U9217 (N_9217,N_9000,N_9014);
or U9218 (N_9218,N_9079,N_9057);
and U9219 (N_9219,N_9045,N_9112);
nand U9220 (N_9220,N_9045,N_9099);
nand U9221 (N_9221,N_9089,N_9086);
nand U9222 (N_9222,N_9063,N_9008);
nand U9223 (N_9223,N_9051,N_9014);
nand U9224 (N_9224,N_9022,N_9027);
xor U9225 (N_9225,N_9044,N_9095);
or U9226 (N_9226,N_9020,N_9039);
nor U9227 (N_9227,N_9081,N_9108);
nor U9228 (N_9228,N_9038,N_9045);
or U9229 (N_9229,N_9036,N_9102);
and U9230 (N_9230,N_9047,N_9039);
nor U9231 (N_9231,N_9073,N_9047);
or U9232 (N_9232,N_9060,N_9021);
nand U9233 (N_9233,N_9061,N_9007);
xor U9234 (N_9234,N_9087,N_9084);
nor U9235 (N_9235,N_9018,N_9102);
nand U9236 (N_9236,N_9101,N_9073);
and U9237 (N_9237,N_9046,N_9112);
nand U9238 (N_9238,N_9031,N_9082);
nor U9239 (N_9239,N_9118,N_9116);
nand U9240 (N_9240,N_9111,N_9090);
nand U9241 (N_9241,N_9007,N_9116);
and U9242 (N_9242,N_9045,N_9120);
nor U9243 (N_9243,N_9029,N_9019);
and U9244 (N_9244,N_9005,N_9032);
nand U9245 (N_9245,N_9118,N_9111);
nand U9246 (N_9246,N_9114,N_9073);
or U9247 (N_9247,N_9089,N_9091);
and U9248 (N_9248,N_9103,N_9018);
nor U9249 (N_9249,N_9064,N_9108);
or U9250 (N_9250,N_9142,N_9177);
and U9251 (N_9251,N_9245,N_9212);
nand U9252 (N_9252,N_9135,N_9173);
and U9253 (N_9253,N_9134,N_9181);
or U9254 (N_9254,N_9143,N_9219);
xor U9255 (N_9255,N_9190,N_9155);
and U9256 (N_9256,N_9202,N_9239);
nand U9257 (N_9257,N_9238,N_9125);
and U9258 (N_9258,N_9211,N_9243);
nand U9259 (N_9259,N_9126,N_9159);
nor U9260 (N_9260,N_9168,N_9178);
or U9261 (N_9261,N_9184,N_9215);
nor U9262 (N_9262,N_9214,N_9217);
nor U9263 (N_9263,N_9166,N_9201);
and U9264 (N_9264,N_9228,N_9207);
or U9265 (N_9265,N_9138,N_9193);
nand U9266 (N_9266,N_9198,N_9236);
and U9267 (N_9267,N_9235,N_9203);
nor U9268 (N_9268,N_9170,N_9226);
or U9269 (N_9269,N_9189,N_9232);
nand U9270 (N_9270,N_9140,N_9146);
and U9271 (N_9271,N_9147,N_9197);
nor U9272 (N_9272,N_9151,N_9231);
nand U9273 (N_9273,N_9164,N_9247);
and U9274 (N_9274,N_9163,N_9233);
nand U9275 (N_9275,N_9162,N_9246);
or U9276 (N_9276,N_9220,N_9185);
nor U9277 (N_9277,N_9175,N_9131);
xnor U9278 (N_9278,N_9136,N_9132);
nand U9279 (N_9279,N_9160,N_9237);
and U9280 (N_9280,N_9172,N_9240);
and U9281 (N_9281,N_9206,N_9204);
nor U9282 (N_9282,N_9199,N_9133);
and U9283 (N_9283,N_9153,N_9210);
nand U9284 (N_9284,N_9249,N_9130);
nand U9285 (N_9285,N_9194,N_9158);
nand U9286 (N_9286,N_9183,N_9169);
nand U9287 (N_9287,N_9174,N_9225);
and U9288 (N_9288,N_9191,N_9187);
nor U9289 (N_9289,N_9221,N_9141);
or U9290 (N_9290,N_9223,N_9139);
or U9291 (N_9291,N_9213,N_9234);
nand U9292 (N_9292,N_9229,N_9152);
and U9293 (N_9293,N_9208,N_9171);
xnor U9294 (N_9294,N_9209,N_9179);
or U9295 (N_9295,N_9230,N_9149);
nor U9296 (N_9296,N_9218,N_9161);
nor U9297 (N_9297,N_9227,N_9205);
nand U9298 (N_9298,N_9154,N_9224);
and U9299 (N_9299,N_9242,N_9248);
or U9300 (N_9300,N_9137,N_9180);
or U9301 (N_9301,N_9165,N_9150);
and U9302 (N_9302,N_9188,N_9157);
and U9303 (N_9303,N_9156,N_9244);
nand U9304 (N_9304,N_9196,N_9195);
and U9305 (N_9305,N_9222,N_9182);
nor U9306 (N_9306,N_9129,N_9176);
nor U9307 (N_9307,N_9241,N_9144);
nand U9308 (N_9308,N_9186,N_9145);
and U9309 (N_9309,N_9127,N_9200);
or U9310 (N_9310,N_9192,N_9216);
nor U9311 (N_9311,N_9148,N_9128);
nand U9312 (N_9312,N_9167,N_9136);
and U9313 (N_9313,N_9171,N_9153);
and U9314 (N_9314,N_9141,N_9229);
nand U9315 (N_9315,N_9183,N_9154);
or U9316 (N_9316,N_9143,N_9211);
nor U9317 (N_9317,N_9207,N_9186);
nor U9318 (N_9318,N_9188,N_9206);
nand U9319 (N_9319,N_9177,N_9146);
or U9320 (N_9320,N_9137,N_9233);
or U9321 (N_9321,N_9131,N_9223);
nor U9322 (N_9322,N_9226,N_9176);
nand U9323 (N_9323,N_9214,N_9247);
nor U9324 (N_9324,N_9151,N_9182);
nor U9325 (N_9325,N_9238,N_9182);
and U9326 (N_9326,N_9180,N_9205);
or U9327 (N_9327,N_9232,N_9180);
and U9328 (N_9328,N_9202,N_9210);
xor U9329 (N_9329,N_9191,N_9229);
nand U9330 (N_9330,N_9139,N_9240);
nor U9331 (N_9331,N_9175,N_9135);
and U9332 (N_9332,N_9240,N_9207);
nor U9333 (N_9333,N_9240,N_9181);
nand U9334 (N_9334,N_9222,N_9249);
nand U9335 (N_9335,N_9232,N_9144);
nor U9336 (N_9336,N_9241,N_9135);
nand U9337 (N_9337,N_9189,N_9209);
and U9338 (N_9338,N_9153,N_9174);
nor U9339 (N_9339,N_9170,N_9219);
and U9340 (N_9340,N_9176,N_9234);
xor U9341 (N_9341,N_9151,N_9247);
or U9342 (N_9342,N_9248,N_9199);
and U9343 (N_9343,N_9158,N_9199);
nand U9344 (N_9344,N_9187,N_9170);
nand U9345 (N_9345,N_9173,N_9129);
nor U9346 (N_9346,N_9156,N_9216);
and U9347 (N_9347,N_9202,N_9174);
nor U9348 (N_9348,N_9140,N_9180);
nor U9349 (N_9349,N_9164,N_9206);
or U9350 (N_9350,N_9161,N_9190);
nand U9351 (N_9351,N_9199,N_9190);
nand U9352 (N_9352,N_9172,N_9146);
nand U9353 (N_9353,N_9247,N_9208);
nand U9354 (N_9354,N_9211,N_9136);
and U9355 (N_9355,N_9223,N_9189);
or U9356 (N_9356,N_9242,N_9198);
xor U9357 (N_9357,N_9172,N_9218);
nand U9358 (N_9358,N_9178,N_9242);
or U9359 (N_9359,N_9182,N_9173);
and U9360 (N_9360,N_9146,N_9171);
or U9361 (N_9361,N_9154,N_9236);
or U9362 (N_9362,N_9134,N_9177);
nand U9363 (N_9363,N_9152,N_9214);
nor U9364 (N_9364,N_9228,N_9203);
or U9365 (N_9365,N_9125,N_9171);
nor U9366 (N_9366,N_9203,N_9156);
nand U9367 (N_9367,N_9159,N_9128);
or U9368 (N_9368,N_9171,N_9188);
nor U9369 (N_9369,N_9144,N_9240);
or U9370 (N_9370,N_9201,N_9217);
nand U9371 (N_9371,N_9199,N_9182);
and U9372 (N_9372,N_9179,N_9213);
nor U9373 (N_9373,N_9143,N_9168);
nand U9374 (N_9374,N_9142,N_9152);
or U9375 (N_9375,N_9281,N_9310);
or U9376 (N_9376,N_9286,N_9250);
nand U9377 (N_9377,N_9313,N_9255);
xor U9378 (N_9378,N_9373,N_9315);
and U9379 (N_9379,N_9321,N_9314);
nand U9380 (N_9380,N_9325,N_9361);
and U9381 (N_9381,N_9324,N_9346);
nand U9382 (N_9382,N_9320,N_9252);
nor U9383 (N_9383,N_9289,N_9351);
and U9384 (N_9384,N_9307,N_9349);
or U9385 (N_9385,N_9344,N_9300);
or U9386 (N_9386,N_9282,N_9279);
nand U9387 (N_9387,N_9273,N_9322);
nor U9388 (N_9388,N_9256,N_9296);
and U9389 (N_9389,N_9330,N_9291);
nor U9390 (N_9390,N_9295,N_9318);
nand U9391 (N_9391,N_9277,N_9357);
nand U9392 (N_9392,N_9323,N_9327);
and U9393 (N_9393,N_9283,N_9259);
nor U9394 (N_9394,N_9334,N_9338);
or U9395 (N_9395,N_9275,N_9303);
nor U9396 (N_9396,N_9294,N_9264);
or U9397 (N_9397,N_9308,N_9305);
xor U9398 (N_9398,N_9358,N_9285);
nand U9399 (N_9399,N_9312,N_9251);
nand U9400 (N_9400,N_9284,N_9272);
or U9401 (N_9401,N_9271,N_9274);
nand U9402 (N_9402,N_9309,N_9262);
xnor U9403 (N_9403,N_9365,N_9288);
nand U9404 (N_9404,N_9298,N_9332);
xor U9405 (N_9405,N_9367,N_9316);
nand U9406 (N_9406,N_9352,N_9311);
or U9407 (N_9407,N_9371,N_9372);
nand U9408 (N_9408,N_9366,N_9268);
or U9409 (N_9409,N_9328,N_9347);
and U9410 (N_9410,N_9269,N_9263);
and U9411 (N_9411,N_9293,N_9292);
and U9412 (N_9412,N_9329,N_9287);
and U9413 (N_9413,N_9260,N_9270);
or U9414 (N_9414,N_9331,N_9374);
and U9415 (N_9415,N_9363,N_9342);
or U9416 (N_9416,N_9345,N_9276);
or U9417 (N_9417,N_9364,N_9267);
xnor U9418 (N_9418,N_9302,N_9258);
nand U9419 (N_9419,N_9353,N_9350);
xor U9420 (N_9420,N_9280,N_9326);
and U9421 (N_9421,N_9337,N_9368);
and U9422 (N_9422,N_9341,N_9278);
xnor U9423 (N_9423,N_9261,N_9266);
nand U9424 (N_9424,N_9336,N_9301);
and U9425 (N_9425,N_9257,N_9253);
or U9426 (N_9426,N_9355,N_9297);
or U9427 (N_9427,N_9317,N_9265);
nand U9428 (N_9428,N_9354,N_9304);
and U9429 (N_9429,N_9343,N_9348);
or U9430 (N_9430,N_9306,N_9254);
nand U9431 (N_9431,N_9335,N_9359);
or U9432 (N_9432,N_9369,N_9340);
xnor U9433 (N_9433,N_9299,N_9333);
and U9434 (N_9434,N_9362,N_9290);
and U9435 (N_9435,N_9370,N_9360);
nand U9436 (N_9436,N_9339,N_9319);
nand U9437 (N_9437,N_9356,N_9300);
and U9438 (N_9438,N_9272,N_9333);
nor U9439 (N_9439,N_9307,N_9268);
xnor U9440 (N_9440,N_9348,N_9256);
or U9441 (N_9441,N_9348,N_9259);
nor U9442 (N_9442,N_9342,N_9338);
and U9443 (N_9443,N_9335,N_9333);
or U9444 (N_9444,N_9325,N_9270);
nor U9445 (N_9445,N_9279,N_9261);
nor U9446 (N_9446,N_9296,N_9341);
nand U9447 (N_9447,N_9269,N_9332);
and U9448 (N_9448,N_9251,N_9278);
and U9449 (N_9449,N_9344,N_9250);
nand U9450 (N_9450,N_9332,N_9364);
or U9451 (N_9451,N_9282,N_9313);
and U9452 (N_9452,N_9320,N_9340);
or U9453 (N_9453,N_9367,N_9270);
and U9454 (N_9454,N_9356,N_9348);
nand U9455 (N_9455,N_9334,N_9364);
nand U9456 (N_9456,N_9264,N_9268);
and U9457 (N_9457,N_9279,N_9277);
nor U9458 (N_9458,N_9303,N_9288);
nand U9459 (N_9459,N_9359,N_9336);
nor U9460 (N_9460,N_9260,N_9327);
nor U9461 (N_9461,N_9287,N_9324);
and U9462 (N_9462,N_9267,N_9274);
xnor U9463 (N_9463,N_9275,N_9339);
and U9464 (N_9464,N_9278,N_9331);
nand U9465 (N_9465,N_9295,N_9282);
nor U9466 (N_9466,N_9304,N_9275);
nand U9467 (N_9467,N_9364,N_9317);
nand U9468 (N_9468,N_9332,N_9319);
and U9469 (N_9469,N_9365,N_9260);
and U9470 (N_9470,N_9337,N_9253);
and U9471 (N_9471,N_9322,N_9339);
nand U9472 (N_9472,N_9348,N_9303);
nor U9473 (N_9473,N_9287,N_9355);
nand U9474 (N_9474,N_9325,N_9280);
and U9475 (N_9475,N_9294,N_9282);
or U9476 (N_9476,N_9334,N_9287);
and U9477 (N_9477,N_9297,N_9251);
nand U9478 (N_9478,N_9316,N_9253);
and U9479 (N_9479,N_9361,N_9348);
and U9480 (N_9480,N_9348,N_9297);
and U9481 (N_9481,N_9345,N_9251);
and U9482 (N_9482,N_9316,N_9333);
nand U9483 (N_9483,N_9259,N_9374);
or U9484 (N_9484,N_9351,N_9288);
nor U9485 (N_9485,N_9295,N_9257);
xor U9486 (N_9486,N_9332,N_9338);
and U9487 (N_9487,N_9287,N_9280);
nor U9488 (N_9488,N_9347,N_9268);
nor U9489 (N_9489,N_9301,N_9250);
or U9490 (N_9490,N_9286,N_9345);
or U9491 (N_9491,N_9365,N_9287);
xor U9492 (N_9492,N_9288,N_9290);
and U9493 (N_9493,N_9371,N_9306);
or U9494 (N_9494,N_9357,N_9370);
and U9495 (N_9495,N_9303,N_9287);
or U9496 (N_9496,N_9335,N_9362);
or U9497 (N_9497,N_9283,N_9293);
and U9498 (N_9498,N_9353,N_9253);
or U9499 (N_9499,N_9327,N_9359);
xnor U9500 (N_9500,N_9407,N_9443);
or U9501 (N_9501,N_9466,N_9440);
and U9502 (N_9502,N_9379,N_9433);
xor U9503 (N_9503,N_9473,N_9403);
or U9504 (N_9504,N_9404,N_9498);
nand U9505 (N_9505,N_9392,N_9401);
nor U9506 (N_9506,N_9406,N_9469);
nor U9507 (N_9507,N_9417,N_9434);
or U9508 (N_9508,N_9429,N_9476);
and U9509 (N_9509,N_9486,N_9412);
or U9510 (N_9510,N_9467,N_9421);
and U9511 (N_9511,N_9432,N_9472);
or U9512 (N_9512,N_9378,N_9376);
nand U9513 (N_9513,N_9449,N_9470);
or U9514 (N_9514,N_9491,N_9451);
nor U9515 (N_9515,N_9471,N_9384);
or U9516 (N_9516,N_9389,N_9456);
nor U9517 (N_9517,N_9454,N_9408);
nor U9518 (N_9518,N_9381,N_9398);
xor U9519 (N_9519,N_9439,N_9446);
or U9520 (N_9520,N_9492,N_9390);
nand U9521 (N_9521,N_9493,N_9444);
and U9522 (N_9522,N_9385,N_9420);
and U9523 (N_9523,N_9416,N_9427);
nor U9524 (N_9524,N_9455,N_9382);
xor U9525 (N_9525,N_9488,N_9490);
nor U9526 (N_9526,N_9463,N_9475);
or U9527 (N_9527,N_9428,N_9448);
nor U9528 (N_9528,N_9410,N_9497);
xor U9529 (N_9529,N_9436,N_9483);
and U9530 (N_9530,N_9468,N_9461);
nand U9531 (N_9531,N_9395,N_9477);
nor U9532 (N_9532,N_9441,N_9437);
nand U9533 (N_9533,N_9481,N_9399);
nand U9534 (N_9534,N_9418,N_9452);
nor U9535 (N_9535,N_9419,N_9377);
nor U9536 (N_9536,N_9414,N_9447);
and U9537 (N_9537,N_9423,N_9430);
nor U9538 (N_9538,N_9453,N_9438);
nand U9539 (N_9539,N_9484,N_9383);
xor U9540 (N_9540,N_9494,N_9499);
and U9541 (N_9541,N_9496,N_9487);
or U9542 (N_9542,N_9445,N_9402);
nand U9543 (N_9543,N_9435,N_9474);
nand U9544 (N_9544,N_9479,N_9397);
and U9545 (N_9545,N_9465,N_9450);
xnor U9546 (N_9546,N_9393,N_9426);
or U9547 (N_9547,N_9460,N_9386);
nor U9548 (N_9548,N_9495,N_9391);
or U9549 (N_9549,N_9380,N_9457);
nand U9550 (N_9550,N_9480,N_9411);
and U9551 (N_9551,N_9387,N_9394);
and U9552 (N_9552,N_9396,N_9422);
nor U9553 (N_9553,N_9425,N_9409);
nor U9554 (N_9554,N_9375,N_9459);
nand U9555 (N_9555,N_9405,N_9442);
nand U9556 (N_9556,N_9464,N_9462);
xor U9557 (N_9557,N_9400,N_9413);
and U9558 (N_9558,N_9485,N_9415);
or U9559 (N_9559,N_9478,N_9458);
nand U9560 (N_9560,N_9489,N_9424);
nand U9561 (N_9561,N_9431,N_9482);
or U9562 (N_9562,N_9388,N_9456);
nand U9563 (N_9563,N_9417,N_9483);
or U9564 (N_9564,N_9396,N_9494);
and U9565 (N_9565,N_9456,N_9401);
and U9566 (N_9566,N_9463,N_9402);
nand U9567 (N_9567,N_9404,N_9422);
nor U9568 (N_9568,N_9461,N_9437);
or U9569 (N_9569,N_9384,N_9492);
or U9570 (N_9570,N_9479,N_9464);
nand U9571 (N_9571,N_9428,N_9493);
xnor U9572 (N_9572,N_9471,N_9400);
nand U9573 (N_9573,N_9408,N_9468);
nor U9574 (N_9574,N_9408,N_9491);
nor U9575 (N_9575,N_9393,N_9388);
or U9576 (N_9576,N_9463,N_9381);
nor U9577 (N_9577,N_9434,N_9478);
or U9578 (N_9578,N_9380,N_9381);
nand U9579 (N_9579,N_9409,N_9464);
xnor U9580 (N_9580,N_9419,N_9385);
nor U9581 (N_9581,N_9381,N_9416);
and U9582 (N_9582,N_9455,N_9478);
or U9583 (N_9583,N_9405,N_9385);
xnor U9584 (N_9584,N_9458,N_9499);
nand U9585 (N_9585,N_9398,N_9412);
or U9586 (N_9586,N_9379,N_9416);
and U9587 (N_9587,N_9384,N_9483);
nand U9588 (N_9588,N_9424,N_9422);
xnor U9589 (N_9589,N_9387,N_9375);
xnor U9590 (N_9590,N_9379,N_9407);
xor U9591 (N_9591,N_9405,N_9452);
nor U9592 (N_9592,N_9479,N_9387);
and U9593 (N_9593,N_9401,N_9496);
and U9594 (N_9594,N_9442,N_9417);
nor U9595 (N_9595,N_9448,N_9417);
or U9596 (N_9596,N_9497,N_9435);
xor U9597 (N_9597,N_9452,N_9477);
or U9598 (N_9598,N_9437,N_9399);
or U9599 (N_9599,N_9426,N_9456);
nor U9600 (N_9600,N_9493,N_9489);
nor U9601 (N_9601,N_9381,N_9426);
nand U9602 (N_9602,N_9432,N_9423);
nand U9603 (N_9603,N_9427,N_9482);
nor U9604 (N_9604,N_9381,N_9377);
nor U9605 (N_9605,N_9494,N_9421);
or U9606 (N_9606,N_9445,N_9422);
nand U9607 (N_9607,N_9426,N_9385);
nand U9608 (N_9608,N_9497,N_9421);
or U9609 (N_9609,N_9448,N_9388);
nor U9610 (N_9610,N_9489,N_9384);
and U9611 (N_9611,N_9413,N_9419);
nand U9612 (N_9612,N_9407,N_9467);
nor U9613 (N_9613,N_9392,N_9424);
nand U9614 (N_9614,N_9495,N_9421);
or U9615 (N_9615,N_9483,N_9459);
or U9616 (N_9616,N_9455,N_9400);
nor U9617 (N_9617,N_9405,N_9409);
xnor U9618 (N_9618,N_9450,N_9471);
or U9619 (N_9619,N_9495,N_9393);
nand U9620 (N_9620,N_9398,N_9479);
xnor U9621 (N_9621,N_9462,N_9404);
nand U9622 (N_9622,N_9388,N_9461);
and U9623 (N_9623,N_9431,N_9447);
xor U9624 (N_9624,N_9418,N_9445);
and U9625 (N_9625,N_9563,N_9618);
or U9626 (N_9626,N_9535,N_9564);
nand U9627 (N_9627,N_9605,N_9551);
nor U9628 (N_9628,N_9504,N_9584);
nand U9629 (N_9629,N_9562,N_9502);
xnor U9630 (N_9630,N_9539,N_9540);
nor U9631 (N_9631,N_9597,N_9506);
or U9632 (N_9632,N_9542,N_9600);
nor U9633 (N_9633,N_9525,N_9585);
nand U9634 (N_9634,N_9617,N_9550);
xor U9635 (N_9635,N_9553,N_9552);
nor U9636 (N_9636,N_9522,N_9521);
and U9637 (N_9637,N_9616,N_9508);
xnor U9638 (N_9638,N_9598,N_9591);
nand U9639 (N_9639,N_9530,N_9558);
and U9640 (N_9640,N_9505,N_9590);
and U9641 (N_9641,N_9538,N_9622);
nor U9642 (N_9642,N_9578,N_9607);
and U9643 (N_9643,N_9599,N_9517);
and U9644 (N_9644,N_9595,N_9609);
nand U9645 (N_9645,N_9601,N_9603);
and U9646 (N_9646,N_9577,N_9531);
and U9647 (N_9647,N_9546,N_9559);
and U9648 (N_9648,N_9586,N_9536);
nor U9649 (N_9649,N_9556,N_9570);
nor U9650 (N_9650,N_9533,N_9526);
nand U9651 (N_9651,N_9520,N_9596);
nor U9652 (N_9652,N_9568,N_9624);
or U9653 (N_9653,N_9614,N_9579);
nor U9654 (N_9654,N_9574,N_9516);
and U9655 (N_9655,N_9602,N_9509);
nand U9656 (N_9656,N_9543,N_9612);
nor U9657 (N_9657,N_9501,N_9593);
and U9658 (N_9658,N_9560,N_9575);
nand U9659 (N_9659,N_9623,N_9512);
nor U9660 (N_9660,N_9583,N_9604);
xnor U9661 (N_9661,N_9519,N_9611);
nand U9662 (N_9662,N_9548,N_9594);
xnor U9663 (N_9663,N_9569,N_9511);
xor U9664 (N_9664,N_9571,N_9606);
and U9665 (N_9665,N_9588,N_9547);
nor U9666 (N_9666,N_9528,N_9544);
or U9667 (N_9667,N_9619,N_9524);
nand U9668 (N_9668,N_9541,N_9561);
nand U9669 (N_9669,N_9518,N_9537);
xor U9670 (N_9670,N_9613,N_9514);
nand U9671 (N_9671,N_9567,N_9581);
or U9672 (N_9672,N_9555,N_9610);
nor U9673 (N_9673,N_9608,N_9589);
or U9674 (N_9674,N_9554,N_9532);
nand U9675 (N_9675,N_9510,N_9566);
nand U9676 (N_9676,N_9592,N_9527);
and U9677 (N_9677,N_9615,N_9534);
or U9678 (N_9678,N_9515,N_9573);
or U9679 (N_9679,N_9500,N_9620);
or U9680 (N_9680,N_9523,N_9545);
nor U9681 (N_9681,N_9529,N_9565);
nand U9682 (N_9682,N_9582,N_9587);
and U9683 (N_9683,N_9507,N_9572);
nor U9684 (N_9684,N_9621,N_9549);
nor U9685 (N_9685,N_9513,N_9576);
nand U9686 (N_9686,N_9557,N_9503);
or U9687 (N_9687,N_9580,N_9505);
nand U9688 (N_9688,N_9621,N_9514);
xor U9689 (N_9689,N_9551,N_9573);
or U9690 (N_9690,N_9567,N_9592);
or U9691 (N_9691,N_9567,N_9602);
or U9692 (N_9692,N_9582,N_9610);
and U9693 (N_9693,N_9596,N_9563);
and U9694 (N_9694,N_9535,N_9571);
xnor U9695 (N_9695,N_9575,N_9530);
or U9696 (N_9696,N_9560,N_9545);
nand U9697 (N_9697,N_9605,N_9539);
and U9698 (N_9698,N_9501,N_9606);
nor U9699 (N_9699,N_9588,N_9504);
nand U9700 (N_9700,N_9538,N_9591);
nand U9701 (N_9701,N_9503,N_9520);
nor U9702 (N_9702,N_9539,N_9595);
nor U9703 (N_9703,N_9509,N_9510);
nor U9704 (N_9704,N_9529,N_9592);
and U9705 (N_9705,N_9527,N_9512);
or U9706 (N_9706,N_9537,N_9578);
and U9707 (N_9707,N_9588,N_9577);
or U9708 (N_9708,N_9529,N_9535);
or U9709 (N_9709,N_9603,N_9512);
nand U9710 (N_9710,N_9571,N_9551);
and U9711 (N_9711,N_9550,N_9506);
xnor U9712 (N_9712,N_9579,N_9527);
nor U9713 (N_9713,N_9569,N_9523);
xor U9714 (N_9714,N_9525,N_9503);
nor U9715 (N_9715,N_9536,N_9558);
xnor U9716 (N_9716,N_9548,N_9595);
nand U9717 (N_9717,N_9590,N_9624);
nand U9718 (N_9718,N_9535,N_9547);
or U9719 (N_9719,N_9585,N_9598);
and U9720 (N_9720,N_9610,N_9559);
and U9721 (N_9721,N_9554,N_9588);
nor U9722 (N_9722,N_9525,N_9589);
nand U9723 (N_9723,N_9602,N_9507);
and U9724 (N_9724,N_9597,N_9586);
and U9725 (N_9725,N_9543,N_9587);
nand U9726 (N_9726,N_9527,N_9624);
nand U9727 (N_9727,N_9572,N_9612);
or U9728 (N_9728,N_9588,N_9619);
nand U9729 (N_9729,N_9605,N_9548);
nand U9730 (N_9730,N_9564,N_9615);
or U9731 (N_9731,N_9551,N_9623);
and U9732 (N_9732,N_9536,N_9554);
nand U9733 (N_9733,N_9513,N_9591);
or U9734 (N_9734,N_9598,N_9546);
xor U9735 (N_9735,N_9505,N_9604);
nor U9736 (N_9736,N_9621,N_9547);
nand U9737 (N_9737,N_9614,N_9521);
nor U9738 (N_9738,N_9552,N_9517);
and U9739 (N_9739,N_9516,N_9517);
or U9740 (N_9740,N_9517,N_9608);
and U9741 (N_9741,N_9573,N_9501);
and U9742 (N_9742,N_9572,N_9546);
xor U9743 (N_9743,N_9620,N_9617);
or U9744 (N_9744,N_9510,N_9622);
nor U9745 (N_9745,N_9501,N_9509);
nand U9746 (N_9746,N_9530,N_9507);
and U9747 (N_9747,N_9558,N_9511);
and U9748 (N_9748,N_9514,N_9614);
nand U9749 (N_9749,N_9528,N_9522);
nand U9750 (N_9750,N_9693,N_9694);
nor U9751 (N_9751,N_9732,N_9703);
or U9752 (N_9752,N_9743,N_9699);
or U9753 (N_9753,N_9634,N_9661);
nand U9754 (N_9754,N_9670,N_9653);
nand U9755 (N_9755,N_9660,N_9726);
nand U9756 (N_9756,N_9705,N_9627);
nand U9757 (N_9757,N_9682,N_9625);
xnor U9758 (N_9758,N_9738,N_9713);
nor U9759 (N_9759,N_9657,N_9636);
xnor U9760 (N_9760,N_9719,N_9700);
nand U9761 (N_9761,N_9720,N_9666);
nand U9762 (N_9762,N_9646,N_9701);
and U9763 (N_9763,N_9638,N_9665);
and U9764 (N_9764,N_9669,N_9731);
and U9765 (N_9765,N_9687,N_9628);
xor U9766 (N_9766,N_9641,N_9640);
nor U9767 (N_9767,N_9671,N_9652);
and U9768 (N_9768,N_9746,N_9741);
or U9769 (N_9769,N_9656,N_9744);
and U9770 (N_9770,N_9698,N_9711);
nor U9771 (N_9771,N_9729,N_9686);
xor U9772 (N_9772,N_9733,N_9736);
xor U9773 (N_9773,N_9675,N_9679);
nand U9774 (N_9774,N_9626,N_9647);
nand U9775 (N_9775,N_9637,N_9667);
and U9776 (N_9776,N_9690,N_9749);
and U9777 (N_9777,N_9704,N_9723);
and U9778 (N_9778,N_9681,N_9632);
and U9779 (N_9779,N_9709,N_9680);
and U9780 (N_9780,N_9644,N_9745);
or U9781 (N_9781,N_9697,N_9737);
nand U9782 (N_9782,N_9714,N_9629);
or U9783 (N_9783,N_9649,N_9663);
and U9784 (N_9784,N_9740,N_9696);
nand U9785 (N_9785,N_9747,N_9708);
nand U9786 (N_9786,N_9710,N_9689);
and U9787 (N_9787,N_9664,N_9662);
or U9788 (N_9788,N_9630,N_9707);
nor U9789 (N_9789,N_9734,N_9706);
nand U9790 (N_9790,N_9742,N_9735);
nor U9791 (N_9791,N_9655,N_9651);
and U9792 (N_9792,N_9721,N_9658);
xnor U9793 (N_9793,N_9648,N_9677);
and U9794 (N_9794,N_9715,N_9685);
and U9795 (N_9795,N_9678,N_9643);
nand U9796 (N_9796,N_9692,N_9672);
nor U9797 (N_9797,N_9730,N_9717);
nor U9798 (N_9798,N_9748,N_9674);
nor U9799 (N_9799,N_9712,N_9673);
xnor U9800 (N_9800,N_9645,N_9725);
nand U9801 (N_9801,N_9688,N_9650);
and U9802 (N_9802,N_9639,N_9739);
or U9803 (N_9803,N_9695,N_9631);
nand U9804 (N_9804,N_9684,N_9728);
nor U9805 (N_9805,N_9691,N_9683);
xnor U9806 (N_9806,N_9633,N_9642);
nand U9807 (N_9807,N_9654,N_9718);
or U9808 (N_9808,N_9635,N_9724);
nor U9809 (N_9809,N_9722,N_9668);
or U9810 (N_9810,N_9676,N_9727);
and U9811 (N_9811,N_9659,N_9716);
nand U9812 (N_9812,N_9702,N_9655);
nor U9813 (N_9813,N_9640,N_9721);
and U9814 (N_9814,N_9635,N_9745);
or U9815 (N_9815,N_9718,N_9711);
nor U9816 (N_9816,N_9669,N_9657);
nand U9817 (N_9817,N_9719,N_9709);
xnor U9818 (N_9818,N_9732,N_9643);
xnor U9819 (N_9819,N_9741,N_9671);
or U9820 (N_9820,N_9692,N_9634);
xor U9821 (N_9821,N_9687,N_9665);
xnor U9822 (N_9822,N_9737,N_9625);
or U9823 (N_9823,N_9670,N_9699);
nand U9824 (N_9824,N_9731,N_9745);
nand U9825 (N_9825,N_9633,N_9720);
xor U9826 (N_9826,N_9703,N_9667);
nand U9827 (N_9827,N_9710,N_9671);
nand U9828 (N_9828,N_9673,N_9710);
xor U9829 (N_9829,N_9671,N_9692);
or U9830 (N_9830,N_9625,N_9749);
nor U9831 (N_9831,N_9643,N_9651);
nor U9832 (N_9832,N_9699,N_9679);
and U9833 (N_9833,N_9681,N_9645);
or U9834 (N_9834,N_9728,N_9713);
and U9835 (N_9835,N_9649,N_9690);
or U9836 (N_9836,N_9712,N_9680);
nor U9837 (N_9837,N_9695,N_9706);
or U9838 (N_9838,N_9687,N_9734);
nand U9839 (N_9839,N_9643,N_9743);
and U9840 (N_9840,N_9685,N_9738);
or U9841 (N_9841,N_9749,N_9660);
nor U9842 (N_9842,N_9743,N_9728);
and U9843 (N_9843,N_9670,N_9675);
and U9844 (N_9844,N_9746,N_9676);
and U9845 (N_9845,N_9701,N_9688);
nor U9846 (N_9846,N_9735,N_9672);
xnor U9847 (N_9847,N_9712,N_9709);
and U9848 (N_9848,N_9725,N_9713);
xor U9849 (N_9849,N_9667,N_9704);
or U9850 (N_9850,N_9725,N_9667);
and U9851 (N_9851,N_9668,N_9716);
nand U9852 (N_9852,N_9647,N_9668);
and U9853 (N_9853,N_9667,N_9636);
nand U9854 (N_9854,N_9740,N_9695);
and U9855 (N_9855,N_9739,N_9714);
nor U9856 (N_9856,N_9744,N_9702);
nand U9857 (N_9857,N_9662,N_9734);
nor U9858 (N_9858,N_9673,N_9631);
and U9859 (N_9859,N_9679,N_9694);
xnor U9860 (N_9860,N_9730,N_9742);
nor U9861 (N_9861,N_9739,N_9679);
xnor U9862 (N_9862,N_9703,N_9697);
and U9863 (N_9863,N_9634,N_9673);
xor U9864 (N_9864,N_9746,N_9639);
or U9865 (N_9865,N_9677,N_9647);
or U9866 (N_9866,N_9632,N_9625);
or U9867 (N_9867,N_9665,N_9712);
or U9868 (N_9868,N_9688,N_9723);
nand U9869 (N_9869,N_9717,N_9736);
nand U9870 (N_9870,N_9666,N_9708);
nor U9871 (N_9871,N_9725,N_9640);
nand U9872 (N_9872,N_9638,N_9661);
nor U9873 (N_9873,N_9746,N_9685);
nor U9874 (N_9874,N_9740,N_9627);
and U9875 (N_9875,N_9869,N_9871);
and U9876 (N_9876,N_9866,N_9841);
or U9877 (N_9877,N_9852,N_9816);
or U9878 (N_9878,N_9834,N_9822);
nor U9879 (N_9879,N_9763,N_9823);
or U9880 (N_9880,N_9828,N_9837);
or U9881 (N_9881,N_9783,N_9795);
nor U9882 (N_9882,N_9799,N_9873);
and U9883 (N_9883,N_9802,N_9808);
and U9884 (N_9884,N_9867,N_9758);
nand U9885 (N_9885,N_9805,N_9851);
nor U9886 (N_9886,N_9835,N_9778);
and U9887 (N_9887,N_9764,N_9820);
nor U9888 (N_9888,N_9840,N_9771);
nor U9889 (N_9889,N_9829,N_9754);
nand U9890 (N_9890,N_9831,N_9847);
or U9891 (N_9891,N_9814,N_9838);
xnor U9892 (N_9892,N_9762,N_9789);
or U9893 (N_9893,N_9865,N_9832);
and U9894 (N_9894,N_9794,N_9845);
nand U9895 (N_9895,N_9830,N_9826);
and U9896 (N_9896,N_9773,N_9797);
and U9897 (N_9897,N_9839,N_9770);
or U9898 (N_9898,N_9853,N_9861);
xnor U9899 (N_9899,N_9872,N_9756);
nand U9900 (N_9900,N_9751,N_9856);
nand U9901 (N_9901,N_9759,N_9760);
nor U9902 (N_9902,N_9786,N_9848);
and U9903 (N_9903,N_9863,N_9806);
nor U9904 (N_9904,N_9874,N_9825);
nor U9905 (N_9905,N_9765,N_9846);
nor U9906 (N_9906,N_9807,N_9821);
nand U9907 (N_9907,N_9870,N_9780);
or U9908 (N_9908,N_9750,N_9819);
nand U9909 (N_9909,N_9793,N_9782);
nand U9910 (N_9910,N_9776,N_9818);
and U9911 (N_9911,N_9864,N_9854);
nand U9912 (N_9912,N_9753,N_9772);
or U9913 (N_9913,N_9801,N_9790);
or U9914 (N_9914,N_9768,N_9796);
or U9915 (N_9915,N_9791,N_9788);
and U9916 (N_9916,N_9809,N_9868);
nor U9917 (N_9917,N_9774,N_9800);
xnor U9918 (N_9918,N_9859,N_9855);
or U9919 (N_9919,N_9824,N_9833);
xor U9920 (N_9920,N_9812,N_9850);
nor U9921 (N_9921,N_9766,N_9785);
or U9922 (N_9922,N_9810,N_9843);
nand U9923 (N_9923,N_9862,N_9767);
nor U9924 (N_9924,N_9757,N_9860);
nor U9925 (N_9925,N_9761,N_9857);
nor U9926 (N_9926,N_9815,N_9804);
nor U9927 (N_9927,N_9842,N_9836);
nor U9928 (N_9928,N_9781,N_9769);
and U9929 (N_9929,N_9784,N_9811);
or U9930 (N_9930,N_9752,N_9775);
nor U9931 (N_9931,N_9787,N_9803);
nor U9932 (N_9932,N_9798,N_9755);
nor U9933 (N_9933,N_9844,N_9849);
or U9934 (N_9934,N_9827,N_9779);
and U9935 (N_9935,N_9858,N_9777);
nor U9936 (N_9936,N_9813,N_9792);
and U9937 (N_9937,N_9817,N_9783);
nand U9938 (N_9938,N_9810,N_9759);
nor U9939 (N_9939,N_9822,N_9752);
nor U9940 (N_9940,N_9813,N_9856);
nor U9941 (N_9941,N_9755,N_9858);
or U9942 (N_9942,N_9821,N_9834);
nor U9943 (N_9943,N_9830,N_9760);
nand U9944 (N_9944,N_9865,N_9841);
nand U9945 (N_9945,N_9788,N_9765);
or U9946 (N_9946,N_9825,N_9797);
nor U9947 (N_9947,N_9754,N_9855);
and U9948 (N_9948,N_9804,N_9849);
and U9949 (N_9949,N_9763,N_9812);
nor U9950 (N_9950,N_9771,N_9865);
or U9951 (N_9951,N_9782,N_9873);
nor U9952 (N_9952,N_9806,N_9760);
nand U9953 (N_9953,N_9810,N_9835);
xnor U9954 (N_9954,N_9789,N_9814);
nand U9955 (N_9955,N_9821,N_9867);
or U9956 (N_9956,N_9782,N_9761);
or U9957 (N_9957,N_9796,N_9818);
and U9958 (N_9958,N_9851,N_9818);
nor U9959 (N_9959,N_9805,N_9773);
nor U9960 (N_9960,N_9829,N_9815);
xor U9961 (N_9961,N_9855,N_9850);
and U9962 (N_9962,N_9769,N_9842);
xnor U9963 (N_9963,N_9751,N_9867);
or U9964 (N_9964,N_9825,N_9842);
nand U9965 (N_9965,N_9863,N_9811);
and U9966 (N_9966,N_9858,N_9764);
or U9967 (N_9967,N_9793,N_9760);
nand U9968 (N_9968,N_9772,N_9861);
or U9969 (N_9969,N_9869,N_9799);
and U9970 (N_9970,N_9873,N_9862);
xor U9971 (N_9971,N_9807,N_9841);
nor U9972 (N_9972,N_9779,N_9772);
or U9973 (N_9973,N_9834,N_9789);
nand U9974 (N_9974,N_9786,N_9859);
and U9975 (N_9975,N_9756,N_9794);
and U9976 (N_9976,N_9824,N_9786);
and U9977 (N_9977,N_9763,N_9854);
and U9978 (N_9978,N_9873,N_9768);
and U9979 (N_9979,N_9783,N_9840);
nor U9980 (N_9980,N_9857,N_9866);
nand U9981 (N_9981,N_9768,N_9823);
and U9982 (N_9982,N_9844,N_9753);
nand U9983 (N_9983,N_9785,N_9863);
xnor U9984 (N_9984,N_9831,N_9771);
nand U9985 (N_9985,N_9801,N_9804);
xnor U9986 (N_9986,N_9812,N_9803);
and U9987 (N_9987,N_9851,N_9819);
nor U9988 (N_9988,N_9840,N_9756);
and U9989 (N_9989,N_9754,N_9767);
nand U9990 (N_9990,N_9852,N_9791);
or U9991 (N_9991,N_9766,N_9802);
or U9992 (N_9992,N_9751,N_9845);
and U9993 (N_9993,N_9801,N_9754);
xnor U9994 (N_9994,N_9753,N_9807);
and U9995 (N_9995,N_9824,N_9814);
xor U9996 (N_9996,N_9833,N_9750);
nand U9997 (N_9997,N_9830,N_9750);
nor U9998 (N_9998,N_9865,N_9799);
and U9999 (N_9999,N_9843,N_9861);
nor U10000 (N_10000,N_9996,N_9977);
xor U10001 (N_10001,N_9981,N_9930);
and U10002 (N_10002,N_9914,N_9921);
nand U10003 (N_10003,N_9960,N_9998);
or U10004 (N_10004,N_9879,N_9915);
nand U10005 (N_10005,N_9988,N_9894);
nor U10006 (N_10006,N_9939,N_9953);
and U10007 (N_10007,N_9893,N_9980);
nor U10008 (N_10008,N_9993,N_9889);
and U10009 (N_10009,N_9878,N_9963);
xnor U10010 (N_10010,N_9931,N_9898);
and U10011 (N_10011,N_9904,N_9932);
nand U10012 (N_10012,N_9936,N_9892);
and U10013 (N_10013,N_9969,N_9947);
or U10014 (N_10014,N_9958,N_9920);
nand U10015 (N_10015,N_9983,N_9948);
nor U10016 (N_10016,N_9916,N_9961);
nand U10017 (N_10017,N_9995,N_9962);
or U10018 (N_10018,N_9917,N_9941);
nand U10019 (N_10019,N_9944,N_9997);
nand U10020 (N_10020,N_9909,N_9940);
or U10021 (N_10021,N_9952,N_9966);
xor U10022 (N_10022,N_9884,N_9986);
nand U10023 (N_10023,N_9888,N_9905);
nor U10024 (N_10024,N_9985,N_9965);
and U10025 (N_10025,N_9938,N_9942);
nor U10026 (N_10026,N_9891,N_9933);
nand U10027 (N_10027,N_9886,N_9912);
nor U10028 (N_10028,N_9970,N_9902);
nand U10029 (N_10029,N_9973,N_9994);
nor U10030 (N_10030,N_9957,N_9964);
or U10031 (N_10031,N_9906,N_9890);
and U10032 (N_10032,N_9918,N_9895);
or U10033 (N_10033,N_9968,N_9927);
nor U10034 (N_10034,N_9946,N_9992);
nor U10035 (N_10035,N_9987,N_9926);
and U10036 (N_10036,N_9950,N_9989);
and U10037 (N_10037,N_9982,N_9922);
and U10038 (N_10038,N_9907,N_9896);
nand U10039 (N_10039,N_9882,N_9876);
or U10040 (N_10040,N_9976,N_9887);
or U10041 (N_10041,N_9974,N_9951);
nand U10042 (N_10042,N_9923,N_9919);
or U10043 (N_10043,N_9978,N_9881);
and U10044 (N_10044,N_9979,N_9910);
nand U10045 (N_10045,N_9911,N_9897);
nor U10046 (N_10046,N_9949,N_9943);
or U10047 (N_10047,N_9913,N_9900);
nand U10048 (N_10048,N_9935,N_9925);
nand U10049 (N_10049,N_9972,N_9984);
nor U10050 (N_10050,N_9899,N_9885);
and U10051 (N_10051,N_9956,N_9959);
nor U10052 (N_10052,N_9875,N_9877);
and U10053 (N_10053,N_9929,N_9880);
or U10054 (N_10054,N_9928,N_9924);
nand U10055 (N_10055,N_9945,N_9954);
xnor U10056 (N_10056,N_9908,N_9990);
nand U10057 (N_10057,N_9975,N_9934);
xnor U10058 (N_10058,N_9991,N_9999);
or U10059 (N_10059,N_9901,N_9883);
nand U10060 (N_10060,N_9971,N_9955);
nand U10061 (N_10061,N_9937,N_9903);
xor U10062 (N_10062,N_9967,N_9887);
nand U10063 (N_10063,N_9968,N_9908);
nand U10064 (N_10064,N_9951,N_9898);
nor U10065 (N_10065,N_9993,N_9935);
xor U10066 (N_10066,N_9948,N_9972);
and U10067 (N_10067,N_9957,N_9987);
nor U10068 (N_10068,N_9919,N_9924);
or U10069 (N_10069,N_9958,N_9979);
nand U10070 (N_10070,N_9945,N_9889);
nand U10071 (N_10071,N_9931,N_9974);
or U10072 (N_10072,N_9901,N_9907);
or U10073 (N_10073,N_9886,N_9952);
xor U10074 (N_10074,N_9896,N_9986);
nand U10075 (N_10075,N_9975,N_9894);
and U10076 (N_10076,N_9889,N_9990);
and U10077 (N_10077,N_9961,N_9907);
nor U10078 (N_10078,N_9906,N_9947);
xnor U10079 (N_10079,N_9927,N_9902);
nor U10080 (N_10080,N_9956,N_9891);
and U10081 (N_10081,N_9894,N_9918);
nor U10082 (N_10082,N_9925,N_9881);
or U10083 (N_10083,N_9996,N_9922);
nand U10084 (N_10084,N_9897,N_9985);
or U10085 (N_10085,N_9881,N_9970);
nand U10086 (N_10086,N_9982,N_9924);
or U10087 (N_10087,N_9916,N_9931);
or U10088 (N_10088,N_9920,N_9941);
nand U10089 (N_10089,N_9907,N_9915);
and U10090 (N_10090,N_9941,N_9940);
or U10091 (N_10091,N_9881,N_9931);
nor U10092 (N_10092,N_9959,N_9881);
and U10093 (N_10093,N_9883,N_9913);
nor U10094 (N_10094,N_9959,N_9967);
and U10095 (N_10095,N_9982,N_9944);
nor U10096 (N_10096,N_9926,N_9937);
and U10097 (N_10097,N_9904,N_9908);
or U10098 (N_10098,N_9964,N_9996);
or U10099 (N_10099,N_9942,N_9979);
nand U10100 (N_10100,N_9921,N_9898);
xor U10101 (N_10101,N_9929,N_9941);
and U10102 (N_10102,N_9917,N_9994);
or U10103 (N_10103,N_9955,N_9915);
and U10104 (N_10104,N_9974,N_9987);
nor U10105 (N_10105,N_9891,N_9978);
and U10106 (N_10106,N_9884,N_9891);
or U10107 (N_10107,N_9940,N_9884);
and U10108 (N_10108,N_9928,N_9918);
or U10109 (N_10109,N_9878,N_9907);
xnor U10110 (N_10110,N_9902,N_9922);
nand U10111 (N_10111,N_9931,N_9937);
or U10112 (N_10112,N_9879,N_9967);
nor U10113 (N_10113,N_9991,N_9922);
nor U10114 (N_10114,N_9958,N_9967);
nor U10115 (N_10115,N_9920,N_9919);
nor U10116 (N_10116,N_9992,N_9887);
and U10117 (N_10117,N_9984,N_9911);
xnor U10118 (N_10118,N_9928,N_9890);
nor U10119 (N_10119,N_9945,N_9897);
nor U10120 (N_10120,N_9924,N_9876);
nand U10121 (N_10121,N_9987,N_9893);
nor U10122 (N_10122,N_9899,N_9894);
xor U10123 (N_10123,N_9878,N_9886);
nor U10124 (N_10124,N_9956,N_9995);
nand U10125 (N_10125,N_10114,N_10111);
xnor U10126 (N_10126,N_10119,N_10122);
nand U10127 (N_10127,N_10056,N_10101);
nor U10128 (N_10128,N_10120,N_10099);
or U10129 (N_10129,N_10094,N_10042);
or U10130 (N_10130,N_10040,N_10096);
and U10131 (N_10131,N_10005,N_10029);
xor U10132 (N_10132,N_10121,N_10009);
or U10133 (N_10133,N_10001,N_10053);
nor U10134 (N_10134,N_10086,N_10062);
nand U10135 (N_10135,N_10065,N_10081);
nor U10136 (N_10136,N_10004,N_10051);
nand U10137 (N_10137,N_10034,N_10061);
nand U10138 (N_10138,N_10017,N_10044);
or U10139 (N_10139,N_10106,N_10124);
nor U10140 (N_10140,N_10075,N_10091);
or U10141 (N_10141,N_10037,N_10104);
or U10142 (N_10142,N_10010,N_10033);
xor U10143 (N_10143,N_10109,N_10048);
and U10144 (N_10144,N_10028,N_10045);
or U10145 (N_10145,N_10107,N_10074);
and U10146 (N_10146,N_10024,N_10082);
or U10147 (N_10147,N_10123,N_10014);
and U10148 (N_10148,N_10026,N_10097);
and U10149 (N_10149,N_10116,N_10043);
xor U10150 (N_10150,N_10023,N_10006);
or U10151 (N_10151,N_10100,N_10118);
nor U10152 (N_10152,N_10018,N_10013);
nor U10153 (N_10153,N_10093,N_10077);
nand U10154 (N_10154,N_10103,N_10021);
or U10155 (N_10155,N_10039,N_10066);
nor U10156 (N_10156,N_10059,N_10000);
and U10157 (N_10157,N_10060,N_10089);
nor U10158 (N_10158,N_10105,N_10079);
xor U10159 (N_10159,N_10041,N_10036);
xnor U10160 (N_10160,N_10072,N_10115);
or U10161 (N_10161,N_10108,N_10069);
and U10162 (N_10162,N_10102,N_10087);
xor U10163 (N_10163,N_10113,N_10070);
xor U10164 (N_10164,N_10085,N_10073);
or U10165 (N_10165,N_10090,N_10052);
nand U10166 (N_10166,N_10031,N_10046);
nand U10167 (N_10167,N_10055,N_10025);
nand U10168 (N_10168,N_10002,N_10088);
nand U10169 (N_10169,N_10110,N_10003);
nand U10170 (N_10170,N_10071,N_10117);
and U10171 (N_10171,N_10080,N_10092);
or U10172 (N_10172,N_10027,N_10032);
nor U10173 (N_10173,N_10016,N_10067);
nand U10174 (N_10174,N_10057,N_10076);
nand U10175 (N_10175,N_10054,N_10022);
nand U10176 (N_10176,N_10019,N_10112);
nand U10177 (N_10177,N_10063,N_10058);
nand U10178 (N_10178,N_10038,N_10012);
nor U10179 (N_10179,N_10015,N_10083);
nand U10180 (N_10180,N_10084,N_10049);
nand U10181 (N_10181,N_10035,N_10064);
and U10182 (N_10182,N_10078,N_10047);
or U10183 (N_10183,N_10098,N_10030);
or U10184 (N_10184,N_10068,N_10050);
nand U10185 (N_10185,N_10095,N_10008);
xor U10186 (N_10186,N_10007,N_10011);
and U10187 (N_10187,N_10020,N_10063);
nor U10188 (N_10188,N_10042,N_10034);
and U10189 (N_10189,N_10078,N_10110);
and U10190 (N_10190,N_10092,N_10017);
or U10191 (N_10191,N_10122,N_10030);
nand U10192 (N_10192,N_10078,N_10057);
and U10193 (N_10193,N_10068,N_10060);
nor U10194 (N_10194,N_10060,N_10026);
nor U10195 (N_10195,N_10005,N_10065);
and U10196 (N_10196,N_10049,N_10002);
nor U10197 (N_10197,N_10043,N_10122);
or U10198 (N_10198,N_10119,N_10103);
nor U10199 (N_10199,N_10033,N_10065);
and U10200 (N_10200,N_10101,N_10114);
or U10201 (N_10201,N_10060,N_10023);
nor U10202 (N_10202,N_10036,N_10004);
nor U10203 (N_10203,N_10013,N_10112);
and U10204 (N_10204,N_10049,N_10124);
and U10205 (N_10205,N_10076,N_10001);
xor U10206 (N_10206,N_10087,N_10004);
or U10207 (N_10207,N_10043,N_10001);
nor U10208 (N_10208,N_10001,N_10035);
and U10209 (N_10209,N_10012,N_10004);
and U10210 (N_10210,N_10078,N_10020);
xnor U10211 (N_10211,N_10072,N_10068);
nand U10212 (N_10212,N_10075,N_10080);
or U10213 (N_10213,N_10087,N_10070);
nor U10214 (N_10214,N_10112,N_10078);
and U10215 (N_10215,N_10076,N_10073);
and U10216 (N_10216,N_10033,N_10046);
or U10217 (N_10217,N_10101,N_10039);
nand U10218 (N_10218,N_10053,N_10111);
and U10219 (N_10219,N_10054,N_10089);
or U10220 (N_10220,N_10070,N_10111);
xor U10221 (N_10221,N_10023,N_10111);
nand U10222 (N_10222,N_10082,N_10027);
and U10223 (N_10223,N_10055,N_10067);
nor U10224 (N_10224,N_10038,N_10057);
or U10225 (N_10225,N_10057,N_10110);
and U10226 (N_10226,N_10080,N_10121);
nor U10227 (N_10227,N_10001,N_10017);
nor U10228 (N_10228,N_10003,N_10114);
or U10229 (N_10229,N_10021,N_10051);
nand U10230 (N_10230,N_10118,N_10083);
nor U10231 (N_10231,N_10092,N_10039);
nor U10232 (N_10232,N_10054,N_10011);
nand U10233 (N_10233,N_10072,N_10051);
nand U10234 (N_10234,N_10039,N_10060);
nor U10235 (N_10235,N_10061,N_10096);
or U10236 (N_10236,N_10059,N_10018);
nand U10237 (N_10237,N_10028,N_10003);
or U10238 (N_10238,N_10070,N_10097);
or U10239 (N_10239,N_10065,N_10109);
nand U10240 (N_10240,N_10054,N_10010);
nand U10241 (N_10241,N_10061,N_10003);
nor U10242 (N_10242,N_10099,N_10023);
nor U10243 (N_10243,N_10070,N_10008);
or U10244 (N_10244,N_10097,N_10121);
and U10245 (N_10245,N_10032,N_10121);
and U10246 (N_10246,N_10038,N_10054);
nand U10247 (N_10247,N_10098,N_10092);
nand U10248 (N_10248,N_10082,N_10045);
and U10249 (N_10249,N_10066,N_10034);
or U10250 (N_10250,N_10246,N_10184);
nor U10251 (N_10251,N_10227,N_10170);
nor U10252 (N_10252,N_10203,N_10174);
nand U10253 (N_10253,N_10139,N_10213);
xnor U10254 (N_10254,N_10209,N_10158);
nor U10255 (N_10255,N_10215,N_10163);
nor U10256 (N_10256,N_10175,N_10191);
and U10257 (N_10257,N_10204,N_10222);
nor U10258 (N_10258,N_10127,N_10199);
or U10259 (N_10259,N_10216,N_10181);
nor U10260 (N_10260,N_10171,N_10176);
or U10261 (N_10261,N_10190,N_10237);
nor U10262 (N_10262,N_10146,N_10224);
nand U10263 (N_10263,N_10189,N_10136);
xnor U10264 (N_10264,N_10148,N_10172);
or U10265 (N_10265,N_10206,N_10161);
nor U10266 (N_10266,N_10233,N_10142);
nand U10267 (N_10267,N_10225,N_10244);
nand U10268 (N_10268,N_10223,N_10128);
xnor U10269 (N_10269,N_10177,N_10143);
nor U10270 (N_10270,N_10135,N_10201);
or U10271 (N_10271,N_10221,N_10141);
nor U10272 (N_10272,N_10238,N_10165);
and U10273 (N_10273,N_10164,N_10229);
nor U10274 (N_10274,N_10182,N_10147);
or U10275 (N_10275,N_10187,N_10242);
or U10276 (N_10276,N_10219,N_10188);
or U10277 (N_10277,N_10228,N_10180);
nand U10278 (N_10278,N_10166,N_10198);
and U10279 (N_10279,N_10160,N_10214);
nand U10280 (N_10280,N_10168,N_10197);
and U10281 (N_10281,N_10193,N_10248);
and U10282 (N_10282,N_10236,N_10153);
nand U10283 (N_10283,N_10235,N_10151);
nand U10284 (N_10284,N_10126,N_10162);
or U10285 (N_10285,N_10167,N_10212);
and U10286 (N_10286,N_10217,N_10230);
xnor U10287 (N_10287,N_10194,N_10226);
xor U10288 (N_10288,N_10132,N_10241);
and U10289 (N_10289,N_10173,N_10149);
nor U10290 (N_10290,N_10155,N_10133);
and U10291 (N_10291,N_10208,N_10239);
nor U10292 (N_10292,N_10131,N_10130);
or U10293 (N_10293,N_10159,N_10178);
xor U10294 (N_10294,N_10210,N_10249);
and U10295 (N_10295,N_10240,N_10137);
nor U10296 (N_10296,N_10156,N_10185);
nor U10297 (N_10297,N_10183,N_10202);
nor U10298 (N_10298,N_10134,N_10231);
and U10299 (N_10299,N_10207,N_10150);
nor U10300 (N_10300,N_10195,N_10218);
nor U10301 (N_10301,N_10234,N_10152);
xor U10302 (N_10302,N_10192,N_10140);
or U10303 (N_10303,N_10196,N_10125);
nor U10304 (N_10304,N_10205,N_10247);
nor U10305 (N_10305,N_10169,N_10145);
or U10306 (N_10306,N_10154,N_10186);
nand U10307 (N_10307,N_10179,N_10138);
or U10308 (N_10308,N_10200,N_10211);
and U10309 (N_10309,N_10243,N_10245);
or U10310 (N_10310,N_10220,N_10129);
nand U10311 (N_10311,N_10157,N_10144);
nor U10312 (N_10312,N_10232,N_10219);
nor U10313 (N_10313,N_10237,N_10231);
nor U10314 (N_10314,N_10174,N_10213);
and U10315 (N_10315,N_10166,N_10183);
or U10316 (N_10316,N_10208,N_10133);
nor U10317 (N_10317,N_10160,N_10236);
nor U10318 (N_10318,N_10140,N_10134);
xor U10319 (N_10319,N_10248,N_10228);
nor U10320 (N_10320,N_10186,N_10222);
and U10321 (N_10321,N_10222,N_10192);
nor U10322 (N_10322,N_10173,N_10147);
and U10323 (N_10323,N_10219,N_10227);
nor U10324 (N_10324,N_10168,N_10145);
nand U10325 (N_10325,N_10225,N_10141);
or U10326 (N_10326,N_10222,N_10151);
nand U10327 (N_10327,N_10136,N_10133);
or U10328 (N_10328,N_10142,N_10167);
nand U10329 (N_10329,N_10246,N_10185);
nor U10330 (N_10330,N_10175,N_10193);
or U10331 (N_10331,N_10206,N_10154);
nand U10332 (N_10332,N_10218,N_10222);
nor U10333 (N_10333,N_10199,N_10225);
or U10334 (N_10334,N_10236,N_10149);
or U10335 (N_10335,N_10202,N_10234);
and U10336 (N_10336,N_10213,N_10225);
and U10337 (N_10337,N_10170,N_10178);
and U10338 (N_10338,N_10156,N_10207);
or U10339 (N_10339,N_10146,N_10186);
nor U10340 (N_10340,N_10210,N_10238);
nor U10341 (N_10341,N_10170,N_10226);
nor U10342 (N_10342,N_10145,N_10214);
nor U10343 (N_10343,N_10170,N_10248);
and U10344 (N_10344,N_10178,N_10206);
and U10345 (N_10345,N_10164,N_10141);
or U10346 (N_10346,N_10243,N_10184);
nand U10347 (N_10347,N_10233,N_10234);
xnor U10348 (N_10348,N_10177,N_10146);
and U10349 (N_10349,N_10148,N_10131);
or U10350 (N_10350,N_10198,N_10171);
nor U10351 (N_10351,N_10154,N_10248);
nand U10352 (N_10352,N_10158,N_10167);
nor U10353 (N_10353,N_10135,N_10202);
nor U10354 (N_10354,N_10247,N_10231);
and U10355 (N_10355,N_10214,N_10236);
and U10356 (N_10356,N_10205,N_10234);
or U10357 (N_10357,N_10125,N_10246);
or U10358 (N_10358,N_10246,N_10137);
nand U10359 (N_10359,N_10140,N_10210);
and U10360 (N_10360,N_10228,N_10158);
nand U10361 (N_10361,N_10239,N_10129);
xnor U10362 (N_10362,N_10154,N_10223);
or U10363 (N_10363,N_10219,N_10144);
or U10364 (N_10364,N_10188,N_10139);
nor U10365 (N_10365,N_10129,N_10167);
nor U10366 (N_10366,N_10176,N_10165);
or U10367 (N_10367,N_10160,N_10163);
xnor U10368 (N_10368,N_10196,N_10178);
or U10369 (N_10369,N_10162,N_10145);
and U10370 (N_10370,N_10195,N_10216);
and U10371 (N_10371,N_10168,N_10211);
nor U10372 (N_10372,N_10169,N_10224);
xnor U10373 (N_10373,N_10246,N_10164);
nand U10374 (N_10374,N_10164,N_10206);
nor U10375 (N_10375,N_10371,N_10343);
or U10376 (N_10376,N_10308,N_10283);
and U10377 (N_10377,N_10270,N_10366);
and U10378 (N_10378,N_10305,N_10304);
nand U10379 (N_10379,N_10265,N_10340);
or U10380 (N_10380,N_10339,N_10361);
or U10381 (N_10381,N_10354,N_10258);
and U10382 (N_10382,N_10275,N_10303);
xor U10383 (N_10383,N_10274,N_10309);
or U10384 (N_10384,N_10373,N_10284);
nand U10385 (N_10385,N_10315,N_10324);
nand U10386 (N_10386,N_10316,N_10319);
nand U10387 (N_10387,N_10286,N_10299);
nor U10388 (N_10388,N_10374,N_10273);
nand U10389 (N_10389,N_10292,N_10328);
nand U10390 (N_10390,N_10297,N_10266);
nor U10391 (N_10391,N_10257,N_10337);
and U10392 (N_10392,N_10254,N_10353);
nor U10393 (N_10393,N_10325,N_10289);
nor U10394 (N_10394,N_10259,N_10296);
and U10395 (N_10395,N_10261,N_10307);
and U10396 (N_10396,N_10322,N_10314);
and U10397 (N_10397,N_10280,N_10278);
or U10398 (N_10398,N_10345,N_10294);
nand U10399 (N_10399,N_10360,N_10341);
or U10400 (N_10400,N_10331,N_10276);
nand U10401 (N_10401,N_10349,N_10302);
or U10402 (N_10402,N_10348,N_10293);
nor U10403 (N_10403,N_10369,N_10277);
and U10404 (N_10404,N_10352,N_10350);
or U10405 (N_10405,N_10312,N_10317);
nor U10406 (N_10406,N_10363,N_10300);
nand U10407 (N_10407,N_10263,N_10272);
nand U10408 (N_10408,N_10368,N_10279);
or U10409 (N_10409,N_10321,N_10344);
and U10410 (N_10410,N_10342,N_10281);
nand U10411 (N_10411,N_10295,N_10268);
and U10412 (N_10412,N_10320,N_10362);
nand U10413 (N_10413,N_10267,N_10359);
nand U10414 (N_10414,N_10327,N_10334);
nand U10415 (N_10415,N_10365,N_10290);
nor U10416 (N_10416,N_10264,N_10330);
nor U10417 (N_10417,N_10333,N_10255);
nor U10418 (N_10418,N_10346,N_10357);
and U10419 (N_10419,N_10311,N_10253);
or U10420 (N_10420,N_10370,N_10262);
xor U10421 (N_10421,N_10351,N_10298);
nor U10422 (N_10422,N_10269,N_10306);
or U10423 (N_10423,N_10271,N_10260);
or U10424 (N_10424,N_10326,N_10358);
and U10425 (N_10425,N_10364,N_10355);
or U10426 (N_10426,N_10313,N_10288);
nor U10427 (N_10427,N_10338,N_10372);
or U10428 (N_10428,N_10282,N_10291);
xnor U10429 (N_10429,N_10251,N_10256);
and U10430 (N_10430,N_10336,N_10332);
xnor U10431 (N_10431,N_10310,N_10285);
or U10432 (N_10432,N_10323,N_10367);
nand U10433 (N_10433,N_10347,N_10250);
nand U10434 (N_10434,N_10329,N_10287);
nand U10435 (N_10435,N_10252,N_10301);
nand U10436 (N_10436,N_10356,N_10335);
and U10437 (N_10437,N_10318,N_10329);
nand U10438 (N_10438,N_10328,N_10290);
nor U10439 (N_10439,N_10291,N_10323);
nand U10440 (N_10440,N_10374,N_10369);
nor U10441 (N_10441,N_10293,N_10281);
or U10442 (N_10442,N_10352,N_10371);
and U10443 (N_10443,N_10278,N_10331);
or U10444 (N_10444,N_10363,N_10370);
xnor U10445 (N_10445,N_10332,N_10309);
or U10446 (N_10446,N_10359,N_10373);
nand U10447 (N_10447,N_10255,N_10263);
or U10448 (N_10448,N_10284,N_10252);
nor U10449 (N_10449,N_10305,N_10354);
nor U10450 (N_10450,N_10366,N_10294);
and U10451 (N_10451,N_10305,N_10348);
and U10452 (N_10452,N_10353,N_10299);
nor U10453 (N_10453,N_10327,N_10306);
and U10454 (N_10454,N_10271,N_10255);
nand U10455 (N_10455,N_10299,N_10289);
or U10456 (N_10456,N_10320,N_10305);
nor U10457 (N_10457,N_10302,N_10347);
xor U10458 (N_10458,N_10295,N_10297);
nor U10459 (N_10459,N_10367,N_10259);
and U10460 (N_10460,N_10262,N_10344);
or U10461 (N_10461,N_10291,N_10260);
nand U10462 (N_10462,N_10269,N_10335);
xnor U10463 (N_10463,N_10300,N_10313);
or U10464 (N_10464,N_10355,N_10350);
or U10465 (N_10465,N_10270,N_10297);
nor U10466 (N_10466,N_10253,N_10290);
xnor U10467 (N_10467,N_10286,N_10348);
nand U10468 (N_10468,N_10274,N_10278);
and U10469 (N_10469,N_10309,N_10271);
or U10470 (N_10470,N_10306,N_10322);
nor U10471 (N_10471,N_10360,N_10299);
nor U10472 (N_10472,N_10296,N_10305);
or U10473 (N_10473,N_10289,N_10275);
and U10474 (N_10474,N_10336,N_10373);
nor U10475 (N_10475,N_10367,N_10355);
nand U10476 (N_10476,N_10252,N_10277);
and U10477 (N_10477,N_10300,N_10352);
nand U10478 (N_10478,N_10310,N_10338);
nor U10479 (N_10479,N_10363,N_10288);
and U10480 (N_10480,N_10326,N_10346);
and U10481 (N_10481,N_10255,N_10342);
nand U10482 (N_10482,N_10359,N_10355);
or U10483 (N_10483,N_10273,N_10303);
nand U10484 (N_10484,N_10366,N_10272);
and U10485 (N_10485,N_10279,N_10316);
and U10486 (N_10486,N_10255,N_10254);
or U10487 (N_10487,N_10337,N_10357);
or U10488 (N_10488,N_10299,N_10293);
and U10489 (N_10489,N_10312,N_10347);
nand U10490 (N_10490,N_10362,N_10250);
nand U10491 (N_10491,N_10339,N_10296);
nor U10492 (N_10492,N_10331,N_10364);
or U10493 (N_10493,N_10346,N_10333);
nor U10494 (N_10494,N_10349,N_10303);
nor U10495 (N_10495,N_10264,N_10312);
nor U10496 (N_10496,N_10294,N_10282);
or U10497 (N_10497,N_10267,N_10358);
and U10498 (N_10498,N_10265,N_10308);
or U10499 (N_10499,N_10300,N_10285);
and U10500 (N_10500,N_10444,N_10474);
and U10501 (N_10501,N_10395,N_10380);
and U10502 (N_10502,N_10403,N_10451);
xnor U10503 (N_10503,N_10399,N_10384);
nand U10504 (N_10504,N_10385,N_10412);
nand U10505 (N_10505,N_10497,N_10437);
nand U10506 (N_10506,N_10475,N_10494);
or U10507 (N_10507,N_10427,N_10450);
and U10508 (N_10508,N_10470,N_10405);
or U10509 (N_10509,N_10484,N_10386);
or U10510 (N_10510,N_10445,N_10432);
or U10511 (N_10511,N_10430,N_10490);
or U10512 (N_10512,N_10415,N_10447);
or U10513 (N_10513,N_10473,N_10413);
and U10514 (N_10514,N_10382,N_10400);
nor U10515 (N_10515,N_10453,N_10376);
xor U10516 (N_10516,N_10377,N_10436);
nor U10517 (N_10517,N_10429,N_10411);
nand U10518 (N_10518,N_10393,N_10493);
nor U10519 (N_10519,N_10379,N_10381);
nor U10520 (N_10520,N_10397,N_10394);
nand U10521 (N_10521,N_10461,N_10407);
and U10522 (N_10522,N_10442,N_10392);
or U10523 (N_10523,N_10398,N_10478);
nor U10524 (N_10524,N_10387,N_10471);
nor U10525 (N_10525,N_10406,N_10479);
xnor U10526 (N_10526,N_10499,N_10454);
and U10527 (N_10527,N_10431,N_10489);
xor U10528 (N_10528,N_10465,N_10464);
or U10529 (N_10529,N_10416,N_10402);
nor U10530 (N_10530,N_10417,N_10375);
and U10531 (N_10531,N_10498,N_10457);
and U10532 (N_10532,N_10423,N_10483);
nor U10533 (N_10533,N_10463,N_10409);
and U10534 (N_10534,N_10396,N_10408);
nor U10535 (N_10535,N_10449,N_10481);
or U10536 (N_10536,N_10389,N_10410);
xor U10537 (N_10537,N_10455,N_10486);
xor U10538 (N_10538,N_10459,N_10462);
or U10539 (N_10539,N_10438,N_10476);
or U10540 (N_10540,N_10440,N_10456);
and U10541 (N_10541,N_10420,N_10448);
or U10542 (N_10542,N_10404,N_10388);
and U10543 (N_10543,N_10466,N_10468);
or U10544 (N_10544,N_10485,N_10428);
nor U10545 (N_10545,N_10458,N_10421);
nand U10546 (N_10546,N_10477,N_10460);
xor U10547 (N_10547,N_10401,N_10414);
nor U10548 (N_10548,N_10433,N_10488);
xor U10549 (N_10549,N_10452,N_10496);
nor U10550 (N_10550,N_10383,N_10441);
and U10551 (N_10551,N_10482,N_10391);
and U10552 (N_10552,N_10434,N_10487);
nand U10553 (N_10553,N_10492,N_10435);
or U10554 (N_10554,N_10467,N_10419);
or U10555 (N_10555,N_10491,N_10469);
nand U10556 (N_10556,N_10426,N_10424);
nor U10557 (N_10557,N_10443,N_10495);
nand U10558 (N_10558,N_10422,N_10418);
and U10559 (N_10559,N_10446,N_10480);
or U10560 (N_10560,N_10378,N_10472);
xnor U10561 (N_10561,N_10425,N_10439);
nand U10562 (N_10562,N_10390,N_10457);
nand U10563 (N_10563,N_10489,N_10403);
nor U10564 (N_10564,N_10402,N_10499);
or U10565 (N_10565,N_10378,N_10469);
nand U10566 (N_10566,N_10451,N_10419);
nor U10567 (N_10567,N_10396,N_10383);
nand U10568 (N_10568,N_10378,N_10459);
nand U10569 (N_10569,N_10490,N_10475);
nand U10570 (N_10570,N_10421,N_10403);
nand U10571 (N_10571,N_10475,N_10467);
and U10572 (N_10572,N_10426,N_10474);
and U10573 (N_10573,N_10484,N_10406);
or U10574 (N_10574,N_10402,N_10428);
and U10575 (N_10575,N_10427,N_10481);
or U10576 (N_10576,N_10440,N_10476);
and U10577 (N_10577,N_10406,N_10489);
or U10578 (N_10578,N_10407,N_10459);
nand U10579 (N_10579,N_10405,N_10450);
nor U10580 (N_10580,N_10467,N_10473);
nor U10581 (N_10581,N_10459,N_10461);
nor U10582 (N_10582,N_10489,N_10392);
or U10583 (N_10583,N_10441,N_10448);
and U10584 (N_10584,N_10461,N_10485);
nor U10585 (N_10585,N_10496,N_10424);
and U10586 (N_10586,N_10459,N_10413);
and U10587 (N_10587,N_10488,N_10384);
nor U10588 (N_10588,N_10390,N_10463);
nand U10589 (N_10589,N_10455,N_10446);
nor U10590 (N_10590,N_10425,N_10410);
nor U10591 (N_10591,N_10495,N_10391);
and U10592 (N_10592,N_10468,N_10473);
nor U10593 (N_10593,N_10470,N_10454);
and U10594 (N_10594,N_10468,N_10487);
nor U10595 (N_10595,N_10388,N_10440);
or U10596 (N_10596,N_10375,N_10394);
nand U10597 (N_10597,N_10474,N_10495);
nand U10598 (N_10598,N_10393,N_10465);
and U10599 (N_10599,N_10437,N_10479);
nor U10600 (N_10600,N_10476,N_10463);
nand U10601 (N_10601,N_10452,N_10376);
nand U10602 (N_10602,N_10430,N_10449);
nand U10603 (N_10603,N_10467,N_10377);
and U10604 (N_10604,N_10433,N_10481);
nand U10605 (N_10605,N_10436,N_10440);
and U10606 (N_10606,N_10400,N_10434);
xor U10607 (N_10607,N_10481,N_10389);
nor U10608 (N_10608,N_10398,N_10402);
nor U10609 (N_10609,N_10466,N_10404);
and U10610 (N_10610,N_10480,N_10407);
and U10611 (N_10611,N_10377,N_10478);
and U10612 (N_10612,N_10433,N_10423);
and U10613 (N_10613,N_10478,N_10397);
and U10614 (N_10614,N_10424,N_10411);
or U10615 (N_10615,N_10408,N_10496);
nand U10616 (N_10616,N_10404,N_10438);
nor U10617 (N_10617,N_10416,N_10400);
or U10618 (N_10618,N_10438,N_10465);
xor U10619 (N_10619,N_10401,N_10424);
nor U10620 (N_10620,N_10377,N_10448);
or U10621 (N_10621,N_10478,N_10449);
xnor U10622 (N_10622,N_10426,N_10400);
and U10623 (N_10623,N_10447,N_10395);
nor U10624 (N_10624,N_10391,N_10457);
nor U10625 (N_10625,N_10521,N_10606);
xor U10626 (N_10626,N_10567,N_10533);
nand U10627 (N_10627,N_10554,N_10578);
or U10628 (N_10628,N_10590,N_10575);
or U10629 (N_10629,N_10559,N_10539);
and U10630 (N_10630,N_10501,N_10582);
nor U10631 (N_10631,N_10502,N_10570);
nand U10632 (N_10632,N_10619,N_10574);
nand U10633 (N_10633,N_10548,N_10523);
nor U10634 (N_10634,N_10584,N_10609);
or U10635 (N_10635,N_10527,N_10618);
nor U10636 (N_10636,N_10563,N_10610);
xor U10637 (N_10637,N_10564,N_10596);
or U10638 (N_10638,N_10576,N_10580);
nand U10639 (N_10639,N_10601,N_10586);
nor U10640 (N_10640,N_10552,N_10566);
nand U10641 (N_10641,N_10506,N_10538);
nor U10642 (N_10642,N_10510,N_10519);
nor U10643 (N_10643,N_10603,N_10540);
nor U10644 (N_10644,N_10617,N_10615);
or U10645 (N_10645,N_10518,N_10534);
nor U10646 (N_10646,N_10505,N_10612);
and U10647 (N_10647,N_10604,N_10543);
nand U10648 (N_10648,N_10551,N_10513);
or U10649 (N_10649,N_10556,N_10550);
and U10650 (N_10650,N_10520,N_10500);
nor U10651 (N_10651,N_10613,N_10600);
and U10652 (N_10652,N_10621,N_10605);
or U10653 (N_10653,N_10542,N_10583);
and U10654 (N_10654,N_10589,N_10591);
or U10655 (N_10655,N_10611,N_10545);
nand U10656 (N_10656,N_10547,N_10560);
nor U10657 (N_10657,N_10561,N_10525);
nor U10658 (N_10658,N_10546,N_10624);
and U10659 (N_10659,N_10515,N_10508);
nand U10660 (N_10660,N_10588,N_10544);
nor U10661 (N_10661,N_10622,N_10562);
or U10662 (N_10662,N_10568,N_10614);
nand U10663 (N_10663,N_10581,N_10524);
or U10664 (N_10664,N_10598,N_10608);
and U10665 (N_10665,N_10503,N_10579);
or U10666 (N_10666,N_10607,N_10577);
nand U10667 (N_10667,N_10587,N_10531);
nor U10668 (N_10668,N_10571,N_10569);
nand U10669 (N_10669,N_10595,N_10592);
or U10670 (N_10670,N_10530,N_10549);
or U10671 (N_10671,N_10529,N_10504);
nor U10672 (N_10672,N_10585,N_10565);
nor U10673 (N_10673,N_10541,N_10537);
or U10674 (N_10674,N_10532,N_10557);
nor U10675 (N_10675,N_10516,N_10616);
or U10676 (N_10676,N_10599,N_10593);
or U10677 (N_10677,N_10558,N_10594);
and U10678 (N_10678,N_10602,N_10522);
nand U10679 (N_10679,N_10511,N_10528);
nor U10680 (N_10680,N_10526,N_10623);
and U10681 (N_10681,N_10535,N_10517);
and U10682 (N_10682,N_10572,N_10536);
nor U10683 (N_10683,N_10514,N_10512);
xnor U10684 (N_10684,N_10573,N_10597);
nand U10685 (N_10685,N_10553,N_10507);
nand U10686 (N_10686,N_10555,N_10509);
nand U10687 (N_10687,N_10620,N_10553);
nor U10688 (N_10688,N_10516,N_10607);
or U10689 (N_10689,N_10614,N_10569);
nand U10690 (N_10690,N_10598,N_10596);
nor U10691 (N_10691,N_10558,N_10623);
and U10692 (N_10692,N_10527,N_10562);
or U10693 (N_10693,N_10621,N_10529);
and U10694 (N_10694,N_10546,N_10510);
nor U10695 (N_10695,N_10602,N_10555);
nand U10696 (N_10696,N_10586,N_10623);
and U10697 (N_10697,N_10506,N_10582);
or U10698 (N_10698,N_10512,N_10607);
or U10699 (N_10699,N_10614,N_10571);
and U10700 (N_10700,N_10512,N_10622);
or U10701 (N_10701,N_10580,N_10568);
or U10702 (N_10702,N_10548,N_10608);
nand U10703 (N_10703,N_10542,N_10500);
nand U10704 (N_10704,N_10529,N_10623);
or U10705 (N_10705,N_10557,N_10597);
nand U10706 (N_10706,N_10563,N_10542);
nand U10707 (N_10707,N_10615,N_10552);
xor U10708 (N_10708,N_10510,N_10544);
and U10709 (N_10709,N_10528,N_10531);
and U10710 (N_10710,N_10521,N_10612);
xnor U10711 (N_10711,N_10604,N_10590);
xnor U10712 (N_10712,N_10555,N_10522);
nand U10713 (N_10713,N_10600,N_10524);
nor U10714 (N_10714,N_10507,N_10543);
nor U10715 (N_10715,N_10505,N_10619);
or U10716 (N_10716,N_10505,N_10608);
and U10717 (N_10717,N_10556,N_10528);
nor U10718 (N_10718,N_10577,N_10586);
or U10719 (N_10719,N_10551,N_10537);
nand U10720 (N_10720,N_10577,N_10515);
xor U10721 (N_10721,N_10555,N_10533);
or U10722 (N_10722,N_10551,N_10561);
nor U10723 (N_10723,N_10500,N_10527);
nor U10724 (N_10724,N_10558,N_10577);
nor U10725 (N_10725,N_10500,N_10579);
and U10726 (N_10726,N_10535,N_10525);
nor U10727 (N_10727,N_10611,N_10539);
or U10728 (N_10728,N_10608,N_10595);
nand U10729 (N_10729,N_10608,N_10559);
or U10730 (N_10730,N_10598,N_10623);
and U10731 (N_10731,N_10569,N_10608);
or U10732 (N_10732,N_10538,N_10622);
and U10733 (N_10733,N_10605,N_10509);
and U10734 (N_10734,N_10617,N_10581);
and U10735 (N_10735,N_10507,N_10583);
xor U10736 (N_10736,N_10576,N_10575);
nand U10737 (N_10737,N_10606,N_10562);
nor U10738 (N_10738,N_10618,N_10607);
xnor U10739 (N_10739,N_10507,N_10547);
xnor U10740 (N_10740,N_10524,N_10556);
xor U10741 (N_10741,N_10595,N_10577);
and U10742 (N_10742,N_10581,N_10555);
nand U10743 (N_10743,N_10567,N_10515);
and U10744 (N_10744,N_10511,N_10620);
and U10745 (N_10745,N_10587,N_10524);
xor U10746 (N_10746,N_10591,N_10550);
nor U10747 (N_10747,N_10557,N_10540);
and U10748 (N_10748,N_10521,N_10503);
and U10749 (N_10749,N_10531,N_10602);
nand U10750 (N_10750,N_10691,N_10637);
and U10751 (N_10751,N_10720,N_10702);
xnor U10752 (N_10752,N_10653,N_10713);
nor U10753 (N_10753,N_10701,N_10655);
or U10754 (N_10754,N_10672,N_10717);
nor U10755 (N_10755,N_10731,N_10658);
nand U10756 (N_10756,N_10721,N_10670);
nor U10757 (N_10757,N_10686,N_10738);
xnor U10758 (N_10758,N_10679,N_10735);
xnor U10759 (N_10759,N_10742,N_10633);
xnor U10760 (N_10760,N_10728,N_10725);
nand U10761 (N_10761,N_10671,N_10740);
nor U10762 (N_10762,N_10675,N_10693);
and U10763 (N_10763,N_10696,N_10643);
and U10764 (N_10764,N_10724,N_10695);
nand U10765 (N_10765,N_10668,N_10642);
or U10766 (N_10766,N_10715,N_10677);
and U10767 (N_10767,N_10688,N_10659);
nor U10768 (N_10768,N_10685,N_10704);
nand U10769 (N_10769,N_10690,N_10714);
nand U10770 (N_10770,N_10698,N_10716);
nand U10771 (N_10771,N_10711,N_10689);
nand U10772 (N_10772,N_10667,N_10710);
nand U10773 (N_10773,N_10629,N_10663);
nor U10774 (N_10774,N_10632,N_10627);
nor U10775 (N_10775,N_10748,N_10648);
xor U10776 (N_10776,N_10645,N_10649);
or U10777 (N_10777,N_10638,N_10626);
nand U10778 (N_10778,N_10640,N_10708);
nor U10779 (N_10779,N_10635,N_10682);
and U10780 (N_10780,N_10683,N_10700);
and U10781 (N_10781,N_10732,N_10630);
nor U10782 (N_10782,N_10674,N_10719);
nor U10783 (N_10783,N_10703,N_10729);
and U10784 (N_10784,N_10747,N_10694);
and U10785 (N_10785,N_10749,N_10644);
or U10786 (N_10786,N_10687,N_10692);
nor U10787 (N_10787,N_10636,N_10722);
and U10788 (N_10788,N_10656,N_10712);
nand U10789 (N_10789,N_10739,N_10718);
and U10790 (N_10790,N_10743,N_10723);
nand U10791 (N_10791,N_10736,N_10662);
or U10792 (N_10792,N_10625,N_10699);
nand U10793 (N_10793,N_10697,N_10706);
nor U10794 (N_10794,N_10661,N_10650);
nand U10795 (N_10795,N_10666,N_10727);
and U10796 (N_10796,N_10664,N_10657);
nand U10797 (N_10797,N_10681,N_10639);
nand U10798 (N_10798,N_10665,N_10654);
nand U10799 (N_10799,N_10646,N_10741);
or U10800 (N_10800,N_10669,N_10745);
or U10801 (N_10801,N_10730,N_10641);
nor U10802 (N_10802,N_10707,N_10734);
nor U10803 (N_10803,N_10746,N_10660);
xor U10804 (N_10804,N_10684,N_10705);
or U10805 (N_10805,N_10652,N_10647);
xor U10806 (N_10806,N_10676,N_10726);
or U10807 (N_10807,N_10634,N_10628);
and U10808 (N_10808,N_10631,N_10733);
and U10809 (N_10809,N_10680,N_10673);
nand U10810 (N_10810,N_10678,N_10737);
nor U10811 (N_10811,N_10651,N_10744);
nand U10812 (N_10812,N_10709,N_10678);
nand U10813 (N_10813,N_10746,N_10730);
and U10814 (N_10814,N_10684,N_10717);
nor U10815 (N_10815,N_10633,N_10685);
and U10816 (N_10816,N_10625,N_10692);
or U10817 (N_10817,N_10674,N_10638);
nor U10818 (N_10818,N_10646,N_10674);
and U10819 (N_10819,N_10676,N_10702);
nand U10820 (N_10820,N_10686,N_10701);
nand U10821 (N_10821,N_10720,N_10649);
and U10822 (N_10822,N_10744,N_10708);
or U10823 (N_10823,N_10673,N_10711);
nand U10824 (N_10824,N_10665,N_10749);
or U10825 (N_10825,N_10712,N_10649);
nand U10826 (N_10826,N_10665,N_10670);
and U10827 (N_10827,N_10670,N_10698);
nand U10828 (N_10828,N_10686,N_10693);
and U10829 (N_10829,N_10656,N_10679);
or U10830 (N_10830,N_10631,N_10696);
or U10831 (N_10831,N_10687,N_10671);
nor U10832 (N_10832,N_10644,N_10728);
nand U10833 (N_10833,N_10670,N_10628);
nand U10834 (N_10834,N_10658,N_10668);
nor U10835 (N_10835,N_10648,N_10650);
xor U10836 (N_10836,N_10677,N_10720);
or U10837 (N_10837,N_10718,N_10654);
nor U10838 (N_10838,N_10698,N_10625);
and U10839 (N_10839,N_10740,N_10634);
nand U10840 (N_10840,N_10655,N_10736);
and U10841 (N_10841,N_10649,N_10641);
xor U10842 (N_10842,N_10718,N_10716);
and U10843 (N_10843,N_10713,N_10647);
or U10844 (N_10844,N_10704,N_10664);
or U10845 (N_10845,N_10681,N_10677);
or U10846 (N_10846,N_10651,N_10643);
and U10847 (N_10847,N_10698,N_10719);
or U10848 (N_10848,N_10740,N_10654);
and U10849 (N_10849,N_10688,N_10684);
nand U10850 (N_10850,N_10746,N_10747);
or U10851 (N_10851,N_10705,N_10722);
nor U10852 (N_10852,N_10692,N_10717);
and U10853 (N_10853,N_10724,N_10732);
and U10854 (N_10854,N_10660,N_10626);
or U10855 (N_10855,N_10740,N_10699);
and U10856 (N_10856,N_10633,N_10640);
nand U10857 (N_10857,N_10709,N_10719);
nand U10858 (N_10858,N_10676,N_10736);
nor U10859 (N_10859,N_10637,N_10712);
nand U10860 (N_10860,N_10746,N_10697);
nor U10861 (N_10861,N_10734,N_10682);
xnor U10862 (N_10862,N_10682,N_10715);
or U10863 (N_10863,N_10741,N_10659);
xnor U10864 (N_10864,N_10729,N_10692);
and U10865 (N_10865,N_10658,N_10718);
nor U10866 (N_10866,N_10662,N_10723);
nand U10867 (N_10867,N_10628,N_10718);
or U10868 (N_10868,N_10664,N_10746);
or U10869 (N_10869,N_10657,N_10681);
or U10870 (N_10870,N_10734,N_10625);
and U10871 (N_10871,N_10679,N_10687);
or U10872 (N_10872,N_10641,N_10711);
or U10873 (N_10873,N_10719,N_10694);
or U10874 (N_10874,N_10646,N_10650);
xnor U10875 (N_10875,N_10842,N_10821);
nand U10876 (N_10876,N_10808,N_10817);
xnor U10877 (N_10877,N_10823,N_10865);
and U10878 (N_10878,N_10784,N_10814);
nand U10879 (N_10879,N_10838,N_10780);
and U10880 (N_10880,N_10802,N_10871);
xnor U10881 (N_10881,N_10854,N_10827);
nand U10882 (N_10882,N_10778,N_10845);
and U10883 (N_10883,N_10757,N_10807);
and U10884 (N_10884,N_10753,N_10806);
or U10885 (N_10885,N_10826,N_10822);
or U10886 (N_10886,N_10825,N_10832);
and U10887 (N_10887,N_10799,N_10750);
nand U10888 (N_10888,N_10766,N_10840);
and U10889 (N_10889,N_10851,N_10794);
nor U10890 (N_10890,N_10834,N_10856);
nor U10891 (N_10891,N_10857,N_10759);
and U10892 (N_10892,N_10755,N_10874);
nand U10893 (N_10893,N_10855,N_10783);
nor U10894 (N_10894,N_10830,N_10764);
xor U10895 (N_10895,N_10828,N_10863);
or U10896 (N_10896,N_10797,N_10824);
and U10897 (N_10897,N_10763,N_10803);
and U10898 (N_10898,N_10793,N_10812);
or U10899 (N_10899,N_10813,N_10758);
or U10900 (N_10900,N_10815,N_10862);
and U10901 (N_10901,N_10770,N_10789);
or U10902 (N_10902,N_10870,N_10831);
and U10903 (N_10903,N_10788,N_10769);
nor U10904 (N_10904,N_10801,N_10833);
nand U10905 (N_10905,N_10752,N_10841);
nor U10906 (N_10906,N_10771,N_10796);
nand U10907 (N_10907,N_10810,N_10787);
or U10908 (N_10908,N_10848,N_10820);
or U10909 (N_10909,N_10775,N_10791);
or U10910 (N_10910,N_10765,N_10835);
nand U10911 (N_10911,N_10819,N_10804);
nor U10912 (N_10912,N_10847,N_10816);
and U10913 (N_10913,N_10768,N_10756);
nand U10914 (N_10914,N_10785,N_10839);
or U10915 (N_10915,N_10850,N_10846);
or U10916 (N_10916,N_10760,N_10761);
or U10917 (N_10917,N_10860,N_10866);
or U10918 (N_10918,N_10776,N_10811);
nor U10919 (N_10919,N_10836,N_10868);
and U10920 (N_10920,N_10782,N_10781);
or U10921 (N_10921,N_10777,N_10798);
and U10922 (N_10922,N_10844,N_10859);
nand U10923 (N_10923,N_10852,N_10861);
xnor U10924 (N_10924,N_10754,N_10867);
nor U10925 (N_10925,N_10790,N_10829);
and U10926 (N_10926,N_10837,N_10818);
or U10927 (N_10927,N_10751,N_10795);
nand U10928 (N_10928,N_10872,N_10772);
nor U10929 (N_10929,N_10805,N_10864);
and U10930 (N_10930,N_10849,N_10843);
nand U10931 (N_10931,N_10762,N_10767);
nor U10932 (N_10932,N_10779,N_10869);
and U10933 (N_10933,N_10786,N_10858);
and U10934 (N_10934,N_10809,N_10774);
nand U10935 (N_10935,N_10800,N_10853);
nor U10936 (N_10936,N_10792,N_10873);
or U10937 (N_10937,N_10773,N_10839);
nand U10938 (N_10938,N_10773,N_10763);
or U10939 (N_10939,N_10792,N_10770);
nor U10940 (N_10940,N_10853,N_10780);
or U10941 (N_10941,N_10776,N_10868);
xnor U10942 (N_10942,N_10776,N_10756);
and U10943 (N_10943,N_10765,N_10799);
and U10944 (N_10944,N_10847,N_10775);
nand U10945 (N_10945,N_10844,N_10760);
xnor U10946 (N_10946,N_10824,N_10802);
or U10947 (N_10947,N_10865,N_10755);
and U10948 (N_10948,N_10785,N_10800);
nor U10949 (N_10949,N_10800,N_10781);
or U10950 (N_10950,N_10784,N_10780);
nand U10951 (N_10951,N_10802,N_10791);
nand U10952 (N_10952,N_10846,N_10849);
and U10953 (N_10953,N_10767,N_10857);
nand U10954 (N_10954,N_10823,N_10824);
or U10955 (N_10955,N_10831,N_10865);
and U10956 (N_10956,N_10821,N_10831);
or U10957 (N_10957,N_10750,N_10856);
nand U10958 (N_10958,N_10867,N_10824);
and U10959 (N_10959,N_10867,N_10870);
or U10960 (N_10960,N_10775,N_10805);
xnor U10961 (N_10961,N_10864,N_10793);
or U10962 (N_10962,N_10868,N_10869);
and U10963 (N_10963,N_10821,N_10813);
or U10964 (N_10964,N_10761,N_10850);
and U10965 (N_10965,N_10867,N_10809);
and U10966 (N_10966,N_10863,N_10864);
and U10967 (N_10967,N_10867,N_10775);
and U10968 (N_10968,N_10858,N_10782);
and U10969 (N_10969,N_10854,N_10843);
xnor U10970 (N_10970,N_10806,N_10758);
nand U10971 (N_10971,N_10825,N_10870);
or U10972 (N_10972,N_10762,N_10755);
xnor U10973 (N_10973,N_10769,N_10822);
nand U10974 (N_10974,N_10784,N_10870);
or U10975 (N_10975,N_10757,N_10784);
or U10976 (N_10976,N_10845,N_10760);
or U10977 (N_10977,N_10778,N_10815);
or U10978 (N_10978,N_10826,N_10813);
and U10979 (N_10979,N_10839,N_10803);
or U10980 (N_10980,N_10843,N_10870);
xor U10981 (N_10981,N_10767,N_10770);
nand U10982 (N_10982,N_10811,N_10784);
nand U10983 (N_10983,N_10785,N_10818);
nor U10984 (N_10984,N_10783,N_10824);
or U10985 (N_10985,N_10782,N_10776);
and U10986 (N_10986,N_10750,N_10798);
nand U10987 (N_10987,N_10764,N_10761);
nand U10988 (N_10988,N_10795,N_10784);
or U10989 (N_10989,N_10789,N_10870);
nand U10990 (N_10990,N_10847,N_10852);
nor U10991 (N_10991,N_10792,N_10777);
xnor U10992 (N_10992,N_10835,N_10800);
or U10993 (N_10993,N_10765,N_10813);
nand U10994 (N_10994,N_10820,N_10823);
nand U10995 (N_10995,N_10839,N_10861);
xnor U10996 (N_10996,N_10763,N_10758);
nor U10997 (N_10997,N_10827,N_10819);
and U10998 (N_10998,N_10795,N_10846);
nand U10999 (N_10999,N_10792,N_10804);
nor U11000 (N_11000,N_10931,N_10966);
xnor U11001 (N_11001,N_10922,N_10996);
nor U11002 (N_11002,N_10921,N_10924);
nor U11003 (N_11003,N_10943,N_10881);
nor U11004 (N_11004,N_10913,N_10889);
or U11005 (N_11005,N_10901,N_10885);
nor U11006 (N_11006,N_10953,N_10884);
or U11007 (N_11007,N_10992,N_10986);
xnor U11008 (N_11008,N_10961,N_10916);
nor U11009 (N_11009,N_10995,N_10982);
and U11010 (N_11010,N_10886,N_10975);
nor U11011 (N_11011,N_10978,N_10910);
nor U11012 (N_11012,N_10907,N_10959);
xnor U11013 (N_11013,N_10951,N_10882);
nor U11014 (N_11014,N_10905,N_10941);
or U11015 (N_11015,N_10896,N_10918);
nor U11016 (N_11016,N_10987,N_10962);
nor U11017 (N_11017,N_10942,N_10970);
nand U11018 (N_11018,N_10993,N_10891);
and U11019 (N_11019,N_10976,N_10912);
or U11020 (N_11020,N_10888,N_10967);
and U11021 (N_11021,N_10906,N_10960);
nand U11022 (N_11022,N_10879,N_10950);
nor U11023 (N_11023,N_10923,N_10973);
or U11024 (N_11024,N_10897,N_10944);
nand U11025 (N_11025,N_10911,N_10964);
nand U11026 (N_11026,N_10955,N_10927);
nand U11027 (N_11027,N_10957,N_10917);
nor U11028 (N_11028,N_10972,N_10904);
and U11029 (N_11029,N_10935,N_10945);
nand U11030 (N_11030,N_10998,N_10877);
or U11031 (N_11031,N_10933,N_10939);
nand U11032 (N_11032,N_10936,N_10937);
and U11033 (N_11033,N_10919,N_10908);
nand U11034 (N_11034,N_10948,N_10974);
and U11035 (N_11035,N_10952,N_10963);
xnor U11036 (N_11036,N_10947,N_10979);
nor U11037 (N_11037,N_10909,N_10938);
or U11038 (N_11038,N_10969,N_10985);
or U11039 (N_11039,N_10893,N_10928);
nor U11040 (N_11040,N_10965,N_10971);
and U11041 (N_11041,N_10956,N_10898);
or U11042 (N_11042,N_10946,N_10954);
nor U11043 (N_11043,N_10929,N_10894);
and U11044 (N_11044,N_10899,N_10988);
and U11045 (N_11045,N_10981,N_10968);
xor U11046 (N_11046,N_10883,N_10925);
or U11047 (N_11047,N_10915,N_10926);
nor U11048 (N_11048,N_10994,N_10876);
nor U11049 (N_11049,N_10991,N_10983);
nor U11050 (N_11050,N_10875,N_10902);
or U11051 (N_11051,N_10890,N_10980);
and U11052 (N_11052,N_10977,N_10895);
nor U11053 (N_11053,N_10990,N_10984);
and U11054 (N_11054,N_10900,N_10940);
and U11055 (N_11055,N_10914,N_10999);
or U11056 (N_11056,N_10903,N_10989);
nor U11057 (N_11057,N_10958,N_10997);
nand U11058 (N_11058,N_10932,N_10920);
nor U11059 (N_11059,N_10949,N_10878);
or U11060 (N_11060,N_10880,N_10930);
or U11061 (N_11061,N_10892,N_10887);
and U11062 (N_11062,N_10934,N_10939);
nor U11063 (N_11063,N_10883,N_10967);
nand U11064 (N_11064,N_10998,N_10960);
and U11065 (N_11065,N_10899,N_10897);
and U11066 (N_11066,N_10989,N_10913);
nor U11067 (N_11067,N_10880,N_10894);
and U11068 (N_11068,N_10969,N_10962);
or U11069 (N_11069,N_10945,N_10968);
or U11070 (N_11070,N_10970,N_10926);
or U11071 (N_11071,N_10901,N_10945);
or U11072 (N_11072,N_10880,N_10952);
nor U11073 (N_11073,N_10903,N_10931);
and U11074 (N_11074,N_10901,N_10962);
nand U11075 (N_11075,N_10964,N_10953);
xor U11076 (N_11076,N_10922,N_10916);
nand U11077 (N_11077,N_10883,N_10914);
or U11078 (N_11078,N_10993,N_10927);
xor U11079 (N_11079,N_10933,N_10877);
nand U11080 (N_11080,N_10986,N_10944);
and U11081 (N_11081,N_10885,N_10928);
nor U11082 (N_11082,N_10903,N_10992);
and U11083 (N_11083,N_10999,N_10972);
and U11084 (N_11084,N_10924,N_10912);
or U11085 (N_11085,N_10913,N_10921);
nor U11086 (N_11086,N_10936,N_10908);
or U11087 (N_11087,N_10953,N_10882);
or U11088 (N_11088,N_10893,N_10938);
nor U11089 (N_11089,N_10972,N_10939);
or U11090 (N_11090,N_10885,N_10921);
and U11091 (N_11091,N_10939,N_10994);
nor U11092 (N_11092,N_10993,N_10896);
xnor U11093 (N_11093,N_10928,N_10917);
and U11094 (N_11094,N_10957,N_10887);
and U11095 (N_11095,N_10896,N_10960);
xor U11096 (N_11096,N_10877,N_10952);
and U11097 (N_11097,N_10882,N_10922);
or U11098 (N_11098,N_10968,N_10925);
nor U11099 (N_11099,N_10950,N_10880);
or U11100 (N_11100,N_10899,N_10880);
nor U11101 (N_11101,N_10978,N_10895);
or U11102 (N_11102,N_10914,N_10910);
nand U11103 (N_11103,N_10981,N_10993);
and U11104 (N_11104,N_10898,N_10912);
nand U11105 (N_11105,N_10956,N_10893);
nand U11106 (N_11106,N_10936,N_10933);
nand U11107 (N_11107,N_10942,N_10902);
or U11108 (N_11108,N_10878,N_10945);
or U11109 (N_11109,N_10965,N_10978);
xor U11110 (N_11110,N_10911,N_10989);
and U11111 (N_11111,N_10987,N_10950);
nand U11112 (N_11112,N_10932,N_10909);
or U11113 (N_11113,N_10919,N_10938);
and U11114 (N_11114,N_10923,N_10898);
nand U11115 (N_11115,N_10910,N_10913);
and U11116 (N_11116,N_10914,N_10944);
and U11117 (N_11117,N_10901,N_10920);
xor U11118 (N_11118,N_10875,N_10948);
nand U11119 (N_11119,N_10981,N_10947);
nand U11120 (N_11120,N_10972,N_10990);
xor U11121 (N_11121,N_10974,N_10895);
nor U11122 (N_11122,N_10985,N_10913);
and U11123 (N_11123,N_10973,N_10900);
or U11124 (N_11124,N_10982,N_10906);
nand U11125 (N_11125,N_11013,N_11026);
and U11126 (N_11126,N_11120,N_11101);
nand U11127 (N_11127,N_11090,N_11031);
nand U11128 (N_11128,N_11053,N_11054);
nor U11129 (N_11129,N_11070,N_11103);
or U11130 (N_11130,N_11020,N_11012);
xnor U11131 (N_11131,N_11046,N_11035);
or U11132 (N_11132,N_11063,N_11061);
or U11133 (N_11133,N_11094,N_11105);
nand U11134 (N_11134,N_11000,N_11009);
nand U11135 (N_11135,N_11047,N_11029);
and U11136 (N_11136,N_11079,N_11051);
and U11137 (N_11137,N_11119,N_11049);
nor U11138 (N_11138,N_11006,N_11030);
or U11139 (N_11139,N_11093,N_11092);
nor U11140 (N_11140,N_11066,N_11077);
xnor U11141 (N_11141,N_11060,N_11067);
nand U11142 (N_11142,N_11068,N_11059);
nor U11143 (N_11143,N_11018,N_11058);
nand U11144 (N_11144,N_11123,N_11087);
xnor U11145 (N_11145,N_11019,N_11042);
and U11146 (N_11146,N_11017,N_11008);
or U11147 (N_11147,N_11034,N_11078);
and U11148 (N_11148,N_11089,N_11082);
and U11149 (N_11149,N_11112,N_11091);
and U11150 (N_11150,N_11002,N_11003);
nor U11151 (N_11151,N_11039,N_11055);
nor U11152 (N_11152,N_11088,N_11022);
and U11153 (N_11153,N_11044,N_11001);
and U11154 (N_11154,N_11116,N_11015);
or U11155 (N_11155,N_11081,N_11076);
and U11156 (N_11156,N_11005,N_11118);
nor U11157 (N_11157,N_11121,N_11033);
nand U11158 (N_11158,N_11071,N_11106);
nand U11159 (N_11159,N_11043,N_11099);
nand U11160 (N_11160,N_11069,N_11027);
and U11161 (N_11161,N_11072,N_11038);
or U11162 (N_11162,N_11037,N_11062);
nor U11163 (N_11163,N_11102,N_11004);
xnor U11164 (N_11164,N_11036,N_11048);
nor U11165 (N_11165,N_11025,N_11023);
nor U11166 (N_11166,N_11056,N_11064);
and U11167 (N_11167,N_11028,N_11040);
nand U11168 (N_11168,N_11085,N_11016);
and U11169 (N_11169,N_11098,N_11114);
nor U11170 (N_11170,N_11075,N_11011);
nor U11171 (N_11171,N_11021,N_11124);
nand U11172 (N_11172,N_11050,N_11045);
nor U11173 (N_11173,N_11041,N_11122);
and U11174 (N_11174,N_11115,N_11111);
or U11175 (N_11175,N_11107,N_11065);
xor U11176 (N_11176,N_11014,N_11109);
nor U11177 (N_11177,N_11117,N_11032);
xor U11178 (N_11178,N_11086,N_11113);
xor U11179 (N_11179,N_11057,N_11110);
and U11180 (N_11180,N_11024,N_11108);
xor U11181 (N_11181,N_11073,N_11074);
nor U11182 (N_11182,N_11097,N_11080);
or U11183 (N_11183,N_11104,N_11052);
nand U11184 (N_11184,N_11083,N_11084);
xor U11185 (N_11185,N_11096,N_11010);
or U11186 (N_11186,N_11100,N_11007);
and U11187 (N_11187,N_11095,N_11101);
nor U11188 (N_11188,N_11108,N_11066);
nor U11189 (N_11189,N_11057,N_11031);
nor U11190 (N_11190,N_11124,N_11068);
nand U11191 (N_11191,N_11000,N_11031);
nor U11192 (N_11192,N_11011,N_11098);
or U11193 (N_11193,N_11017,N_11093);
nor U11194 (N_11194,N_11069,N_11084);
nor U11195 (N_11195,N_11064,N_11100);
and U11196 (N_11196,N_11113,N_11109);
and U11197 (N_11197,N_11121,N_11093);
xnor U11198 (N_11198,N_11057,N_11074);
nor U11199 (N_11199,N_11108,N_11117);
or U11200 (N_11200,N_11001,N_11037);
nand U11201 (N_11201,N_11021,N_11017);
or U11202 (N_11202,N_11043,N_11119);
nand U11203 (N_11203,N_11001,N_11041);
and U11204 (N_11204,N_11053,N_11077);
and U11205 (N_11205,N_11022,N_11029);
or U11206 (N_11206,N_11011,N_11095);
or U11207 (N_11207,N_11119,N_11079);
or U11208 (N_11208,N_11085,N_11012);
nand U11209 (N_11209,N_11068,N_11108);
and U11210 (N_11210,N_11062,N_11105);
or U11211 (N_11211,N_11084,N_11090);
nand U11212 (N_11212,N_11017,N_11025);
xnor U11213 (N_11213,N_11012,N_11069);
and U11214 (N_11214,N_11027,N_11007);
nor U11215 (N_11215,N_11010,N_11042);
nand U11216 (N_11216,N_11026,N_11039);
and U11217 (N_11217,N_11000,N_11044);
and U11218 (N_11218,N_11108,N_11032);
nand U11219 (N_11219,N_11022,N_11090);
xor U11220 (N_11220,N_11051,N_11124);
nand U11221 (N_11221,N_11024,N_11123);
or U11222 (N_11222,N_11021,N_11033);
or U11223 (N_11223,N_11123,N_11013);
nor U11224 (N_11224,N_11081,N_11114);
xnor U11225 (N_11225,N_11019,N_11076);
or U11226 (N_11226,N_11056,N_11086);
nand U11227 (N_11227,N_11117,N_11056);
and U11228 (N_11228,N_11043,N_11015);
nor U11229 (N_11229,N_11124,N_11083);
or U11230 (N_11230,N_11047,N_11107);
nor U11231 (N_11231,N_11021,N_11043);
or U11232 (N_11232,N_11118,N_11097);
nand U11233 (N_11233,N_11103,N_11068);
or U11234 (N_11234,N_11109,N_11006);
xnor U11235 (N_11235,N_11123,N_11100);
and U11236 (N_11236,N_11001,N_11110);
and U11237 (N_11237,N_11034,N_11059);
xor U11238 (N_11238,N_11074,N_11004);
and U11239 (N_11239,N_11099,N_11065);
and U11240 (N_11240,N_11074,N_11055);
or U11241 (N_11241,N_11103,N_11005);
nor U11242 (N_11242,N_11058,N_11106);
or U11243 (N_11243,N_11005,N_11008);
and U11244 (N_11244,N_11049,N_11001);
nor U11245 (N_11245,N_11054,N_11014);
or U11246 (N_11246,N_11093,N_11088);
and U11247 (N_11247,N_11109,N_11047);
nand U11248 (N_11248,N_11093,N_11041);
and U11249 (N_11249,N_11032,N_11087);
and U11250 (N_11250,N_11183,N_11174);
and U11251 (N_11251,N_11210,N_11162);
or U11252 (N_11252,N_11240,N_11129);
and U11253 (N_11253,N_11181,N_11152);
nand U11254 (N_11254,N_11226,N_11232);
or U11255 (N_11255,N_11182,N_11191);
nand U11256 (N_11256,N_11139,N_11206);
nand U11257 (N_11257,N_11216,N_11133);
and U11258 (N_11258,N_11211,N_11235);
or U11259 (N_11259,N_11153,N_11179);
nor U11260 (N_11260,N_11198,N_11178);
nor U11261 (N_11261,N_11195,N_11230);
and U11262 (N_11262,N_11202,N_11138);
nor U11263 (N_11263,N_11228,N_11249);
xor U11264 (N_11264,N_11194,N_11215);
or U11265 (N_11265,N_11187,N_11165);
or U11266 (N_11266,N_11164,N_11171);
nor U11267 (N_11267,N_11213,N_11192);
nor U11268 (N_11268,N_11144,N_11239);
or U11269 (N_11269,N_11220,N_11125);
or U11270 (N_11270,N_11203,N_11214);
or U11271 (N_11271,N_11247,N_11238);
nor U11272 (N_11272,N_11147,N_11177);
or U11273 (N_11273,N_11205,N_11222);
nand U11274 (N_11274,N_11224,N_11172);
nand U11275 (N_11275,N_11150,N_11180);
or U11276 (N_11276,N_11188,N_11126);
and U11277 (N_11277,N_11175,N_11176);
nand U11278 (N_11278,N_11169,N_11151);
or U11279 (N_11279,N_11209,N_11130);
and U11280 (N_11280,N_11199,N_11231);
and U11281 (N_11281,N_11170,N_11167);
nand U11282 (N_11282,N_11166,N_11248);
and U11283 (N_11283,N_11207,N_11156);
and U11284 (N_11284,N_11173,N_11223);
and U11285 (N_11285,N_11157,N_11160);
and U11286 (N_11286,N_11140,N_11189);
nor U11287 (N_11287,N_11149,N_11135);
or U11288 (N_11288,N_11168,N_11148);
xnor U11289 (N_11289,N_11145,N_11159);
xnor U11290 (N_11290,N_11142,N_11141);
or U11291 (N_11291,N_11217,N_11234);
and U11292 (N_11292,N_11212,N_11218);
or U11293 (N_11293,N_11163,N_11155);
nor U11294 (N_11294,N_11201,N_11184);
nand U11295 (N_11295,N_11244,N_11245);
or U11296 (N_11296,N_11134,N_11193);
and U11297 (N_11297,N_11208,N_11186);
nor U11298 (N_11298,N_11225,N_11219);
xnor U11299 (N_11299,N_11127,N_11154);
nor U11300 (N_11300,N_11146,N_11221);
xor U11301 (N_11301,N_11185,N_11229);
and U11302 (N_11302,N_11246,N_11241);
or U11303 (N_11303,N_11227,N_11243);
nand U11304 (N_11304,N_11143,N_11204);
nor U11305 (N_11305,N_11233,N_11196);
nor U11306 (N_11306,N_11161,N_11137);
and U11307 (N_11307,N_11158,N_11197);
nand U11308 (N_11308,N_11131,N_11136);
and U11309 (N_11309,N_11190,N_11128);
or U11310 (N_11310,N_11132,N_11200);
nand U11311 (N_11311,N_11237,N_11242);
or U11312 (N_11312,N_11236,N_11226);
nor U11313 (N_11313,N_11210,N_11228);
and U11314 (N_11314,N_11214,N_11134);
nor U11315 (N_11315,N_11246,N_11130);
nand U11316 (N_11316,N_11177,N_11231);
nor U11317 (N_11317,N_11153,N_11236);
nand U11318 (N_11318,N_11174,N_11220);
xnor U11319 (N_11319,N_11173,N_11146);
nand U11320 (N_11320,N_11249,N_11244);
and U11321 (N_11321,N_11129,N_11241);
xor U11322 (N_11322,N_11164,N_11150);
or U11323 (N_11323,N_11230,N_11219);
and U11324 (N_11324,N_11184,N_11157);
nand U11325 (N_11325,N_11242,N_11136);
nor U11326 (N_11326,N_11236,N_11210);
or U11327 (N_11327,N_11164,N_11228);
xor U11328 (N_11328,N_11136,N_11151);
or U11329 (N_11329,N_11171,N_11193);
and U11330 (N_11330,N_11184,N_11235);
nand U11331 (N_11331,N_11235,N_11164);
or U11332 (N_11332,N_11246,N_11240);
nor U11333 (N_11333,N_11200,N_11134);
nand U11334 (N_11334,N_11190,N_11185);
or U11335 (N_11335,N_11235,N_11156);
or U11336 (N_11336,N_11192,N_11235);
xnor U11337 (N_11337,N_11198,N_11230);
and U11338 (N_11338,N_11222,N_11231);
and U11339 (N_11339,N_11154,N_11138);
nor U11340 (N_11340,N_11181,N_11147);
nand U11341 (N_11341,N_11160,N_11191);
nand U11342 (N_11342,N_11192,N_11171);
and U11343 (N_11343,N_11198,N_11183);
and U11344 (N_11344,N_11216,N_11183);
nand U11345 (N_11345,N_11248,N_11187);
nand U11346 (N_11346,N_11139,N_11157);
nand U11347 (N_11347,N_11222,N_11217);
nand U11348 (N_11348,N_11226,N_11205);
nand U11349 (N_11349,N_11173,N_11152);
nor U11350 (N_11350,N_11226,N_11131);
or U11351 (N_11351,N_11152,N_11131);
xor U11352 (N_11352,N_11143,N_11164);
nand U11353 (N_11353,N_11132,N_11210);
nor U11354 (N_11354,N_11242,N_11129);
and U11355 (N_11355,N_11145,N_11188);
xor U11356 (N_11356,N_11175,N_11181);
nand U11357 (N_11357,N_11220,N_11221);
and U11358 (N_11358,N_11194,N_11133);
nand U11359 (N_11359,N_11177,N_11144);
or U11360 (N_11360,N_11144,N_11178);
nand U11361 (N_11361,N_11221,N_11169);
or U11362 (N_11362,N_11148,N_11130);
or U11363 (N_11363,N_11161,N_11201);
nor U11364 (N_11364,N_11138,N_11200);
and U11365 (N_11365,N_11184,N_11176);
nand U11366 (N_11366,N_11168,N_11130);
nor U11367 (N_11367,N_11180,N_11220);
and U11368 (N_11368,N_11139,N_11165);
nand U11369 (N_11369,N_11196,N_11169);
and U11370 (N_11370,N_11244,N_11131);
and U11371 (N_11371,N_11157,N_11207);
or U11372 (N_11372,N_11146,N_11132);
xor U11373 (N_11373,N_11184,N_11205);
nor U11374 (N_11374,N_11223,N_11126);
or U11375 (N_11375,N_11307,N_11350);
nor U11376 (N_11376,N_11330,N_11265);
and U11377 (N_11377,N_11341,N_11275);
or U11378 (N_11378,N_11348,N_11313);
or U11379 (N_11379,N_11329,N_11273);
nor U11380 (N_11380,N_11328,N_11262);
nor U11381 (N_11381,N_11346,N_11349);
and U11382 (N_11382,N_11356,N_11304);
and U11383 (N_11383,N_11272,N_11312);
and U11384 (N_11384,N_11267,N_11368);
nand U11385 (N_11385,N_11343,N_11309);
nand U11386 (N_11386,N_11296,N_11334);
and U11387 (N_11387,N_11289,N_11354);
nand U11388 (N_11388,N_11365,N_11351);
or U11389 (N_11389,N_11308,N_11323);
nor U11390 (N_11390,N_11285,N_11250);
nor U11391 (N_11391,N_11251,N_11276);
xor U11392 (N_11392,N_11255,N_11305);
or U11393 (N_11393,N_11266,N_11352);
nand U11394 (N_11394,N_11331,N_11299);
nor U11395 (N_11395,N_11288,N_11342);
nand U11396 (N_11396,N_11319,N_11291);
or U11397 (N_11397,N_11298,N_11340);
or U11398 (N_11398,N_11306,N_11283);
and U11399 (N_11399,N_11336,N_11301);
nor U11400 (N_11400,N_11269,N_11254);
nand U11401 (N_11401,N_11360,N_11315);
or U11402 (N_11402,N_11324,N_11322);
nor U11403 (N_11403,N_11345,N_11370);
and U11404 (N_11404,N_11292,N_11253);
or U11405 (N_11405,N_11290,N_11282);
xnor U11406 (N_11406,N_11261,N_11325);
nand U11407 (N_11407,N_11357,N_11277);
and U11408 (N_11408,N_11372,N_11311);
nor U11409 (N_11409,N_11271,N_11338);
and U11410 (N_11410,N_11326,N_11344);
nor U11411 (N_11411,N_11362,N_11317);
or U11412 (N_11412,N_11264,N_11327);
nor U11413 (N_11413,N_11318,N_11335);
or U11414 (N_11414,N_11355,N_11310);
or U11415 (N_11415,N_11337,N_11314);
and U11416 (N_11416,N_11302,N_11286);
nand U11417 (N_11417,N_11258,N_11366);
or U11418 (N_11418,N_11371,N_11297);
or U11419 (N_11419,N_11364,N_11293);
nor U11420 (N_11420,N_11295,N_11270);
nor U11421 (N_11421,N_11316,N_11361);
or U11422 (N_11422,N_11287,N_11279);
nor U11423 (N_11423,N_11367,N_11280);
or U11424 (N_11424,N_11263,N_11358);
nor U11425 (N_11425,N_11347,N_11256);
nor U11426 (N_11426,N_11281,N_11294);
nor U11427 (N_11427,N_11257,N_11284);
and U11428 (N_11428,N_11369,N_11374);
and U11429 (N_11429,N_11303,N_11259);
and U11430 (N_11430,N_11373,N_11278);
and U11431 (N_11431,N_11363,N_11274);
nor U11432 (N_11432,N_11300,N_11268);
nor U11433 (N_11433,N_11320,N_11333);
or U11434 (N_11434,N_11359,N_11332);
and U11435 (N_11435,N_11321,N_11339);
or U11436 (N_11436,N_11252,N_11353);
nand U11437 (N_11437,N_11260,N_11311);
and U11438 (N_11438,N_11367,N_11357);
and U11439 (N_11439,N_11330,N_11264);
nand U11440 (N_11440,N_11344,N_11327);
and U11441 (N_11441,N_11295,N_11293);
or U11442 (N_11442,N_11364,N_11353);
and U11443 (N_11443,N_11323,N_11312);
nor U11444 (N_11444,N_11358,N_11267);
or U11445 (N_11445,N_11276,N_11278);
or U11446 (N_11446,N_11291,N_11253);
or U11447 (N_11447,N_11338,N_11266);
and U11448 (N_11448,N_11281,N_11288);
or U11449 (N_11449,N_11294,N_11254);
or U11450 (N_11450,N_11336,N_11293);
or U11451 (N_11451,N_11329,N_11270);
and U11452 (N_11452,N_11316,N_11282);
xnor U11453 (N_11453,N_11349,N_11265);
nor U11454 (N_11454,N_11292,N_11373);
and U11455 (N_11455,N_11263,N_11344);
and U11456 (N_11456,N_11251,N_11303);
and U11457 (N_11457,N_11294,N_11264);
and U11458 (N_11458,N_11312,N_11319);
nor U11459 (N_11459,N_11279,N_11344);
nor U11460 (N_11460,N_11328,N_11285);
nor U11461 (N_11461,N_11257,N_11320);
nor U11462 (N_11462,N_11342,N_11319);
and U11463 (N_11463,N_11284,N_11368);
nor U11464 (N_11464,N_11282,N_11338);
or U11465 (N_11465,N_11313,N_11285);
nor U11466 (N_11466,N_11283,N_11295);
and U11467 (N_11467,N_11285,N_11372);
nand U11468 (N_11468,N_11353,N_11322);
nor U11469 (N_11469,N_11285,N_11257);
and U11470 (N_11470,N_11323,N_11256);
and U11471 (N_11471,N_11293,N_11289);
and U11472 (N_11472,N_11372,N_11336);
nor U11473 (N_11473,N_11328,N_11352);
nor U11474 (N_11474,N_11275,N_11340);
nor U11475 (N_11475,N_11323,N_11368);
nand U11476 (N_11476,N_11283,N_11360);
nand U11477 (N_11477,N_11276,N_11362);
xnor U11478 (N_11478,N_11273,N_11314);
and U11479 (N_11479,N_11290,N_11291);
and U11480 (N_11480,N_11260,N_11358);
and U11481 (N_11481,N_11343,N_11278);
nand U11482 (N_11482,N_11290,N_11364);
and U11483 (N_11483,N_11274,N_11289);
nor U11484 (N_11484,N_11329,N_11292);
xor U11485 (N_11485,N_11327,N_11306);
nor U11486 (N_11486,N_11356,N_11300);
xnor U11487 (N_11487,N_11281,N_11372);
nand U11488 (N_11488,N_11250,N_11267);
nor U11489 (N_11489,N_11286,N_11346);
or U11490 (N_11490,N_11300,N_11342);
nor U11491 (N_11491,N_11257,N_11331);
or U11492 (N_11492,N_11256,N_11320);
xnor U11493 (N_11493,N_11332,N_11274);
nand U11494 (N_11494,N_11255,N_11362);
nor U11495 (N_11495,N_11363,N_11267);
nand U11496 (N_11496,N_11271,N_11367);
nor U11497 (N_11497,N_11253,N_11339);
and U11498 (N_11498,N_11369,N_11326);
nor U11499 (N_11499,N_11357,N_11341);
or U11500 (N_11500,N_11441,N_11393);
nor U11501 (N_11501,N_11426,N_11478);
and U11502 (N_11502,N_11488,N_11483);
nor U11503 (N_11503,N_11388,N_11400);
xnor U11504 (N_11504,N_11406,N_11474);
and U11505 (N_11505,N_11435,N_11427);
nor U11506 (N_11506,N_11377,N_11477);
or U11507 (N_11507,N_11476,N_11376);
nor U11508 (N_11508,N_11461,N_11450);
nor U11509 (N_11509,N_11385,N_11496);
xor U11510 (N_11510,N_11495,N_11492);
and U11511 (N_11511,N_11459,N_11463);
and U11512 (N_11512,N_11472,N_11456);
or U11513 (N_11513,N_11432,N_11468);
nor U11514 (N_11514,N_11402,N_11454);
and U11515 (N_11515,N_11487,N_11493);
nor U11516 (N_11516,N_11405,N_11413);
xnor U11517 (N_11517,N_11378,N_11455);
and U11518 (N_11518,N_11437,N_11382);
nand U11519 (N_11519,N_11448,N_11384);
xor U11520 (N_11520,N_11375,N_11479);
and U11521 (N_11521,N_11480,N_11423);
nor U11522 (N_11522,N_11458,N_11482);
or U11523 (N_11523,N_11439,N_11445);
nor U11524 (N_11524,N_11491,N_11412);
or U11525 (N_11525,N_11396,N_11490);
or U11526 (N_11526,N_11415,N_11418);
nand U11527 (N_11527,N_11414,N_11484);
nor U11528 (N_11528,N_11410,N_11436);
nand U11529 (N_11529,N_11386,N_11430);
and U11530 (N_11530,N_11409,N_11449);
and U11531 (N_11531,N_11420,N_11411);
or U11532 (N_11532,N_11447,N_11391);
and U11533 (N_11533,N_11422,N_11408);
or U11534 (N_11534,N_11387,N_11471);
xor U11535 (N_11535,N_11417,N_11407);
or U11536 (N_11536,N_11380,N_11404);
and U11537 (N_11537,N_11416,N_11440);
nand U11538 (N_11538,N_11444,N_11453);
and U11539 (N_11539,N_11419,N_11475);
or U11540 (N_11540,N_11381,N_11433);
nand U11541 (N_11541,N_11379,N_11442);
nor U11542 (N_11542,N_11431,N_11438);
or U11543 (N_11543,N_11428,N_11486);
and U11544 (N_11544,N_11434,N_11394);
nand U11545 (N_11545,N_11429,N_11443);
or U11546 (N_11546,N_11481,N_11470);
nor U11547 (N_11547,N_11494,N_11457);
nand U11548 (N_11548,N_11424,N_11467);
xnor U11549 (N_11549,N_11460,N_11465);
nand U11550 (N_11550,N_11469,N_11398);
nor U11551 (N_11551,N_11399,N_11403);
xnor U11552 (N_11552,N_11473,N_11446);
and U11553 (N_11553,N_11395,N_11392);
or U11554 (N_11554,N_11421,N_11425);
and U11555 (N_11555,N_11466,N_11401);
and U11556 (N_11556,N_11498,N_11452);
nand U11557 (N_11557,N_11397,N_11497);
nor U11558 (N_11558,N_11485,N_11383);
or U11559 (N_11559,N_11451,N_11462);
or U11560 (N_11560,N_11489,N_11464);
xor U11561 (N_11561,N_11390,N_11499);
xnor U11562 (N_11562,N_11389,N_11469);
nand U11563 (N_11563,N_11414,N_11427);
and U11564 (N_11564,N_11393,N_11410);
nor U11565 (N_11565,N_11476,N_11484);
or U11566 (N_11566,N_11477,N_11446);
nor U11567 (N_11567,N_11499,N_11461);
nand U11568 (N_11568,N_11431,N_11376);
nor U11569 (N_11569,N_11379,N_11396);
xnor U11570 (N_11570,N_11377,N_11412);
nand U11571 (N_11571,N_11452,N_11467);
nor U11572 (N_11572,N_11404,N_11417);
nor U11573 (N_11573,N_11428,N_11409);
nor U11574 (N_11574,N_11433,N_11457);
or U11575 (N_11575,N_11478,N_11401);
or U11576 (N_11576,N_11493,N_11409);
nand U11577 (N_11577,N_11468,N_11423);
xor U11578 (N_11578,N_11375,N_11389);
and U11579 (N_11579,N_11473,N_11448);
and U11580 (N_11580,N_11450,N_11453);
xnor U11581 (N_11581,N_11441,N_11389);
nand U11582 (N_11582,N_11403,N_11458);
xor U11583 (N_11583,N_11475,N_11444);
or U11584 (N_11584,N_11410,N_11456);
or U11585 (N_11585,N_11451,N_11413);
and U11586 (N_11586,N_11488,N_11473);
and U11587 (N_11587,N_11462,N_11463);
or U11588 (N_11588,N_11485,N_11411);
and U11589 (N_11589,N_11391,N_11426);
and U11590 (N_11590,N_11485,N_11418);
nor U11591 (N_11591,N_11416,N_11470);
xnor U11592 (N_11592,N_11402,N_11469);
nand U11593 (N_11593,N_11460,N_11488);
and U11594 (N_11594,N_11404,N_11436);
xor U11595 (N_11595,N_11427,N_11379);
nor U11596 (N_11596,N_11466,N_11480);
nor U11597 (N_11597,N_11389,N_11450);
nand U11598 (N_11598,N_11451,N_11419);
nand U11599 (N_11599,N_11469,N_11425);
nor U11600 (N_11600,N_11491,N_11437);
nand U11601 (N_11601,N_11381,N_11431);
or U11602 (N_11602,N_11417,N_11446);
or U11603 (N_11603,N_11390,N_11483);
nor U11604 (N_11604,N_11411,N_11397);
nand U11605 (N_11605,N_11430,N_11465);
or U11606 (N_11606,N_11426,N_11456);
nand U11607 (N_11607,N_11465,N_11411);
or U11608 (N_11608,N_11445,N_11449);
nand U11609 (N_11609,N_11419,N_11462);
xor U11610 (N_11610,N_11498,N_11474);
or U11611 (N_11611,N_11450,N_11485);
nand U11612 (N_11612,N_11388,N_11463);
and U11613 (N_11613,N_11391,N_11381);
nor U11614 (N_11614,N_11455,N_11416);
nor U11615 (N_11615,N_11441,N_11450);
nand U11616 (N_11616,N_11476,N_11427);
nand U11617 (N_11617,N_11470,N_11401);
nor U11618 (N_11618,N_11416,N_11376);
and U11619 (N_11619,N_11465,N_11392);
nand U11620 (N_11620,N_11401,N_11495);
nand U11621 (N_11621,N_11388,N_11403);
nand U11622 (N_11622,N_11469,N_11480);
and U11623 (N_11623,N_11450,N_11381);
nor U11624 (N_11624,N_11409,N_11489);
or U11625 (N_11625,N_11623,N_11591);
xor U11626 (N_11626,N_11570,N_11620);
xor U11627 (N_11627,N_11535,N_11606);
nand U11628 (N_11628,N_11546,N_11515);
nand U11629 (N_11629,N_11588,N_11552);
and U11630 (N_11630,N_11581,N_11509);
nand U11631 (N_11631,N_11560,N_11564);
nand U11632 (N_11632,N_11542,N_11503);
and U11633 (N_11633,N_11558,N_11506);
and U11634 (N_11634,N_11602,N_11579);
and U11635 (N_11635,N_11599,N_11565);
or U11636 (N_11636,N_11583,N_11527);
xnor U11637 (N_11637,N_11607,N_11510);
nor U11638 (N_11638,N_11541,N_11621);
nor U11639 (N_11639,N_11594,N_11593);
or U11640 (N_11640,N_11538,N_11573);
nand U11641 (N_11641,N_11531,N_11590);
nor U11642 (N_11642,N_11596,N_11556);
or U11643 (N_11643,N_11574,N_11504);
xor U11644 (N_11644,N_11547,N_11601);
or U11645 (N_11645,N_11605,N_11608);
or U11646 (N_11646,N_11572,N_11536);
nand U11647 (N_11647,N_11603,N_11550);
nor U11648 (N_11648,N_11568,N_11569);
xnor U11649 (N_11649,N_11537,N_11559);
xnor U11650 (N_11650,N_11511,N_11554);
or U11651 (N_11651,N_11539,N_11571);
or U11652 (N_11652,N_11600,N_11530);
nor U11653 (N_11653,N_11529,N_11614);
or U11654 (N_11654,N_11540,N_11501);
or U11655 (N_11655,N_11533,N_11580);
nand U11656 (N_11656,N_11544,N_11520);
nor U11657 (N_11657,N_11616,N_11589);
nand U11658 (N_11658,N_11584,N_11523);
nand U11659 (N_11659,N_11609,N_11519);
nor U11660 (N_11660,N_11563,N_11545);
nand U11661 (N_11661,N_11577,N_11543);
nand U11662 (N_11662,N_11582,N_11553);
or U11663 (N_11663,N_11517,N_11551);
and U11664 (N_11664,N_11549,N_11528);
nor U11665 (N_11665,N_11557,N_11514);
nand U11666 (N_11666,N_11562,N_11567);
or U11667 (N_11667,N_11587,N_11522);
nand U11668 (N_11668,N_11622,N_11507);
nand U11669 (N_11669,N_11598,N_11513);
nor U11670 (N_11670,N_11586,N_11595);
or U11671 (N_11671,N_11585,N_11526);
nor U11672 (N_11672,N_11561,N_11613);
and U11673 (N_11673,N_11512,N_11576);
nand U11674 (N_11674,N_11604,N_11617);
nor U11675 (N_11675,N_11500,N_11612);
xnor U11676 (N_11676,N_11516,N_11597);
nand U11677 (N_11677,N_11534,N_11508);
nor U11678 (N_11678,N_11555,N_11532);
nand U11679 (N_11679,N_11524,N_11525);
or U11680 (N_11680,N_11624,N_11615);
xnor U11681 (N_11681,N_11502,N_11610);
nand U11682 (N_11682,N_11578,N_11518);
or U11683 (N_11683,N_11521,N_11548);
nor U11684 (N_11684,N_11566,N_11618);
and U11685 (N_11685,N_11575,N_11611);
and U11686 (N_11686,N_11505,N_11619);
nor U11687 (N_11687,N_11592,N_11520);
or U11688 (N_11688,N_11568,N_11540);
nand U11689 (N_11689,N_11609,N_11525);
nand U11690 (N_11690,N_11619,N_11568);
and U11691 (N_11691,N_11547,N_11595);
xnor U11692 (N_11692,N_11608,N_11557);
nor U11693 (N_11693,N_11616,N_11547);
and U11694 (N_11694,N_11521,N_11534);
nand U11695 (N_11695,N_11519,N_11583);
or U11696 (N_11696,N_11618,N_11536);
or U11697 (N_11697,N_11620,N_11621);
nor U11698 (N_11698,N_11533,N_11510);
nor U11699 (N_11699,N_11503,N_11618);
xor U11700 (N_11700,N_11538,N_11623);
and U11701 (N_11701,N_11549,N_11599);
and U11702 (N_11702,N_11590,N_11521);
xor U11703 (N_11703,N_11613,N_11507);
and U11704 (N_11704,N_11500,N_11512);
nor U11705 (N_11705,N_11602,N_11505);
or U11706 (N_11706,N_11602,N_11614);
or U11707 (N_11707,N_11534,N_11591);
nor U11708 (N_11708,N_11584,N_11598);
nand U11709 (N_11709,N_11601,N_11570);
nor U11710 (N_11710,N_11552,N_11600);
nand U11711 (N_11711,N_11610,N_11519);
nor U11712 (N_11712,N_11518,N_11540);
and U11713 (N_11713,N_11564,N_11582);
xor U11714 (N_11714,N_11502,N_11579);
or U11715 (N_11715,N_11513,N_11602);
nand U11716 (N_11716,N_11518,N_11507);
or U11717 (N_11717,N_11525,N_11500);
nand U11718 (N_11718,N_11515,N_11614);
and U11719 (N_11719,N_11514,N_11512);
or U11720 (N_11720,N_11608,N_11537);
and U11721 (N_11721,N_11599,N_11526);
and U11722 (N_11722,N_11529,N_11540);
and U11723 (N_11723,N_11535,N_11619);
and U11724 (N_11724,N_11594,N_11565);
and U11725 (N_11725,N_11551,N_11526);
nor U11726 (N_11726,N_11623,N_11506);
or U11727 (N_11727,N_11517,N_11561);
nand U11728 (N_11728,N_11620,N_11550);
and U11729 (N_11729,N_11576,N_11500);
and U11730 (N_11730,N_11540,N_11602);
and U11731 (N_11731,N_11604,N_11522);
nand U11732 (N_11732,N_11524,N_11547);
or U11733 (N_11733,N_11560,N_11524);
and U11734 (N_11734,N_11554,N_11559);
and U11735 (N_11735,N_11574,N_11538);
or U11736 (N_11736,N_11619,N_11538);
and U11737 (N_11737,N_11573,N_11519);
xor U11738 (N_11738,N_11607,N_11571);
nor U11739 (N_11739,N_11534,N_11601);
nor U11740 (N_11740,N_11621,N_11572);
xnor U11741 (N_11741,N_11530,N_11544);
or U11742 (N_11742,N_11603,N_11618);
nand U11743 (N_11743,N_11523,N_11612);
nand U11744 (N_11744,N_11597,N_11514);
and U11745 (N_11745,N_11541,N_11576);
nand U11746 (N_11746,N_11623,N_11556);
nor U11747 (N_11747,N_11591,N_11547);
nand U11748 (N_11748,N_11526,N_11591);
or U11749 (N_11749,N_11588,N_11621);
nand U11750 (N_11750,N_11633,N_11717);
nand U11751 (N_11751,N_11709,N_11658);
or U11752 (N_11752,N_11646,N_11742);
nand U11753 (N_11753,N_11643,N_11644);
nand U11754 (N_11754,N_11728,N_11712);
nor U11755 (N_11755,N_11698,N_11677);
and U11756 (N_11756,N_11744,N_11674);
or U11757 (N_11757,N_11720,N_11669);
nor U11758 (N_11758,N_11727,N_11738);
nand U11759 (N_11759,N_11707,N_11635);
nand U11760 (N_11760,N_11630,N_11697);
or U11761 (N_11761,N_11684,N_11650);
and U11762 (N_11762,N_11631,N_11637);
nor U11763 (N_11763,N_11719,N_11670);
or U11764 (N_11764,N_11691,N_11743);
and U11765 (N_11765,N_11652,N_11722);
and U11766 (N_11766,N_11649,N_11626);
and U11767 (N_11767,N_11628,N_11714);
or U11768 (N_11768,N_11662,N_11676);
nor U11769 (N_11769,N_11745,N_11664);
and U11770 (N_11770,N_11700,N_11640);
and U11771 (N_11771,N_11681,N_11715);
or U11772 (N_11772,N_11659,N_11716);
nor U11773 (N_11773,N_11696,N_11747);
and U11774 (N_11774,N_11648,N_11735);
nor U11775 (N_11775,N_11656,N_11686);
xor U11776 (N_11776,N_11653,N_11704);
nand U11777 (N_11777,N_11737,N_11671);
nand U11778 (N_11778,N_11729,N_11663);
nand U11779 (N_11779,N_11636,N_11741);
nand U11780 (N_11780,N_11642,N_11645);
and U11781 (N_11781,N_11693,N_11748);
or U11782 (N_11782,N_11634,N_11713);
and U11783 (N_11783,N_11705,N_11695);
nor U11784 (N_11784,N_11710,N_11721);
nand U11785 (N_11785,N_11655,N_11673);
or U11786 (N_11786,N_11657,N_11647);
nor U11787 (N_11787,N_11725,N_11660);
nor U11788 (N_11788,N_11724,N_11672);
nand U11789 (N_11789,N_11732,N_11638);
nand U11790 (N_11790,N_11665,N_11723);
nand U11791 (N_11791,N_11685,N_11701);
and U11792 (N_11792,N_11739,N_11678);
nor U11793 (N_11793,N_11702,N_11651);
and U11794 (N_11794,N_11688,N_11682);
and U11795 (N_11795,N_11749,N_11746);
nand U11796 (N_11796,N_11703,N_11692);
xor U11797 (N_11797,N_11641,N_11711);
nor U11798 (N_11798,N_11675,N_11632);
and U11799 (N_11799,N_11683,N_11679);
and U11800 (N_11800,N_11680,N_11687);
or U11801 (N_11801,N_11730,N_11668);
xnor U11802 (N_11802,N_11654,N_11706);
xor U11803 (N_11803,N_11718,N_11625);
nor U11804 (N_11804,N_11734,N_11666);
or U11805 (N_11805,N_11667,N_11708);
nor U11806 (N_11806,N_11661,N_11627);
or U11807 (N_11807,N_11733,N_11726);
xnor U11808 (N_11808,N_11689,N_11740);
nand U11809 (N_11809,N_11699,N_11731);
and U11810 (N_11810,N_11629,N_11639);
nand U11811 (N_11811,N_11736,N_11694);
nand U11812 (N_11812,N_11690,N_11727);
nor U11813 (N_11813,N_11631,N_11673);
xnor U11814 (N_11814,N_11686,N_11709);
xor U11815 (N_11815,N_11673,N_11684);
nor U11816 (N_11816,N_11684,N_11706);
nor U11817 (N_11817,N_11672,N_11704);
nand U11818 (N_11818,N_11691,N_11687);
nor U11819 (N_11819,N_11710,N_11643);
nand U11820 (N_11820,N_11668,N_11733);
nand U11821 (N_11821,N_11674,N_11676);
and U11822 (N_11822,N_11668,N_11746);
and U11823 (N_11823,N_11684,N_11724);
and U11824 (N_11824,N_11711,N_11650);
or U11825 (N_11825,N_11677,N_11627);
nand U11826 (N_11826,N_11749,N_11641);
or U11827 (N_11827,N_11670,N_11686);
nor U11828 (N_11828,N_11652,N_11654);
nor U11829 (N_11829,N_11703,N_11629);
and U11830 (N_11830,N_11723,N_11679);
or U11831 (N_11831,N_11650,N_11661);
and U11832 (N_11832,N_11631,N_11748);
nand U11833 (N_11833,N_11717,N_11714);
nor U11834 (N_11834,N_11743,N_11670);
or U11835 (N_11835,N_11661,N_11707);
or U11836 (N_11836,N_11633,N_11628);
or U11837 (N_11837,N_11652,N_11695);
or U11838 (N_11838,N_11671,N_11633);
nand U11839 (N_11839,N_11747,N_11658);
nor U11840 (N_11840,N_11711,N_11748);
nor U11841 (N_11841,N_11635,N_11633);
nor U11842 (N_11842,N_11640,N_11627);
or U11843 (N_11843,N_11747,N_11713);
and U11844 (N_11844,N_11714,N_11733);
nand U11845 (N_11845,N_11746,N_11700);
nor U11846 (N_11846,N_11648,N_11654);
nor U11847 (N_11847,N_11719,N_11626);
nand U11848 (N_11848,N_11654,N_11736);
nor U11849 (N_11849,N_11645,N_11716);
nand U11850 (N_11850,N_11692,N_11683);
and U11851 (N_11851,N_11659,N_11731);
and U11852 (N_11852,N_11674,N_11694);
xnor U11853 (N_11853,N_11729,N_11713);
and U11854 (N_11854,N_11747,N_11635);
xor U11855 (N_11855,N_11691,N_11700);
or U11856 (N_11856,N_11747,N_11677);
nor U11857 (N_11857,N_11695,N_11665);
and U11858 (N_11858,N_11748,N_11699);
nor U11859 (N_11859,N_11642,N_11707);
nand U11860 (N_11860,N_11730,N_11695);
or U11861 (N_11861,N_11718,N_11719);
nor U11862 (N_11862,N_11694,N_11633);
and U11863 (N_11863,N_11637,N_11687);
nand U11864 (N_11864,N_11683,N_11639);
and U11865 (N_11865,N_11711,N_11642);
nand U11866 (N_11866,N_11733,N_11627);
nor U11867 (N_11867,N_11749,N_11662);
nor U11868 (N_11868,N_11666,N_11745);
nor U11869 (N_11869,N_11679,N_11625);
or U11870 (N_11870,N_11703,N_11644);
and U11871 (N_11871,N_11667,N_11668);
nand U11872 (N_11872,N_11700,N_11631);
nor U11873 (N_11873,N_11634,N_11627);
nand U11874 (N_11874,N_11684,N_11654);
and U11875 (N_11875,N_11756,N_11852);
nand U11876 (N_11876,N_11796,N_11781);
and U11877 (N_11877,N_11859,N_11855);
or U11878 (N_11878,N_11785,N_11820);
or U11879 (N_11879,N_11846,N_11798);
nand U11880 (N_11880,N_11829,N_11828);
nor U11881 (N_11881,N_11772,N_11821);
xor U11882 (N_11882,N_11816,N_11815);
and U11883 (N_11883,N_11766,N_11865);
nor U11884 (N_11884,N_11843,N_11770);
nand U11885 (N_11885,N_11805,N_11804);
and U11886 (N_11886,N_11838,N_11834);
nor U11887 (N_11887,N_11755,N_11773);
or U11888 (N_11888,N_11873,N_11863);
nor U11889 (N_11889,N_11810,N_11813);
xnor U11890 (N_11890,N_11845,N_11836);
and U11891 (N_11891,N_11868,N_11819);
nand U11892 (N_11892,N_11854,N_11814);
nor U11893 (N_11893,N_11817,N_11860);
nor U11894 (N_11894,N_11753,N_11870);
xnor U11895 (N_11895,N_11786,N_11835);
nand U11896 (N_11896,N_11752,N_11856);
nand U11897 (N_11897,N_11808,N_11827);
nor U11898 (N_11898,N_11837,N_11787);
nand U11899 (N_11899,N_11750,N_11830);
and U11900 (N_11900,N_11761,N_11826);
or U11901 (N_11901,N_11763,N_11867);
nand U11902 (N_11902,N_11809,N_11825);
and U11903 (N_11903,N_11754,N_11800);
nand U11904 (N_11904,N_11822,N_11840);
nor U11905 (N_11905,N_11769,N_11789);
and U11906 (N_11906,N_11765,N_11775);
and U11907 (N_11907,N_11782,N_11801);
xnor U11908 (N_11908,N_11759,N_11818);
nor U11909 (N_11909,N_11803,N_11866);
nor U11910 (N_11910,N_11788,N_11832);
or U11911 (N_11911,N_11774,N_11812);
and U11912 (N_11912,N_11794,N_11771);
and U11913 (N_11913,N_11760,N_11851);
nand U11914 (N_11914,N_11793,N_11831);
nand U11915 (N_11915,N_11777,N_11833);
and U11916 (N_11916,N_11807,N_11849);
and U11917 (N_11917,N_11758,N_11762);
nor U11918 (N_11918,N_11874,N_11792);
or U11919 (N_11919,N_11767,N_11857);
and U11920 (N_11920,N_11848,N_11776);
or U11921 (N_11921,N_11797,N_11757);
nor U11922 (N_11922,N_11872,N_11799);
and U11923 (N_11923,N_11802,N_11751);
nand U11924 (N_11924,N_11780,N_11847);
or U11925 (N_11925,N_11823,N_11824);
nor U11926 (N_11926,N_11861,N_11764);
nand U11927 (N_11927,N_11783,N_11784);
xnor U11928 (N_11928,N_11842,N_11778);
nor U11929 (N_11929,N_11791,N_11858);
nand U11930 (N_11930,N_11779,N_11864);
nor U11931 (N_11931,N_11795,N_11844);
or U11932 (N_11932,N_11850,N_11862);
or U11933 (N_11933,N_11806,N_11869);
and U11934 (N_11934,N_11839,N_11871);
nand U11935 (N_11935,N_11841,N_11811);
or U11936 (N_11936,N_11853,N_11790);
and U11937 (N_11937,N_11768,N_11764);
and U11938 (N_11938,N_11779,N_11832);
or U11939 (N_11939,N_11854,N_11758);
xor U11940 (N_11940,N_11855,N_11856);
or U11941 (N_11941,N_11806,N_11829);
nor U11942 (N_11942,N_11811,N_11821);
xor U11943 (N_11943,N_11837,N_11805);
and U11944 (N_11944,N_11833,N_11836);
nand U11945 (N_11945,N_11790,N_11874);
nand U11946 (N_11946,N_11845,N_11868);
or U11947 (N_11947,N_11763,N_11794);
xor U11948 (N_11948,N_11781,N_11816);
xor U11949 (N_11949,N_11861,N_11806);
and U11950 (N_11950,N_11859,N_11751);
and U11951 (N_11951,N_11811,N_11772);
xor U11952 (N_11952,N_11848,N_11835);
or U11953 (N_11953,N_11816,N_11801);
nor U11954 (N_11954,N_11870,N_11817);
nand U11955 (N_11955,N_11797,N_11753);
nor U11956 (N_11956,N_11819,N_11801);
and U11957 (N_11957,N_11813,N_11773);
and U11958 (N_11958,N_11792,N_11830);
xor U11959 (N_11959,N_11801,N_11788);
nand U11960 (N_11960,N_11859,N_11806);
nor U11961 (N_11961,N_11751,N_11843);
and U11962 (N_11962,N_11750,N_11777);
or U11963 (N_11963,N_11759,N_11839);
nand U11964 (N_11964,N_11830,N_11873);
nor U11965 (N_11965,N_11858,N_11802);
and U11966 (N_11966,N_11856,N_11861);
nand U11967 (N_11967,N_11763,N_11872);
xor U11968 (N_11968,N_11829,N_11765);
xnor U11969 (N_11969,N_11839,N_11765);
and U11970 (N_11970,N_11821,N_11765);
and U11971 (N_11971,N_11789,N_11816);
nor U11972 (N_11972,N_11842,N_11804);
nand U11973 (N_11973,N_11853,N_11846);
or U11974 (N_11974,N_11829,N_11752);
and U11975 (N_11975,N_11809,N_11773);
and U11976 (N_11976,N_11821,N_11762);
xor U11977 (N_11977,N_11759,N_11762);
and U11978 (N_11978,N_11859,N_11773);
nand U11979 (N_11979,N_11785,N_11765);
and U11980 (N_11980,N_11836,N_11843);
nor U11981 (N_11981,N_11846,N_11815);
nor U11982 (N_11982,N_11791,N_11788);
nand U11983 (N_11983,N_11780,N_11778);
or U11984 (N_11984,N_11838,N_11858);
nor U11985 (N_11985,N_11794,N_11864);
nand U11986 (N_11986,N_11785,N_11758);
nand U11987 (N_11987,N_11828,N_11783);
or U11988 (N_11988,N_11780,N_11851);
or U11989 (N_11989,N_11805,N_11771);
nor U11990 (N_11990,N_11780,N_11754);
nand U11991 (N_11991,N_11834,N_11808);
and U11992 (N_11992,N_11858,N_11831);
nand U11993 (N_11993,N_11802,N_11769);
nand U11994 (N_11994,N_11834,N_11846);
and U11995 (N_11995,N_11872,N_11855);
nor U11996 (N_11996,N_11769,N_11871);
and U11997 (N_11997,N_11812,N_11849);
or U11998 (N_11998,N_11757,N_11753);
xnor U11999 (N_11999,N_11842,N_11850);
nor U12000 (N_12000,N_11991,N_11969);
nor U12001 (N_12001,N_11979,N_11896);
and U12002 (N_12002,N_11974,N_11955);
and U12003 (N_12003,N_11928,N_11883);
nor U12004 (N_12004,N_11993,N_11886);
nor U12005 (N_12005,N_11909,N_11983);
and U12006 (N_12006,N_11953,N_11878);
or U12007 (N_12007,N_11908,N_11984);
xor U12008 (N_12008,N_11950,N_11893);
and U12009 (N_12009,N_11990,N_11949);
and U12010 (N_12010,N_11923,N_11916);
nand U12011 (N_12011,N_11876,N_11946);
nor U12012 (N_12012,N_11941,N_11880);
and U12013 (N_12013,N_11890,N_11943);
xnor U12014 (N_12014,N_11898,N_11910);
nor U12015 (N_12015,N_11989,N_11912);
nor U12016 (N_12016,N_11954,N_11970);
xor U12017 (N_12017,N_11963,N_11988);
nand U12018 (N_12018,N_11975,N_11951);
nand U12019 (N_12019,N_11957,N_11921);
and U12020 (N_12020,N_11967,N_11927);
nor U12021 (N_12021,N_11884,N_11906);
or U12022 (N_12022,N_11971,N_11892);
nor U12023 (N_12023,N_11877,N_11997);
nand U12024 (N_12024,N_11960,N_11897);
nand U12025 (N_12025,N_11885,N_11964);
xor U12026 (N_12026,N_11930,N_11899);
xnor U12027 (N_12027,N_11956,N_11891);
nor U12028 (N_12028,N_11879,N_11942);
nand U12029 (N_12029,N_11959,N_11980);
or U12030 (N_12030,N_11933,N_11962);
or U12031 (N_12031,N_11925,N_11976);
or U12032 (N_12032,N_11895,N_11924);
or U12033 (N_12033,N_11945,N_11913);
or U12034 (N_12034,N_11985,N_11935);
or U12035 (N_12035,N_11995,N_11926);
nor U12036 (N_12036,N_11948,N_11972);
or U12037 (N_12037,N_11952,N_11958);
nor U12038 (N_12038,N_11996,N_11937);
nand U12039 (N_12039,N_11987,N_11911);
nand U12040 (N_12040,N_11966,N_11986);
and U12041 (N_12041,N_11982,N_11875);
or U12042 (N_12042,N_11938,N_11904);
or U12043 (N_12043,N_11961,N_11901);
and U12044 (N_12044,N_11929,N_11905);
nor U12045 (N_12045,N_11903,N_11914);
and U12046 (N_12046,N_11931,N_11940);
nor U12047 (N_12047,N_11947,N_11889);
xnor U12048 (N_12048,N_11882,N_11902);
or U12049 (N_12049,N_11894,N_11919);
or U12050 (N_12050,N_11978,N_11887);
nand U12051 (N_12051,N_11968,N_11973);
or U12052 (N_12052,N_11932,N_11939);
or U12053 (N_12053,N_11981,N_11918);
nand U12054 (N_12054,N_11965,N_11977);
xor U12055 (N_12055,N_11936,N_11992);
and U12056 (N_12056,N_11922,N_11881);
and U12057 (N_12057,N_11917,N_11944);
or U12058 (N_12058,N_11998,N_11994);
nand U12059 (N_12059,N_11920,N_11934);
and U12060 (N_12060,N_11900,N_11907);
and U12061 (N_12061,N_11888,N_11915);
nor U12062 (N_12062,N_11999,N_11978);
and U12063 (N_12063,N_11888,N_11961);
or U12064 (N_12064,N_11937,N_11900);
nor U12065 (N_12065,N_11908,N_11959);
and U12066 (N_12066,N_11938,N_11888);
or U12067 (N_12067,N_11884,N_11915);
nor U12068 (N_12068,N_11926,N_11886);
or U12069 (N_12069,N_11988,N_11994);
or U12070 (N_12070,N_11960,N_11978);
xnor U12071 (N_12071,N_11946,N_11993);
or U12072 (N_12072,N_11933,N_11945);
or U12073 (N_12073,N_11961,N_11880);
nand U12074 (N_12074,N_11948,N_11947);
nand U12075 (N_12075,N_11975,N_11968);
nor U12076 (N_12076,N_11915,N_11982);
nand U12077 (N_12077,N_11895,N_11941);
xnor U12078 (N_12078,N_11915,N_11976);
or U12079 (N_12079,N_11987,N_11958);
nand U12080 (N_12080,N_11924,N_11992);
and U12081 (N_12081,N_11938,N_11927);
or U12082 (N_12082,N_11889,N_11900);
nand U12083 (N_12083,N_11993,N_11876);
nor U12084 (N_12084,N_11913,N_11903);
nand U12085 (N_12085,N_11888,N_11966);
nand U12086 (N_12086,N_11970,N_11889);
and U12087 (N_12087,N_11947,N_11883);
or U12088 (N_12088,N_11897,N_11915);
nand U12089 (N_12089,N_11986,N_11997);
nand U12090 (N_12090,N_11905,N_11881);
nand U12091 (N_12091,N_11898,N_11892);
nand U12092 (N_12092,N_11930,N_11932);
or U12093 (N_12093,N_11932,N_11968);
nor U12094 (N_12094,N_11902,N_11968);
and U12095 (N_12095,N_11879,N_11920);
nor U12096 (N_12096,N_11885,N_11945);
nor U12097 (N_12097,N_11984,N_11950);
xnor U12098 (N_12098,N_11928,N_11945);
and U12099 (N_12099,N_11909,N_11981);
xnor U12100 (N_12100,N_11976,N_11998);
nor U12101 (N_12101,N_11978,N_11876);
nand U12102 (N_12102,N_11942,N_11951);
nor U12103 (N_12103,N_11940,N_11929);
nor U12104 (N_12104,N_11939,N_11884);
nand U12105 (N_12105,N_11967,N_11931);
xnor U12106 (N_12106,N_11959,N_11987);
nor U12107 (N_12107,N_11963,N_11934);
nor U12108 (N_12108,N_11979,N_11914);
and U12109 (N_12109,N_11982,N_11938);
or U12110 (N_12110,N_11963,N_11929);
nand U12111 (N_12111,N_11936,N_11998);
and U12112 (N_12112,N_11924,N_11961);
xnor U12113 (N_12113,N_11986,N_11917);
nand U12114 (N_12114,N_11998,N_11904);
nor U12115 (N_12115,N_11929,N_11948);
nand U12116 (N_12116,N_11954,N_11877);
and U12117 (N_12117,N_11917,N_11966);
nor U12118 (N_12118,N_11881,N_11956);
nor U12119 (N_12119,N_11892,N_11976);
nor U12120 (N_12120,N_11916,N_11957);
nor U12121 (N_12121,N_11994,N_11957);
and U12122 (N_12122,N_11961,N_11968);
or U12123 (N_12123,N_11928,N_11902);
or U12124 (N_12124,N_11995,N_11949);
or U12125 (N_12125,N_12031,N_12038);
xor U12126 (N_12126,N_12001,N_12082);
and U12127 (N_12127,N_12026,N_12025);
and U12128 (N_12128,N_12118,N_12097);
or U12129 (N_12129,N_12047,N_12071);
or U12130 (N_12130,N_12006,N_12003);
nor U12131 (N_12131,N_12049,N_12043);
xnor U12132 (N_12132,N_12119,N_12014);
nor U12133 (N_12133,N_12040,N_12028);
xnor U12134 (N_12134,N_12112,N_12117);
and U12135 (N_12135,N_12116,N_12017);
or U12136 (N_12136,N_12042,N_12090);
or U12137 (N_12137,N_12104,N_12093);
and U12138 (N_12138,N_12019,N_12011);
and U12139 (N_12139,N_12109,N_12056);
xor U12140 (N_12140,N_12048,N_12085);
nor U12141 (N_12141,N_12106,N_12076);
nand U12142 (N_12142,N_12012,N_12100);
xnor U12143 (N_12143,N_12078,N_12075);
and U12144 (N_12144,N_12115,N_12121);
or U12145 (N_12145,N_12059,N_12002);
and U12146 (N_12146,N_12023,N_12051);
and U12147 (N_12147,N_12092,N_12033);
nor U12148 (N_12148,N_12105,N_12089);
and U12149 (N_12149,N_12102,N_12039);
or U12150 (N_12150,N_12009,N_12060);
and U12151 (N_12151,N_12122,N_12058);
or U12152 (N_12152,N_12000,N_12063);
nand U12153 (N_12153,N_12084,N_12065);
or U12154 (N_12154,N_12101,N_12062);
or U12155 (N_12155,N_12054,N_12016);
nor U12156 (N_12156,N_12096,N_12073);
nor U12157 (N_12157,N_12007,N_12015);
and U12158 (N_12158,N_12052,N_12021);
or U12159 (N_12159,N_12067,N_12079);
nor U12160 (N_12160,N_12044,N_12055);
or U12161 (N_12161,N_12103,N_12066);
or U12162 (N_12162,N_12108,N_12050);
or U12163 (N_12163,N_12114,N_12037);
xor U12164 (N_12164,N_12029,N_12094);
nand U12165 (N_12165,N_12086,N_12091);
and U12166 (N_12166,N_12036,N_12041);
or U12167 (N_12167,N_12074,N_12099);
nand U12168 (N_12168,N_12005,N_12020);
nand U12169 (N_12169,N_12070,N_12080);
and U12170 (N_12170,N_12083,N_12095);
nand U12171 (N_12171,N_12087,N_12045);
and U12172 (N_12172,N_12123,N_12098);
nor U12173 (N_12173,N_12077,N_12004);
and U12174 (N_12174,N_12030,N_12034);
and U12175 (N_12175,N_12018,N_12113);
or U12176 (N_12176,N_12072,N_12081);
nand U12177 (N_12177,N_12061,N_12064);
or U12178 (N_12178,N_12022,N_12013);
and U12179 (N_12179,N_12111,N_12027);
and U12180 (N_12180,N_12032,N_12107);
xnor U12181 (N_12181,N_12008,N_12053);
nor U12182 (N_12182,N_12024,N_12010);
nor U12183 (N_12183,N_12110,N_12035);
nor U12184 (N_12184,N_12057,N_12046);
or U12185 (N_12185,N_12069,N_12124);
xnor U12186 (N_12186,N_12068,N_12120);
nand U12187 (N_12187,N_12088,N_12027);
nor U12188 (N_12188,N_12078,N_12013);
or U12189 (N_12189,N_12079,N_12020);
xnor U12190 (N_12190,N_12034,N_12002);
or U12191 (N_12191,N_12085,N_12007);
or U12192 (N_12192,N_12017,N_12073);
and U12193 (N_12193,N_12019,N_12001);
and U12194 (N_12194,N_12067,N_12068);
or U12195 (N_12195,N_12124,N_12021);
xnor U12196 (N_12196,N_12066,N_12078);
nand U12197 (N_12197,N_12106,N_12098);
xnor U12198 (N_12198,N_12103,N_12084);
nand U12199 (N_12199,N_12095,N_12047);
nand U12200 (N_12200,N_12090,N_12103);
nor U12201 (N_12201,N_12121,N_12049);
nand U12202 (N_12202,N_12047,N_12124);
or U12203 (N_12203,N_12107,N_12078);
or U12204 (N_12204,N_12065,N_12094);
or U12205 (N_12205,N_12092,N_12098);
nand U12206 (N_12206,N_12048,N_12040);
nand U12207 (N_12207,N_12003,N_12085);
nand U12208 (N_12208,N_12073,N_12064);
nand U12209 (N_12209,N_12108,N_12016);
nor U12210 (N_12210,N_12120,N_12032);
and U12211 (N_12211,N_12068,N_12051);
xnor U12212 (N_12212,N_12001,N_12062);
nand U12213 (N_12213,N_12000,N_12103);
nor U12214 (N_12214,N_12040,N_12060);
and U12215 (N_12215,N_12044,N_12024);
or U12216 (N_12216,N_12111,N_12064);
nor U12217 (N_12217,N_12008,N_12024);
nand U12218 (N_12218,N_12036,N_12111);
or U12219 (N_12219,N_12065,N_12048);
nand U12220 (N_12220,N_12120,N_12072);
nor U12221 (N_12221,N_12038,N_12115);
or U12222 (N_12222,N_12002,N_12101);
or U12223 (N_12223,N_12124,N_12119);
or U12224 (N_12224,N_12120,N_12100);
nor U12225 (N_12225,N_12005,N_12109);
nor U12226 (N_12226,N_12098,N_12020);
nand U12227 (N_12227,N_12052,N_12016);
or U12228 (N_12228,N_12013,N_12016);
or U12229 (N_12229,N_12103,N_12060);
or U12230 (N_12230,N_12094,N_12071);
and U12231 (N_12231,N_12076,N_12071);
and U12232 (N_12232,N_12100,N_12037);
and U12233 (N_12233,N_12085,N_12124);
and U12234 (N_12234,N_12020,N_12071);
or U12235 (N_12235,N_12094,N_12022);
nand U12236 (N_12236,N_12107,N_12065);
and U12237 (N_12237,N_12034,N_12107);
nand U12238 (N_12238,N_12093,N_12083);
nor U12239 (N_12239,N_12057,N_12018);
nor U12240 (N_12240,N_12004,N_12047);
nand U12241 (N_12241,N_12096,N_12038);
and U12242 (N_12242,N_12033,N_12004);
nand U12243 (N_12243,N_12086,N_12026);
xnor U12244 (N_12244,N_12003,N_12047);
xnor U12245 (N_12245,N_12076,N_12018);
nand U12246 (N_12246,N_12095,N_12092);
and U12247 (N_12247,N_12096,N_12100);
xnor U12248 (N_12248,N_12076,N_12080);
nor U12249 (N_12249,N_12015,N_12116);
nor U12250 (N_12250,N_12201,N_12199);
and U12251 (N_12251,N_12210,N_12225);
or U12252 (N_12252,N_12243,N_12179);
or U12253 (N_12253,N_12197,N_12186);
nor U12254 (N_12254,N_12168,N_12219);
nor U12255 (N_12255,N_12145,N_12165);
nand U12256 (N_12256,N_12154,N_12233);
nor U12257 (N_12257,N_12190,N_12188);
nand U12258 (N_12258,N_12142,N_12237);
or U12259 (N_12259,N_12182,N_12224);
nand U12260 (N_12260,N_12139,N_12152);
nand U12261 (N_12261,N_12126,N_12157);
or U12262 (N_12262,N_12235,N_12241);
nor U12263 (N_12263,N_12202,N_12140);
and U12264 (N_12264,N_12147,N_12208);
and U12265 (N_12265,N_12158,N_12153);
and U12266 (N_12266,N_12213,N_12159);
nor U12267 (N_12267,N_12227,N_12212);
or U12268 (N_12268,N_12178,N_12209);
and U12269 (N_12269,N_12217,N_12249);
xnor U12270 (N_12270,N_12170,N_12207);
and U12271 (N_12271,N_12143,N_12148);
nor U12272 (N_12272,N_12163,N_12183);
and U12273 (N_12273,N_12155,N_12185);
or U12274 (N_12274,N_12223,N_12176);
xnor U12275 (N_12275,N_12220,N_12222);
nand U12276 (N_12276,N_12229,N_12129);
nand U12277 (N_12277,N_12181,N_12133);
and U12278 (N_12278,N_12127,N_12128);
nor U12279 (N_12279,N_12138,N_12205);
nand U12280 (N_12280,N_12172,N_12156);
xnor U12281 (N_12281,N_12193,N_12211);
or U12282 (N_12282,N_12231,N_12134);
nand U12283 (N_12283,N_12184,N_12204);
or U12284 (N_12284,N_12232,N_12141);
nor U12285 (N_12285,N_12160,N_12162);
nor U12286 (N_12286,N_12161,N_12151);
and U12287 (N_12287,N_12203,N_12215);
nor U12288 (N_12288,N_12239,N_12131);
xor U12289 (N_12289,N_12144,N_12200);
nor U12290 (N_12290,N_12130,N_12171);
or U12291 (N_12291,N_12247,N_12173);
or U12292 (N_12292,N_12149,N_12180);
nand U12293 (N_12293,N_12221,N_12167);
xnor U12294 (N_12294,N_12192,N_12206);
and U12295 (N_12295,N_12146,N_12135);
or U12296 (N_12296,N_12191,N_12125);
xnor U12297 (N_12297,N_12150,N_12242);
and U12298 (N_12298,N_12226,N_12164);
and U12299 (N_12299,N_12174,N_12240);
or U12300 (N_12300,N_12244,N_12216);
nand U12301 (N_12301,N_12214,N_12132);
and U12302 (N_12302,N_12248,N_12245);
nand U12303 (N_12303,N_12228,N_12234);
nor U12304 (N_12304,N_12175,N_12196);
or U12305 (N_12305,N_12230,N_12198);
nand U12306 (N_12306,N_12189,N_12169);
xnor U12307 (N_12307,N_12195,N_12236);
nand U12308 (N_12308,N_12136,N_12238);
nand U12309 (N_12309,N_12194,N_12218);
nand U12310 (N_12310,N_12187,N_12246);
nor U12311 (N_12311,N_12177,N_12137);
nor U12312 (N_12312,N_12166,N_12197);
or U12313 (N_12313,N_12238,N_12186);
nor U12314 (N_12314,N_12202,N_12166);
nor U12315 (N_12315,N_12141,N_12151);
or U12316 (N_12316,N_12175,N_12188);
nor U12317 (N_12317,N_12238,N_12245);
and U12318 (N_12318,N_12231,N_12190);
nor U12319 (N_12319,N_12134,N_12191);
nand U12320 (N_12320,N_12248,N_12188);
nor U12321 (N_12321,N_12208,N_12238);
and U12322 (N_12322,N_12197,N_12160);
nand U12323 (N_12323,N_12146,N_12125);
nand U12324 (N_12324,N_12140,N_12166);
or U12325 (N_12325,N_12241,N_12186);
and U12326 (N_12326,N_12157,N_12223);
or U12327 (N_12327,N_12209,N_12128);
xor U12328 (N_12328,N_12189,N_12245);
nand U12329 (N_12329,N_12135,N_12163);
nand U12330 (N_12330,N_12175,N_12209);
and U12331 (N_12331,N_12247,N_12230);
nor U12332 (N_12332,N_12178,N_12179);
nand U12333 (N_12333,N_12140,N_12213);
nor U12334 (N_12334,N_12242,N_12186);
nor U12335 (N_12335,N_12237,N_12165);
or U12336 (N_12336,N_12189,N_12203);
nor U12337 (N_12337,N_12242,N_12154);
and U12338 (N_12338,N_12225,N_12131);
nor U12339 (N_12339,N_12190,N_12172);
nand U12340 (N_12340,N_12137,N_12148);
nor U12341 (N_12341,N_12214,N_12128);
or U12342 (N_12342,N_12232,N_12145);
and U12343 (N_12343,N_12177,N_12240);
and U12344 (N_12344,N_12198,N_12221);
xor U12345 (N_12345,N_12147,N_12162);
or U12346 (N_12346,N_12156,N_12129);
nor U12347 (N_12347,N_12199,N_12237);
nor U12348 (N_12348,N_12142,N_12185);
and U12349 (N_12349,N_12212,N_12170);
or U12350 (N_12350,N_12186,N_12224);
nor U12351 (N_12351,N_12201,N_12234);
or U12352 (N_12352,N_12170,N_12204);
nand U12353 (N_12353,N_12203,N_12221);
nand U12354 (N_12354,N_12192,N_12151);
or U12355 (N_12355,N_12173,N_12153);
nand U12356 (N_12356,N_12159,N_12148);
nor U12357 (N_12357,N_12239,N_12207);
nand U12358 (N_12358,N_12186,N_12219);
nor U12359 (N_12359,N_12141,N_12181);
or U12360 (N_12360,N_12217,N_12155);
or U12361 (N_12361,N_12233,N_12208);
nand U12362 (N_12362,N_12156,N_12133);
nand U12363 (N_12363,N_12144,N_12172);
nor U12364 (N_12364,N_12191,N_12178);
nor U12365 (N_12365,N_12166,N_12237);
and U12366 (N_12366,N_12142,N_12248);
and U12367 (N_12367,N_12147,N_12139);
or U12368 (N_12368,N_12209,N_12199);
and U12369 (N_12369,N_12179,N_12228);
and U12370 (N_12370,N_12215,N_12134);
and U12371 (N_12371,N_12149,N_12227);
xor U12372 (N_12372,N_12243,N_12185);
nand U12373 (N_12373,N_12156,N_12154);
xor U12374 (N_12374,N_12193,N_12225);
nand U12375 (N_12375,N_12357,N_12283);
nor U12376 (N_12376,N_12342,N_12358);
and U12377 (N_12377,N_12368,N_12351);
nor U12378 (N_12378,N_12317,N_12349);
nor U12379 (N_12379,N_12307,N_12279);
xor U12380 (N_12380,N_12327,N_12353);
xnor U12381 (N_12381,N_12336,N_12274);
and U12382 (N_12382,N_12295,N_12289);
nor U12383 (N_12383,N_12303,N_12263);
or U12384 (N_12384,N_12277,N_12280);
or U12385 (N_12385,N_12372,N_12286);
nor U12386 (N_12386,N_12276,N_12294);
or U12387 (N_12387,N_12281,N_12373);
nor U12388 (N_12388,N_12270,N_12313);
nor U12389 (N_12389,N_12254,N_12311);
nand U12390 (N_12390,N_12297,N_12370);
nand U12391 (N_12391,N_12366,N_12331);
nor U12392 (N_12392,N_12359,N_12258);
nor U12393 (N_12393,N_12324,N_12361);
and U12394 (N_12394,N_12339,N_12255);
nand U12395 (N_12395,N_12347,N_12329);
and U12396 (N_12396,N_12323,N_12367);
nand U12397 (N_12397,N_12287,N_12371);
xor U12398 (N_12398,N_12320,N_12321);
or U12399 (N_12399,N_12266,N_12262);
nor U12400 (N_12400,N_12344,N_12340);
nor U12401 (N_12401,N_12374,N_12291);
and U12402 (N_12402,N_12345,N_12253);
nor U12403 (N_12403,N_12284,N_12304);
or U12404 (N_12404,N_12306,N_12332);
or U12405 (N_12405,N_12292,N_12363);
xnor U12406 (N_12406,N_12278,N_12328);
and U12407 (N_12407,N_12298,N_12290);
nor U12408 (N_12408,N_12348,N_12350);
or U12409 (N_12409,N_12265,N_12264);
nand U12410 (N_12410,N_12275,N_12296);
nand U12411 (N_12411,N_12326,N_12337);
and U12412 (N_12412,N_12256,N_12354);
nand U12413 (N_12413,N_12260,N_12316);
xor U12414 (N_12414,N_12355,N_12305);
or U12415 (N_12415,N_12318,N_12314);
nand U12416 (N_12416,N_12302,N_12356);
and U12417 (N_12417,N_12273,N_12250);
or U12418 (N_12418,N_12338,N_12301);
or U12419 (N_12419,N_12312,N_12362);
or U12420 (N_12420,N_12300,N_12315);
nand U12421 (N_12421,N_12272,N_12308);
and U12422 (N_12422,N_12360,N_12288);
and U12423 (N_12423,N_12267,N_12269);
nor U12424 (N_12424,N_12346,N_12251);
nand U12425 (N_12425,N_12325,N_12330);
and U12426 (N_12426,N_12268,N_12352);
and U12427 (N_12427,N_12259,N_12334);
and U12428 (N_12428,N_12343,N_12335);
and U12429 (N_12429,N_12293,N_12261);
or U12430 (N_12430,N_12341,N_12309);
xnor U12431 (N_12431,N_12299,N_12285);
xnor U12432 (N_12432,N_12365,N_12310);
nor U12433 (N_12433,N_12319,N_12282);
nor U12434 (N_12434,N_12271,N_12252);
nor U12435 (N_12435,N_12369,N_12322);
nor U12436 (N_12436,N_12257,N_12364);
and U12437 (N_12437,N_12333,N_12356);
or U12438 (N_12438,N_12258,N_12259);
nand U12439 (N_12439,N_12314,N_12355);
xor U12440 (N_12440,N_12287,N_12342);
or U12441 (N_12441,N_12311,N_12250);
nor U12442 (N_12442,N_12287,N_12289);
or U12443 (N_12443,N_12258,N_12311);
nand U12444 (N_12444,N_12266,N_12299);
nand U12445 (N_12445,N_12287,N_12293);
nand U12446 (N_12446,N_12304,N_12322);
and U12447 (N_12447,N_12265,N_12281);
nand U12448 (N_12448,N_12309,N_12374);
and U12449 (N_12449,N_12342,N_12339);
and U12450 (N_12450,N_12352,N_12266);
nand U12451 (N_12451,N_12303,N_12359);
or U12452 (N_12452,N_12345,N_12357);
nor U12453 (N_12453,N_12306,N_12261);
nor U12454 (N_12454,N_12314,N_12269);
or U12455 (N_12455,N_12317,N_12270);
nor U12456 (N_12456,N_12318,N_12347);
nand U12457 (N_12457,N_12263,N_12261);
nand U12458 (N_12458,N_12267,N_12307);
nand U12459 (N_12459,N_12331,N_12370);
and U12460 (N_12460,N_12358,N_12309);
xnor U12461 (N_12461,N_12266,N_12291);
nand U12462 (N_12462,N_12269,N_12260);
nor U12463 (N_12463,N_12345,N_12333);
or U12464 (N_12464,N_12351,N_12344);
and U12465 (N_12465,N_12301,N_12274);
nor U12466 (N_12466,N_12269,N_12358);
nor U12467 (N_12467,N_12343,N_12283);
or U12468 (N_12468,N_12371,N_12276);
or U12469 (N_12469,N_12321,N_12328);
or U12470 (N_12470,N_12293,N_12366);
and U12471 (N_12471,N_12333,N_12297);
nand U12472 (N_12472,N_12347,N_12334);
xor U12473 (N_12473,N_12302,N_12251);
nor U12474 (N_12474,N_12317,N_12373);
or U12475 (N_12475,N_12334,N_12263);
or U12476 (N_12476,N_12259,N_12296);
nor U12477 (N_12477,N_12309,N_12307);
and U12478 (N_12478,N_12342,N_12361);
and U12479 (N_12479,N_12282,N_12336);
nor U12480 (N_12480,N_12280,N_12351);
xnor U12481 (N_12481,N_12316,N_12357);
and U12482 (N_12482,N_12330,N_12256);
and U12483 (N_12483,N_12321,N_12276);
xor U12484 (N_12484,N_12304,N_12359);
nor U12485 (N_12485,N_12320,N_12284);
xor U12486 (N_12486,N_12258,N_12263);
or U12487 (N_12487,N_12337,N_12340);
xor U12488 (N_12488,N_12283,N_12332);
xnor U12489 (N_12489,N_12274,N_12299);
nor U12490 (N_12490,N_12263,N_12341);
and U12491 (N_12491,N_12275,N_12363);
or U12492 (N_12492,N_12269,N_12326);
nand U12493 (N_12493,N_12330,N_12302);
and U12494 (N_12494,N_12274,N_12344);
or U12495 (N_12495,N_12264,N_12325);
and U12496 (N_12496,N_12328,N_12279);
or U12497 (N_12497,N_12296,N_12302);
nand U12498 (N_12498,N_12258,N_12343);
or U12499 (N_12499,N_12306,N_12358);
nor U12500 (N_12500,N_12393,N_12450);
and U12501 (N_12501,N_12477,N_12487);
nor U12502 (N_12502,N_12389,N_12400);
nand U12503 (N_12503,N_12474,N_12440);
nand U12504 (N_12504,N_12432,N_12498);
nor U12505 (N_12505,N_12484,N_12426);
and U12506 (N_12506,N_12475,N_12408);
or U12507 (N_12507,N_12434,N_12442);
and U12508 (N_12508,N_12468,N_12390);
and U12509 (N_12509,N_12378,N_12418);
and U12510 (N_12510,N_12382,N_12394);
xnor U12511 (N_12511,N_12470,N_12424);
and U12512 (N_12512,N_12377,N_12490);
and U12513 (N_12513,N_12401,N_12419);
or U12514 (N_12514,N_12412,N_12464);
nand U12515 (N_12515,N_12427,N_12443);
nand U12516 (N_12516,N_12482,N_12485);
and U12517 (N_12517,N_12472,N_12465);
nand U12518 (N_12518,N_12410,N_12491);
or U12519 (N_12519,N_12456,N_12460);
xor U12520 (N_12520,N_12461,N_12481);
nand U12521 (N_12521,N_12435,N_12420);
and U12522 (N_12522,N_12488,N_12494);
nor U12523 (N_12523,N_12396,N_12391);
or U12524 (N_12524,N_12411,N_12478);
nand U12525 (N_12525,N_12399,N_12387);
nand U12526 (N_12526,N_12406,N_12462);
nand U12527 (N_12527,N_12433,N_12455);
and U12528 (N_12528,N_12495,N_12376);
xor U12529 (N_12529,N_12421,N_12476);
or U12530 (N_12530,N_12398,N_12414);
or U12531 (N_12531,N_12445,N_12422);
and U12532 (N_12532,N_12452,N_12417);
or U12533 (N_12533,N_12453,N_12496);
nor U12534 (N_12534,N_12405,N_12431);
or U12535 (N_12535,N_12441,N_12499);
and U12536 (N_12536,N_12459,N_12380);
nand U12537 (N_12537,N_12386,N_12429);
xnor U12538 (N_12538,N_12454,N_12409);
nor U12539 (N_12539,N_12448,N_12388);
and U12540 (N_12540,N_12402,N_12446);
xor U12541 (N_12541,N_12497,N_12449);
and U12542 (N_12542,N_12457,N_12395);
nand U12543 (N_12543,N_12384,N_12416);
or U12544 (N_12544,N_12379,N_12413);
nand U12545 (N_12545,N_12439,N_12473);
or U12546 (N_12546,N_12415,N_12404);
nand U12547 (N_12547,N_12407,N_12451);
or U12548 (N_12548,N_12430,N_12489);
xor U12549 (N_12549,N_12438,N_12425);
nor U12550 (N_12550,N_12423,N_12493);
nand U12551 (N_12551,N_12492,N_12483);
xnor U12552 (N_12552,N_12480,N_12486);
nand U12553 (N_12553,N_12436,N_12467);
nor U12554 (N_12554,N_12392,N_12383);
nand U12555 (N_12555,N_12381,N_12479);
or U12556 (N_12556,N_12428,N_12444);
nand U12557 (N_12557,N_12385,N_12375);
nor U12558 (N_12558,N_12466,N_12471);
nand U12559 (N_12559,N_12458,N_12447);
nand U12560 (N_12560,N_12463,N_12469);
or U12561 (N_12561,N_12437,N_12397);
nor U12562 (N_12562,N_12403,N_12420);
and U12563 (N_12563,N_12414,N_12494);
nor U12564 (N_12564,N_12385,N_12450);
and U12565 (N_12565,N_12424,N_12467);
nor U12566 (N_12566,N_12396,N_12384);
or U12567 (N_12567,N_12436,N_12391);
xnor U12568 (N_12568,N_12450,N_12399);
nand U12569 (N_12569,N_12461,N_12393);
nor U12570 (N_12570,N_12462,N_12474);
xor U12571 (N_12571,N_12461,N_12430);
xnor U12572 (N_12572,N_12455,N_12438);
and U12573 (N_12573,N_12428,N_12431);
nand U12574 (N_12574,N_12489,N_12493);
nand U12575 (N_12575,N_12434,N_12477);
nand U12576 (N_12576,N_12417,N_12407);
nand U12577 (N_12577,N_12433,N_12486);
and U12578 (N_12578,N_12426,N_12400);
nand U12579 (N_12579,N_12385,N_12410);
or U12580 (N_12580,N_12469,N_12442);
and U12581 (N_12581,N_12482,N_12447);
or U12582 (N_12582,N_12389,N_12464);
nand U12583 (N_12583,N_12391,N_12419);
and U12584 (N_12584,N_12450,N_12493);
nand U12585 (N_12585,N_12439,N_12405);
or U12586 (N_12586,N_12378,N_12485);
nand U12587 (N_12587,N_12377,N_12441);
and U12588 (N_12588,N_12417,N_12497);
and U12589 (N_12589,N_12493,N_12424);
nand U12590 (N_12590,N_12443,N_12474);
nor U12591 (N_12591,N_12457,N_12419);
and U12592 (N_12592,N_12461,N_12425);
and U12593 (N_12593,N_12402,N_12380);
or U12594 (N_12594,N_12447,N_12452);
nand U12595 (N_12595,N_12461,N_12451);
nor U12596 (N_12596,N_12424,N_12376);
and U12597 (N_12597,N_12422,N_12388);
nor U12598 (N_12598,N_12474,N_12442);
and U12599 (N_12599,N_12466,N_12422);
nor U12600 (N_12600,N_12496,N_12455);
or U12601 (N_12601,N_12400,N_12488);
nand U12602 (N_12602,N_12497,N_12390);
nor U12603 (N_12603,N_12382,N_12415);
nand U12604 (N_12604,N_12451,N_12421);
or U12605 (N_12605,N_12383,N_12490);
nand U12606 (N_12606,N_12429,N_12378);
nand U12607 (N_12607,N_12499,N_12497);
or U12608 (N_12608,N_12478,N_12491);
nand U12609 (N_12609,N_12444,N_12401);
and U12610 (N_12610,N_12495,N_12445);
and U12611 (N_12611,N_12498,N_12421);
xor U12612 (N_12612,N_12408,N_12426);
nor U12613 (N_12613,N_12499,N_12425);
nand U12614 (N_12614,N_12478,N_12428);
nand U12615 (N_12615,N_12474,N_12451);
and U12616 (N_12616,N_12400,N_12391);
and U12617 (N_12617,N_12459,N_12485);
or U12618 (N_12618,N_12439,N_12475);
and U12619 (N_12619,N_12414,N_12463);
and U12620 (N_12620,N_12433,N_12488);
nor U12621 (N_12621,N_12381,N_12484);
and U12622 (N_12622,N_12495,N_12493);
nand U12623 (N_12623,N_12491,N_12460);
xnor U12624 (N_12624,N_12404,N_12440);
and U12625 (N_12625,N_12562,N_12602);
nand U12626 (N_12626,N_12567,N_12592);
xor U12627 (N_12627,N_12623,N_12510);
xor U12628 (N_12628,N_12601,N_12524);
and U12629 (N_12629,N_12546,N_12563);
nor U12630 (N_12630,N_12608,N_12509);
nor U12631 (N_12631,N_12518,N_12568);
nor U12632 (N_12632,N_12534,N_12599);
nor U12633 (N_12633,N_12588,N_12538);
nand U12634 (N_12634,N_12532,N_12522);
and U12635 (N_12635,N_12583,N_12580);
nand U12636 (N_12636,N_12615,N_12593);
nand U12637 (N_12637,N_12561,N_12515);
nor U12638 (N_12638,N_12519,N_12566);
and U12639 (N_12639,N_12545,N_12527);
nor U12640 (N_12640,N_12556,N_12500);
nor U12641 (N_12641,N_12511,N_12528);
nor U12642 (N_12642,N_12570,N_12598);
xor U12643 (N_12643,N_12620,N_12557);
nor U12644 (N_12644,N_12517,N_12604);
and U12645 (N_12645,N_12520,N_12572);
nand U12646 (N_12646,N_12617,N_12558);
xor U12647 (N_12647,N_12578,N_12603);
nor U12648 (N_12648,N_12573,N_12609);
nand U12649 (N_12649,N_12612,N_12569);
xnor U12650 (N_12650,N_12614,N_12514);
or U12651 (N_12651,N_12513,N_12553);
nor U12652 (N_12652,N_12536,N_12516);
and U12653 (N_12653,N_12574,N_12531);
nand U12654 (N_12654,N_12548,N_12539);
and U12655 (N_12655,N_12564,N_12611);
or U12656 (N_12656,N_12523,N_12547);
nand U12657 (N_12657,N_12624,N_12610);
nand U12658 (N_12658,N_12560,N_12576);
nand U12659 (N_12659,N_12542,N_12622);
xnor U12660 (N_12660,N_12571,N_12587);
nand U12661 (N_12661,N_12596,N_12521);
and U12662 (N_12662,N_12579,N_12541);
and U12663 (N_12663,N_12607,N_12543);
nor U12664 (N_12664,N_12591,N_12585);
nand U12665 (N_12665,N_12575,N_12577);
nand U12666 (N_12666,N_12594,N_12530);
or U12667 (N_12667,N_12606,N_12526);
nor U12668 (N_12668,N_12529,N_12605);
nor U12669 (N_12669,N_12590,N_12555);
or U12670 (N_12670,N_12559,N_12503);
xnor U12671 (N_12671,N_12597,N_12586);
nor U12672 (N_12672,N_12619,N_12600);
nor U12673 (N_12673,N_12505,N_12613);
nor U12674 (N_12674,N_12554,N_12501);
nand U12675 (N_12675,N_12535,N_12581);
nor U12676 (N_12676,N_12616,N_12525);
and U12677 (N_12677,N_12595,N_12506);
or U12678 (N_12678,N_12507,N_12550);
nor U12679 (N_12679,N_12537,N_12504);
nor U12680 (N_12680,N_12621,N_12618);
and U12681 (N_12681,N_12540,N_12584);
or U12682 (N_12682,N_12589,N_12582);
nor U12683 (N_12683,N_12508,N_12552);
nor U12684 (N_12684,N_12533,N_12544);
and U12685 (N_12685,N_12565,N_12551);
nand U12686 (N_12686,N_12512,N_12549);
nand U12687 (N_12687,N_12502,N_12623);
or U12688 (N_12688,N_12565,N_12574);
and U12689 (N_12689,N_12598,N_12535);
nor U12690 (N_12690,N_12516,N_12598);
nand U12691 (N_12691,N_12598,N_12504);
and U12692 (N_12692,N_12579,N_12573);
or U12693 (N_12693,N_12591,N_12608);
nor U12694 (N_12694,N_12501,N_12610);
or U12695 (N_12695,N_12555,N_12606);
and U12696 (N_12696,N_12599,N_12607);
or U12697 (N_12697,N_12554,N_12557);
and U12698 (N_12698,N_12553,N_12510);
xnor U12699 (N_12699,N_12565,N_12569);
or U12700 (N_12700,N_12600,N_12610);
nand U12701 (N_12701,N_12589,N_12512);
or U12702 (N_12702,N_12587,N_12596);
or U12703 (N_12703,N_12509,N_12622);
nor U12704 (N_12704,N_12585,N_12594);
nand U12705 (N_12705,N_12536,N_12599);
and U12706 (N_12706,N_12557,N_12540);
nand U12707 (N_12707,N_12576,N_12500);
nor U12708 (N_12708,N_12568,N_12613);
nor U12709 (N_12709,N_12592,N_12588);
and U12710 (N_12710,N_12580,N_12527);
and U12711 (N_12711,N_12548,N_12584);
nand U12712 (N_12712,N_12525,N_12563);
or U12713 (N_12713,N_12613,N_12555);
or U12714 (N_12714,N_12515,N_12591);
nor U12715 (N_12715,N_12577,N_12618);
or U12716 (N_12716,N_12615,N_12555);
xnor U12717 (N_12717,N_12534,N_12612);
or U12718 (N_12718,N_12592,N_12536);
and U12719 (N_12719,N_12537,N_12623);
nand U12720 (N_12720,N_12582,N_12524);
and U12721 (N_12721,N_12512,N_12538);
nor U12722 (N_12722,N_12621,N_12508);
nand U12723 (N_12723,N_12531,N_12553);
nor U12724 (N_12724,N_12617,N_12618);
nand U12725 (N_12725,N_12501,N_12580);
nor U12726 (N_12726,N_12528,N_12575);
xnor U12727 (N_12727,N_12587,N_12594);
nand U12728 (N_12728,N_12624,N_12614);
or U12729 (N_12729,N_12622,N_12570);
or U12730 (N_12730,N_12601,N_12596);
nand U12731 (N_12731,N_12586,N_12595);
or U12732 (N_12732,N_12590,N_12585);
or U12733 (N_12733,N_12553,N_12505);
and U12734 (N_12734,N_12607,N_12512);
or U12735 (N_12735,N_12597,N_12513);
and U12736 (N_12736,N_12550,N_12509);
nor U12737 (N_12737,N_12619,N_12576);
and U12738 (N_12738,N_12592,N_12624);
or U12739 (N_12739,N_12590,N_12616);
and U12740 (N_12740,N_12572,N_12553);
xnor U12741 (N_12741,N_12603,N_12515);
and U12742 (N_12742,N_12535,N_12555);
nor U12743 (N_12743,N_12594,N_12520);
nand U12744 (N_12744,N_12593,N_12609);
nand U12745 (N_12745,N_12624,N_12622);
nor U12746 (N_12746,N_12620,N_12601);
xnor U12747 (N_12747,N_12608,N_12508);
xnor U12748 (N_12748,N_12528,N_12609);
nor U12749 (N_12749,N_12599,N_12517);
nor U12750 (N_12750,N_12637,N_12715);
or U12751 (N_12751,N_12639,N_12649);
nand U12752 (N_12752,N_12712,N_12628);
nand U12753 (N_12753,N_12659,N_12691);
nor U12754 (N_12754,N_12685,N_12731);
nand U12755 (N_12755,N_12702,N_12713);
and U12756 (N_12756,N_12666,N_12723);
or U12757 (N_12757,N_12737,N_12650);
or U12758 (N_12758,N_12646,N_12665);
and U12759 (N_12759,N_12658,N_12726);
nand U12760 (N_12760,N_12745,N_12724);
xor U12761 (N_12761,N_12682,N_12652);
nand U12762 (N_12762,N_12667,N_12684);
nand U12763 (N_12763,N_12630,N_12670);
nor U12764 (N_12764,N_12641,N_12674);
nor U12765 (N_12765,N_12678,N_12743);
nand U12766 (N_12766,N_12662,N_12734);
nor U12767 (N_12767,N_12632,N_12676);
nor U12768 (N_12768,N_12717,N_12697);
or U12769 (N_12769,N_12720,N_12625);
nand U12770 (N_12770,N_12725,N_12675);
and U12771 (N_12771,N_12738,N_12729);
nor U12772 (N_12772,N_12681,N_12648);
nor U12773 (N_12773,N_12741,N_12704);
xnor U12774 (N_12774,N_12740,N_12739);
or U12775 (N_12775,N_12696,N_12672);
nor U12776 (N_12776,N_12644,N_12626);
or U12777 (N_12777,N_12703,N_12688);
xor U12778 (N_12778,N_12690,N_12645);
and U12779 (N_12779,N_12627,N_12653);
nand U12780 (N_12780,N_12719,N_12669);
and U12781 (N_12781,N_12749,N_12705);
nor U12782 (N_12782,N_12656,N_12742);
and U12783 (N_12783,N_12636,N_12699);
or U12784 (N_12784,N_12747,N_12660);
nor U12785 (N_12785,N_12709,N_12651);
nand U12786 (N_12786,N_12683,N_12668);
or U12787 (N_12787,N_12647,N_12654);
and U12788 (N_12788,N_12689,N_12708);
nand U12789 (N_12789,N_12694,N_12728);
and U12790 (N_12790,N_12707,N_12693);
nand U12791 (N_12791,N_12730,N_12714);
and U12792 (N_12792,N_12695,N_12687);
and U12793 (N_12793,N_12677,N_12711);
nand U12794 (N_12794,N_12679,N_12643);
nor U12795 (N_12795,N_12718,N_12706);
xor U12796 (N_12796,N_12727,N_12680);
nand U12797 (N_12797,N_12657,N_12716);
xnor U12798 (N_12798,N_12701,N_12640);
or U12799 (N_12799,N_12686,N_12635);
nor U12800 (N_12800,N_12746,N_12655);
and U12801 (N_12801,N_12733,N_12710);
or U12802 (N_12802,N_12629,N_12673);
or U12803 (N_12803,N_12721,N_12735);
nor U12804 (N_12804,N_12642,N_12671);
or U12805 (N_12805,N_12736,N_12700);
xnor U12806 (N_12806,N_12748,N_12631);
nand U12807 (N_12807,N_12692,N_12633);
nand U12808 (N_12808,N_12661,N_12698);
nand U12809 (N_12809,N_12732,N_12744);
or U12810 (N_12810,N_12663,N_12722);
nand U12811 (N_12811,N_12664,N_12638);
nor U12812 (N_12812,N_12634,N_12670);
nand U12813 (N_12813,N_12742,N_12730);
nor U12814 (N_12814,N_12749,N_12678);
and U12815 (N_12815,N_12674,N_12721);
nor U12816 (N_12816,N_12732,N_12676);
nand U12817 (N_12817,N_12725,N_12705);
or U12818 (N_12818,N_12666,N_12681);
nand U12819 (N_12819,N_12749,N_12644);
nand U12820 (N_12820,N_12648,N_12633);
nand U12821 (N_12821,N_12692,N_12739);
nand U12822 (N_12822,N_12643,N_12705);
and U12823 (N_12823,N_12657,N_12740);
nand U12824 (N_12824,N_12661,N_12747);
and U12825 (N_12825,N_12671,N_12685);
or U12826 (N_12826,N_12656,N_12695);
and U12827 (N_12827,N_12633,N_12720);
or U12828 (N_12828,N_12708,N_12739);
nand U12829 (N_12829,N_12638,N_12741);
nand U12830 (N_12830,N_12672,N_12722);
nor U12831 (N_12831,N_12631,N_12651);
and U12832 (N_12832,N_12704,N_12718);
or U12833 (N_12833,N_12749,N_12698);
and U12834 (N_12834,N_12744,N_12632);
nand U12835 (N_12835,N_12640,N_12693);
nand U12836 (N_12836,N_12640,N_12692);
nand U12837 (N_12837,N_12655,N_12709);
nand U12838 (N_12838,N_12649,N_12689);
or U12839 (N_12839,N_12646,N_12712);
or U12840 (N_12840,N_12747,N_12634);
nand U12841 (N_12841,N_12663,N_12716);
nor U12842 (N_12842,N_12684,N_12649);
nor U12843 (N_12843,N_12683,N_12636);
nand U12844 (N_12844,N_12733,N_12640);
or U12845 (N_12845,N_12682,N_12728);
nand U12846 (N_12846,N_12712,N_12736);
or U12847 (N_12847,N_12728,N_12644);
nor U12848 (N_12848,N_12745,N_12728);
and U12849 (N_12849,N_12645,N_12633);
nand U12850 (N_12850,N_12681,N_12739);
or U12851 (N_12851,N_12734,N_12649);
nor U12852 (N_12852,N_12711,N_12659);
nor U12853 (N_12853,N_12694,N_12748);
and U12854 (N_12854,N_12721,N_12649);
and U12855 (N_12855,N_12626,N_12654);
or U12856 (N_12856,N_12691,N_12724);
or U12857 (N_12857,N_12705,N_12669);
and U12858 (N_12858,N_12704,N_12686);
xnor U12859 (N_12859,N_12698,N_12696);
or U12860 (N_12860,N_12727,N_12699);
xor U12861 (N_12861,N_12671,N_12679);
nor U12862 (N_12862,N_12686,N_12647);
and U12863 (N_12863,N_12669,N_12728);
or U12864 (N_12864,N_12733,N_12730);
and U12865 (N_12865,N_12718,N_12684);
and U12866 (N_12866,N_12650,N_12686);
xnor U12867 (N_12867,N_12740,N_12632);
or U12868 (N_12868,N_12628,N_12657);
nand U12869 (N_12869,N_12684,N_12694);
or U12870 (N_12870,N_12627,N_12727);
nand U12871 (N_12871,N_12693,N_12747);
or U12872 (N_12872,N_12746,N_12701);
nand U12873 (N_12873,N_12749,N_12740);
xor U12874 (N_12874,N_12744,N_12627);
and U12875 (N_12875,N_12807,N_12873);
and U12876 (N_12876,N_12841,N_12772);
or U12877 (N_12877,N_12770,N_12760);
xnor U12878 (N_12878,N_12803,N_12805);
and U12879 (N_12879,N_12780,N_12872);
nand U12880 (N_12880,N_12863,N_12777);
nor U12881 (N_12881,N_12858,N_12857);
and U12882 (N_12882,N_12845,N_12806);
or U12883 (N_12883,N_12825,N_12787);
and U12884 (N_12884,N_12862,N_12768);
and U12885 (N_12885,N_12759,N_12784);
nor U12886 (N_12886,N_12752,N_12824);
or U12887 (N_12887,N_12814,N_12812);
nor U12888 (N_12888,N_12838,N_12800);
or U12889 (N_12889,N_12765,N_12843);
nor U12890 (N_12890,N_12793,N_12860);
nand U12891 (N_12891,N_12855,N_12785);
nand U12892 (N_12892,N_12775,N_12783);
nor U12893 (N_12893,N_12864,N_12767);
nor U12894 (N_12894,N_12868,N_12782);
xor U12895 (N_12895,N_12833,N_12790);
or U12896 (N_12896,N_12854,N_12773);
and U12897 (N_12897,N_12842,N_12828);
nor U12898 (N_12898,N_12786,N_12789);
xnor U12899 (N_12899,N_12820,N_12850);
nor U12900 (N_12900,N_12844,N_12761);
or U12901 (N_12901,N_12769,N_12758);
or U12902 (N_12902,N_12778,N_12836);
nor U12903 (N_12903,N_12874,N_12818);
xor U12904 (N_12904,N_12822,N_12791);
and U12905 (N_12905,N_12856,N_12830);
or U12906 (N_12906,N_12870,N_12799);
or U12907 (N_12907,N_12766,N_12861);
or U12908 (N_12908,N_12846,N_12817);
xor U12909 (N_12909,N_12788,N_12832);
nand U12910 (N_12910,N_12802,N_12827);
nor U12911 (N_12911,N_12853,N_12859);
xnor U12912 (N_12912,N_12819,N_12792);
and U12913 (N_12913,N_12837,N_12751);
and U12914 (N_12914,N_12829,N_12750);
or U12915 (N_12915,N_12811,N_12795);
nor U12916 (N_12916,N_12794,N_12756);
nor U12917 (N_12917,N_12779,N_12848);
or U12918 (N_12918,N_12849,N_12757);
and U12919 (N_12919,N_12776,N_12867);
nor U12920 (N_12920,N_12852,N_12835);
and U12921 (N_12921,N_12771,N_12804);
nand U12922 (N_12922,N_12831,N_12816);
nor U12923 (N_12923,N_12810,N_12809);
or U12924 (N_12924,N_12865,N_12764);
nand U12925 (N_12925,N_12834,N_12753);
nand U12926 (N_12926,N_12866,N_12826);
nand U12927 (N_12927,N_12871,N_12808);
or U12928 (N_12928,N_12763,N_12840);
xnor U12929 (N_12929,N_12839,N_12851);
and U12930 (N_12930,N_12754,N_12762);
nand U12931 (N_12931,N_12781,N_12801);
nor U12932 (N_12932,N_12813,N_12847);
nor U12933 (N_12933,N_12755,N_12869);
xor U12934 (N_12934,N_12815,N_12774);
xnor U12935 (N_12935,N_12821,N_12796);
or U12936 (N_12936,N_12823,N_12798);
nor U12937 (N_12937,N_12797,N_12793);
and U12938 (N_12938,N_12855,N_12763);
or U12939 (N_12939,N_12775,N_12796);
xnor U12940 (N_12940,N_12761,N_12872);
nor U12941 (N_12941,N_12860,N_12854);
nor U12942 (N_12942,N_12839,N_12785);
nor U12943 (N_12943,N_12758,N_12855);
and U12944 (N_12944,N_12811,N_12870);
or U12945 (N_12945,N_12834,N_12849);
or U12946 (N_12946,N_12824,N_12774);
nor U12947 (N_12947,N_12772,N_12750);
xor U12948 (N_12948,N_12770,N_12843);
or U12949 (N_12949,N_12774,N_12773);
xor U12950 (N_12950,N_12840,N_12761);
xor U12951 (N_12951,N_12775,N_12832);
nand U12952 (N_12952,N_12818,N_12789);
nand U12953 (N_12953,N_12857,N_12790);
and U12954 (N_12954,N_12874,N_12834);
xor U12955 (N_12955,N_12853,N_12803);
and U12956 (N_12956,N_12853,N_12826);
and U12957 (N_12957,N_12767,N_12769);
and U12958 (N_12958,N_12840,N_12821);
xnor U12959 (N_12959,N_12816,N_12798);
and U12960 (N_12960,N_12863,N_12855);
or U12961 (N_12961,N_12810,N_12754);
nor U12962 (N_12962,N_12827,N_12850);
xor U12963 (N_12963,N_12857,N_12865);
and U12964 (N_12964,N_12828,N_12768);
nand U12965 (N_12965,N_12821,N_12841);
and U12966 (N_12966,N_12764,N_12753);
or U12967 (N_12967,N_12812,N_12855);
nand U12968 (N_12968,N_12819,N_12871);
or U12969 (N_12969,N_12801,N_12871);
or U12970 (N_12970,N_12799,N_12805);
xor U12971 (N_12971,N_12855,N_12766);
or U12972 (N_12972,N_12810,N_12759);
or U12973 (N_12973,N_12860,N_12763);
and U12974 (N_12974,N_12856,N_12789);
nand U12975 (N_12975,N_12832,N_12755);
nor U12976 (N_12976,N_12764,N_12808);
xor U12977 (N_12977,N_12865,N_12759);
nand U12978 (N_12978,N_12839,N_12772);
nand U12979 (N_12979,N_12808,N_12779);
and U12980 (N_12980,N_12793,N_12845);
or U12981 (N_12981,N_12776,N_12851);
or U12982 (N_12982,N_12837,N_12789);
or U12983 (N_12983,N_12789,N_12795);
and U12984 (N_12984,N_12754,N_12855);
and U12985 (N_12985,N_12851,N_12750);
nor U12986 (N_12986,N_12764,N_12850);
or U12987 (N_12987,N_12857,N_12839);
or U12988 (N_12988,N_12789,N_12757);
or U12989 (N_12989,N_12781,N_12750);
and U12990 (N_12990,N_12821,N_12827);
or U12991 (N_12991,N_12785,N_12866);
and U12992 (N_12992,N_12771,N_12765);
and U12993 (N_12993,N_12864,N_12762);
nand U12994 (N_12994,N_12771,N_12760);
and U12995 (N_12995,N_12790,N_12819);
and U12996 (N_12996,N_12813,N_12775);
or U12997 (N_12997,N_12812,N_12846);
nand U12998 (N_12998,N_12808,N_12807);
or U12999 (N_12999,N_12758,N_12751);
or U13000 (N_13000,N_12966,N_12896);
nand U13001 (N_13001,N_12969,N_12994);
nand U13002 (N_13002,N_12892,N_12991);
nor U13003 (N_13003,N_12986,N_12940);
xnor U13004 (N_13004,N_12888,N_12919);
xor U13005 (N_13005,N_12886,N_12895);
and U13006 (N_13006,N_12973,N_12877);
or U13007 (N_13007,N_12914,N_12974);
or U13008 (N_13008,N_12908,N_12988);
xnor U13009 (N_13009,N_12944,N_12875);
or U13010 (N_13010,N_12931,N_12906);
nand U13011 (N_13011,N_12976,N_12900);
nor U13012 (N_13012,N_12992,N_12916);
nand U13013 (N_13013,N_12987,N_12893);
xnor U13014 (N_13014,N_12977,N_12975);
nand U13015 (N_13015,N_12881,N_12962);
or U13016 (N_13016,N_12964,N_12955);
nand U13017 (N_13017,N_12938,N_12998);
and U13018 (N_13018,N_12928,N_12949);
xnor U13019 (N_13019,N_12915,N_12985);
nand U13020 (N_13020,N_12960,N_12958);
or U13021 (N_13021,N_12945,N_12910);
nor U13022 (N_13022,N_12954,N_12909);
nand U13023 (N_13023,N_12927,N_12924);
or U13024 (N_13024,N_12882,N_12980);
and U13025 (N_13025,N_12995,N_12929);
and U13026 (N_13026,N_12903,N_12942);
or U13027 (N_13027,N_12965,N_12901);
nand U13028 (N_13028,N_12936,N_12887);
nor U13029 (N_13029,N_12939,N_12951);
or U13030 (N_13030,N_12913,N_12898);
nand U13031 (N_13031,N_12993,N_12884);
and U13032 (N_13032,N_12918,N_12921);
nor U13033 (N_13033,N_12970,N_12922);
nand U13034 (N_13034,N_12885,N_12935);
or U13035 (N_13035,N_12943,N_12997);
nand U13036 (N_13036,N_12934,N_12996);
xnor U13037 (N_13037,N_12968,N_12981);
or U13038 (N_13038,N_12947,N_12982);
xor U13039 (N_13039,N_12999,N_12990);
or U13040 (N_13040,N_12983,N_12889);
and U13041 (N_13041,N_12946,N_12907);
or U13042 (N_13042,N_12880,N_12937);
nand U13043 (N_13043,N_12899,N_12894);
xor U13044 (N_13044,N_12890,N_12878);
nand U13045 (N_13045,N_12952,N_12930);
xor U13046 (N_13046,N_12926,N_12971);
nand U13047 (N_13047,N_12917,N_12963);
or U13048 (N_13048,N_12961,N_12933);
nor U13049 (N_13049,N_12905,N_12959);
nand U13050 (N_13050,N_12984,N_12879);
and U13051 (N_13051,N_12948,N_12972);
and U13052 (N_13052,N_12912,N_12932);
nand U13053 (N_13053,N_12904,N_12923);
nor U13054 (N_13054,N_12957,N_12891);
and U13055 (N_13055,N_12902,N_12989);
xor U13056 (N_13056,N_12967,N_12911);
nand U13057 (N_13057,N_12925,N_12941);
nand U13058 (N_13058,N_12920,N_12950);
or U13059 (N_13059,N_12897,N_12979);
and U13060 (N_13060,N_12978,N_12956);
and U13061 (N_13061,N_12883,N_12953);
nand U13062 (N_13062,N_12876,N_12962);
xor U13063 (N_13063,N_12994,N_12914);
or U13064 (N_13064,N_12922,N_12982);
or U13065 (N_13065,N_12929,N_12924);
and U13066 (N_13066,N_12910,N_12957);
or U13067 (N_13067,N_12923,N_12879);
or U13068 (N_13068,N_12991,N_12948);
nand U13069 (N_13069,N_12891,N_12921);
or U13070 (N_13070,N_12948,N_12945);
nor U13071 (N_13071,N_12932,N_12977);
nand U13072 (N_13072,N_12920,N_12961);
nand U13073 (N_13073,N_12916,N_12970);
nor U13074 (N_13074,N_12889,N_12928);
or U13075 (N_13075,N_12983,N_12950);
or U13076 (N_13076,N_12885,N_12978);
nor U13077 (N_13077,N_12939,N_12929);
xnor U13078 (N_13078,N_12917,N_12914);
nor U13079 (N_13079,N_12912,N_12879);
nand U13080 (N_13080,N_12882,N_12957);
nor U13081 (N_13081,N_12975,N_12943);
or U13082 (N_13082,N_12973,N_12983);
nand U13083 (N_13083,N_12974,N_12987);
and U13084 (N_13084,N_12991,N_12963);
or U13085 (N_13085,N_12961,N_12938);
and U13086 (N_13086,N_12957,N_12908);
or U13087 (N_13087,N_12926,N_12986);
and U13088 (N_13088,N_12972,N_12980);
nand U13089 (N_13089,N_12899,N_12910);
nor U13090 (N_13090,N_12877,N_12970);
and U13091 (N_13091,N_12953,N_12962);
and U13092 (N_13092,N_12953,N_12887);
or U13093 (N_13093,N_12920,N_12973);
nor U13094 (N_13094,N_12985,N_12913);
nor U13095 (N_13095,N_12945,N_12903);
nand U13096 (N_13096,N_12926,N_12991);
nor U13097 (N_13097,N_12940,N_12915);
and U13098 (N_13098,N_12969,N_12914);
and U13099 (N_13099,N_12959,N_12894);
nand U13100 (N_13100,N_12896,N_12934);
xnor U13101 (N_13101,N_12885,N_12944);
nand U13102 (N_13102,N_12908,N_12934);
nand U13103 (N_13103,N_12930,N_12971);
or U13104 (N_13104,N_12954,N_12928);
and U13105 (N_13105,N_12983,N_12906);
or U13106 (N_13106,N_12882,N_12903);
nand U13107 (N_13107,N_12968,N_12958);
or U13108 (N_13108,N_12948,N_12891);
and U13109 (N_13109,N_12996,N_12951);
and U13110 (N_13110,N_12983,N_12962);
nor U13111 (N_13111,N_12911,N_12934);
nand U13112 (N_13112,N_12891,N_12975);
xnor U13113 (N_13113,N_12904,N_12892);
or U13114 (N_13114,N_12876,N_12927);
and U13115 (N_13115,N_12929,N_12962);
and U13116 (N_13116,N_12971,N_12906);
or U13117 (N_13117,N_12979,N_12927);
nor U13118 (N_13118,N_12941,N_12964);
nand U13119 (N_13119,N_12954,N_12923);
xnor U13120 (N_13120,N_12977,N_12961);
and U13121 (N_13121,N_12900,N_12942);
or U13122 (N_13122,N_12938,N_12899);
nand U13123 (N_13123,N_12989,N_12993);
or U13124 (N_13124,N_12976,N_12968);
xnor U13125 (N_13125,N_13045,N_13066);
or U13126 (N_13126,N_13088,N_13112);
nor U13127 (N_13127,N_13059,N_13113);
nand U13128 (N_13128,N_13015,N_13019);
nand U13129 (N_13129,N_13091,N_13014);
and U13130 (N_13130,N_13024,N_13122);
xor U13131 (N_13131,N_13077,N_13079);
nand U13132 (N_13132,N_13038,N_13053);
or U13133 (N_13133,N_13050,N_13008);
nand U13134 (N_13134,N_13090,N_13076);
xor U13135 (N_13135,N_13099,N_13089);
nor U13136 (N_13136,N_13114,N_13057);
and U13137 (N_13137,N_13051,N_13106);
or U13138 (N_13138,N_13036,N_13069);
or U13139 (N_13139,N_13073,N_13103);
nand U13140 (N_13140,N_13060,N_13100);
xor U13141 (N_13141,N_13072,N_13124);
or U13142 (N_13142,N_13062,N_13006);
nor U13143 (N_13143,N_13041,N_13118);
nand U13144 (N_13144,N_13013,N_13116);
nand U13145 (N_13145,N_13095,N_13035);
nand U13146 (N_13146,N_13007,N_13009);
and U13147 (N_13147,N_13012,N_13052);
xnor U13148 (N_13148,N_13110,N_13056);
or U13149 (N_13149,N_13055,N_13028);
nor U13150 (N_13150,N_13084,N_13031);
and U13151 (N_13151,N_13064,N_13032);
nor U13152 (N_13152,N_13115,N_13104);
xor U13153 (N_13153,N_13033,N_13087);
nor U13154 (N_13154,N_13111,N_13107);
and U13155 (N_13155,N_13034,N_13094);
nor U13156 (N_13156,N_13044,N_13023);
or U13157 (N_13157,N_13080,N_13098);
nand U13158 (N_13158,N_13030,N_13119);
or U13159 (N_13159,N_13074,N_13049);
nor U13160 (N_13160,N_13071,N_13065);
or U13161 (N_13161,N_13000,N_13018);
and U13162 (N_13162,N_13054,N_13063);
and U13163 (N_13163,N_13026,N_13017);
nand U13164 (N_13164,N_13011,N_13085);
and U13165 (N_13165,N_13037,N_13003);
xnor U13166 (N_13166,N_13046,N_13042);
or U13167 (N_13167,N_13120,N_13086);
nand U13168 (N_13168,N_13097,N_13121);
nor U13169 (N_13169,N_13029,N_13082);
and U13170 (N_13170,N_13070,N_13016);
nand U13171 (N_13171,N_13002,N_13047);
xnor U13172 (N_13172,N_13078,N_13061);
nor U13173 (N_13173,N_13004,N_13048);
nor U13174 (N_13174,N_13096,N_13092);
or U13175 (N_13175,N_13068,N_13010);
nand U13176 (N_13176,N_13067,N_13001);
xnor U13177 (N_13177,N_13025,N_13093);
nand U13178 (N_13178,N_13108,N_13043);
nor U13179 (N_13179,N_13027,N_13040);
nand U13180 (N_13180,N_13123,N_13022);
nand U13181 (N_13181,N_13109,N_13039);
nand U13182 (N_13182,N_13102,N_13058);
and U13183 (N_13183,N_13105,N_13075);
nand U13184 (N_13184,N_13005,N_13117);
and U13185 (N_13185,N_13020,N_13083);
nand U13186 (N_13186,N_13101,N_13081);
or U13187 (N_13187,N_13021,N_13117);
nand U13188 (N_13188,N_13124,N_13030);
nor U13189 (N_13189,N_13057,N_13064);
nor U13190 (N_13190,N_13069,N_13119);
and U13191 (N_13191,N_13021,N_13085);
or U13192 (N_13192,N_13074,N_13064);
or U13193 (N_13193,N_13040,N_13045);
or U13194 (N_13194,N_13104,N_13004);
and U13195 (N_13195,N_13035,N_13036);
nand U13196 (N_13196,N_13123,N_13028);
and U13197 (N_13197,N_13122,N_13006);
nor U13198 (N_13198,N_13043,N_13007);
or U13199 (N_13199,N_13064,N_13029);
nand U13200 (N_13200,N_13076,N_13096);
nand U13201 (N_13201,N_13030,N_13019);
and U13202 (N_13202,N_13093,N_13019);
nand U13203 (N_13203,N_13080,N_13124);
and U13204 (N_13204,N_13077,N_13012);
or U13205 (N_13205,N_13105,N_13004);
and U13206 (N_13206,N_13069,N_13016);
nor U13207 (N_13207,N_13087,N_13122);
nand U13208 (N_13208,N_13005,N_13036);
and U13209 (N_13209,N_13074,N_13039);
xor U13210 (N_13210,N_13011,N_13114);
nand U13211 (N_13211,N_13072,N_13037);
nor U13212 (N_13212,N_13002,N_13113);
xor U13213 (N_13213,N_13120,N_13124);
or U13214 (N_13214,N_13058,N_13112);
nor U13215 (N_13215,N_13028,N_13104);
xor U13216 (N_13216,N_13065,N_13112);
or U13217 (N_13217,N_13040,N_13024);
nand U13218 (N_13218,N_13021,N_13095);
and U13219 (N_13219,N_13109,N_13102);
nand U13220 (N_13220,N_13068,N_13079);
nor U13221 (N_13221,N_13110,N_13102);
nor U13222 (N_13222,N_13026,N_13041);
or U13223 (N_13223,N_13048,N_13081);
nor U13224 (N_13224,N_13018,N_13059);
nor U13225 (N_13225,N_13049,N_13032);
nor U13226 (N_13226,N_13090,N_13070);
and U13227 (N_13227,N_13001,N_13071);
nand U13228 (N_13228,N_13011,N_13022);
xnor U13229 (N_13229,N_13002,N_13115);
nor U13230 (N_13230,N_13020,N_13055);
nor U13231 (N_13231,N_13034,N_13121);
or U13232 (N_13232,N_13032,N_13094);
or U13233 (N_13233,N_13087,N_13002);
nand U13234 (N_13234,N_13000,N_13086);
or U13235 (N_13235,N_13124,N_13077);
and U13236 (N_13236,N_13030,N_13099);
or U13237 (N_13237,N_13048,N_13006);
nand U13238 (N_13238,N_13028,N_13017);
nand U13239 (N_13239,N_13070,N_13068);
or U13240 (N_13240,N_13002,N_13093);
nand U13241 (N_13241,N_13025,N_13105);
nand U13242 (N_13242,N_13119,N_13061);
xor U13243 (N_13243,N_13044,N_13109);
and U13244 (N_13244,N_13104,N_13061);
nor U13245 (N_13245,N_13059,N_13095);
and U13246 (N_13246,N_13072,N_13019);
or U13247 (N_13247,N_13045,N_13054);
nor U13248 (N_13248,N_13077,N_13028);
and U13249 (N_13249,N_13092,N_13086);
nor U13250 (N_13250,N_13156,N_13188);
and U13251 (N_13251,N_13157,N_13205);
and U13252 (N_13252,N_13190,N_13246);
nand U13253 (N_13253,N_13221,N_13192);
nor U13254 (N_13254,N_13159,N_13141);
or U13255 (N_13255,N_13230,N_13220);
or U13256 (N_13256,N_13134,N_13152);
nor U13257 (N_13257,N_13158,N_13129);
nand U13258 (N_13258,N_13136,N_13216);
nor U13259 (N_13259,N_13199,N_13201);
and U13260 (N_13260,N_13154,N_13163);
xnor U13261 (N_13261,N_13182,N_13247);
nand U13262 (N_13262,N_13242,N_13166);
or U13263 (N_13263,N_13168,N_13193);
and U13264 (N_13264,N_13240,N_13236);
nand U13265 (N_13265,N_13126,N_13237);
nand U13266 (N_13266,N_13231,N_13146);
nor U13267 (N_13267,N_13248,N_13191);
nor U13268 (N_13268,N_13180,N_13172);
nand U13269 (N_13269,N_13208,N_13243);
and U13270 (N_13270,N_13198,N_13167);
nor U13271 (N_13271,N_13127,N_13171);
and U13272 (N_13272,N_13140,N_13249);
nor U13273 (N_13273,N_13227,N_13148);
or U13274 (N_13274,N_13133,N_13215);
nor U13275 (N_13275,N_13226,N_13209);
and U13276 (N_13276,N_13204,N_13229);
nor U13277 (N_13277,N_13149,N_13144);
xor U13278 (N_13278,N_13125,N_13153);
xor U13279 (N_13279,N_13225,N_13165);
nand U13280 (N_13280,N_13161,N_13181);
nor U13281 (N_13281,N_13241,N_13183);
nor U13282 (N_13282,N_13235,N_13160);
and U13283 (N_13283,N_13150,N_13164);
and U13284 (N_13284,N_13234,N_13155);
nand U13285 (N_13285,N_13194,N_13137);
and U13286 (N_13286,N_13186,N_13214);
nand U13287 (N_13287,N_13210,N_13173);
nand U13288 (N_13288,N_13218,N_13245);
and U13289 (N_13289,N_13200,N_13202);
xor U13290 (N_13290,N_13130,N_13207);
nand U13291 (N_13291,N_13211,N_13195);
nor U13292 (N_13292,N_13178,N_13228);
nand U13293 (N_13293,N_13176,N_13232);
nand U13294 (N_13294,N_13222,N_13169);
or U13295 (N_13295,N_13162,N_13187);
and U13296 (N_13296,N_13184,N_13239);
and U13297 (N_13297,N_13174,N_13170);
or U13298 (N_13298,N_13224,N_13142);
nor U13299 (N_13299,N_13145,N_13138);
or U13300 (N_13300,N_13128,N_13233);
nor U13301 (N_13301,N_13203,N_13132);
nor U13302 (N_13302,N_13177,N_13213);
and U13303 (N_13303,N_13206,N_13175);
or U13304 (N_13304,N_13135,N_13238);
nor U13305 (N_13305,N_13131,N_13179);
or U13306 (N_13306,N_13219,N_13139);
or U13307 (N_13307,N_13217,N_13196);
and U13308 (N_13308,N_13223,N_13151);
xor U13309 (N_13309,N_13197,N_13212);
nor U13310 (N_13310,N_13143,N_13244);
and U13311 (N_13311,N_13147,N_13185);
or U13312 (N_13312,N_13189,N_13179);
or U13313 (N_13313,N_13137,N_13241);
xnor U13314 (N_13314,N_13174,N_13202);
or U13315 (N_13315,N_13160,N_13233);
nor U13316 (N_13316,N_13188,N_13131);
nand U13317 (N_13317,N_13153,N_13204);
nor U13318 (N_13318,N_13231,N_13148);
nor U13319 (N_13319,N_13202,N_13162);
or U13320 (N_13320,N_13164,N_13204);
or U13321 (N_13321,N_13209,N_13190);
nand U13322 (N_13322,N_13208,N_13152);
nor U13323 (N_13323,N_13186,N_13196);
nand U13324 (N_13324,N_13126,N_13148);
and U13325 (N_13325,N_13126,N_13240);
nor U13326 (N_13326,N_13186,N_13133);
nor U13327 (N_13327,N_13212,N_13142);
or U13328 (N_13328,N_13226,N_13157);
xor U13329 (N_13329,N_13147,N_13132);
xor U13330 (N_13330,N_13235,N_13205);
and U13331 (N_13331,N_13162,N_13211);
nand U13332 (N_13332,N_13178,N_13174);
and U13333 (N_13333,N_13145,N_13239);
xor U13334 (N_13334,N_13190,N_13249);
or U13335 (N_13335,N_13195,N_13200);
and U13336 (N_13336,N_13212,N_13208);
or U13337 (N_13337,N_13154,N_13200);
and U13338 (N_13338,N_13181,N_13144);
nand U13339 (N_13339,N_13186,N_13135);
nor U13340 (N_13340,N_13194,N_13155);
and U13341 (N_13341,N_13246,N_13227);
or U13342 (N_13342,N_13229,N_13199);
nand U13343 (N_13343,N_13174,N_13193);
or U13344 (N_13344,N_13234,N_13196);
and U13345 (N_13345,N_13213,N_13223);
nand U13346 (N_13346,N_13239,N_13207);
nor U13347 (N_13347,N_13180,N_13186);
nand U13348 (N_13348,N_13181,N_13166);
nand U13349 (N_13349,N_13247,N_13150);
xor U13350 (N_13350,N_13247,N_13242);
nor U13351 (N_13351,N_13165,N_13171);
and U13352 (N_13352,N_13134,N_13163);
or U13353 (N_13353,N_13184,N_13154);
xor U13354 (N_13354,N_13156,N_13239);
nor U13355 (N_13355,N_13125,N_13245);
nand U13356 (N_13356,N_13176,N_13162);
or U13357 (N_13357,N_13181,N_13198);
or U13358 (N_13358,N_13237,N_13143);
and U13359 (N_13359,N_13170,N_13242);
and U13360 (N_13360,N_13194,N_13186);
or U13361 (N_13361,N_13185,N_13127);
and U13362 (N_13362,N_13153,N_13220);
or U13363 (N_13363,N_13217,N_13239);
or U13364 (N_13364,N_13180,N_13201);
and U13365 (N_13365,N_13172,N_13157);
or U13366 (N_13366,N_13193,N_13189);
or U13367 (N_13367,N_13136,N_13220);
xor U13368 (N_13368,N_13182,N_13213);
xnor U13369 (N_13369,N_13149,N_13228);
xor U13370 (N_13370,N_13175,N_13166);
xnor U13371 (N_13371,N_13233,N_13159);
nor U13372 (N_13372,N_13192,N_13234);
or U13373 (N_13373,N_13168,N_13196);
xor U13374 (N_13374,N_13236,N_13224);
and U13375 (N_13375,N_13286,N_13368);
nor U13376 (N_13376,N_13322,N_13315);
nor U13377 (N_13377,N_13280,N_13357);
nand U13378 (N_13378,N_13262,N_13270);
nand U13379 (N_13379,N_13316,N_13365);
nand U13380 (N_13380,N_13367,N_13308);
nand U13381 (N_13381,N_13320,N_13331);
nand U13382 (N_13382,N_13341,N_13272);
and U13383 (N_13383,N_13283,N_13345);
nand U13384 (N_13384,N_13285,N_13327);
nand U13385 (N_13385,N_13264,N_13259);
and U13386 (N_13386,N_13353,N_13348);
and U13387 (N_13387,N_13271,N_13266);
nor U13388 (N_13388,N_13276,N_13310);
or U13389 (N_13389,N_13332,N_13294);
nand U13390 (N_13390,N_13299,N_13343);
or U13391 (N_13391,N_13251,N_13347);
or U13392 (N_13392,N_13307,N_13319);
nand U13393 (N_13393,N_13328,N_13371);
nor U13394 (N_13394,N_13370,N_13363);
nand U13395 (N_13395,N_13335,N_13301);
xnor U13396 (N_13396,N_13290,N_13306);
or U13397 (N_13397,N_13333,N_13289);
xor U13398 (N_13398,N_13253,N_13252);
nor U13399 (N_13399,N_13336,N_13351);
and U13400 (N_13400,N_13324,N_13258);
or U13401 (N_13401,N_13267,N_13275);
xor U13402 (N_13402,N_13366,N_13274);
nand U13403 (N_13403,N_13288,N_13372);
or U13404 (N_13404,N_13250,N_13293);
xor U13405 (N_13405,N_13300,N_13263);
nand U13406 (N_13406,N_13282,N_13309);
and U13407 (N_13407,N_13321,N_13281);
nor U13408 (N_13408,N_13304,N_13361);
nand U13409 (N_13409,N_13305,N_13296);
xor U13410 (N_13410,N_13325,N_13342);
nor U13411 (N_13411,N_13323,N_13355);
or U13412 (N_13412,N_13273,N_13279);
nor U13413 (N_13413,N_13356,N_13314);
nand U13414 (N_13414,N_13256,N_13261);
or U13415 (N_13415,N_13268,N_13265);
nor U13416 (N_13416,N_13297,N_13362);
nor U13417 (N_13417,N_13330,N_13364);
or U13418 (N_13418,N_13302,N_13360);
nand U13419 (N_13419,N_13313,N_13350);
nand U13420 (N_13420,N_13255,N_13374);
nand U13421 (N_13421,N_13334,N_13295);
nor U13422 (N_13422,N_13269,N_13287);
or U13423 (N_13423,N_13292,N_13284);
nand U13424 (N_13424,N_13329,N_13278);
nor U13425 (N_13425,N_13277,N_13318);
xnor U13426 (N_13426,N_13358,N_13337);
and U13427 (N_13427,N_13298,N_13312);
nand U13428 (N_13428,N_13344,N_13291);
or U13429 (N_13429,N_13257,N_13338);
nor U13430 (N_13430,N_13349,N_13311);
and U13431 (N_13431,N_13373,N_13346);
and U13432 (N_13432,N_13354,N_13339);
and U13433 (N_13433,N_13303,N_13352);
and U13434 (N_13434,N_13340,N_13369);
or U13435 (N_13435,N_13317,N_13260);
and U13436 (N_13436,N_13359,N_13326);
or U13437 (N_13437,N_13254,N_13315);
and U13438 (N_13438,N_13319,N_13365);
or U13439 (N_13439,N_13364,N_13251);
and U13440 (N_13440,N_13343,N_13270);
or U13441 (N_13441,N_13268,N_13297);
and U13442 (N_13442,N_13352,N_13272);
xnor U13443 (N_13443,N_13324,N_13266);
or U13444 (N_13444,N_13374,N_13295);
nor U13445 (N_13445,N_13327,N_13324);
nand U13446 (N_13446,N_13335,N_13313);
nand U13447 (N_13447,N_13336,N_13277);
and U13448 (N_13448,N_13292,N_13351);
and U13449 (N_13449,N_13347,N_13300);
or U13450 (N_13450,N_13339,N_13277);
or U13451 (N_13451,N_13360,N_13260);
nor U13452 (N_13452,N_13291,N_13349);
nor U13453 (N_13453,N_13347,N_13331);
nor U13454 (N_13454,N_13333,N_13290);
nor U13455 (N_13455,N_13289,N_13263);
xor U13456 (N_13456,N_13264,N_13336);
nand U13457 (N_13457,N_13316,N_13278);
and U13458 (N_13458,N_13362,N_13353);
nor U13459 (N_13459,N_13305,N_13338);
and U13460 (N_13460,N_13360,N_13371);
and U13461 (N_13461,N_13262,N_13365);
or U13462 (N_13462,N_13352,N_13274);
xnor U13463 (N_13463,N_13291,N_13356);
nand U13464 (N_13464,N_13278,N_13305);
nor U13465 (N_13465,N_13352,N_13320);
nand U13466 (N_13466,N_13283,N_13274);
nand U13467 (N_13467,N_13374,N_13358);
and U13468 (N_13468,N_13370,N_13265);
or U13469 (N_13469,N_13285,N_13282);
and U13470 (N_13470,N_13340,N_13320);
or U13471 (N_13471,N_13342,N_13308);
and U13472 (N_13472,N_13321,N_13324);
or U13473 (N_13473,N_13254,N_13352);
and U13474 (N_13474,N_13252,N_13362);
xor U13475 (N_13475,N_13293,N_13254);
xnor U13476 (N_13476,N_13259,N_13343);
nand U13477 (N_13477,N_13280,N_13366);
or U13478 (N_13478,N_13311,N_13251);
nor U13479 (N_13479,N_13267,N_13326);
and U13480 (N_13480,N_13261,N_13311);
or U13481 (N_13481,N_13268,N_13345);
xor U13482 (N_13482,N_13336,N_13327);
and U13483 (N_13483,N_13314,N_13283);
nand U13484 (N_13484,N_13329,N_13330);
and U13485 (N_13485,N_13302,N_13336);
nor U13486 (N_13486,N_13270,N_13259);
or U13487 (N_13487,N_13269,N_13285);
or U13488 (N_13488,N_13318,N_13257);
nand U13489 (N_13489,N_13335,N_13348);
nand U13490 (N_13490,N_13301,N_13263);
and U13491 (N_13491,N_13340,N_13307);
nor U13492 (N_13492,N_13319,N_13333);
and U13493 (N_13493,N_13264,N_13335);
nor U13494 (N_13494,N_13308,N_13302);
nand U13495 (N_13495,N_13278,N_13373);
nand U13496 (N_13496,N_13342,N_13265);
nand U13497 (N_13497,N_13302,N_13250);
nor U13498 (N_13498,N_13302,N_13283);
nor U13499 (N_13499,N_13351,N_13302);
or U13500 (N_13500,N_13398,N_13466);
or U13501 (N_13501,N_13432,N_13392);
or U13502 (N_13502,N_13409,N_13449);
nand U13503 (N_13503,N_13375,N_13403);
and U13504 (N_13504,N_13378,N_13470);
and U13505 (N_13505,N_13483,N_13425);
nand U13506 (N_13506,N_13438,N_13469);
and U13507 (N_13507,N_13499,N_13455);
nor U13508 (N_13508,N_13411,N_13468);
xnor U13509 (N_13509,N_13384,N_13421);
or U13510 (N_13510,N_13493,N_13451);
and U13511 (N_13511,N_13498,N_13408);
and U13512 (N_13512,N_13400,N_13404);
nand U13513 (N_13513,N_13423,N_13475);
nand U13514 (N_13514,N_13387,N_13386);
or U13515 (N_13515,N_13389,N_13485);
and U13516 (N_13516,N_13431,N_13406);
or U13517 (N_13517,N_13477,N_13418);
or U13518 (N_13518,N_13481,N_13494);
or U13519 (N_13519,N_13454,N_13401);
and U13520 (N_13520,N_13445,N_13462);
or U13521 (N_13521,N_13480,N_13473);
and U13522 (N_13522,N_13453,N_13441);
xor U13523 (N_13523,N_13381,N_13417);
xnor U13524 (N_13524,N_13490,N_13376);
nand U13525 (N_13525,N_13399,N_13457);
or U13526 (N_13526,N_13491,N_13434);
nor U13527 (N_13527,N_13396,N_13393);
xor U13528 (N_13528,N_13489,N_13492);
nor U13529 (N_13529,N_13428,N_13420);
and U13530 (N_13530,N_13419,N_13383);
and U13531 (N_13531,N_13458,N_13443);
or U13532 (N_13532,N_13380,N_13474);
or U13533 (N_13533,N_13397,N_13437);
nand U13534 (N_13534,N_13479,N_13388);
nand U13535 (N_13535,N_13382,N_13448);
nor U13536 (N_13536,N_13433,N_13414);
xor U13537 (N_13537,N_13460,N_13467);
and U13538 (N_13538,N_13461,N_13436);
nor U13539 (N_13539,N_13395,N_13472);
and U13540 (N_13540,N_13464,N_13426);
or U13541 (N_13541,N_13405,N_13478);
and U13542 (N_13542,N_13444,N_13412);
or U13543 (N_13543,N_13463,N_13422);
or U13544 (N_13544,N_13410,N_13450);
and U13545 (N_13545,N_13391,N_13402);
nand U13546 (N_13546,N_13390,N_13476);
xor U13547 (N_13547,N_13484,N_13413);
and U13548 (N_13548,N_13459,N_13447);
nand U13549 (N_13549,N_13430,N_13488);
and U13550 (N_13550,N_13471,N_13452);
xnor U13551 (N_13551,N_13394,N_13495);
and U13552 (N_13552,N_13456,N_13487);
or U13553 (N_13553,N_13429,N_13465);
nor U13554 (N_13554,N_13486,N_13497);
and U13555 (N_13555,N_13446,N_13439);
or U13556 (N_13556,N_13427,N_13424);
and U13557 (N_13557,N_13482,N_13379);
nand U13558 (N_13558,N_13407,N_13377);
nor U13559 (N_13559,N_13385,N_13416);
nor U13560 (N_13560,N_13440,N_13415);
and U13561 (N_13561,N_13442,N_13496);
or U13562 (N_13562,N_13435,N_13430);
nor U13563 (N_13563,N_13497,N_13402);
nor U13564 (N_13564,N_13462,N_13416);
and U13565 (N_13565,N_13437,N_13380);
nand U13566 (N_13566,N_13429,N_13419);
nand U13567 (N_13567,N_13454,N_13476);
nor U13568 (N_13568,N_13471,N_13473);
or U13569 (N_13569,N_13469,N_13427);
xnor U13570 (N_13570,N_13378,N_13408);
nand U13571 (N_13571,N_13476,N_13473);
nand U13572 (N_13572,N_13443,N_13379);
or U13573 (N_13573,N_13494,N_13489);
or U13574 (N_13574,N_13431,N_13462);
nor U13575 (N_13575,N_13407,N_13391);
nor U13576 (N_13576,N_13479,N_13422);
xor U13577 (N_13577,N_13376,N_13391);
nor U13578 (N_13578,N_13405,N_13451);
or U13579 (N_13579,N_13447,N_13440);
or U13580 (N_13580,N_13378,N_13456);
and U13581 (N_13581,N_13396,N_13377);
xor U13582 (N_13582,N_13479,N_13442);
or U13583 (N_13583,N_13493,N_13401);
or U13584 (N_13584,N_13447,N_13462);
nand U13585 (N_13585,N_13437,N_13426);
nand U13586 (N_13586,N_13445,N_13439);
or U13587 (N_13587,N_13376,N_13452);
xor U13588 (N_13588,N_13494,N_13413);
nor U13589 (N_13589,N_13472,N_13425);
or U13590 (N_13590,N_13486,N_13428);
nand U13591 (N_13591,N_13378,N_13413);
nand U13592 (N_13592,N_13408,N_13454);
and U13593 (N_13593,N_13411,N_13447);
or U13594 (N_13594,N_13490,N_13497);
and U13595 (N_13595,N_13497,N_13463);
nand U13596 (N_13596,N_13434,N_13414);
and U13597 (N_13597,N_13475,N_13470);
nor U13598 (N_13598,N_13447,N_13420);
and U13599 (N_13599,N_13387,N_13379);
nand U13600 (N_13600,N_13399,N_13423);
and U13601 (N_13601,N_13380,N_13425);
nand U13602 (N_13602,N_13390,N_13380);
and U13603 (N_13603,N_13429,N_13409);
and U13604 (N_13604,N_13468,N_13464);
or U13605 (N_13605,N_13425,N_13463);
or U13606 (N_13606,N_13460,N_13409);
xnor U13607 (N_13607,N_13486,N_13401);
nand U13608 (N_13608,N_13410,N_13417);
and U13609 (N_13609,N_13479,N_13444);
and U13610 (N_13610,N_13480,N_13472);
xnor U13611 (N_13611,N_13494,N_13469);
nor U13612 (N_13612,N_13470,N_13432);
and U13613 (N_13613,N_13433,N_13390);
or U13614 (N_13614,N_13393,N_13485);
or U13615 (N_13615,N_13458,N_13415);
nor U13616 (N_13616,N_13482,N_13381);
nor U13617 (N_13617,N_13406,N_13381);
and U13618 (N_13618,N_13407,N_13466);
or U13619 (N_13619,N_13390,N_13464);
xor U13620 (N_13620,N_13411,N_13459);
nand U13621 (N_13621,N_13390,N_13430);
nand U13622 (N_13622,N_13493,N_13458);
or U13623 (N_13623,N_13427,N_13492);
or U13624 (N_13624,N_13405,N_13470);
xnor U13625 (N_13625,N_13597,N_13562);
or U13626 (N_13626,N_13532,N_13622);
and U13627 (N_13627,N_13584,N_13550);
nand U13628 (N_13628,N_13580,N_13610);
nand U13629 (N_13629,N_13567,N_13524);
nand U13630 (N_13630,N_13545,N_13611);
and U13631 (N_13631,N_13557,N_13608);
nor U13632 (N_13632,N_13559,N_13548);
and U13633 (N_13633,N_13506,N_13566);
or U13634 (N_13634,N_13589,N_13521);
and U13635 (N_13635,N_13515,N_13501);
nor U13636 (N_13636,N_13514,N_13538);
or U13637 (N_13637,N_13573,N_13549);
and U13638 (N_13638,N_13556,N_13587);
nand U13639 (N_13639,N_13537,N_13596);
xnor U13640 (N_13640,N_13565,N_13583);
or U13641 (N_13641,N_13551,N_13531);
xnor U13642 (N_13642,N_13623,N_13560);
and U13643 (N_13643,N_13511,N_13547);
nor U13644 (N_13644,N_13602,N_13525);
nor U13645 (N_13645,N_13503,N_13618);
and U13646 (N_13646,N_13609,N_13542);
and U13647 (N_13647,N_13568,N_13605);
and U13648 (N_13648,N_13510,N_13512);
nor U13649 (N_13649,N_13607,N_13535);
nor U13650 (N_13650,N_13561,N_13523);
xnor U13651 (N_13651,N_13553,N_13571);
or U13652 (N_13652,N_13533,N_13544);
and U13653 (N_13653,N_13513,N_13519);
and U13654 (N_13654,N_13601,N_13613);
or U13655 (N_13655,N_13590,N_13575);
xnor U13656 (N_13656,N_13517,N_13558);
nand U13657 (N_13657,N_13586,N_13563);
or U13658 (N_13658,N_13620,N_13619);
or U13659 (N_13659,N_13509,N_13522);
or U13660 (N_13660,N_13536,N_13520);
or U13661 (N_13661,N_13529,N_13572);
or U13662 (N_13662,N_13615,N_13508);
xnor U13663 (N_13663,N_13616,N_13530);
nand U13664 (N_13664,N_13526,N_13500);
nand U13665 (N_13665,N_13541,N_13574);
and U13666 (N_13666,N_13600,N_13624);
or U13667 (N_13667,N_13516,N_13576);
or U13668 (N_13668,N_13579,N_13504);
nor U13669 (N_13669,N_13578,N_13505);
nor U13670 (N_13670,N_13527,N_13507);
nor U13671 (N_13671,N_13569,N_13588);
or U13672 (N_13672,N_13604,N_13552);
nand U13673 (N_13673,N_13534,N_13621);
nor U13674 (N_13674,N_13592,N_13540);
xor U13675 (N_13675,N_13606,N_13570);
and U13676 (N_13676,N_13502,N_13581);
and U13677 (N_13677,N_13598,N_13614);
nand U13678 (N_13678,N_13518,N_13582);
nand U13679 (N_13679,N_13543,N_13546);
or U13680 (N_13680,N_13593,N_13555);
nand U13681 (N_13681,N_13539,N_13617);
nand U13682 (N_13682,N_13528,N_13564);
xor U13683 (N_13683,N_13603,N_13585);
nor U13684 (N_13684,N_13612,N_13554);
nor U13685 (N_13685,N_13595,N_13594);
and U13686 (N_13686,N_13591,N_13599);
nor U13687 (N_13687,N_13577,N_13544);
or U13688 (N_13688,N_13593,N_13590);
and U13689 (N_13689,N_13624,N_13538);
or U13690 (N_13690,N_13589,N_13514);
or U13691 (N_13691,N_13530,N_13525);
nand U13692 (N_13692,N_13591,N_13529);
nor U13693 (N_13693,N_13605,N_13598);
nand U13694 (N_13694,N_13587,N_13511);
nand U13695 (N_13695,N_13585,N_13582);
or U13696 (N_13696,N_13568,N_13582);
nand U13697 (N_13697,N_13569,N_13531);
and U13698 (N_13698,N_13615,N_13585);
nor U13699 (N_13699,N_13527,N_13554);
xnor U13700 (N_13700,N_13603,N_13572);
nand U13701 (N_13701,N_13602,N_13565);
nor U13702 (N_13702,N_13588,N_13519);
and U13703 (N_13703,N_13588,N_13587);
and U13704 (N_13704,N_13525,N_13555);
nand U13705 (N_13705,N_13519,N_13547);
and U13706 (N_13706,N_13554,N_13538);
nand U13707 (N_13707,N_13620,N_13609);
nand U13708 (N_13708,N_13505,N_13520);
and U13709 (N_13709,N_13620,N_13582);
nand U13710 (N_13710,N_13503,N_13541);
or U13711 (N_13711,N_13530,N_13619);
nor U13712 (N_13712,N_13574,N_13544);
nand U13713 (N_13713,N_13618,N_13512);
and U13714 (N_13714,N_13556,N_13607);
nand U13715 (N_13715,N_13580,N_13506);
and U13716 (N_13716,N_13566,N_13569);
xnor U13717 (N_13717,N_13546,N_13612);
nand U13718 (N_13718,N_13525,N_13541);
nand U13719 (N_13719,N_13535,N_13553);
or U13720 (N_13720,N_13529,N_13609);
nand U13721 (N_13721,N_13553,N_13540);
nand U13722 (N_13722,N_13621,N_13591);
nor U13723 (N_13723,N_13593,N_13584);
nand U13724 (N_13724,N_13536,N_13575);
and U13725 (N_13725,N_13521,N_13544);
xnor U13726 (N_13726,N_13613,N_13503);
nor U13727 (N_13727,N_13506,N_13619);
or U13728 (N_13728,N_13598,N_13591);
nand U13729 (N_13729,N_13533,N_13546);
nor U13730 (N_13730,N_13554,N_13562);
nor U13731 (N_13731,N_13505,N_13605);
nand U13732 (N_13732,N_13617,N_13558);
nand U13733 (N_13733,N_13582,N_13614);
nor U13734 (N_13734,N_13504,N_13563);
or U13735 (N_13735,N_13613,N_13508);
nor U13736 (N_13736,N_13556,N_13559);
nor U13737 (N_13737,N_13521,N_13585);
xnor U13738 (N_13738,N_13509,N_13556);
and U13739 (N_13739,N_13568,N_13580);
and U13740 (N_13740,N_13571,N_13547);
or U13741 (N_13741,N_13531,N_13580);
or U13742 (N_13742,N_13576,N_13573);
and U13743 (N_13743,N_13567,N_13589);
or U13744 (N_13744,N_13505,N_13543);
or U13745 (N_13745,N_13565,N_13576);
or U13746 (N_13746,N_13589,N_13591);
nor U13747 (N_13747,N_13596,N_13501);
nor U13748 (N_13748,N_13589,N_13593);
and U13749 (N_13749,N_13512,N_13565);
nand U13750 (N_13750,N_13648,N_13715);
nand U13751 (N_13751,N_13744,N_13655);
xnor U13752 (N_13752,N_13743,N_13675);
xnor U13753 (N_13753,N_13651,N_13630);
nor U13754 (N_13754,N_13684,N_13678);
xor U13755 (N_13755,N_13668,N_13665);
or U13756 (N_13756,N_13736,N_13674);
xor U13757 (N_13757,N_13720,N_13659);
or U13758 (N_13758,N_13693,N_13628);
or U13759 (N_13759,N_13647,N_13725);
and U13760 (N_13760,N_13731,N_13676);
and U13761 (N_13761,N_13639,N_13726);
or U13762 (N_13762,N_13664,N_13702);
or U13763 (N_13763,N_13633,N_13735);
xor U13764 (N_13764,N_13646,N_13727);
nor U13765 (N_13765,N_13708,N_13716);
nand U13766 (N_13766,N_13696,N_13687);
nand U13767 (N_13767,N_13714,N_13653);
xor U13768 (N_13768,N_13719,N_13748);
or U13769 (N_13769,N_13652,N_13667);
and U13770 (N_13770,N_13732,N_13711);
nand U13771 (N_13771,N_13683,N_13643);
nor U13772 (N_13772,N_13697,N_13631);
and U13773 (N_13773,N_13635,N_13691);
nand U13774 (N_13774,N_13728,N_13707);
nand U13775 (N_13775,N_13699,N_13689);
xnor U13776 (N_13776,N_13679,N_13723);
and U13777 (N_13777,N_13681,N_13644);
nand U13778 (N_13778,N_13645,N_13680);
nand U13779 (N_13779,N_13749,N_13673);
nand U13780 (N_13780,N_13705,N_13671);
nor U13781 (N_13781,N_13729,N_13704);
nor U13782 (N_13782,N_13656,N_13740);
and U13783 (N_13783,N_13654,N_13746);
nand U13784 (N_13784,N_13692,N_13739);
or U13785 (N_13785,N_13730,N_13661);
nor U13786 (N_13786,N_13698,N_13706);
and U13787 (N_13787,N_13636,N_13741);
nand U13788 (N_13788,N_13629,N_13733);
nor U13789 (N_13789,N_13627,N_13747);
nor U13790 (N_13790,N_13721,N_13717);
xnor U13791 (N_13791,N_13626,N_13637);
and U13792 (N_13792,N_13742,N_13738);
and U13793 (N_13793,N_13657,N_13724);
nand U13794 (N_13794,N_13718,N_13701);
or U13795 (N_13795,N_13695,N_13722);
nor U13796 (N_13796,N_13663,N_13658);
and U13797 (N_13797,N_13666,N_13682);
nor U13798 (N_13798,N_13734,N_13625);
xor U13799 (N_13799,N_13677,N_13690);
nor U13800 (N_13800,N_13670,N_13641);
xnor U13801 (N_13801,N_13703,N_13694);
nor U13802 (N_13802,N_13660,N_13686);
nor U13803 (N_13803,N_13745,N_13634);
nor U13804 (N_13804,N_13638,N_13685);
or U13805 (N_13805,N_13710,N_13672);
nor U13806 (N_13806,N_13713,N_13632);
nor U13807 (N_13807,N_13662,N_13640);
nor U13808 (N_13808,N_13709,N_13650);
or U13809 (N_13809,N_13642,N_13649);
nand U13810 (N_13810,N_13700,N_13669);
nor U13811 (N_13811,N_13712,N_13688);
and U13812 (N_13812,N_13737,N_13627);
xnor U13813 (N_13813,N_13721,N_13635);
and U13814 (N_13814,N_13715,N_13679);
or U13815 (N_13815,N_13685,N_13719);
and U13816 (N_13816,N_13685,N_13656);
or U13817 (N_13817,N_13713,N_13697);
nand U13818 (N_13818,N_13705,N_13735);
nand U13819 (N_13819,N_13657,N_13660);
and U13820 (N_13820,N_13748,N_13664);
nand U13821 (N_13821,N_13700,N_13626);
nand U13822 (N_13822,N_13709,N_13711);
nor U13823 (N_13823,N_13739,N_13646);
nand U13824 (N_13824,N_13649,N_13625);
and U13825 (N_13825,N_13678,N_13677);
nor U13826 (N_13826,N_13710,N_13711);
nand U13827 (N_13827,N_13641,N_13729);
xor U13828 (N_13828,N_13677,N_13700);
nand U13829 (N_13829,N_13691,N_13633);
xnor U13830 (N_13830,N_13664,N_13719);
nand U13831 (N_13831,N_13736,N_13632);
nor U13832 (N_13832,N_13668,N_13726);
nand U13833 (N_13833,N_13677,N_13704);
and U13834 (N_13834,N_13637,N_13675);
or U13835 (N_13835,N_13641,N_13744);
or U13836 (N_13836,N_13690,N_13649);
nor U13837 (N_13837,N_13719,N_13747);
or U13838 (N_13838,N_13657,N_13737);
or U13839 (N_13839,N_13662,N_13730);
or U13840 (N_13840,N_13675,N_13739);
and U13841 (N_13841,N_13681,N_13692);
nor U13842 (N_13842,N_13745,N_13708);
nor U13843 (N_13843,N_13664,N_13626);
xor U13844 (N_13844,N_13684,N_13743);
or U13845 (N_13845,N_13689,N_13656);
or U13846 (N_13846,N_13664,N_13647);
nand U13847 (N_13847,N_13649,N_13661);
xor U13848 (N_13848,N_13689,N_13736);
nand U13849 (N_13849,N_13712,N_13640);
nor U13850 (N_13850,N_13702,N_13626);
nand U13851 (N_13851,N_13626,N_13672);
or U13852 (N_13852,N_13732,N_13697);
nand U13853 (N_13853,N_13653,N_13718);
nand U13854 (N_13854,N_13697,N_13626);
xnor U13855 (N_13855,N_13650,N_13688);
and U13856 (N_13856,N_13715,N_13642);
and U13857 (N_13857,N_13724,N_13675);
nand U13858 (N_13858,N_13663,N_13693);
xnor U13859 (N_13859,N_13679,N_13659);
nor U13860 (N_13860,N_13685,N_13710);
or U13861 (N_13861,N_13697,N_13730);
nand U13862 (N_13862,N_13720,N_13691);
nand U13863 (N_13863,N_13686,N_13736);
xnor U13864 (N_13864,N_13633,N_13625);
or U13865 (N_13865,N_13670,N_13677);
nand U13866 (N_13866,N_13631,N_13647);
nor U13867 (N_13867,N_13700,N_13730);
xnor U13868 (N_13868,N_13673,N_13722);
and U13869 (N_13869,N_13628,N_13749);
or U13870 (N_13870,N_13698,N_13746);
xnor U13871 (N_13871,N_13647,N_13637);
nor U13872 (N_13872,N_13674,N_13726);
nor U13873 (N_13873,N_13724,N_13648);
xnor U13874 (N_13874,N_13735,N_13728);
and U13875 (N_13875,N_13816,N_13813);
or U13876 (N_13876,N_13776,N_13854);
nor U13877 (N_13877,N_13822,N_13836);
nor U13878 (N_13878,N_13852,N_13859);
xor U13879 (N_13879,N_13796,N_13824);
and U13880 (N_13880,N_13857,N_13868);
xor U13881 (N_13881,N_13787,N_13837);
or U13882 (N_13882,N_13825,N_13773);
and U13883 (N_13883,N_13811,N_13841);
nor U13884 (N_13884,N_13842,N_13874);
nand U13885 (N_13885,N_13761,N_13869);
nand U13886 (N_13886,N_13834,N_13871);
xor U13887 (N_13887,N_13753,N_13750);
xor U13888 (N_13888,N_13872,N_13778);
nand U13889 (N_13889,N_13823,N_13829);
and U13890 (N_13890,N_13850,N_13858);
nand U13891 (N_13891,N_13832,N_13848);
and U13892 (N_13892,N_13846,N_13751);
and U13893 (N_13893,N_13767,N_13774);
nor U13894 (N_13894,N_13768,N_13769);
nand U13895 (N_13895,N_13764,N_13840);
nand U13896 (N_13896,N_13808,N_13772);
nand U13897 (N_13897,N_13843,N_13798);
and U13898 (N_13898,N_13828,N_13788);
nor U13899 (N_13899,N_13819,N_13826);
xor U13900 (N_13900,N_13851,N_13756);
nor U13901 (N_13901,N_13831,N_13783);
or U13902 (N_13902,N_13835,N_13805);
nor U13903 (N_13903,N_13817,N_13771);
xnor U13904 (N_13904,N_13833,N_13814);
nand U13905 (N_13905,N_13847,N_13807);
and U13906 (N_13906,N_13866,N_13789);
xor U13907 (N_13907,N_13856,N_13804);
and U13908 (N_13908,N_13797,N_13755);
and U13909 (N_13909,N_13766,N_13827);
nor U13910 (N_13910,N_13795,N_13777);
and U13911 (N_13911,N_13862,N_13820);
or U13912 (N_13912,N_13792,N_13867);
xor U13913 (N_13913,N_13861,N_13803);
and U13914 (N_13914,N_13765,N_13809);
nor U13915 (N_13915,N_13784,N_13810);
xnor U13916 (N_13916,N_13806,N_13863);
nor U13917 (N_13917,N_13791,N_13865);
and U13918 (N_13918,N_13752,N_13821);
and U13919 (N_13919,N_13802,N_13782);
nand U13920 (N_13920,N_13754,N_13758);
and U13921 (N_13921,N_13794,N_13785);
nor U13922 (N_13922,N_13775,N_13799);
or U13923 (N_13923,N_13779,N_13757);
or U13924 (N_13924,N_13786,N_13873);
nor U13925 (N_13925,N_13853,N_13830);
nand U13926 (N_13926,N_13759,N_13793);
xnor U13927 (N_13927,N_13763,N_13849);
nand U13928 (N_13928,N_13801,N_13762);
or U13929 (N_13929,N_13812,N_13860);
or U13930 (N_13930,N_13800,N_13770);
or U13931 (N_13931,N_13844,N_13790);
and U13932 (N_13932,N_13838,N_13839);
or U13933 (N_13933,N_13781,N_13864);
and U13934 (N_13934,N_13818,N_13870);
nor U13935 (N_13935,N_13760,N_13855);
or U13936 (N_13936,N_13780,N_13845);
nand U13937 (N_13937,N_13815,N_13842);
nand U13938 (N_13938,N_13788,N_13863);
xor U13939 (N_13939,N_13856,N_13758);
and U13940 (N_13940,N_13822,N_13771);
nor U13941 (N_13941,N_13807,N_13757);
or U13942 (N_13942,N_13823,N_13771);
and U13943 (N_13943,N_13784,N_13795);
nand U13944 (N_13944,N_13851,N_13762);
nor U13945 (N_13945,N_13854,N_13783);
or U13946 (N_13946,N_13789,N_13750);
nor U13947 (N_13947,N_13872,N_13811);
nor U13948 (N_13948,N_13791,N_13817);
nand U13949 (N_13949,N_13826,N_13789);
or U13950 (N_13950,N_13778,N_13809);
xnor U13951 (N_13951,N_13785,N_13806);
nand U13952 (N_13952,N_13855,N_13840);
nor U13953 (N_13953,N_13830,N_13813);
or U13954 (N_13954,N_13822,N_13802);
and U13955 (N_13955,N_13843,N_13803);
nand U13956 (N_13956,N_13767,N_13750);
xnor U13957 (N_13957,N_13819,N_13802);
nor U13958 (N_13958,N_13796,N_13769);
and U13959 (N_13959,N_13779,N_13776);
xor U13960 (N_13960,N_13776,N_13783);
and U13961 (N_13961,N_13753,N_13854);
or U13962 (N_13962,N_13759,N_13831);
nand U13963 (N_13963,N_13813,N_13867);
and U13964 (N_13964,N_13752,N_13784);
xnor U13965 (N_13965,N_13843,N_13870);
nor U13966 (N_13966,N_13780,N_13859);
nor U13967 (N_13967,N_13846,N_13849);
nand U13968 (N_13968,N_13854,N_13795);
or U13969 (N_13969,N_13874,N_13790);
or U13970 (N_13970,N_13790,N_13783);
or U13971 (N_13971,N_13808,N_13859);
nand U13972 (N_13972,N_13850,N_13784);
and U13973 (N_13973,N_13858,N_13814);
nand U13974 (N_13974,N_13871,N_13797);
and U13975 (N_13975,N_13809,N_13818);
nand U13976 (N_13976,N_13765,N_13805);
or U13977 (N_13977,N_13821,N_13814);
nand U13978 (N_13978,N_13785,N_13783);
nand U13979 (N_13979,N_13804,N_13754);
and U13980 (N_13980,N_13829,N_13763);
nand U13981 (N_13981,N_13775,N_13793);
or U13982 (N_13982,N_13834,N_13830);
nand U13983 (N_13983,N_13841,N_13752);
and U13984 (N_13984,N_13832,N_13793);
and U13985 (N_13985,N_13750,N_13804);
nor U13986 (N_13986,N_13829,N_13837);
or U13987 (N_13987,N_13855,N_13826);
xor U13988 (N_13988,N_13786,N_13773);
nand U13989 (N_13989,N_13802,N_13776);
nor U13990 (N_13990,N_13761,N_13815);
or U13991 (N_13991,N_13765,N_13755);
nand U13992 (N_13992,N_13804,N_13768);
or U13993 (N_13993,N_13797,N_13823);
nor U13994 (N_13994,N_13821,N_13794);
nand U13995 (N_13995,N_13771,N_13848);
nor U13996 (N_13996,N_13820,N_13858);
xor U13997 (N_13997,N_13780,N_13796);
or U13998 (N_13998,N_13766,N_13825);
nand U13999 (N_13999,N_13836,N_13778);
or U14000 (N_14000,N_13927,N_13939);
nand U14001 (N_14001,N_13890,N_13967);
nor U14002 (N_14002,N_13973,N_13885);
or U14003 (N_14003,N_13914,N_13907);
and U14004 (N_14004,N_13974,N_13984);
or U14005 (N_14005,N_13883,N_13954);
xnor U14006 (N_14006,N_13886,N_13986);
and U14007 (N_14007,N_13922,N_13978);
or U14008 (N_14008,N_13906,N_13944);
and U14009 (N_14009,N_13992,N_13930);
or U14010 (N_14010,N_13904,N_13879);
nand U14011 (N_14011,N_13937,N_13892);
xor U14012 (N_14012,N_13915,N_13898);
nor U14013 (N_14013,N_13989,N_13962);
or U14014 (N_14014,N_13920,N_13982);
nand U14015 (N_14015,N_13884,N_13887);
nand U14016 (N_14016,N_13932,N_13903);
nand U14017 (N_14017,N_13924,N_13919);
nor U14018 (N_14018,N_13899,N_13936);
or U14019 (N_14019,N_13999,N_13947);
nand U14020 (N_14020,N_13926,N_13900);
xor U14021 (N_14021,N_13923,N_13993);
nand U14022 (N_14022,N_13979,N_13935);
nor U14023 (N_14023,N_13975,N_13961);
and U14024 (N_14024,N_13888,N_13971);
nor U14025 (N_14025,N_13946,N_13902);
nand U14026 (N_14026,N_13988,N_13896);
nor U14027 (N_14027,N_13951,N_13889);
nand U14028 (N_14028,N_13983,N_13997);
nor U14029 (N_14029,N_13916,N_13928);
and U14030 (N_14030,N_13945,N_13948);
or U14031 (N_14031,N_13880,N_13878);
nand U14032 (N_14032,N_13912,N_13969);
and U14033 (N_14033,N_13980,N_13933);
nand U14034 (N_14034,N_13970,N_13996);
xor U14035 (N_14035,N_13958,N_13905);
nor U14036 (N_14036,N_13968,N_13911);
nor U14037 (N_14037,N_13882,N_13908);
and U14038 (N_14038,N_13942,N_13965);
nand U14039 (N_14039,N_13985,N_13918);
nor U14040 (N_14040,N_13894,N_13925);
nand U14041 (N_14041,N_13949,N_13929);
or U14042 (N_14042,N_13893,N_13991);
nor U14043 (N_14043,N_13960,N_13963);
and U14044 (N_14044,N_13909,N_13897);
or U14045 (N_14045,N_13994,N_13881);
nand U14046 (N_14046,N_13895,N_13959);
nand U14047 (N_14047,N_13952,N_13901);
nand U14048 (N_14048,N_13977,N_13876);
xor U14049 (N_14049,N_13938,N_13910);
nor U14050 (N_14050,N_13957,N_13956);
nand U14051 (N_14051,N_13972,N_13998);
and U14052 (N_14052,N_13875,N_13877);
or U14053 (N_14053,N_13934,N_13943);
and U14054 (N_14054,N_13950,N_13955);
xor U14055 (N_14055,N_13941,N_13953);
nand U14056 (N_14056,N_13921,N_13931);
nor U14057 (N_14057,N_13917,N_13990);
nor U14058 (N_14058,N_13891,N_13964);
nand U14059 (N_14059,N_13966,N_13981);
nand U14060 (N_14060,N_13940,N_13913);
nor U14061 (N_14061,N_13995,N_13987);
and U14062 (N_14062,N_13976,N_13919);
xnor U14063 (N_14063,N_13978,N_13976);
nor U14064 (N_14064,N_13928,N_13881);
nand U14065 (N_14065,N_13919,N_13916);
and U14066 (N_14066,N_13914,N_13923);
xnor U14067 (N_14067,N_13879,N_13911);
nand U14068 (N_14068,N_13932,N_13955);
nor U14069 (N_14069,N_13915,N_13990);
nor U14070 (N_14070,N_13988,N_13936);
or U14071 (N_14071,N_13896,N_13976);
or U14072 (N_14072,N_13938,N_13911);
nand U14073 (N_14073,N_13986,N_13990);
and U14074 (N_14074,N_13990,N_13885);
nor U14075 (N_14075,N_13932,N_13884);
nor U14076 (N_14076,N_13900,N_13995);
and U14077 (N_14077,N_13952,N_13925);
or U14078 (N_14078,N_13954,N_13970);
nor U14079 (N_14079,N_13948,N_13938);
or U14080 (N_14080,N_13893,N_13958);
nor U14081 (N_14081,N_13930,N_13957);
nor U14082 (N_14082,N_13968,N_13912);
or U14083 (N_14083,N_13992,N_13877);
nand U14084 (N_14084,N_13895,N_13886);
or U14085 (N_14085,N_13993,N_13970);
nor U14086 (N_14086,N_13981,N_13892);
nor U14087 (N_14087,N_13896,N_13970);
nor U14088 (N_14088,N_13875,N_13976);
nor U14089 (N_14089,N_13979,N_13944);
nand U14090 (N_14090,N_13927,N_13996);
nand U14091 (N_14091,N_13932,N_13992);
and U14092 (N_14092,N_13900,N_13940);
xor U14093 (N_14093,N_13973,N_13929);
nand U14094 (N_14094,N_13920,N_13964);
or U14095 (N_14095,N_13896,N_13981);
or U14096 (N_14096,N_13932,N_13966);
nor U14097 (N_14097,N_13943,N_13880);
xor U14098 (N_14098,N_13985,N_13968);
or U14099 (N_14099,N_13965,N_13945);
or U14100 (N_14100,N_13981,N_13977);
nor U14101 (N_14101,N_13997,N_13968);
nor U14102 (N_14102,N_13999,N_13968);
or U14103 (N_14103,N_13981,N_13914);
and U14104 (N_14104,N_13887,N_13988);
and U14105 (N_14105,N_13923,N_13958);
nor U14106 (N_14106,N_13990,N_13919);
and U14107 (N_14107,N_13920,N_13977);
or U14108 (N_14108,N_13896,N_13958);
or U14109 (N_14109,N_13899,N_13938);
nand U14110 (N_14110,N_13963,N_13996);
or U14111 (N_14111,N_13894,N_13935);
nor U14112 (N_14112,N_13965,N_13895);
nor U14113 (N_14113,N_13995,N_13911);
xnor U14114 (N_14114,N_13998,N_13985);
nand U14115 (N_14115,N_13956,N_13907);
and U14116 (N_14116,N_13945,N_13976);
nor U14117 (N_14117,N_13907,N_13904);
nor U14118 (N_14118,N_13900,N_13996);
nand U14119 (N_14119,N_13983,N_13934);
or U14120 (N_14120,N_13917,N_13891);
xnor U14121 (N_14121,N_13877,N_13970);
nand U14122 (N_14122,N_13889,N_13987);
nand U14123 (N_14123,N_13927,N_13974);
and U14124 (N_14124,N_13950,N_13997);
nor U14125 (N_14125,N_14103,N_14097);
nand U14126 (N_14126,N_14062,N_14016);
nand U14127 (N_14127,N_14115,N_14109);
xor U14128 (N_14128,N_14034,N_14106);
nor U14129 (N_14129,N_14091,N_14041);
and U14130 (N_14130,N_14068,N_14019);
xor U14131 (N_14131,N_14110,N_14027);
xnor U14132 (N_14132,N_14064,N_14018);
and U14133 (N_14133,N_14122,N_14032);
nor U14134 (N_14134,N_14071,N_14111);
xnor U14135 (N_14135,N_14120,N_14118);
nand U14136 (N_14136,N_14093,N_14038);
or U14137 (N_14137,N_14114,N_14099);
nand U14138 (N_14138,N_14050,N_14024);
nor U14139 (N_14139,N_14045,N_14107);
or U14140 (N_14140,N_14026,N_14025);
xor U14141 (N_14141,N_14040,N_14084);
or U14142 (N_14142,N_14117,N_14073);
xor U14143 (N_14143,N_14011,N_14044);
and U14144 (N_14144,N_14076,N_14029);
nor U14145 (N_14145,N_14004,N_14092);
xor U14146 (N_14146,N_14089,N_14047);
nand U14147 (N_14147,N_14102,N_14082);
and U14148 (N_14148,N_14055,N_14023);
nor U14149 (N_14149,N_14009,N_14095);
nand U14150 (N_14150,N_14070,N_14061);
nor U14151 (N_14151,N_14066,N_14035);
nand U14152 (N_14152,N_14077,N_14020);
nor U14153 (N_14153,N_14087,N_14048);
nand U14154 (N_14154,N_14058,N_14037);
and U14155 (N_14155,N_14031,N_14005);
xnor U14156 (N_14156,N_14078,N_14052);
nor U14157 (N_14157,N_14022,N_14013);
xnor U14158 (N_14158,N_14051,N_14079);
xnor U14159 (N_14159,N_14039,N_14049);
and U14160 (N_14160,N_14123,N_14081);
and U14161 (N_14161,N_14003,N_14060);
or U14162 (N_14162,N_14083,N_14059);
xor U14163 (N_14163,N_14053,N_14065);
and U14164 (N_14164,N_14014,N_14119);
nand U14165 (N_14165,N_14012,N_14021);
or U14166 (N_14166,N_14057,N_14124);
nor U14167 (N_14167,N_14063,N_14086);
and U14168 (N_14168,N_14056,N_14108);
xnor U14169 (N_14169,N_14088,N_14094);
xor U14170 (N_14170,N_14054,N_14098);
nand U14171 (N_14171,N_14030,N_14067);
and U14172 (N_14172,N_14100,N_14043);
nand U14173 (N_14173,N_14015,N_14006);
nand U14174 (N_14174,N_14002,N_14036);
xnor U14175 (N_14175,N_14080,N_14001);
and U14176 (N_14176,N_14069,N_14105);
or U14177 (N_14177,N_14121,N_14112);
or U14178 (N_14178,N_14116,N_14046);
xnor U14179 (N_14179,N_14104,N_14028);
or U14180 (N_14180,N_14096,N_14010);
and U14181 (N_14181,N_14113,N_14008);
nor U14182 (N_14182,N_14074,N_14000);
and U14183 (N_14183,N_14090,N_14042);
or U14184 (N_14184,N_14075,N_14072);
and U14185 (N_14185,N_14101,N_14033);
nor U14186 (N_14186,N_14017,N_14085);
and U14187 (N_14187,N_14007,N_14051);
nor U14188 (N_14188,N_14069,N_14039);
nor U14189 (N_14189,N_14012,N_14033);
or U14190 (N_14190,N_14068,N_14094);
nor U14191 (N_14191,N_14102,N_14120);
or U14192 (N_14192,N_14040,N_14114);
and U14193 (N_14193,N_14001,N_14021);
nor U14194 (N_14194,N_14053,N_14117);
nand U14195 (N_14195,N_14080,N_14023);
and U14196 (N_14196,N_14066,N_14067);
xor U14197 (N_14197,N_14056,N_14033);
xnor U14198 (N_14198,N_14100,N_14119);
nor U14199 (N_14199,N_14001,N_14048);
nand U14200 (N_14200,N_14075,N_14049);
nand U14201 (N_14201,N_14088,N_14098);
or U14202 (N_14202,N_14022,N_14085);
nand U14203 (N_14203,N_14004,N_14107);
or U14204 (N_14204,N_14066,N_14074);
xnor U14205 (N_14205,N_14046,N_14091);
nor U14206 (N_14206,N_14029,N_14019);
nor U14207 (N_14207,N_14073,N_14098);
or U14208 (N_14208,N_14055,N_14109);
nor U14209 (N_14209,N_14099,N_14083);
or U14210 (N_14210,N_14103,N_14082);
nand U14211 (N_14211,N_14099,N_14120);
or U14212 (N_14212,N_14056,N_14070);
nor U14213 (N_14213,N_14091,N_14106);
nor U14214 (N_14214,N_14100,N_14118);
and U14215 (N_14215,N_14120,N_14058);
and U14216 (N_14216,N_14079,N_14058);
nor U14217 (N_14217,N_14031,N_14094);
and U14218 (N_14218,N_14121,N_14082);
nand U14219 (N_14219,N_14061,N_14099);
nand U14220 (N_14220,N_14000,N_14021);
xnor U14221 (N_14221,N_14023,N_14083);
xor U14222 (N_14222,N_14120,N_14072);
and U14223 (N_14223,N_14060,N_14032);
or U14224 (N_14224,N_14029,N_14010);
nor U14225 (N_14225,N_14095,N_14033);
nor U14226 (N_14226,N_14053,N_14036);
nand U14227 (N_14227,N_14068,N_14077);
nor U14228 (N_14228,N_14117,N_14123);
and U14229 (N_14229,N_14098,N_14124);
or U14230 (N_14230,N_14066,N_14123);
nor U14231 (N_14231,N_14053,N_14091);
and U14232 (N_14232,N_14040,N_14032);
nand U14233 (N_14233,N_14032,N_14039);
nand U14234 (N_14234,N_14051,N_14068);
nor U14235 (N_14235,N_14122,N_14036);
nor U14236 (N_14236,N_14053,N_14095);
nor U14237 (N_14237,N_14065,N_14117);
nand U14238 (N_14238,N_14090,N_14054);
nor U14239 (N_14239,N_14095,N_14104);
nor U14240 (N_14240,N_14077,N_14084);
nor U14241 (N_14241,N_14040,N_14011);
and U14242 (N_14242,N_14115,N_14049);
or U14243 (N_14243,N_14032,N_14094);
or U14244 (N_14244,N_14103,N_14020);
or U14245 (N_14245,N_14062,N_14081);
nand U14246 (N_14246,N_14074,N_14027);
or U14247 (N_14247,N_14031,N_14101);
nand U14248 (N_14248,N_14031,N_14043);
or U14249 (N_14249,N_14000,N_14081);
xor U14250 (N_14250,N_14145,N_14213);
and U14251 (N_14251,N_14203,N_14158);
or U14252 (N_14252,N_14177,N_14232);
nand U14253 (N_14253,N_14241,N_14208);
nand U14254 (N_14254,N_14166,N_14162);
nor U14255 (N_14255,N_14134,N_14170);
nor U14256 (N_14256,N_14180,N_14228);
nor U14257 (N_14257,N_14181,N_14136);
nor U14258 (N_14258,N_14186,N_14164);
and U14259 (N_14259,N_14163,N_14195);
xnor U14260 (N_14260,N_14210,N_14242);
xnor U14261 (N_14261,N_14233,N_14201);
and U14262 (N_14262,N_14128,N_14167);
or U14263 (N_14263,N_14248,N_14187);
nor U14264 (N_14264,N_14159,N_14178);
nor U14265 (N_14265,N_14196,N_14146);
and U14266 (N_14266,N_14182,N_14194);
and U14267 (N_14267,N_14174,N_14227);
nand U14268 (N_14268,N_14173,N_14131);
nor U14269 (N_14269,N_14153,N_14230);
nand U14270 (N_14270,N_14239,N_14204);
and U14271 (N_14271,N_14135,N_14175);
and U14272 (N_14272,N_14165,N_14217);
and U14273 (N_14273,N_14150,N_14246);
and U14274 (N_14274,N_14176,N_14224);
or U14275 (N_14275,N_14190,N_14144);
or U14276 (N_14276,N_14151,N_14193);
xor U14277 (N_14277,N_14185,N_14189);
nand U14278 (N_14278,N_14125,N_14222);
or U14279 (N_14279,N_14245,N_14212);
nor U14280 (N_14280,N_14142,N_14140);
nand U14281 (N_14281,N_14179,N_14155);
nand U14282 (N_14282,N_14215,N_14234);
nand U14283 (N_14283,N_14199,N_14126);
nor U14284 (N_14284,N_14138,N_14130);
or U14285 (N_14285,N_14188,N_14243);
and U14286 (N_14286,N_14127,N_14211);
or U14287 (N_14287,N_14191,N_14198);
and U14288 (N_14288,N_14148,N_14236);
xor U14289 (N_14289,N_14218,N_14220);
nand U14290 (N_14290,N_14247,N_14139);
and U14291 (N_14291,N_14160,N_14226);
nor U14292 (N_14292,N_14157,N_14221);
xnor U14293 (N_14293,N_14152,N_14214);
nand U14294 (N_14294,N_14183,N_14161);
or U14295 (N_14295,N_14133,N_14172);
xnor U14296 (N_14296,N_14184,N_14237);
and U14297 (N_14297,N_14156,N_14229);
xor U14298 (N_14298,N_14240,N_14147);
nand U14299 (N_14299,N_14200,N_14149);
nor U14300 (N_14300,N_14249,N_14143);
nand U14301 (N_14301,N_14171,N_14192);
and U14302 (N_14302,N_14205,N_14206);
nor U14303 (N_14303,N_14168,N_14141);
nor U14304 (N_14304,N_14238,N_14223);
and U14305 (N_14305,N_14202,N_14132);
nand U14306 (N_14306,N_14216,N_14207);
and U14307 (N_14307,N_14244,N_14137);
nand U14308 (N_14308,N_14169,N_14219);
and U14309 (N_14309,N_14225,N_14235);
or U14310 (N_14310,N_14129,N_14231);
or U14311 (N_14311,N_14154,N_14197);
or U14312 (N_14312,N_14209,N_14225);
nand U14313 (N_14313,N_14183,N_14186);
nand U14314 (N_14314,N_14154,N_14213);
and U14315 (N_14315,N_14162,N_14219);
or U14316 (N_14316,N_14197,N_14237);
nor U14317 (N_14317,N_14148,N_14134);
nor U14318 (N_14318,N_14136,N_14167);
or U14319 (N_14319,N_14206,N_14130);
or U14320 (N_14320,N_14249,N_14206);
nor U14321 (N_14321,N_14205,N_14193);
or U14322 (N_14322,N_14235,N_14135);
xnor U14323 (N_14323,N_14227,N_14212);
and U14324 (N_14324,N_14175,N_14147);
xnor U14325 (N_14325,N_14128,N_14195);
or U14326 (N_14326,N_14211,N_14163);
or U14327 (N_14327,N_14167,N_14212);
nor U14328 (N_14328,N_14164,N_14181);
nor U14329 (N_14329,N_14170,N_14173);
and U14330 (N_14330,N_14177,N_14183);
and U14331 (N_14331,N_14216,N_14139);
or U14332 (N_14332,N_14162,N_14209);
xor U14333 (N_14333,N_14140,N_14165);
nand U14334 (N_14334,N_14213,N_14152);
or U14335 (N_14335,N_14181,N_14208);
xor U14336 (N_14336,N_14146,N_14226);
xor U14337 (N_14337,N_14209,N_14187);
nand U14338 (N_14338,N_14193,N_14247);
nand U14339 (N_14339,N_14232,N_14242);
nor U14340 (N_14340,N_14156,N_14172);
and U14341 (N_14341,N_14194,N_14241);
nand U14342 (N_14342,N_14178,N_14149);
nand U14343 (N_14343,N_14223,N_14198);
or U14344 (N_14344,N_14210,N_14223);
nand U14345 (N_14345,N_14155,N_14190);
nor U14346 (N_14346,N_14178,N_14179);
nor U14347 (N_14347,N_14198,N_14244);
or U14348 (N_14348,N_14160,N_14181);
nand U14349 (N_14349,N_14208,N_14197);
nor U14350 (N_14350,N_14183,N_14187);
nor U14351 (N_14351,N_14191,N_14142);
nand U14352 (N_14352,N_14192,N_14143);
or U14353 (N_14353,N_14212,N_14196);
nand U14354 (N_14354,N_14134,N_14146);
nor U14355 (N_14355,N_14234,N_14210);
nand U14356 (N_14356,N_14143,N_14247);
nand U14357 (N_14357,N_14234,N_14194);
or U14358 (N_14358,N_14167,N_14147);
nand U14359 (N_14359,N_14199,N_14226);
and U14360 (N_14360,N_14188,N_14134);
nand U14361 (N_14361,N_14165,N_14152);
nor U14362 (N_14362,N_14245,N_14236);
or U14363 (N_14363,N_14194,N_14229);
xnor U14364 (N_14364,N_14167,N_14141);
or U14365 (N_14365,N_14193,N_14222);
xnor U14366 (N_14366,N_14198,N_14159);
nand U14367 (N_14367,N_14185,N_14201);
or U14368 (N_14368,N_14244,N_14232);
or U14369 (N_14369,N_14185,N_14225);
or U14370 (N_14370,N_14149,N_14181);
or U14371 (N_14371,N_14180,N_14229);
or U14372 (N_14372,N_14231,N_14145);
and U14373 (N_14373,N_14168,N_14146);
xor U14374 (N_14374,N_14240,N_14241);
nand U14375 (N_14375,N_14335,N_14307);
nand U14376 (N_14376,N_14305,N_14344);
nor U14377 (N_14377,N_14345,N_14313);
nand U14378 (N_14378,N_14269,N_14341);
and U14379 (N_14379,N_14353,N_14322);
or U14380 (N_14380,N_14360,N_14281);
or U14381 (N_14381,N_14336,N_14290);
nor U14382 (N_14382,N_14348,N_14359);
and U14383 (N_14383,N_14321,N_14351);
and U14384 (N_14384,N_14352,N_14284);
nand U14385 (N_14385,N_14320,N_14273);
xor U14386 (N_14386,N_14283,N_14308);
and U14387 (N_14387,N_14347,N_14274);
and U14388 (N_14388,N_14267,N_14319);
or U14389 (N_14389,N_14298,N_14311);
and U14390 (N_14390,N_14303,N_14255);
nand U14391 (N_14391,N_14357,N_14349);
and U14392 (N_14392,N_14369,N_14265);
nor U14393 (N_14393,N_14314,N_14302);
and U14394 (N_14394,N_14330,N_14374);
nor U14395 (N_14395,N_14340,N_14306);
nor U14396 (N_14396,N_14364,N_14292);
and U14397 (N_14397,N_14342,N_14291);
xnor U14398 (N_14398,N_14337,N_14272);
nor U14399 (N_14399,N_14263,N_14296);
xnor U14400 (N_14400,N_14331,N_14316);
and U14401 (N_14401,N_14278,N_14301);
or U14402 (N_14402,N_14268,N_14312);
nor U14403 (N_14403,N_14294,N_14275);
nand U14404 (N_14404,N_14354,N_14258);
xnor U14405 (N_14405,N_14363,N_14355);
nand U14406 (N_14406,N_14356,N_14270);
nand U14407 (N_14407,N_14260,N_14257);
nor U14408 (N_14408,N_14261,N_14367);
nand U14409 (N_14409,N_14343,N_14280);
and U14410 (N_14410,N_14323,N_14372);
nand U14411 (N_14411,N_14373,N_14339);
and U14412 (N_14412,N_14333,N_14289);
and U14413 (N_14413,N_14318,N_14338);
and U14414 (N_14414,N_14288,N_14362);
or U14415 (N_14415,N_14287,N_14285);
nand U14416 (N_14416,N_14276,N_14368);
xor U14417 (N_14417,N_14334,N_14371);
and U14418 (N_14418,N_14295,N_14262);
or U14419 (N_14419,N_14325,N_14350);
xnor U14420 (N_14420,N_14315,N_14332);
nand U14421 (N_14421,N_14361,N_14286);
and U14422 (N_14422,N_14304,N_14259);
nand U14423 (N_14423,N_14366,N_14252);
nand U14424 (N_14424,N_14253,N_14254);
nor U14425 (N_14425,N_14282,N_14358);
nand U14426 (N_14426,N_14370,N_14328);
and U14427 (N_14427,N_14324,N_14277);
or U14428 (N_14428,N_14326,N_14329);
nand U14429 (N_14429,N_14293,N_14365);
or U14430 (N_14430,N_14264,N_14327);
nor U14431 (N_14431,N_14256,N_14251);
or U14432 (N_14432,N_14266,N_14279);
or U14433 (N_14433,N_14309,N_14300);
nand U14434 (N_14434,N_14271,N_14317);
or U14435 (N_14435,N_14346,N_14250);
nor U14436 (N_14436,N_14299,N_14310);
nor U14437 (N_14437,N_14297,N_14318);
nand U14438 (N_14438,N_14294,N_14355);
nand U14439 (N_14439,N_14283,N_14303);
or U14440 (N_14440,N_14329,N_14317);
nand U14441 (N_14441,N_14350,N_14250);
nand U14442 (N_14442,N_14261,N_14346);
and U14443 (N_14443,N_14344,N_14250);
nor U14444 (N_14444,N_14299,N_14254);
and U14445 (N_14445,N_14354,N_14256);
or U14446 (N_14446,N_14266,N_14257);
nand U14447 (N_14447,N_14296,N_14250);
and U14448 (N_14448,N_14273,N_14325);
and U14449 (N_14449,N_14289,N_14351);
nor U14450 (N_14450,N_14306,N_14347);
or U14451 (N_14451,N_14366,N_14282);
xnor U14452 (N_14452,N_14281,N_14287);
or U14453 (N_14453,N_14284,N_14252);
nor U14454 (N_14454,N_14303,N_14314);
nand U14455 (N_14455,N_14319,N_14289);
and U14456 (N_14456,N_14267,N_14332);
xor U14457 (N_14457,N_14335,N_14250);
nor U14458 (N_14458,N_14361,N_14288);
nor U14459 (N_14459,N_14357,N_14291);
and U14460 (N_14460,N_14266,N_14322);
nand U14461 (N_14461,N_14298,N_14268);
and U14462 (N_14462,N_14307,N_14330);
and U14463 (N_14463,N_14337,N_14293);
nand U14464 (N_14464,N_14307,N_14287);
and U14465 (N_14465,N_14313,N_14334);
or U14466 (N_14466,N_14374,N_14326);
nor U14467 (N_14467,N_14332,N_14334);
or U14468 (N_14468,N_14259,N_14269);
or U14469 (N_14469,N_14269,N_14359);
or U14470 (N_14470,N_14331,N_14312);
xnor U14471 (N_14471,N_14312,N_14368);
nor U14472 (N_14472,N_14277,N_14368);
nand U14473 (N_14473,N_14266,N_14325);
xor U14474 (N_14474,N_14264,N_14346);
nand U14475 (N_14475,N_14342,N_14255);
xnor U14476 (N_14476,N_14360,N_14295);
nand U14477 (N_14477,N_14343,N_14266);
and U14478 (N_14478,N_14322,N_14336);
xor U14479 (N_14479,N_14279,N_14270);
xor U14480 (N_14480,N_14316,N_14341);
and U14481 (N_14481,N_14314,N_14372);
nor U14482 (N_14482,N_14361,N_14370);
and U14483 (N_14483,N_14330,N_14324);
and U14484 (N_14484,N_14358,N_14274);
and U14485 (N_14485,N_14293,N_14280);
and U14486 (N_14486,N_14352,N_14298);
and U14487 (N_14487,N_14325,N_14321);
or U14488 (N_14488,N_14304,N_14349);
and U14489 (N_14489,N_14339,N_14297);
nand U14490 (N_14490,N_14302,N_14334);
nand U14491 (N_14491,N_14293,N_14312);
nor U14492 (N_14492,N_14318,N_14361);
and U14493 (N_14493,N_14293,N_14313);
nor U14494 (N_14494,N_14346,N_14265);
nor U14495 (N_14495,N_14365,N_14345);
or U14496 (N_14496,N_14279,N_14370);
or U14497 (N_14497,N_14303,N_14297);
nor U14498 (N_14498,N_14286,N_14293);
nand U14499 (N_14499,N_14256,N_14335);
nor U14500 (N_14500,N_14492,N_14457);
nor U14501 (N_14501,N_14440,N_14463);
or U14502 (N_14502,N_14389,N_14441);
nand U14503 (N_14503,N_14453,N_14445);
or U14504 (N_14504,N_14444,N_14380);
nand U14505 (N_14505,N_14491,N_14442);
and U14506 (N_14506,N_14426,N_14438);
nand U14507 (N_14507,N_14414,N_14377);
nand U14508 (N_14508,N_14425,N_14412);
and U14509 (N_14509,N_14406,N_14488);
nor U14510 (N_14510,N_14472,N_14481);
nor U14511 (N_14511,N_14400,N_14385);
and U14512 (N_14512,N_14449,N_14468);
nand U14513 (N_14513,N_14421,N_14387);
or U14514 (N_14514,N_14404,N_14430);
and U14515 (N_14515,N_14479,N_14458);
nand U14516 (N_14516,N_14375,N_14474);
or U14517 (N_14517,N_14465,N_14420);
nand U14518 (N_14518,N_14390,N_14388);
xor U14519 (N_14519,N_14396,N_14408);
nand U14520 (N_14520,N_14478,N_14436);
nand U14521 (N_14521,N_14427,N_14428);
nand U14522 (N_14522,N_14464,N_14394);
and U14523 (N_14523,N_14423,N_14376);
xor U14524 (N_14524,N_14486,N_14471);
xor U14525 (N_14525,N_14413,N_14470);
and U14526 (N_14526,N_14397,N_14455);
nor U14527 (N_14527,N_14477,N_14494);
nor U14528 (N_14528,N_14392,N_14405);
nor U14529 (N_14529,N_14498,N_14482);
nor U14530 (N_14530,N_14429,N_14381);
nor U14531 (N_14531,N_14434,N_14424);
nand U14532 (N_14532,N_14462,N_14487);
and U14533 (N_14533,N_14411,N_14393);
or U14534 (N_14534,N_14459,N_14456);
nand U14535 (N_14535,N_14485,N_14416);
nand U14536 (N_14536,N_14435,N_14379);
and U14537 (N_14537,N_14410,N_14446);
or U14538 (N_14538,N_14447,N_14418);
nor U14539 (N_14539,N_14461,N_14496);
nand U14540 (N_14540,N_14489,N_14386);
and U14541 (N_14541,N_14460,N_14450);
nand U14542 (N_14542,N_14402,N_14454);
or U14543 (N_14543,N_14433,N_14495);
and U14544 (N_14544,N_14493,N_14409);
nor U14545 (N_14545,N_14419,N_14437);
nand U14546 (N_14546,N_14497,N_14407);
nor U14547 (N_14547,N_14399,N_14443);
or U14548 (N_14548,N_14499,N_14467);
nor U14549 (N_14549,N_14417,N_14384);
nand U14550 (N_14550,N_14452,N_14490);
and U14551 (N_14551,N_14401,N_14415);
and U14552 (N_14552,N_14378,N_14439);
or U14553 (N_14553,N_14475,N_14448);
xor U14554 (N_14554,N_14395,N_14451);
and U14555 (N_14555,N_14391,N_14466);
nor U14556 (N_14556,N_14382,N_14431);
or U14557 (N_14557,N_14473,N_14403);
and U14558 (N_14558,N_14398,N_14484);
or U14559 (N_14559,N_14422,N_14476);
nor U14560 (N_14560,N_14383,N_14432);
or U14561 (N_14561,N_14480,N_14469);
xnor U14562 (N_14562,N_14483,N_14408);
or U14563 (N_14563,N_14417,N_14404);
nor U14564 (N_14564,N_14419,N_14455);
and U14565 (N_14565,N_14447,N_14483);
or U14566 (N_14566,N_14407,N_14400);
or U14567 (N_14567,N_14451,N_14495);
and U14568 (N_14568,N_14473,N_14490);
or U14569 (N_14569,N_14383,N_14435);
or U14570 (N_14570,N_14468,N_14458);
nand U14571 (N_14571,N_14409,N_14473);
nor U14572 (N_14572,N_14385,N_14446);
or U14573 (N_14573,N_14489,N_14483);
or U14574 (N_14574,N_14481,N_14470);
nor U14575 (N_14575,N_14487,N_14417);
nor U14576 (N_14576,N_14470,N_14433);
nor U14577 (N_14577,N_14397,N_14469);
nor U14578 (N_14578,N_14485,N_14421);
xnor U14579 (N_14579,N_14420,N_14382);
or U14580 (N_14580,N_14456,N_14407);
nor U14581 (N_14581,N_14377,N_14455);
and U14582 (N_14582,N_14476,N_14421);
nor U14583 (N_14583,N_14443,N_14424);
nor U14584 (N_14584,N_14382,N_14447);
nor U14585 (N_14585,N_14415,N_14419);
nor U14586 (N_14586,N_14389,N_14394);
nor U14587 (N_14587,N_14480,N_14413);
nor U14588 (N_14588,N_14475,N_14410);
or U14589 (N_14589,N_14495,N_14463);
nand U14590 (N_14590,N_14443,N_14498);
and U14591 (N_14591,N_14415,N_14409);
or U14592 (N_14592,N_14381,N_14421);
nand U14593 (N_14593,N_14468,N_14463);
and U14594 (N_14594,N_14416,N_14470);
nand U14595 (N_14595,N_14389,N_14410);
xnor U14596 (N_14596,N_14422,N_14427);
and U14597 (N_14597,N_14405,N_14395);
and U14598 (N_14598,N_14416,N_14481);
or U14599 (N_14599,N_14479,N_14489);
nor U14600 (N_14600,N_14421,N_14395);
or U14601 (N_14601,N_14383,N_14496);
nor U14602 (N_14602,N_14415,N_14390);
xor U14603 (N_14603,N_14389,N_14474);
and U14604 (N_14604,N_14413,N_14494);
nand U14605 (N_14605,N_14490,N_14423);
nor U14606 (N_14606,N_14436,N_14434);
and U14607 (N_14607,N_14419,N_14377);
nand U14608 (N_14608,N_14495,N_14431);
or U14609 (N_14609,N_14432,N_14465);
nand U14610 (N_14610,N_14467,N_14474);
or U14611 (N_14611,N_14403,N_14410);
nor U14612 (N_14612,N_14382,N_14390);
and U14613 (N_14613,N_14432,N_14403);
and U14614 (N_14614,N_14414,N_14479);
nor U14615 (N_14615,N_14487,N_14485);
and U14616 (N_14616,N_14440,N_14405);
and U14617 (N_14617,N_14461,N_14442);
and U14618 (N_14618,N_14415,N_14414);
nor U14619 (N_14619,N_14388,N_14450);
and U14620 (N_14620,N_14464,N_14396);
nand U14621 (N_14621,N_14488,N_14385);
nor U14622 (N_14622,N_14460,N_14488);
and U14623 (N_14623,N_14479,N_14390);
or U14624 (N_14624,N_14457,N_14453);
nor U14625 (N_14625,N_14559,N_14606);
nand U14626 (N_14626,N_14580,N_14536);
and U14627 (N_14627,N_14568,N_14616);
nor U14628 (N_14628,N_14507,N_14570);
and U14629 (N_14629,N_14511,N_14541);
or U14630 (N_14630,N_14590,N_14592);
nand U14631 (N_14631,N_14600,N_14596);
nor U14632 (N_14632,N_14529,N_14573);
and U14633 (N_14633,N_14502,N_14619);
and U14634 (N_14634,N_14516,N_14604);
or U14635 (N_14635,N_14553,N_14578);
nand U14636 (N_14636,N_14587,N_14607);
nor U14637 (N_14637,N_14555,N_14566);
nand U14638 (N_14638,N_14543,N_14564);
nor U14639 (N_14639,N_14610,N_14591);
nand U14640 (N_14640,N_14582,N_14581);
nor U14641 (N_14641,N_14585,N_14532);
xnor U14642 (N_14642,N_14574,N_14533);
or U14643 (N_14643,N_14542,N_14557);
xnor U14644 (N_14644,N_14618,N_14534);
nor U14645 (N_14645,N_14593,N_14563);
xnor U14646 (N_14646,N_14520,N_14551);
xor U14647 (N_14647,N_14550,N_14558);
xnor U14648 (N_14648,N_14548,N_14514);
nor U14649 (N_14649,N_14560,N_14524);
and U14650 (N_14650,N_14565,N_14526);
nor U14651 (N_14651,N_14584,N_14523);
nor U14652 (N_14652,N_14579,N_14544);
or U14653 (N_14653,N_14594,N_14562);
nand U14654 (N_14654,N_14556,N_14515);
or U14655 (N_14655,N_14513,N_14521);
and U14656 (N_14656,N_14576,N_14567);
and U14657 (N_14657,N_14595,N_14611);
nand U14658 (N_14658,N_14569,N_14539);
or U14659 (N_14659,N_14612,N_14598);
nand U14660 (N_14660,N_14608,N_14602);
and U14661 (N_14661,N_14503,N_14624);
nand U14662 (N_14662,N_14561,N_14522);
and U14663 (N_14663,N_14583,N_14510);
nor U14664 (N_14664,N_14538,N_14501);
and U14665 (N_14665,N_14530,N_14535);
nand U14666 (N_14666,N_14575,N_14609);
nor U14667 (N_14667,N_14571,N_14577);
and U14668 (N_14668,N_14603,N_14601);
nor U14669 (N_14669,N_14552,N_14527);
nand U14670 (N_14670,N_14588,N_14540);
and U14671 (N_14671,N_14572,N_14525);
nand U14672 (N_14672,N_14531,N_14554);
and U14673 (N_14673,N_14614,N_14597);
nor U14674 (N_14674,N_14599,N_14621);
nand U14675 (N_14675,N_14613,N_14615);
nor U14676 (N_14676,N_14512,N_14617);
nand U14677 (N_14677,N_14605,N_14589);
nand U14678 (N_14678,N_14623,N_14549);
nor U14679 (N_14679,N_14506,N_14537);
and U14680 (N_14680,N_14622,N_14620);
or U14681 (N_14681,N_14519,N_14586);
nand U14682 (N_14682,N_14528,N_14504);
nand U14683 (N_14683,N_14546,N_14545);
xnor U14684 (N_14684,N_14547,N_14508);
or U14685 (N_14685,N_14517,N_14500);
or U14686 (N_14686,N_14509,N_14505);
or U14687 (N_14687,N_14518,N_14536);
and U14688 (N_14688,N_14607,N_14523);
xnor U14689 (N_14689,N_14611,N_14623);
and U14690 (N_14690,N_14544,N_14547);
or U14691 (N_14691,N_14569,N_14545);
nand U14692 (N_14692,N_14571,N_14518);
nand U14693 (N_14693,N_14515,N_14571);
nand U14694 (N_14694,N_14500,N_14519);
or U14695 (N_14695,N_14539,N_14514);
and U14696 (N_14696,N_14547,N_14532);
nand U14697 (N_14697,N_14571,N_14608);
nor U14698 (N_14698,N_14603,N_14529);
nor U14699 (N_14699,N_14533,N_14576);
nand U14700 (N_14700,N_14550,N_14526);
or U14701 (N_14701,N_14584,N_14617);
nor U14702 (N_14702,N_14550,N_14556);
and U14703 (N_14703,N_14546,N_14622);
xor U14704 (N_14704,N_14552,N_14592);
and U14705 (N_14705,N_14607,N_14591);
or U14706 (N_14706,N_14534,N_14568);
or U14707 (N_14707,N_14517,N_14571);
nor U14708 (N_14708,N_14597,N_14588);
and U14709 (N_14709,N_14578,N_14597);
nand U14710 (N_14710,N_14603,N_14564);
nor U14711 (N_14711,N_14542,N_14621);
or U14712 (N_14712,N_14563,N_14542);
nand U14713 (N_14713,N_14557,N_14507);
and U14714 (N_14714,N_14562,N_14573);
nand U14715 (N_14715,N_14616,N_14549);
nor U14716 (N_14716,N_14552,N_14513);
xor U14717 (N_14717,N_14611,N_14503);
nor U14718 (N_14718,N_14604,N_14526);
and U14719 (N_14719,N_14570,N_14624);
nor U14720 (N_14720,N_14621,N_14526);
and U14721 (N_14721,N_14560,N_14604);
or U14722 (N_14722,N_14593,N_14569);
nand U14723 (N_14723,N_14605,N_14521);
or U14724 (N_14724,N_14612,N_14503);
xor U14725 (N_14725,N_14580,N_14616);
nor U14726 (N_14726,N_14606,N_14554);
xnor U14727 (N_14727,N_14591,N_14535);
nor U14728 (N_14728,N_14557,N_14585);
nand U14729 (N_14729,N_14524,N_14562);
and U14730 (N_14730,N_14526,N_14505);
and U14731 (N_14731,N_14608,N_14578);
nand U14732 (N_14732,N_14547,N_14604);
or U14733 (N_14733,N_14595,N_14574);
nand U14734 (N_14734,N_14573,N_14581);
xnor U14735 (N_14735,N_14575,N_14607);
and U14736 (N_14736,N_14526,N_14560);
or U14737 (N_14737,N_14516,N_14579);
nor U14738 (N_14738,N_14572,N_14571);
nand U14739 (N_14739,N_14563,N_14535);
nor U14740 (N_14740,N_14541,N_14563);
or U14741 (N_14741,N_14545,N_14598);
nand U14742 (N_14742,N_14511,N_14590);
and U14743 (N_14743,N_14527,N_14550);
nor U14744 (N_14744,N_14619,N_14580);
nor U14745 (N_14745,N_14518,N_14573);
xnor U14746 (N_14746,N_14515,N_14514);
and U14747 (N_14747,N_14555,N_14558);
and U14748 (N_14748,N_14606,N_14587);
nand U14749 (N_14749,N_14502,N_14607);
and U14750 (N_14750,N_14627,N_14660);
or U14751 (N_14751,N_14738,N_14673);
or U14752 (N_14752,N_14672,N_14631);
or U14753 (N_14753,N_14657,N_14732);
and U14754 (N_14754,N_14739,N_14716);
nand U14755 (N_14755,N_14712,N_14649);
xor U14756 (N_14756,N_14715,N_14636);
or U14757 (N_14757,N_14705,N_14640);
nor U14758 (N_14758,N_14727,N_14670);
or U14759 (N_14759,N_14734,N_14721);
xor U14760 (N_14760,N_14639,N_14730);
and U14761 (N_14761,N_14629,N_14676);
and U14762 (N_14762,N_14625,N_14725);
and U14763 (N_14763,N_14644,N_14637);
or U14764 (N_14764,N_14747,N_14749);
and U14765 (N_14765,N_14736,N_14680);
or U14766 (N_14766,N_14646,N_14742);
or U14767 (N_14767,N_14662,N_14684);
nand U14768 (N_14768,N_14709,N_14686);
nand U14769 (N_14769,N_14677,N_14681);
and U14770 (N_14770,N_14710,N_14665);
and U14771 (N_14771,N_14645,N_14641);
nand U14772 (N_14772,N_14702,N_14669);
and U14773 (N_14773,N_14723,N_14746);
or U14774 (N_14774,N_14743,N_14722);
and U14775 (N_14775,N_14691,N_14648);
or U14776 (N_14776,N_14713,N_14714);
or U14777 (N_14777,N_14666,N_14628);
nand U14778 (N_14778,N_14697,N_14695);
or U14779 (N_14779,N_14682,N_14748);
nand U14780 (N_14780,N_14653,N_14688);
nor U14781 (N_14781,N_14675,N_14708);
nor U14782 (N_14782,N_14663,N_14652);
nand U14783 (N_14783,N_14683,N_14651);
or U14784 (N_14784,N_14679,N_14699);
xnor U14785 (N_14785,N_14706,N_14731);
and U14786 (N_14786,N_14647,N_14737);
nand U14787 (N_14787,N_14701,N_14724);
nand U14788 (N_14788,N_14728,N_14704);
and U14789 (N_14789,N_14741,N_14693);
nor U14790 (N_14790,N_14642,N_14685);
nand U14791 (N_14791,N_14720,N_14745);
and U14792 (N_14792,N_14671,N_14719);
xor U14793 (N_14793,N_14698,N_14678);
nor U14794 (N_14794,N_14696,N_14726);
nor U14795 (N_14795,N_14650,N_14664);
or U14796 (N_14796,N_14733,N_14633);
nand U14797 (N_14797,N_14735,N_14703);
or U14798 (N_14798,N_14707,N_14638);
nand U14799 (N_14799,N_14689,N_14668);
nor U14800 (N_14800,N_14674,N_14655);
and U14801 (N_14801,N_14626,N_14692);
nor U14802 (N_14802,N_14740,N_14729);
nand U14803 (N_14803,N_14635,N_14718);
and U14804 (N_14804,N_14687,N_14656);
or U14805 (N_14805,N_14717,N_14744);
and U14806 (N_14806,N_14690,N_14634);
nor U14807 (N_14807,N_14643,N_14654);
xor U14808 (N_14808,N_14658,N_14694);
nor U14809 (N_14809,N_14630,N_14700);
xnor U14810 (N_14810,N_14659,N_14632);
nor U14811 (N_14811,N_14661,N_14667);
and U14812 (N_14812,N_14711,N_14736);
and U14813 (N_14813,N_14734,N_14733);
nor U14814 (N_14814,N_14749,N_14736);
nor U14815 (N_14815,N_14710,N_14716);
nor U14816 (N_14816,N_14741,N_14666);
nand U14817 (N_14817,N_14642,N_14725);
nor U14818 (N_14818,N_14705,N_14748);
and U14819 (N_14819,N_14632,N_14692);
or U14820 (N_14820,N_14636,N_14740);
nor U14821 (N_14821,N_14626,N_14730);
or U14822 (N_14822,N_14690,N_14712);
or U14823 (N_14823,N_14700,N_14701);
nor U14824 (N_14824,N_14665,N_14676);
nand U14825 (N_14825,N_14634,N_14658);
nor U14826 (N_14826,N_14710,N_14726);
and U14827 (N_14827,N_14748,N_14691);
nor U14828 (N_14828,N_14715,N_14627);
nor U14829 (N_14829,N_14637,N_14683);
and U14830 (N_14830,N_14673,N_14646);
nand U14831 (N_14831,N_14626,N_14665);
nor U14832 (N_14832,N_14689,N_14702);
and U14833 (N_14833,N_14728,N_14662);
or U14834 (N_14834,N_14704,N_14678);
and U14835 (N_14835,N_14629,N_14731);
or U14836 (N_14836,N_14714,N_14668);
nor U14837 (N_14837,N_14688,N_14657);
and U14838 (N_14838,N_14694,N_14719);
and U14839 (N_14839,N_14718,N_14631);
or U14840 (N_14840,N_14683,N_14684);
nand U14841 (N_14841,N_14700,N_14741);
nand U14842 (N_14842,N_14682,N_14684);
xnor U14843 (N_14843,N_14703,N_14656);
and U14844 (N_14844,N_14690,N_14721);
or U14845 (N_14845,N_14710,N_14653);
and U14846 (N_14846,N_14717,N_14630);
or U14847 (N_14847,N_14627,N_14731);
or U14848 (N_14848,N_14626,N_14703);
nand U14849 (N_14849,N_14739,N_14712);
nor U14850 (N_14850,N_14679,N_14648);
and U14851 (N_14851,N_14695,N_14645);
and U14852 (N_14852,N_14712,N_14738);
and U14853 (N_14853,N_14645,N_14711);
nand U14854 (N_14854,N_14705,N_14724);
and U14855 (N_14855,N_14640,N_14696);
or U14856 (N_14856,N_14640,N_14661);
nor U14857 (N_14857,N_14706,N_14742);
or U14858 (N_14858,N_14693,N_14662);
nand U14859 (N_14859,N_14710,N_14678);
or U14860 (N_14860,N_14669,N_14695);
nand U14861 (N_14861,N_14638,N_14629);
and U14862 (N_14862,N_14681,N_14708);
or U14863 (N_14863,N_14666,N_14707);
xnor U14864 (N_14864,N_14721,N_14727);
nand U14865 (N_14865,N_14716,N_14732);
nor U14866 (N_14866,N_14656,N_14735);
nor U14867 (N_14867,N_14739,N_14683);
nor U14868 (N_14868,N_14672,N_14711);
xnor U14869 (N_14869,N_14743,N_14663);
or U14870 (N_14870,N_14710,N_14709);
xor U14871 (N_14871,N_14692,N_14645);
xor U14872 (N_14872,N_14630,N_14748);
nor U14873 (N_14873,N_14699,N_14682);
and U14874 (N_14874,N_14664,N_14709);
nand U14875 (N_14875,N_14832,N_14792);
or U14876 (N_14876,N_14776,N_14755);
nor U14877 (N_14877,N_14871,N_14816);
or U14878 (N_14878,N_14851,N_14825);
nand U14879 (N_14879,N_14759,N_14762);
or U14880 (N_14880,N_14778,N_14829);
or U14881 (N_14881,N_14847,N_14783);
nand U14882 (N_14882,N_14752,N_14794);
or U14883 (N_14883,N_14804,N_14838);
nand U14884 (N_14884,N_14814,N_14820);
or U14885 (N_14885,N_14809,N_14860);
or U14886 (N_14886,N_14786,N_14826);
nor U14887 (N_14887,N_14761,N_14780);
nand U14888 (N_14888,N_14782,N_14754);
xnor U14889 (N_14889,N_14864,N_14787);
or U14890 (N_14890,N_14823,N_14846);
nand U14891 (N_14891,N_14779,N_14859);
nand U14892 (N_14892,N_14800,N_14768);
and U14893 (N_14893,N_14837,N_14751);
nand U14894 (N_14894,N_14750,N_14839);
xnor U14895 (N_14895,N_14843,N_14812);
or U14896 (N_14896,N_14848,N_14852);
or U14897 (N_14897,N_14835,N_14865);
nor U14898 (N_14898,N_14840,N_14856);
xor U14899 (N_14899,N_14874,N_14867);
xor U14900 (N_14900,N_14857,N_14811);
and U14901 (N_14901,N_14789,N_14788);
nor U14902 (N_14902,N_14819,N_14756);
nand U14903 (N_14903,N_14773,N_14868);
nor U14904 (N_14904,N_14767,N_14869);
nand U14905 (N_14905,N_14836,N_14763);
nand U14906 (N_14906,N_14790,N_14870);
xor U14907 (N_14907,N_14791,N_14769);
and U14908 (N_14908,N_14797,N_14760);
and U14909 (N_14909,N_14785,N_14861);
nand U14910 (N_14910,N_14845,N_14822);
and U14911 (N_14911,N_14858,N_14862);
nand U14912 (N_14912,N_14774,N_14841);
xor U14913 (N_14913,N_14834,N_14855);
xnor U14914 (N_14914,N_14771,N_14753);
nor U14915 (N_14915,N_14805,N_14799);
or U14916 (N_14916,N_14830,N_14758);
nand U14917 (N_14917,N_14849,N_14850);
and U14918 (N_14918,N_14833,N_14781);
and U14919 (N_14919,N_14777,N_14775);
nor U14920 (N_14920,N_14807,N_14818);
xnor U14921 (N_14921,N_14824,N_14863);
xor U14922 (N_14922,N_14827,N_14765);
nor U14923 (N_14923,N_14793,N_14803);
nand U14924 (N_14924,N_14764,N_14854);
nor U14925 (N_14925,N_14813,N_14766);
nor U14926 (N_14926,N_14784,N_14844);
nand U14927 (N_14927,N_14796,N_14866);
nand U14928 (N_14928,N_14801,N_14873);
nor U14929 (N_14929,N_14815,N_14810);
nor U14930 (N_14930,N_14821,N_14828);
nand U14931 (N_14931,N_14772,N_14770);
nand U14932 (N_14932,N_14808,N_14842);
or U14933 (N_14933,N_14802,N_14853);
nand U14934 (N_14934,N_14817,N_14757);
and U14935 (N_14935,N_14831,N_14795);
nor U14936 (N_14936,N_14798,N_14872);
or U14937 (N_14937,N_14806,N_14765);
nand U14938 (N_14938,N_14825,N_14783);
and U14939 (N_14939,N_14758,N_14812);
and U14940 (N_14940,N_14861,N_14754);
or U14941 (N_14941,N_14771,N_14855);
nand U14942 (N_14942,N_14815,N_14823);
or U14943 (N_14943,N_14764,N_14776);
nand U14944 (N_14944,N_14775,N_14797);
and U14945 (N_14945,N_14836,N_14835);
nor U14946 (N_14946,N_14845,N_14828);
nand U14947 (N_14947,N_14796,N_14785);
or U14948 (N_14948,N_14845,N_14807);
nand U14949 (N_14949,N_14861,N_14852);
nand U14950 (N_14950,N_14841,N_14827);
and U14951 (N_14951,N_14759,N_14868);
nand U14952 (N_14952,N_14793,N_14867);
nor U14953 (N_14953,N_14828,N_14762);
and U14954 (N_14954,N_14823,N_14820);
nor U14955 (N_14955,N_14824,N_14762);
nor U14956 (N_14956,N_14751,N_14865);
nor U14957 (N_14957,N_14767,N_14768);
nor U14958 (N_14958,N_14798,N_14818);
nand U14959 (N_14959,N_14858,N_14803);
nand U14960 (N_14960,N_14755,N_14826);
or U14961 (N_14961,N_14772,N_14801);
or U14962 (N_14962,N_14800,N_14839);
nor U14963 (N_14963,N_14856,N_14817);
xor U14964 (N_14964,N_14826,N_14764);
and U14965 (N_14965,N_14755,N_14754);
or U14966 (N_14966,N_14792,N_14852);
nor U14967 (N_14967,N_14822,N_14828);
nor U14968 (N_14968,N_14781,N_14822);
or U14969 (N_14969,N_14840,N_14823);
nand U14970 (N_14970,N_14808,N_14854);
or U14971 (N_14971,N_14763,N_14788);
and U14972 (N_14972,N_14838,N_14758);
nor U14973 (N_14973,N_14866,N_14867);
or U14974 (N_14974,N_14780,N_14874);
nand U14975 (N_14975,N_14812,N_14849);
nor U14976 (N_14976,N_14767,N_14844);
and U14977 (N_14977,N_14766,N_14791);
and U14978 (N_14978,N_14792,N_14773);
nand U14979 (N_14979,N_14753,N_14798);
nand U14980 (N_14980,N_14812,N_14778);
nand U14981 (N_14981,N_14789,N_14795);
nor U14982 (N_14982,N_14845,N_14780);
xor U14983 (N_14983,N_14774,N_14796);
nand U14984 (N_14984,N_14767,N_14850);
or U14985 (N_14985,N_14754,N_14862);
or U14986 (N_14986,N_14771,N_14825);
and U14987 (N_14987,N_14824,N_14788);
nor U14988 (N_14988,N_14846,N_14851);
or U14989 (N_14989,N_14859,N_14812);
or U14990 (N_14990,N_14809,N_14847);
nor U14991 (N_14991,N_14817,N_14789);
and U14992 (N_14992,N_14840,N_14836);
and U14993 (N_14993,N_14841,N_14755);
and U14994 (N_14994,N_14844,N_14859);
and U14995 (N_14995,N_14824,N_14774);
and U14996 (N_14996,N_14851,N_14750);
and U14997 (N_14997,N_14769,N_14797);
or U14998 (N_14998,N_14828,N_14755);
nor U14999 (N_14999,N_14767,N_14831);
and UO_0 (O_0,N_14876,N_14942);
nand UO_1 (O_1,N_14902,N_14933);
nand UO_2 (O_2,N_14934,N_14915);
or UO_3 (O_3,N_14940,N_14922);
or UO_4 (O_4,N_14875,N_14980);
xor UO_5 (O_5,N_14919,N_14981);
nor UO_6 (O_6,N_14959,N_14968);
nor UO_7 (O_7,N_14932,N_14889);
nand UO_8 (O_8,N_14900,N_14991);
xnor UO_9 (O_9,N_14949,N_14951);
and UO_10 (O_10,N_14917,N_14995);
nor UO_11 (O_11,N_14946,N_14975);
nand UO_12 (O_12,N_14903,N_14910);
nand UO_13 (O_13,N_14924,N_14978);
and UO_14 (O_14,N_14996,N_14888);
or UO_15 (O_15,N_14967,N_14935);
xnor UO_16 (O_16,N_14882,N_14918);
and UO_17 (O_17,N_14899,N_14971);
and UO_18 (O_18,N_14984,N_14986);
nand UO_19 (O_19,N_14947,N_14972);
nor UO_20 (O_20,N_14927,N_14916);
nor UO_21 (O_21,N_14963,N_14880);
nor UO_22 (O_22,N_14988,N_14878);
nor UO_23 (O_23,N_14923,N_14952);
xnor UO_24 (O_24,N_14944,N_14969);
xor UO_25 (O_25,N_14936,N_14964);
nor UO_26 (O_26,N_14974,N_14904);
or UO_27 (O_27,N_14913,N_14891);
or UO_28 (O_28,N_14905,N_14877);
nor UO_29 (O_29,N_14911,N_14901);
nor UO_30 (O_30,N_14983,N_14896);
nand UO_31 (O_31,N_14884,N_14937);
or UO_32 (O_32,N_14982,N_14973);
and UO_33 (O_33,N_14998,N_14907);
or UO_34 (O_34,N_14939,N_14997);
nor UO_35 (O_35,N_14914,N_14926);
or UO_36 (O_36,N_14931,N_14925);
and UO_37 (O_37,N_14886,N_14881);
nand UO_38 (O_38,N_14883,N_14938);
or UO_39 (O_39,N_14885,N_14989);
or UO_40 (O_40,N_14957,N_14950);
nand UO_41 (O_41,N_14943,N_14999);
or UO_42 (O_42,N_14893,N_14992);
xnor UO_43 (O_43,N_14953,N_14956);
nand UO_44 (O_44,N_14928,N_14894);
and UO_45 (O_45,N_14908,N_14929);
or UO_46 (O_46,N_14898,N_14993);
and UO_47 (O_47,N_14948,N_14909);
and UO_48 (O_48,N_14990,N_14945);
or UO_49 (O_49,N_14892,N_14890);
and UO_50 (O_50,N_14895,N_14958);
xnor UO_51 (O_51,N_14961,N_14977);
or UO_52 (O_52,N_14930,N_14954);
or UO_53 (O_53,N_14912,N_14960);
nor UO_54 (O_54,N_14966,N_14906);
or UO_55 (O_55,N_14920,N_14941);
nor UO_56 (O_56,N_14987,N_14985);
and UO_57 (O_57,N_14965,N_14979);
or UO_58 (O_58,N_14887,N_14970);
nand UO_59 (O_59,N_14955,N_14879);
nor UO_60 (O_60,N_14921,N_14994);
nor UO_61 (O_61,N_14897,N_14976);
and UO_62 (O_62,N_14962,N_14954);
nor UO_63 (O_63,N_14961,N_14893);
nor UO_64 (O_64,N_14936,N_14960);
nand UO_65 (O_65,N_14880,N_14986);
xor UO_66 (O_66,N_14971,N_14998);
nor UO_67 (O_67,N_14890,N_14920);
nand UO_68 (O_68,N_14887,N_14917);
nand UO_69 (O_69,N_14964,N_14891);
nand UO_70 (O_70,N_14965,N_14924);
xnor UO_71 (O_71,N_14931,N_14949);
nor UO_72 (O_72,N_14963,N_14943);
nor UO_73 (O_73,N_14887,N_14928);
nand UO_74 (O_74,N_14979,N_14926);
xnor UO_75 (O_75,N_14942,N_14991);
nor UO_76 (O_76,N_14994,N_14918);
and UO_77 (O_77,N_14949,N_14984);
or UO_78 (O_78,N_14910,N_14899);
nand UO_79 (O_79,N_14943,N_14972);
nand UO_80 (O_80,N_14931,N_14932);
and UO_81 (O_81,N_14905,N_14895);
or UO_82 (O_82,N_14906,N_14902);
nand UO_83 (O_83,N_14951,N_14995);
nor UO_84 (O_84,N_14994,N_14931);
nand UO_85 (O_85,N_14890,N_14996);
and UO_86 (O_86,N_14992,N_14920);
nor UO_87 (O_87,N_14900,N_14883);
xnor UO_88 (O_88,N_14883,N_14917);
nor UO_89 (O_89,N_14938,N_14954);
and UO_90 (O_90,N_14985,N_14974);
nor UO_91 (O_91,N_14875,N_14878);
nor UO_92 (O_92,N_14895,N_14998);
xor UO_93 (O_93,N_14951,N_14983);
or UO_94 (O_94,N_14921,N_14961);
nor UO_95 (O_95,N_14919,N_14949);
nor UO_96 (O_96,N_14988,N_14970);
and UO_97 (O_97,N_14928,N_14893);
nor UO_98 (O_98,N_14987,N_14888);
nor UO_99 (O_99,N_14904,N_14921);
or UO_100 (O_100,N_14937,N_14878);
xor UO_101 (O_101,N_14927,N_14906);
xor UO_102 (O_102,N_14933,N_14934);
and UO_103 (O_103,N_14975,N_14889);
nand UO_104 (O_104,N_14942,N_14984);
nor UO_105 (O_105,N_14896,N_14987);
and UO_106 (O_106,N_14880,N_14878);
or UO_107 (O_107,N_14936,N_14968);
and UO_108 (O_108,N_14901,N_14915);
xnor UO_109 (O_109,N_14969,N_14991);
nand UO_110 (O_110,N_14961,N_14887);
nand UO_111 (O_111,N_14891,N_14980);
or UO_112 (O_112,N_14961,N_14938);
nor UO_113 (O_113,N_14930,N_14903);
and UO_114 (O_114,N_14898,N_14881);
nor UO_115 (O_115,N_14989,N_14882);
nand UO_116 (O_116,N_14900,N_14945);
or UO_117 (O_117,N_14952,N_14877);
or UO_118 (O_118,N_14887,N_14888);
and UO_119 (O_119,N_14875,N_14992);
nand UO_120 (O_120,N_14914,N_14995);
and UO_121 (O_121,N_14965,N_14878);
xnor UO_122 (O_122,N_14899,N_14905);
nor UO_123 (O_123,N_14953,N_14972);
nor UO_124 (O_124,N_14905,N_14988);
and UO_125 (O_125,N_14899,N_14978);
or UO_126 (O_126,N_14975,N_14971);
nor UO_127 (O_127,N_14887,N_14923);
xor UO_128 (O_128,N_14972,N_14882);
nand UO_129 (O_129,N_14978,N_14931);
and UO_130 (O_130,N_14914,N_14886);
and UO_131 (O_131,N_14876,N_14930);
nor UO_132 (O_132,N_14910,N_14889);
nor UO_133 (O_133,N_14877,N_14919);
nand UO_134 (O_134,N_14912,N_14994);
nand UO_135 (O_135,N_14953,N_14917);
xnor UO_136 (O_136,N_14939,N_14975);
nor UO_137 (O_137,N_14878,N_14978);
and UO_138 (O_138,N_14979,N_14992);
nor UO_139 (O_139,N_14905,N_14898);
nor UO_140 (O_140,N_14980,N_14913);
or UO_141 (O_141,N_14979,N_14959);
or UO_142 (O_142,N_14903,N_14885);
nand UO_143 (O_143,N_14956,N_14919);
or UO_144 (O_144,N_14909,N_14913);
nor UO_145 (O_145,N_14931,N_14980);
xnor UO_146 (O_146,N_14920,N_14931);
and UO_147 (O_147,N_14990,N_14919);
xor UO_148 (O_148,N_14902,N_14934);
nand UO_149 (O_149,N_14936,N_14975);
nand UO_150 (O_150,N_14918,N_14877);
xor UO_151 (O_151,N_14982,N_14988);
nand UO_152 (O_152,N_14888,N_14983);
or UO_153 (O_153,N_14986,N_14875);
nand UO_154 (O_154,N_14985,N_14941);
and UO_155 (O_155,N_14932,N_14958);
and UO_156 (O_156,N_14978,N_14894);
nand UO_157 (O_157,N_14941,N_14970);
nand UO_158 (O_158,N_14900,N_14997);
nor UO_159 (O_159,N_14879,N_14953);
and UO_160 (O_160,N_14938,N_14902);
xor UO_161 (O_161,N_14877,N_14907);
xor UO_162 (O_162,N_14941,N_14950);
xnor UO_163 (O_163,N_14971,N_14923);
nor UO_164 (O_164,N_14972,N_14924);
and UO_165 (O_165,N_14990,N_14940);
and UO_166 (O_166,N_14997,N_14975);
nand UO_167 (O_167,N_14971,N_14977);
xor UO_168 (O_168,N_14991,N_14923);
nand UO_169 (O_169,N_14979,N_14970);
or UO_170 (O_170,N_14989,N_14915);
nor UO_171 (O_171,N_14934,N_14955);
and UO_172 (O_172,N_14892,N_14938);
and UO_173 (O_173,N_14938,N_14987);
nand UO_174 (O_174,N_14889,N_14880);
nand UO_175 (O_175,N_14921,N_14938);
nand UO_176 (O_176,N_14981,N_14933);
nand UO_177 (O_177,N_14895,N_14976);
or UO_178 (O_178,N_14889,N_14973);
xor UO_179 (O_179,N_14971,N_14937);
nor UO_180 (O_180,N_14944,N_14906);
xnor UO_181 (O_181,N_14930,N_14938);
nor UO_182 (O_182,N_14953,N_14944);
or UO_183 (O_183,N_14881,N_14944);
or UO_184 (O_184,N_14987,N_14892);
nor UO_185 (O_185,N_14879,N_14905);
and UO_186 (O_186,N_14882,N_14925);
and UO_187 (O_187,N_14930,N_14936);
nor UO_188 (O_188,N_14938,N_14996);
or UO_189 (O_189,N_14930,N_14996);
nand UO_190 (O_190,N_14925,N_14988);
or UO_191 (O_191,N_14965,N_14977);
and UO_192 (O_192,N_14886,N_14976);
nand UO_193 (O_193,N_14888,N_14884);
nor UO_194 (O_194,N_14983,N_14958);
nor UO_195 (O_195,N_14901,N_14954);
and UO_196 (O_196,N_14901,N_14877);
and UO_197 (O_197,N_14895,N_14962);
nor UO_198 (O_198,N_14974,N_14925);
and UO_199 (O_199,N_14896,N_14966);
nor UO_200 (O_200,N_14896,N_14995);
nand UO_201 (O_201,N_14973,N_14922);
or UO_202 (O_202,N_14892,N_14976);
or UO_203 (O_203,N_14993,N_14962);
xnor UO_204 (O_204,N_14995,N_14877);
nand UO_205 (O_205,N_14949,N_14945);
nand UO_206 (O_206,N_14929,N_14996);
nand UO_207 (O_207,N_14917,N_14928);
or UO_208 (O_208,N_14977,N_14988);
nand UO_209 (O_209,N_14917,N_14973);
nand UO_210 (O_210,N_14897,N_14931);
nand UO_211 (O_211,N_14887,N_14994);
and UO_212 (O_212,N_14877,N_14902);
xnor UO_213 (O_213,N_14893,N_14906);
or UO_214 (O_214,N_14879,N_14907);
or UO_215 (O_215,N_14996,N_14993);
nor UO_216 (O_216,N_14947,N_14895);
and UO_217 (O_217,N_14940,N_14929);
and UO_218 (O_218,N_14923,N_14960);
and UO_219 (O_219,N_14942,N_14900);
and UO_220 (O_220,N_14987,N_14893);
nor UO_221 (O_221,N_14954,N_14885);
nor UO_222 (O_222,N_14916,N_14948);
nand UO_223 (O_223,N_14877,N_14981);
nor UO_224 (O_224,N_14978,N_14919);
and UO_225 (O_225,N_14954,N_14948);
xnor UO_226 (O_226,N_14963,N_14906);
nand UO_227 (O_227,N_14878,N_14920);
nor UO_228 (O_228,N_14946,N_14905);
nor UO_229 (O_229,N_14947,N_14990);
and UO_230 (O_230,N_14962,N_14997);
or UO_231 (O_231,N_14953,N_14886);
nand UO_232 (O_232,N_14910,N_14911);
or UO_233 (O_233,N_14975,N_14965);
nand UO_234 (O_234,N_14884,N_14971);
xnor UO_235 (O_235,N_14900,N_14932);
and UO_236 (O_236,N_14890,N_14917);
or UO_237 (O_237,N_14989,N_14955);
nor UO_238 (O_238,N_14911,N_14947);
xor UO_239 (O_239,N_14933,N_14901);
xnor UO_240 (O_240,N_14966,N_14935);
nor UO_241 (O_241,N_14960,N_14980);
nor UO_242 (O_242,N_14974,N_14989);
nor UO_243 (O_243,N_14984,N_14963);
or UO_244 (O_244,N_14931,N_14884);
xnor UO_245 (O_245,N_14877,N_14931);
nand UO_246 (O_246,N_14917,N_14974);
nand UO_247 (O_247,N_14901,N_14913);
nor UO_248 (O_248,N_14953,N_14991);
nor UO_249 (O_249,N_14970,N_14956);
nand UO_250 (O_250,N_14958,N_14927);
nand UO_251 (O_251,N_14916,N_14984);
nand UO_252 (O_252,N_14913,N_14967);
nor UO_253 (O_253,N_14991,N_14908);
and UO_254 (O_254,N_14983,N_14915);
and UO_255 (O_255,N_14988,N_14944);
or UO_256 (O_256,N_14904,N_14945);
and UO_257 (O_257,N_14963,N_14925);
and UO_258 (O_258,N_14891,N_14941);
nand UO_259 (O_259,N_14905,N_14976);
nor UO_260 (O_260,N_14879,N_14903);
and UO_261 (O_261,N_14938,N_14878);
nand UO_262 (O_262,N_14934,N_14939);
or UO_263 (O_263,N_14945,N_14991);
and UO_264 (O_264,N_14963,N_14875);
xor UO_265 (O_265,N_14941,N_14885);
nor UO_266 (O_266,N_14961,N_14900);
and UO_267 (O_267,N_14989,N_14904);
and UO_268 (O_268,N_14966,N_14984);
or UO_269 (O_269,N_14921,N_14876);
and UO_270 (O_270,N_14889,N_14928);
or UO_271 (O_271,N_14907,N_14881);
or UO_272 (O_272,N_14948,N_14985);
nand UO_273 (O_273,N_14931,N_14957);
and UO_274 (O_274,N_14914,N_14887);
nor UO_275 (O_275,N_14912,N_14983);
nand UO_276 (O_276,N_14981,N_14948);
or UO_277 (O_277,N_14920,N_14928);
or UO_278 (O_278,N_14877,N_14994);
or UO_279 (O_279,N_14896,N_14917);
and UO_280 (O_280,N_14909,N_14995);
or UO_281 (O_281,N_14991,N_14903);
nor UO_282 (O_282,N_14917,N_14879);
nor UO_283 (O_283,N_14906,N_14881);
nand UO_284 (O_284,N_14898,N_14988);
nor UO_285 (O_285,N_14993,N_14938);
xnor UO_286 (O_286,N_14900,N_14933);
and UO_287 (O_287,N_14908,N_14900);
xnor UO_288 (O_288,N_14948,N_14999);
or UO_289 (O_289,N_14901,N_14918);
nand UO_290 (O_290,N_14919,N_14915);
nor UO_291 (O_291,N_14889,N_14884);
nor UO_292 (O_292,N_14950,N_14877);
nand UO_293 (O_293,N_14935,N_14949);
nor UO_294 (O_294,N_14943,N_14975);
or UO_295 (O_295,N_14937,N_14963);
and UO_296 (O_296,N_14911,N_14921);
nand UO_297 (O_297,N_14996,N_14947);
or UO_298 (O_298,N_14930,N_14922);
and UO_299 (O_299,N_14955,N_14976);
nand UO_300 (O_300,N_14947,N_14899);
nor UO_301 (O_301,N_14970,N_14908);
and UO_302 (O_302,N_14942,N_14914);
xor UO_303 (O_303,N_14951,N_14880);
or UO_304 (O_304,N_14896,N_14877);
or UO_305 (O_305,N_14898,N_14915);
nor UO_306 (O_306,N_14956,N_14982);
and UO_307 (O_307,N_14886,N_14929);
or UO_308 (O_308,N_14938,N_14884);
xor UO_309 (O_309,N_14875,N_14964);
and UO_310 (O_310,N_14911,N_14889);
nand UO_311 (O_311,N_14958,N_14898);
or UO_312 (O_312,N_14930,N_14940);
or UO_313 (O_313,N_14979,N_14925);
and UO_314 (O_314,N_14988,N_14909);
or UO_315 (O_315,N_14990,N_14910);
nand UO_316 (O_316,N_14990,N_14892);
and UO_317 (O_317,N_14968,N_14942);
and UO_318 (O_318,N_14929,N_14914);
xor UO_319 (O_319,N_14905,N_14920);
and UO_320 (O_320,N_14929,N_14972);
xnor UO_321 (O_321,N_14883,N_14902);
and UO_322 (O_322,N_14935,N_14917);
nand UO_323 (O_323,N_14929,N_14976);
and UO_324 (O_324,N_14882,N_14963);
nor UO_325 (O_325,N_14982,N_14942);
or UO_326 (O_326,N_14934,N_14974);
or UO_327 (O_327,N_14978,N_14965);
nor UO_328 (O_328,N_14971,N_14913);
nand UO_329 (O_329,N_14921,N_14883);
nand UO_330 (O_330,N_14917,N_14940);
and UO_331 (O_331,N_14963,N_14964);
or UO_332 (O_332,N_14940,N_14881);
or UO_333 (O_333,N_14946,N_14972);
nor UO_334 (O_334,N_14985,N_14906);
nand UO_335 (O_335,N_14913,N_14894);
and UO_336 (O_336,N_14927,N_14903);
and UO_337 (O_337,N_14908,N_14982);
nand UO_338 (O_338,N_14942,N_14954);
nor UO_339 (O_339,N_14885,N_14876);
nand UO_340 (O_340,N_14983,N_14909);
and UO_341 (O_341,N_14912,N_14891);
nand UO_342 (O_342,N_14973,N_14956);
or UO_343 (O_343,N_14919,N_14955);
nand UO_344 (O_344,N_14932,N_14892);
xor UO_345 (O_345,N_14993,N_14909);
nand UO_346 (O_346,N_14950,N_14948);
nand UO_347 (O_347,N_14953,N_14955);
nor UO_348 (O_348,N_14965,N_14959);
nor UO_349 (O_349,N_14957,N_14973);
or UO_350 (O_350,N_14895,N_14900);
nand UO_351 (O_351,N_14907,N_14950);
and UO_352 (O_352,N_14928,N_14921);
and UO_353 (O_353,N_14905,N_14979);
xor UO_354 (O_354,N_14898,N_14883);
or UO_355 (O_355,N_14875,N_14945);
nor UO_356 (O_356,N_14937,N_14981);
and UO_357 (O_357,N_14940,N_14877);
and UO_358 (O_358,N_14988,N_14959);
nor UO_359 (O_359,N_14965,N_14905);
or UO_360 (O_360,N_14954,N_14900);
and UO_361 (O_361,N_14907,N_14957);
nor UO_362 (O_362,N_14990,N_14904);
and UO_363 (O_363,N_14883,N_14907);
nor UO_364 (O_364,N_14917,N_14913);
or UO_365 (O_365,N_14908,N_14896);
nor UO_366 (O_366,N_14918,N_14897);
and UO_367 (O_367,N_14920,N_14975);
xor UO_368 (O_368,N_14944,N_14937);
nor UO_369 (O_369,N_14967,N_14920);
and UO_370 (O_370,N_14958,N_14940);
xnor UO_371 (O_371,N_14947,N_14956);
and UO_372 (O_372,N_14893,N_14927);
or UO_373 (O_373,N_14918,N_14931);
nand UO_374 (O_374,N_14928,N_14924);
nand UO_375 (O_375,N_14875,N_14895);
nor UO_376 (O_376,N_14942,N_14979);
or UO_377 (O_377,N_14892,N_14921);
nor UO_378 (O_378,N_14992,N_14901);
and UO_379 (O_379,N_14880,N_14920);
and UO_380 (O_380,N_14945,N_14962);
nand UO_381 (O_381,N_14939,N_14936);
nand UO_382 (O_382,N_14995,N_14993);
xor UO_383 (O_383,N_14914,N_14978);
xor UO_384 (O_384,N_14932,N_14904);
or UO_385 (O_385,N_14967,N_14888);
or UO_386 (O_386,N_14907,N_14956);
nor UO_387 (O_387,N_14946,N_14983);
nand UO_388 (O_388,N_14910,N_14992);
or UO_389 (O_389,N_14954,N_14979);
or UO_390 (O_390,N_14948,N_14932);
and UO_391 (O_391,N_14878,N_14971);
and UO_392 (O_392,N_14898,N_14951);
and UO_393 (O_393,N_14963,N_14987);
and UO_394 (O_394,N_14990,N_14961);
and UO_395 (O_395,N_14995,N_14999);
or UO_396 (O_396,N_14974,N_14967);
nor UO_397 (O_397,N_14946,N_14979);
or UO_398 (O_398,N_14922,N_14915);
nor UO_399 (O_399,N_14925,N_14908);
or UO_400 (O_400,N_14949,N_14987);
or UO_401 (O_401,N_14954,N_14925);
nand UO_402 (O_402,N_14899,N_14962);
nand UO_403 (O_403,N_14926,N_14909);
and UO_404 (O_404,N_14934,N_14908);
nand UO_405 (O_405,N_14937,N_14975);
xnor UO_406 (O_406,N_14882,N_14941);
and UO_407 (O_407,N_14906,N_14939);
and UO_408 (O_408,N_14981,N_14954);
nor UO_409 (O_409,N_14912,N_14986);
nor UO_410 (O_410,N_14993,N_14900);
and UO_411 (O_411,N_14920,N_14997);
or UO_412 (O_412,N_14976,N_14946);
nor UO_413 (O_413,N_14953,N_14911);
nand UO_414 (O_414,N_14926,N_14975);
nor UO_415 (O_415,N_14954,N_14991);
nand UO_416 (O_416,N_14885,N_14913);
and UO_417 (O_417,N_14921,N_14924);
nor UO_418 (O_418,N_14944,N_14934);
and UO_419 (O_419,N_14968,N_14991);
or UO_420 (O_420,N_14910,N_14912);
xor UO_421 (O_421,N_14976,N_14896);
xnor UO_422 (O_422,N_14906,N_14924);
nand UO_423 (O_423,N_14956,N_14955);
xor UO_424 (O_424,N_14906,N_14992);
or UO_425 (O_425,N_14936,N_14927);
and UO_426 (O_426,N_14933,N_14951);
or UO_427 (O_427,N_14986,N_14955);
or UO_428 (O_428,N_14982,N_14921);
nand UO_429 (O_429,N_14985,N_14953);
nand UO_430 (O_430,N_14974,N_14994);
and UO_431 (O_431,N_14921,N_14905);
or UO_432 (O_432,N_14987,N_14881);
or UO_433 (O_433,N_14954,N_14933);
nand UO_434 (O_434,N_14953,N_14934);
or UO_435 (O_435,N_14921,N_14912);
or UO_436 (O_436,N_14967,N_14879);
nor UO_437 (O_437,N_14953,N_14951);
and UO_438 (O_438,N_14948,N_14886);
or UO_439 (O_439,N_14922,N_14955);
nand UO_440 (O_440,N_14935,N_14989);
xnor UO_441 (O_441,N_14919,N_14909);
nor UO_442 (O_442,N_14922,N_14954);
and UO_443 (O_443,N_14979,N_14975);
xor UO_444 (O_444,N_14914,N_14960);
xnor UO_445 (O_445,N_14942,N_14970);
xnor UO_446 (O_446,N_14943,N_14944);
nand UO_447 (O_447,N_14944,N_14931);
nand UO_448 (O_448,N_14999,N_14897);
nor UO_449 (O_449,N_14956,N_14978);
nor UO_450 (O_450,N_14908,N_14950);
and UO_451 (O_451,N_14944,N_14933);
nor UO_452 (O_452,N_14949,N_14926);
xor UO_453 (O_453,N_14968,N_14963);
nand UO_454 (O_454,N_14942,N_14929);
nand UO_455 (O_455,N_14991,N_14997);
and UO_456 (O_456,N_14988,N_14973);
nand UO_457 (O_457,N_14907,N_14886);
and UO_458 (O_458,N_14932,N_14911);
nand UO_459 (O_459,N_14966,N_14949);
or UO_460 (O_460,N_14949,N_14886);
or UO_461 (O_461,N_14961,N_14927);
xnor UO_462 (O_462,N_14921,N_14887);
nor UO_463 (O_463,N_14989,N_14961);
nor UO_464 (O_464,N_14999,N_14985);
nand UO_465 (O_465,N_14993,N_14896);
nand UO_466 (O_466,N_14916,N_14898);
or UO_467 (O_467,N_14934,N_14935);
and UO_468 (O_468,N_14985,N_14950);
and UO_469 (O_469,N_14951,N_14972);
or UO_470 (O_470,N_14915,N_14914);
nor UO_471 (O_471,N_14931,N_14876);
or UO_472 (O_472,N_14898,N_14908);
and UO_473 (O_473,N_14968,N_14920);
and UO_474 (O_474,N_14902,N_14901);
and UO_475 (O_475,N_14904,N_14957);
nand UO_476 (O_476,N_14995,N_14972);
nor UO_477 (O_477,N_14977,N_14889);
nor UO_478 (O_478,N_14909,N_14887);
nand UO_479 (O_479,N_14978,N_14964);
nor UO_480 (O_480,N_14920,N_14907);
or UO_481 (O_481,N_14903,N_14875);
and UO_482 (O_482,N_14887,N_14999);
nor UO_483 (O_483,N_14973,N_14897);
and UO_484 (O_484,N_14979,N_14939);
xnor UO_485 (O_485,N_14951,N_14942);
nand UO_486 (O_486,N_14914,N_14893);
or UO_487 (O_487,N_14977,N_14985);
and UO_488 (O_488,N_14932,N_14908);
and UO_489 (O_489,N_14964,N_14948);
and UO_490 (O_490,N_14935,N_14971);
nor UO_491 (O_491,N_14991,N_14964);
nor UO_492 (O_492,N_14971,N_14896);
nor UO_493 (O_493,N_14936,N_14894);
or UO_494 (O_494,N_14890,N_14919);
or UO_495 (O_495,N_14885,N_14924);
nor UO_496 (O_496,N_14999,N_14883);
or UO_497 (O_497,N_14940,N_14969);
or UO_498 (O_498,N_14943,N_14947);
and UO_499 (O_499,N_14884,N_14985);
nor UO_500 (O_500,N_14988,N_14961);
or UO_501 (O_501,N_14902,N_14981);
and UO_502 (O_502,N_14895,N_14925);
nand UO_503 (O_503,N_14949,N_14906);
and UO_504 (O_504,N_14945,N_14973);
xor UO_505 (O_505,N_14882,N_14947);
nor UO_506 (O_506,N_14908,N_14892);
nor UO_507 (O_507,N_14897,N_14990);
and UO_508 (O_508,N_14940,N_14882);
nor UO_509 (O_509,N_14973,N_14993);
nand UO_510 (O_510,N_14956,N_14975);
nand UO_511 (O_511,N_14931,N_14987);
nand UO_512 (O_512,N_14996,N_14988);
and UO_513 (O_513,N_14951,N_14895);
nor UO_514 (O_514,N_14972,N_14923);
or UO_515 (O_515,N_14900,N_14949);
nand UO_516 (O_516,N_14944,N_14985);
nor UO_517 (O_517,N_14959,N_14904);
nand UO_518 (O_518,N_14952,N_14958);
nor UO_519 (O_519,N_14936,N_14971);
nor UO_520 (O_520,N_14901,N_14912);
nor UO_521 (O_521,N_14928,N_14910);
nand UO_522 (O_522,N_14877,N_14897);
or UO_523 (O_523,N_14971,N_14942);
and UO_524 (O_524,N_14930,N_14935);
or UO_525 (O_525,N_14934,N_14975);
nor UO_526 (O_526,N_14992,N_14879);
nand UO_527 (O_527,N_14879,N_14901);
and UO_528 (O_528,N_14883,N_14880);
nand UO_529 (O_529,N_14976,N_14888);
or UO_530 (O_530,N_14941,N_14957);
nand UO_531 (O_531,N_14927,N_14922);
and UO_532 (O_532,N_14891,N_14928);
nand UO_533 (O_533,N_14998,N_14920);
nor UO_534 (O_534,N_14993,N_14985);
or UO_535 (O_535,N_14892,N_14933);
or UO_536 (O_536,N_14881,N_14885);
and UO_537 (O_537,N_14888,N_14878);
nand UO_538 (O_538,N_14877,N_14921);
nand UO_539 (O_539,N_14956,N_14897);
and UO_540 (O_540,N_14991,N_14905);
or UO_541 (O_541,N_14956,N_14985);
and UO_542 (O_542,N_14876,N_14974);
or UO_543 (O_543,N_14985,N_14980);
or UO_544 (O_544,N_14938,N_14978);
nor UO_545 (O_545,N_14959,N_14946);
nand UO_546 (O_546,N_14946,N_14895);
nor UO_547 (O_547,N_14924,N_14976);
or UO_548 (O_548,N_14885,N_14877);
nand UO_549 (O_549,N_14924,N_14999);
or UO_550 (O_550,N_14996,N_14990);
and UO_551 (O_551,N_14984,N_14894);
nor UO_552 (O_552,N_14944,N_14940);
or UO_553 (O_553,N_14992,N_14961);
and UO_554 (O_554,N_14967,N_14948);
nand UO_555 (O_555,N_14957,N_14939);
nand UO_556 (O_556,N_14982,N_14984);
nor UO_557 (O_557,N_14882,N_14945);
and UO_558 (O_558,N_14969,N_14989);
nand UO_559 (O_559,N_14986,N_14964);
nor UO_560 (O_560,N_14948,N_14955);
or UO_561 (O_561,N_14875,N_14987);
or UO_562 (O_562,N_14886,N_14883);
and UO_563 (O_563,N_14987,N_14955);
and UO_564 (O_564,N_14962,N_14938);
nor UO_565 (O_565,N_14947,N_14930);
nor UO_566 (O_566,N_14940,N_14945);
nand UO_567 (O_567,N_14922,N_14942);
xnor UO_568 (O_568,N_14907,N_14909);
xor UO_569 (O_569,N_14926,N_14970);
nor UO_570 (O_570,N_14948,N_14976);
and UO_571 (O_571,N_14895,N_14943);
nand UO_572 (O_572,N_14985,N_14925);
nor UO_573 (O_573,N_14923,N_14883);
nand UO_574 (O_574,N_14903,N_14977);
and UO_575 (O_575,N_14966,N_14964);
and UO_576 (O_576,N_14919,N_14953);
or UO_577 (O_577,N_14980,N_14984);
nor UO_578 (O_578,N_14982,N_14912);
xor UO_579 (O_579,N_14954,N_14943);
nand UO_580 (O_580,N_14976,N_14925);
and UO_581 (O_581,N_14980,N_14879);
nor UO_582 (O_582,N_14946,N_14893);
or UO_583 (O_583,N_14987,N_14921);
and UO_584 (O_584,N_14890,N_14979);
or UO_585 (O_585,N_14915,N_14953);
and UO_586 (O_586,N_14957,N_14975);
or UO_587 (O_587,N_14924,N_14995);
nor UO_588 (O_588,N_14997,N_14937);
nand UO_589 (O_589,N_14923,N_14921);
nand UO_590 (O_590,N_14998,N_14988);
nand UO_591 (O_591,N_14955,N_14890);
nor UO_592 (O_592,N_14892,N_14942);
nor UO_593 (O_593,N_14976,N_14876);
nor UO_594 (O_594,N_14943,N_14909);
nor UO_595 (O_595,N_14949,N_14928);
xor UO_596 (O_596,N_14893,N_14976);
nor UO_597 (O_597,N_14971,N_14890);
and UO_598 (O_598,N_14877,N_14963);
nand UO_599 (O_599,N_14958,N_14992);
or UO_600 (O_600,N_14992,N_14956);
nand UO_601 (O_601,N_14992,N_14997);
or UO_602 (O_602,N_14958,N_14994);
nor UO_603 (O_603,N_14962,N_14977);
and UO_604 (O_604,N_14967,N_14956);
nand UO_605 (O_605,N_14905,N_14978);
and UO_606 (O_606,N_14899,N_14995);
nor UO_607 (O_607,N_14960,N_14939);
and UO_608 (O_608,N_14927,N_14971);
nor UO_609 (O_609,N_14902,N_14912);
or UO_610 (O_610,N_14978,N_14927);
and UO_611 (O_611,N_14902,N_14882);
nor UO_612 (O_612,N_14953,N_14950);
or UO_613 (O_613,N_14890,N_14930);
and UO_614 (O_614,N_14972,N_14954);
nor UO_615 (O_615,N_14939,N_14897);
or UO_616 (O_616,N_14952,N_14928);
nor UO_617 (O_617,N_14935,N_14927);
nand UO_618 (O_618,N_14943,N_14969);
nand UO_619 (O_619,N_14925,N_14929);
and UO_620 (O_620,N_14902,N_14961);
xnor UO_621 (O_621,N_14882,N_14890);
nand UO_622 (O_622,N_14987,N_14953);
and UO_623 (O_623,N_14889,N_14965);
xnor UO_624 (O_624,N_14886,N_14969);
nor UO_625 (O_625,N_14918,N_14915);
nand UO_626 (O_626,N_14910,N_14896);
xor UO_627 (O_627,N_14919,N_14928);
nand UO_628 (O_628,N_14882,N_14891);
nand UO_629 (O_629,N_14971,N_14898);
nand UO_630 (O_630,N_14997,N_14924);
nor UO_631 (O_631,N_14898,N_14944);
xor UO_632 (O_632,N_14992,N_14938);
or UO_633 (O_633,N_14883,N_14929);
xor UO_634 (O_634,N_14939,N_14933);
nor UO_635 (O_635,N_14944,N_14907);
and UO_636 (O_636,N_14922,N_14963);
nand UO_637 (O_637,N_14910,N_14930);
or UO_638 (O_638,N_14972,N_14997);
nand UO_639 (O_639,N_14918,N_14907);
xor UO_640 (O_640,N_14986,N_14946);
and UO_641 (O_641,N_14895,N_14940);
or UO_642 (O_642,N_14912,N_14877);
and UO_643 (O_643,N_14893,N_14985);
nor UO_644 (O_644,N_14951,N_14943);
xor UO_645 (O_645,N_14905,N_14930);
or UO_646 (O_646,N_14937,N_14914);
nand UO_647 (O_647,N_14931,N_14955);
nand UO_648 (O_648,N_14968,N_14997);
or UO_649 (O_649,N_14960,N_14985);
and UO_650 (O_650,N_14996,N_14967);
nand UO_651 (O_651,N_14898,N_14899);
or UO_652 (O_652,N_14966,N_14940);
nand UO_653 (O_653,N_14959,N_14985);
nand UO_654 (O_654,N_14980,N_14896);
xnor UO_655 (O_655,N_14897,N_14919);
xor UO_656 (O_656,N_14899,N_14933);
xor UO_657 (O_657,N_14901,N_14888);
nand UO_658 (O_658,N_14971,N_14966);
nand UO_659 (O_659,N_14945,N_14902);
and UO_660 (O_660,N_14888,N_14998);
nand UO_661 (O_661,N_14920,N_14945);
nor UO_662 (O_662,N_14900,N_14947);
nor UO_663 (O_663,N_14968,N_14930);
xnor UO_664 (O_664,N_14902,N_14878);
xor UO_665 (O_665,N_14965,N_14972);
or UO_666 (O_666,N_14911,N_14998);
nand UO_667 (O_667,N_14888,N_14897);
and UO_668 (O_668,N_14996,N_14985);
xor UO_669 (O_669,N_14948,N_14891);
nand UO_670 (O_670,N_14995,N_14987);
nor UO_671 (O_671,N_14945,N_14935);
and UO_672 (O_672,N_14996,N_14926);
and UO_673 (O_673,N_14961,N_14916);
and UO_674 (O_674,N_14932,N_14947);
and UO_675 (O_675,N_14953,N_14909);
or UO_676 (O_676,N_14916,N_14892);
nand UO_677 (O_677,N_14989,N_14975);
and UO_678 (O_678,N_14916,N_14938);
nor UO_679 (O_679,N_14890,N_14964);
or UO_680 (O_680,N_14929,N_14902);
nor UO_681 (O_681,N_14985,N_14936);
xnor UO_682 (O_682,N_14878,N_14882);
or UO_683 (O_683,N_14897,N_14986);
nand UO_684 (O_684,N_14963,N_14891);
nand UO_685 (O_685,N_14913,N_14915);
or UO_686 (O_686,N_14991,N_14902);
nand UO_687 (O_687,N_14890,N_14877);
and UO_688 (O_688,N_14875,N_14877);
nand UO_689 (O_689,N_14964,N_14980);
or UO_690 (O_690,N_14892,N_14876);
nor UO_691 (O_691,N_14906,N_14876);
or UO_692 (O_692,N_14974,N_14998);
nand UO_693 (O_693,N_14977,N_14919);
nand UO_694 (O_694,N_14891,N_14937);
nand UO_695 (O_695,N_14942,N_14956);
nor UO_696 (O_696,N_14941,N_14932);
or UO_697 (O_697,N_14980,N_14967);
or UO_698 (O_698,N_14958,N_14919);
and UO_699 (O_699,N_14992,N_14981);
nand UO_700 (O_700,N_14960,N_14957);
nand UO_701 (O_701,N_14908,N_14922);
and UO_702 (O_702,N_14966,N_14977);
or UO_703 (O_703,N_14932,N_14980);
nand UO_704 (O_704,N_14932,N_14966);
or UO_705 (O_705,N_14962,N_14990);
nand UO_706 (O_706,N_14941,N_14971);
or UO_707 (O_707,N_14979,N_14931);
nor UO_708 (O_708,N_14890,N_14936);
nand UO_709 (O_709,N_14995,N_14998);
nand UO_710 (O_710,N_14984,N_14914);
nor UO_711 (O_711,N_14948,N_14958);
xor UO_712 (O_712,N_14923,N_14979);
and UO_713 (O_713,N_14954,N_14940);
or UO_714 (O_714,N_14878,N_14926);
nand UO_715 (O_715,N_14885,N_14953);
nand UO_716 (O_716,N_14907,N_14888);
or UO_717 (O_717,N_14924,N_14877);
nor UO_718 (O_718,N_14918,N_14928);
and UO_719 (O_719,N_14930,N_14960);
nor UO_720 (O_720,N_14963,N_14915);
or UO_721 (O_721,N_14885,N_14948);
nand UO_722 (O_722,N_14891,N_14956);
nand UO_723 (O_723,N_14977,N_14973);
nor UO_724 (O_724,N_14904,N_14924);
or UO_725 (O_725,N_14968,N_14993);
xor UO_726 (O_726,N_14988,N_14933);
or UO_727 (O_727,N_14990,N_14976);
nand UO_728 (O_728,N_14892,N_14997);
nand UO_729 (O_729,N_14921,N_14988);
xor UO_730 (O_730,N_14970,N_14995);
nor UO_731 (O_731,N_14934,N_14977);
and UO_732 (O_732,N_14879,N_14887);
nor UO_733 (O_733,N_14991,N_14987);
nor UO_734 (O_734,N_14998,N_14882);
nand UO_735 (O_735,N_14956,N_14911);
and UO_736 (O_736,N_14965,N_14944);
and UO_737 (O_737,N_14906,N_14970);
nor UO_738 (O_738,N_14973,N_14906);
xnor UO_739 (O_739,N_14907,N_14938);
xnor UO_740 (O_740,N_14999,N_14879);
nand UO_741 (O_741,N_14923,N_14963);
nor UO_742 (O_742,N_14959,N_14954);
nor UO_743 (O_743,N_14940,N_14889);
or UO_744 (O_744,N_14894,N_14897);
nand UO_745 (O_745,N_14953,N_14913);
nand UO_746 (O_746,N_14884,N_14921);
nand UO_747 (O_747,N_14918,N_14985);
nor UO_748 (O_748,N_14909,N_14981);
or UO_749 (O_749,N_14962,N_14910);
nor UO_750 (O_750,N_14998,N_14973);
nor UO_751 (O_751,N_14994,N_14911);
nand UO_752 (O_752,N_14920,N_14909);
or UO_753 (O_753,N_14964,N_14888);
xnor UO_754 (O_754,N_14952,N_14926);
xnor UO_755 (O_755,N_14897,N_14968);
or UO_756 (O_756,N_14893,N_14991);
or UO_757 (O_757,N_14948,N_14941);
and UO_758 (O_758,N_14924,N_14991);
or UO_759 (O_759,N_14888,N_14963);
nor UO_760 (O_760,N_14892,N_14963);
or UO_761 (O_761,N_14924,N_14907);
or UO_762 (O_762,N_14939,N_14991);
and UO_763 (O_763,N_14977,N_14883);
nand UO_764 (O_764,N_14911,N_14986);
and UO_765 (O_765,N_14913,N_14962);
and UO_766 (O_766,N_14924,N_14903);
and UO_767 (O_767,N_14987,N_14998);
nand UO_768 (O_768,N_14999,N_14962);
nand UO_769 (O_769,N_14978,N_14882);
or UO_770 (O_770,N_14955,N_14876);
nor UO_771 (O_771,N_14964,N_14922);
and UO_772 (O_772,N_14889,N_14885);
or UO_773 (O_773,N_14947,N_14944);
and UO_774 (O_774,N_14981,N_14926);
nor UO_775 (O_775,N_14902,N_14918);
and UO_776 (O_776,N_14897,N_14937);
nor UO_777 (O_777,N_14945,N_14943);
or UO_778 (O_778,N_14915,N_14892);
nor UO_779 (O_779,N_14880,N_14914);
and UO_780 (O_780,N_14946,N_14919);
and UO_781 (O_781,N_14909,N_14878);
or UO_782 (O_782,N_14939,N_14989);
or UO_783 (O_783,N_14997,N_14952);
and UO_784 (O_784,N_14880,N_14926);
nand UO_785 (O_785,N_14994,N_14998);
nand UO_786 (O_786,N_14885,N_14909);
nand UO_787 (O_787,N_14924,N_14974);
and UO_788 (O_788,N_14931,N_14907);
nor UO_789 (O_789,N_14977,N_14990);
xor UO_790 (O_790,N_14929,N_14921);
or UO_791 (O_791,N_14945,N_14890);
nor UO_792 (O_792,N_14992,N_14882);
or UO_793 (O_793,N_14892,N_14980);
nand UO_794 (O_794,N_14995,N_14920);
nand UO_795 (O_795,N_14955,N_14927);
nor UO_796 (O_796,N_14907,N_14910);
nand UO_797 (O_797,N_14918,N_14938);
or UO_798 (O_798,N_14898,N_14946);
nand UO_799 (O_799,N_14946,N_14917);
nor UO_800 (O_800,N_14907,N_14884);
nand UO_801 (O_801,N_14902,N_14899);
nor UO_802 (O_802,N_14901,N_14927);
or UO_803 (O_803,N_14880,N_14915);
nand UO_804 (O_804,N_14889,N_14899);
or UO_805 (O_805,N_14933,N_14986);
xnor UO_806 (O_806,N_14937,N_14955);
or UO_807 (O_807,N_14929,N_14954);
or UO_808 (O_808,N_14938,N_14997);
nor UO_809 (O_809,N_14896,N_14923);
and UO_810 (O_810,N_14934,N_14883);
or UO_811 (O_811,N_14978,N_14901);
nand UO_812 (O_812,N_14971,N_14918);
nor UO_813 (O_813,N_14987,N_14890);
or UO_814 (O_814,N_14916,N_14895);
and UO_815 (O_815,N_14971,N_14879);
and UO_816 (O_816,N_14939,N_14926);
and UO_817 (O_817,N_14945,N_14972);
and UO_818 (O_818,N_14944,N_14886);
nand UO_819 (O_819,N_14903,N_14936);
and UO_820 (O_820,N_14927,N_14945);
and UO_821 (O_821,N_14925,N_14957);
nand UO_822 (O_822,N_14983,N_14989);
nor UO_823 (O_823,N_14989,N_14937);
or UO_824 (O_824,N_14985,N_14975);
nor UO_825 (O_825,N_14996,N_14881);
and UO_826 (O_826,N_14960,N_14900);
nand UO_827 (O_827,N_14990,N_14885);
or UO_828 (O_828,N_14941,N_14919);
nor UO_829 (O_829,N_14914,N_14894);
or UO_830 (O_830,N_14960,N_14894);
and UO_831 (O_831,N_14980,N_14979);
nand UO_832 (O_832,N_14910,N_14898);
and UO_833 (O_833,N_14946,N_14921);
nor UO_834 (O_834,N_14896,N_14913);
nand UO_835 (O_835,N_14936,N_14879);
nand UO_836 (O_836,N_14982,N_14878);
nor UO_837 (O_837,N_14895,N_14937);
nand UO_838 (O_838,N_14917,N_14916);
and UO_839 (O_839,N_14954,N_14983);
nand UO_840 (O_840,N_14952,N_14880);
nor UO_841 (O_841,N_14980,N_14917);
or UO_842 (O_842,N_14929,N_14892);
and UO_843 (O_843,N_14908,N_14907);
or UO_844 (O_844,N_14934,N_14954);
nor UO_845 (O_845,N_14894,N_14945);
nor UO_846 (O_846,N_14897,N_14930);
or UO_847 (O_847,N_14894,N_14878);
or UO_848 (O_848,N_14935,N_14900);
nand UO_849 (O_849,N_14915,N_14957);
nor UO_850 (O_850,N_14973,N_14899);
or UO_851 (O_851,N_14939,N_14970);
and UO_852 (O_852,N_14882,N_14926);
nand UO_853 (O_853,N_14900,N_14995);
xor UO_854 (O_854,N_14917,N_14923);
nor UO_855 (O_855,N_14947,N_14890);
nand UO_856 (O_856,N_14984,N_14943);
and UO_857 (O_857,N_14982,N_14884);
nor UO_858 (O_858,N_14922,N_14980);
or UO_859 (O_859,N_14887,N_14952);
nand UO_860 (O_860,N_14902,N_14962);
nor UO_861 (O_861,N_14877,N_14937);
and UO_862 (O_862,N_14879,N_14932);
nor UO_863 (O_863,N_14985,N_14897);
nor UO_864 (O_864,N_14919,N_14988);
nand UO_865 (O_865,N_14903,N_14908);
or UO_866 (O_866,N_14958,N_14982);
and UO_867 (O_867,N_14986,N_14977);
and UO_868 (O_868,N_14963,N_14999);
or UO_869 (O_869,N_14971,N_14949);
and UO_870 (O_870,N_14889,N_14920);
and UO_871 (O_871,N_14919,N_14959);
or UO_872 (O_872,N_14983,N_14905);
or UO_873 (O_873,N_14974,N_14893);
and UO_874 (O_874,N_14935,N_14947);
nor UO_875 (O_875,N_14912,N_14913);
nor UO_876 (O_876,N_14911,N_14996);
and UO_877 (O_877,N_14923,N_14973);
and UO_878 (O_878,N_14950,N_14883);
nand UO_879 (O_879,N_14978,N_14910);
nor UO_880 (O_880,N_14886,N_14936);
xor UO_881 (O_881,N_14983,N_14987);
nand UO_882 (O_882,N_14999,N_14940);
nand UO_883 (O_883,N_14954,N_14936);
nor UO_884 (O_884,N_14896,N_14943);
xnor UO_885 (O_885,N_14989,N_14913);
and UO_886 (O_886,N_14991,N_14999);
nand UO_887 (O_887,N_14994,N_14955);
and UO_888 (O_888,N_14959,N_14948);
and UO_889 (O_889,N_14935,N_14923);
nand UO_890 (O_890,N_14935,N_14881);
or UO_891 (O_891,N_14894,N_14966);
or UO_892 (O_892,N_14943,N_14904);
nor UO_893 (O_893,N_14999,N_14959);
nor UO_894 (O_894,N_14928,N_14913);
and UO_895 (O_895,N_14961,N_14918);
or UO_896 (O_896,N_14983,N_14984);
nand UO_897 (O_897,N_14921,N_14958);
nor UO_898 (O_898,N_14965,N_14998);
nand UO_899 (O_899,N_14919,N_14975);
or UO_900 (O_900,N_14983,N_14969);
or UO_901 (O_901,N_14903,N_14972);
nor UO_902 (O_902,N_14967,N_14893);
nor UO_903 (O_903,N_14915,N_14982);
nor UO_904 (O_904,N_14960,N_14976);
or UO_905 (O_905,N_14914,N_14997);
or UO_906 (O_906,N_14965,N_14888);
nand UO_907 (O_907,N_14975,N_14885);
nand UO_908 (O_908,N_14911,N_14912);
nand UO_909 (O_909,N_14991,N_14915);
xnor UO_910 (O_910,N_14921,N_14980);
or UO_911 (O_911,N_14957,N_14905);
xnor UO_912 (O_912,N_14876,N_14970);
nand UO_913 (O_913,N_14945,N_14924);
nand UO_914 (O_914,N_14959,N_14892);
nor UO_915 (O_915,N_14954,N_14880);
nor UO_916 (O_916,N_14887,N_14933);
nor UO_917 (O_917,N_14879,N_14900);
nor UO_918 (O_918,N_14880,N_14958);
xor UO_919 (O_919,N_14923,N_14982);
nand UO_920 (O_920,N_14976,N_14982);
or UO_921 (O_921,N_14952,N_14956);
nor UO_922 (O_922,N_14920,N_14923);
nand UO_923 (O_923,N_14973,N_14910);
or UO_924 (O_924,N_14955,N_14963);
nand UO_925 (O_925,N_14881,N_14903);
and UO_926 (O_926,N_14966,N_14900);
or UO_927 (O_927,N_14898,N_14889);
and UO_928 (O_928,N_14991,N_14888);
and UO_929 (O_929,N_14910,N_14975);
or UO_930 (O_930,N_14937,N_14964);
and UO_931 (O_931,N_14915,N_14965);
nand UO_932 (O_932,N_14891,N_14927);
and UO_933 (O_933,N_14948,N_14889);
nand UO_934 (O_934,N_14911,N_14938);
nor UO_935 (O_935,N_14976,N_14903);
nand UO_936 (O_936,N_14891,N_14879);
or UO_937 (O_937,N_14933,N_14903);
nor UO_938 (O_938,N_14924,N_14966);
xor UO_939 (O_939,N_14921,N_14914);
nor UO_940 (O_940,N_14966,N_14953);
nand UO_941 (O_941,N_14943,N_14932);
xor UO_942 (O_942,N_14996,N_14899);
or UO_943 (O_943,N_14968,N_14918);
or UO_944 (O_944,N_14948,N_14974);
or UO_945 (O_945,N_14964,N_14926);
or UO_946 (O_946,N_14937,N_14976);
nor UO_947 (O_947,N_14945,N_14963);
or UO_948 (O_948,N_14984,N_14890);
nor UO_949 (O_949,N_14899,N_14943);
and UO_950 (O_950,N_14906,N_14956);
or UO_951 (O_951,N_14875,N_14911);
and UO_952 (O_952,N_14928,N_14946);
nor UO_953 (O_953,N_14992,N_14888);
nor UO_954 (O_954,N_14882,N_14919);
or UO_955 (O_955,N_14890,N_14952);
or UO_956 (O_956,N_14904,N_14998);
nand UO_957 (O_957,N_14999,N_14938);
or UO_958 (O_958,N_14938,N_14937);
and UO_959 (O_959,N_14977,N_14943);
or UO_960 (O_960,N_14992,N_14914);
and UO_961 (O_961,N_14888,N_14985);
and UO_962 (O_962,N_14923,N_14897);
xor UO_963 (O_963,N_14940,N_14901);
nor UO_964 (O_964,N_14965,N_14932);
and UO_965 (O_965,N_14927,N_14918);
nand UO_966 (O_966,N_14949,N_14910);
or UO_967 (O_967,N_14987,N_14947);
nor UO_968 (O_968,N_14921,N_14991);
nand UO_969 (O_969,N_14893,N_14905);
nor UO_970 (O_970,N_14926,N_14941);
nand UO_971 (O_971,N_14893,N_14983);
nor UO_972 (O_972,N_14987,N_14954);
and UO_973 (O_973,N_14906,N_14960);
or UO_974 (O_974,N_14985,N_14943);
nor UO_975 (O_975,N_14894,N_14906);
nand UO_976 (O_976,N_14993,N_14965);
and UO_977 (O_977,N_14952,N_14881);
nor UO_978 (O_978,N_14997,N_14928);
or UO_979 (O_979,N_14909,N_14886);
xnor UO_980 (O_980,N_14916,N_14931);
nand UO_981 (O_981,N_14906,N_14958);
nand UO_982 (O_982,N_14905,N_14972);
nor UO_983 (O_983,N_14899,N_14956);
or UO_984 (O_984,N_14959,N_14935);
or UO_985 (O_985,N_14997,N_14886);
nor UO_986 (O_986,N_14885,N_14910);
and UO_987 (O_987,N_14957,N_14902);
or UO_988 (O_988,N_14963,N_14901);
and UO_989 (O_989,N_14920,N_14921);
nand UO_990 (O_990,N_14975,N_14890);
xnor UO_991 (O_991,N_14949,N_14985);
and UO_992 (O_992,N_14896,N_14926);
xnor UO_993 (O_993,N_14892,N_14996);
nand UO_994 (O_994,N_14935,N_14914);
nand UO_995 (O_995,N_14910,N_14985);
nand UO_996 (O_996,N_14986,N_14915);
xor UO_997 (O_997,N_14999,N_14926);
xor UO_998 (O_998,N_14908,N_14958);
or UO_999 (O_999,N_14947,N_14923);
xor UO_1000 (O_1000,N_14969,N_14904);
or UO_1001 (O_1001,N_14924,N_14884);
or UO_1002 (O_1002,N_14952,N_14946);
nor UO_1003 (O_1003,N_14979,N_14986);
nand UO_1004 (O_1004,N_14901,N_14982);
nand UO_1005 (O_1005,N_14977,N_14912);
and UO_1006 (O_1006,N_14949,N_14975);
or UO_1007 (O_1007,N_14996,N_14928);
or UO_1008 (O_1008,N_14994,N_14925);
nor UO_1009 (O_1009,N_14901,N_14997);
nor UO_1010 (O_1010,N_14950,N_14958);
nand UO_1011 (O_1011,N_14951,N_14990);
xor UO_1012 (O_1012,N_14990,N_14878);
and UO_1013 (O_1013,N_14941,N_14881);
nor UO_1014 (O_1014,N_14899,N_14931);
nand UO_1015 (O_1015,N_14964,N_14887);
nand UO_1016 (O_1016,N_14920,N_14994);
or UO_1017 (O_1017,N_14912,N_14972);
or UO_1018 (O_1018,N_14923,N_14882);
xnor UO_1019 (O_1019,N_14960,N_14941);
or UO_1020 (O_1020,N_14962,N_14951);
nor UO_1021 (O_1021,N_14981,N_14940);
nand UO_1022 (O_1022,N_14912,N_14951);
nand UO_1023 (O_1023,N_14924,N_14880);
and UO_1024 (O_1024,N_14973,N_14951);
nor UO_1025 (O_1025,N_14889,N_14903);
or UO_1026 (O_1026,N_14893,N_14956);
and UO_1027 (O_1027,N_14943,N_14901);
and UO_1028 (O_1028,N_14921,N_14965);
nand UO_1029 (O_1029,N_14903,N_14880);
nor UO_1030 (O_1030,N_14960,N_14886);
nor UO_1031 (O_1031,N_14984,N_14926);
nor UO_1032 (O_1032,N_14893,N_14993);
or UO_1033 (O_1033,N_14889,N_14955);
and UO_1034 (O_1034,N_14994,N_14899);
nor UO_1035 (O_1035,N_14894,N_14983);
and UO_1036 (O_1036,N_14953,N_14931);
and UO_1037 (O_1037,N_14943,N_14957);
xor UO_1038 (O_1038,N_14940,N_14902);
nand UO_1039 (O_1039,N_14952,N_14917);
nand UO_1040 (O_1040,N_14877,N_14951);
nand UO_1041 (O_1041,N_14960,N_14910);
nand UO_1042 (O_1042,N_14921,N_14959);
or UO_1043 (O_1043,N_14957,N_14948);
nand UO_1044 (O_1044,N_14997,N_14933);
nor UO_1045 (O_1045,N_14926,N_14890);
nand UO_1046 (O_1046,N_14945,N_14983);
or UO_1047 (O_1047,N_14992,N_14939);
nand UO_1048 (O_1048,N_14937,N_14960);
nor UO_1049 (O_1049,N_14948,N_14961);
nor UO_1050 (O_1050,N_14898,N_14925);
nand UO_1051 (O_1051,N_14959,N_14966);
xor UO_1052 (O_1052,N_14966,N_14970);
nor UO_1053 (O_1053,N_14934,N_14928);
nor UO_1054 (O_1054,N_14910,N_14876);
nor UO_1055 (O_1055,N_14969,N_14937);
nand UO_1056 (O_1056,N_14929,N_14909);
or UO_1057 (O_1057,N_14915,N_14917);
or UO_1058 (O_1058,N_14886,N_14942);
nor UO_1059 (O_1059,N_14950,N_14887);
xor UO_1060 (O_1060,N_14982,N_14925);
or UO_1061 (O_1061,N_14933,N_14961);
nand UO_1062 (O_1062,N_14950,N_14942);
nor UO_1063 (O_1063,N_14917,N_14939);
or UO_1064 (O_1064,N_14963,N_14950);
or UO_1065 (O_1065,N_14978,N_14987);
nand UO_1066 (O_1066,N_14936,N_14951);
xnor UO_1067 (O_1067,N_14929,N_14920);
and UO_1068 (O_1068,N_14926,N_14918);
nor UO_1069 (O_1069,N_14903,N_14893);
and UO_1070 (O_1070,N_14923,N_14986);
and UO_1071 (O_1071,N_14907,N_14911);
and UO_1072 (O_1072,N_14990,N_14924);
nor UO_1073 (O_1073,N_14980,N_14962);
xnor UO_1074 (O_1074,N_14995,N_14910);
nor UO_1075 (O_1075,N_14916,N_14947);
nor UO_1076 (O_1076,N_14910,N_14953);
and UO_1077 (O_1077,N_14978,N_14959);
nand UO_1078 (O_1078,N_14951,N_14970);
nor UO_1079 (O_1079,N_14990,N_14916);
xor UO_1080 (O_1080,N_14975,N_14917);
nor UO_1081 (O_1081,N_14972,N_14890);
nor UO_1082 (O_1082,N_14921,N_14993);
or UO_1083 (O_1083,N_14993,N_14925);
nand UO_1084 (O_1084,N_14988,N_14989);
nand UO_1085 (O_1085,N_14956,N_14976);
nand UO_1086 (O_1086,N_14884,N_14912);
nor UO_1087 (O_1087,N_14900,N_14886);
or UO_1088 (O_1088,N_14938,N_14895);
nand UO_1089 (O_1089,N_14989,N_14970);
nand UO_1090 (O_1090,N_14943,N_14931);
or UO_1091 (O_1091,N_14889,N_14982);
nand UO_1092 (O_1092,N_14985,N_14989);
nor UO_1093 (O_1093,N_14883,N_14958);
nand UO_1094 (O_1094,N_14947,N_14915);
nor UO_1095 (O_1095,N_14946,N_14911);
and UO_1096 (O_1096,N_14932,N_14977);
nor UO_1097 (O_1097,N_14944,N_14899);
and UO_1098 (O_1098,N_14961,N_14935);
xor UO_1099 (O_1099,N_14952,N_14961);
nor UO_1100 (O_1100,N_14896,N_14875);
nand UO_1101 (O_1101,N_14906,N_14998);
or UO_1102 (O_1102,N_14945,N_14887);
and UO_1103 (O_1103,N_14920,N_14876);
or UO_1104 (O_1104,N_14948,N_14994);
nor UO_1105 (O_1105,N_14900,N_14937);
nor UO_1106 (O_1106,N_14971,N_14932);
or UO_1107 (O_1107,N_14894,N_14900);
nor UO_1108 (O_1108,N_14885,N_14878);
and UO_1109 (O_1109,N_14898,N_14892);
nor UO_1110 (O_1110,N_14947,N_14925);
xor UO_1111 (O_1111,N_14890,N_14911);
or UO_1112 (O_1112,N_14990,N_14913);
xnor UO_1113 (O_1113,N_14969,N_14942);
nand UO_1114 (O_1114,N_14893,N_14997);
nor UO_1115 (O_1115,N_14878,N_14955);
nor UO_1116 (O_1116,N_14981,N_14912);
or UO_1117 (O_1117,N_14983,N_14974);
or UO_1118 (O_1118,N_14952,N_14959);
or UO_1119 (O_1119,N_14960,N_14997);
nand UO_1120 (O_1120,N_14962,N_14946);
or UO_1121 (O_1121,N_14976,N_14920);
nand UO_1122 (O_1122,N_14997,N_14965);
and UO_1123 (O_1123,N_14978,N_14912);
and UO_1124 (O_1124,N_14969,N_14910);
or UO_1125 (O_1125,N_14979,N_14933);
nor UO_1126 (O_1126,N_14997,N_14951);
and UO_1127 (O_1127,N_14898,N_14943);
and UO_1128 (O_1128,N_14910,N_14923);
nor UO_1129 (O_1129,N_14964,N_14972);
or UO_1130 (O_1130,N_14888,N_14889);
nand UO_1131 (O_1131,N_14905,N_14926);
or UO_1132 (O_1132,N_14946,N_14920);
nand UO_1133 (O_1133,N_14901,N_14929);
or UO_1134 (O_1134,N_14983,N_14902);
and UO_1135 (O_1135,N_14875,N_14943);
nand UO_1136 (O_1136,N_14980,N_14953);
xnor UO_1137 (O_1137,N_14934,N_14926);
xor UO_1138 (O_1138,N_14928,N_14931);
nand UO_1139 (O_1139,N_14921,N_14976);
nor UO_1140 (O_1140,N_14882,N_14952);
and UO_1141 (O_1141,N_14996,N_14949);
and UO_1142 (O_1142,N_14949,N_14982);
and UO_1143 (O_1143,N_14972,N_14963);
xnor UO_1144 (O_1144,N_14892,N_14943);
or UO_1145 (O_1145,N_14904,N_14906);
and UO_1146 (O_1146,N_14911,N_14964);
and UO_1147 (O_1147,N_14966,N_14955);
nor UO_1148 (O_1148,N_14973,N_14925);
and UO_1149 (O_1149,N_14938,N_14966);
nand UO_1150 (O_1150,N_14890,N_14937);
nor UO_1151 (O_1151,N_14888,N_14926);
xnor UO_1152 (O_1152,N_14992,N_14900);
and UO_1153 (O_1153,N_14888,N_14911);
and UO_1154 (O_1154,N_14932,N_14992);
and UO_1155 (O_1155,N_14934,N_14930);
or UO_1156 (O_1156,N_14884,N_14878);
nand UO_1157 (O_1157,N_14922,N_14992);
and UO_1158 (O_1158,N_14888,N_14940);
or UO_1159 (O_1159,N_14961,N_14926);
nor UO_1160 (O_1160,N_14968,N_14980);
xor UO_1161 (O_1161,N_14933,N_14877);
nand UO_1162 (O_1162,N_14992,N_14890);
and UO_1163 (O_1163,N_14913,N_14988);
and UO_1164 (O_1164,N_14907,N_14970);
and UO_1165 (O_1165,N_14997,N_14963);
nor UO_1166 (O_1166,N_14964,N_14976);
nor UO_1167 (O_1167,N_14939,N_14913);
and UO_1168 (O_1168,N_14965,N_14967);
nor UO_1169 (O_1169,N_14880,N_14919);
or UO_1170 (O_1170,N_14967,N_14924);
and UO_1171 (O_1171,N_14925,N_14909);
or UO_1172 (O_1172,N_14875,N_14998);
or UO_1173 (O_1173,N_14957,N_14982);
or UO_1174 (O_1174,N_14980,N_14949);
and UO_1175 (O_1175,N_14976,N_14980);
nand UO_1176 (O_1176,N_14944,N_14957);
or UO_1177 (O_1177,N_14977,N_14959);
and UO_1178 (O_1178,N_14897,N_14967);
or UO_1179 (O_1179,N_14949,N_14914);
nand UO_1180 (O_1180,N_14981,N_14929);
and UO_1181 (O_1181,N_14986,N_14958);
nor UO_1182 (O_1182,N_14968,N_14904);
nand UO_1183 (O_1183,N_14973,N_14938);
and UO_1184 (O_1184,N_14930,N_14886);
xnor UO_1185 (O_1185,N_14982,N_14897);
nor UO_1186 (O_1186,N_14912,N_14947);
nand UO_1187 (O_1187,N_14911,N_14960);
nand UO_1188 (O_1188,N_14889,N_14981);
xor UO_1189 (O_1189,N_14986,N_14884);
and UO_1190 (O_1190,N_14924,N_14918);
or UO_1191 (O_1191,N_14960,N_14899);
nand UO_1192 (O_1192,N_14938,N_14882);
or UO_1193 (O_1193,N_14981,N_14952);
nand UO_1194 (O_1194,N_14937,N_14949);
or UO_1195 (O_1195,N_14920,N_14947);
nor UO_1196 (O_1196,N_14902,N_14925);
and UO_1197 (O_1197,N_14932,N_14987);
or UO_1198 (O_1198,N_14884,N_14989);
nor UO_1199 (O_1199,N_14931,N_14942);
nor UO_1200 (O_1200,N_14969,N_14996);
or UO_1201 (O_1201,N_14952,N_14934);
nor UO_1202 (O_1202,N_14973,N_14970);
nand UO_1203 (O_1203,N_14931,N_14889);
or UO_1204 (O_1204,N_14978,N_14922);
or UO_1205 (O_1205,N_14885,N_14891);
nor UO_1206 (O_1206,N_14979,N_14964);
nor UO_1207 (O_1207,N_14950,N_14899);
or UO_1208 (O_1208,N_14942,N_14924);
xnor UO_1209 (O_1209,N_14933,N_14958);
and UO_1210 (O_1210,N_14988,N_14987);
nor UO_1211 (O_1211,N_14951,N_14890);
or UO_1212 (O_1212,N_14964,N_14901);
nand UO_1213 (O_1213,N_14947,N_14927);
nand UO_1214 (O_1214,N_14936,N_14937);
or UO_1215 (O_1215,N_14903,N_14996);
nor UO_1216 (O_1216,N_14983,N_14950);
nor UO_1217 (O_1217,N_14985,N_14938);
and UO_1218 (O_1218,N_14928,N_14925);
or UO_1219 (O_1219,N_14906,N_14909);
nor UO_1220 (O_1220,N_14938,N_14879);
nor UO_1221 (O_1221,N_14984,N_14875);
xnor UO_1222 (O_1222,N_14935,N_14918);
nor UO_1223 (O_1223,N_14947,N_14939);
and UO_1224 (O_1224,N_14955,N_14944);
and UO_1225 (O_1225,N_14911,N_14944);
nor UO_1226 (O_1226,N_14939,N_14875);
and UO_1227 (O_1227,N_14946,N_14947);
or UO_1228 (O_1228,N_14962,N_14926);
or UO_1229 (O_1229,N_14886,N_14940);
or UO_1230 (O_1230,N_14915,N_14940);
nand UO_1231 (O_1231,N_14977,N_14880);
nor UO_1232 (O_1232,N_14951,N_14960);
nor UO_1233 (O_1233,N_14875,N_14881);
nor UO_1234 (O_1234,N_14915,N_14932);
xnor UO_1235 (O_1235,N_14978,N_14947);
nand UO_1236 (O_1236,N_14896,N_14960);
or UO_1237 (O_1237,N_14958,N_14894);
nand UO_1238 (O_1238,N_14984,N_14917);
or UO_1239 (O_1239,N_14907,N_14927);
nor UO_1240 (O_1240,N_14933,N_14888);
nand UO_1241 (O_1241,N_14925,N_14987);
nand UO_1242 (O_1242,N_14888,N_14900);
or UO_1243 (O_1243,N_14889,N_14914);
xnor UO_1244 (O_1244,N_14908,N_14891);
nand UO_1245 (O_1245,N_14884,N_14959);
or UO_1246 (O_1246,N_14994,N_14950);
nand UO_1247 (O_1247,N_14890,N_14990);
xor UO_1248 (O_1248,N_14911,N_14897);
nand UO_1249 (O_1249,N_14953,N_14947);
nand UO_1250 (O_1250,N_14950,N_14924);
or UO_1251 (O_1251,N_14991,N_14909);
or UO_1252 (O_1252,N_14925,N_14904);
nor UO_1253 (O_1253,N_14998,N_14992);
and UO_1254 (O_1254,N_14926,N_14884);
or UO_1255 (O_1255,N_14897,N_14885);
xnor UO_1256 (O_1256,N_14972,N_14934);
nand UO_1257 (O_1257,N_14902,N_14970);
or UO_1258 (O_1258,N_14879,N_14892);
or UO_1259 (O_1259,N_14985,N_14991);
nand UO_1260 (O_1260,N_14988,N_14985);
nor UO_1261 (O_1261,N_14957,N_14969);
nand UO_1262 (O_1262,N_14971,N_14881);
nand UO_1263 (O_1263,N_14948,N_14940);
and UO_1264 (O_1264,N_14969,N_14988);
or UO_1265 (O_1265,N_14961,N_14951);
nand UO_1266 (O_1266,N_14957,N_14953);
or UO_1267 (O_1267,N_14885,N_14923);
xor UO_1268 (O_1268,N_14903,N_14892);
nand UO_1269 (O_1269,N_14974,N_14990);
and UO_1270 (O_1270,N_14922,N_14923);
and UO_1271 (O_1271,N_14980,N_14992);
nand UO_1272 (O_1272,N_14937,N_14885);
or UO_1273 (O_1273,N_14970,N_14944);
nand UO_1274 (O_1274,N_14888,N_14956);
nor UO_1275 (O_1275,N_14913,N_14877);
and UO_1276 (O_1276,N_14883,N_14972);
xnor UO_1277 (O_1277,N_14921,N_14909);
nor UO_1278 (O_1278,N_14988,N_14911);
or UO_1279 (O_1279,N_14889,N_14999);
nand UO_1280 (O_1280,N_14908,N_14983);
xnor UO_1281 (O_1281,N_14946,N_14906);
and UO_1282 (O_1282,N_14923,N_14879);
xnor UO_1283 (O_1283,N_14950,N_14995);
and UO_1284 (O_1284,N_14951,N_14977);
nand UO_1285 (O_1285,N_14962,N_14987);
and UO_1286 (O_1286,N_14994,N_14943);
and UO_1287 (O_1287,N_14977,N_14877);
xor UO_1288 (O_1288,N_14890,N_14941);
nand UO_1289 (O_1289,N_14995,N_14949);
nand UO_1290 (O_1290,N_14896,N_14899);
and UO_1291 (O_1291,N_14916,N_14945);
xnor UO_1292 (O_1292,N_14932,N_14970);
nand UO_1293 (O_1293,N_14921,N_14986);
or UO_1294 (O_1294,N_14977,N_14895);
nor UO_1295 (O_1295,N_14989,N_14971);
nand UO_1296 (O_1296,N_14971,N_14903);
and UO_1297 (O_1297,N_14924,N_14959);
nand UO_1298 (O_1298,N_14919,N_14918);
and UO_1299 (O_1299,N_14947,N_14951);
nand UO_1300 (O_1300,N_14968,N_14877);
nand UO_1301 (O_1301,N_14902,N_14903);
nand UO_1302 (O_1302,N_14972,N_14975);
and UO_1303 (O_1303,N_14936,N_14980);
nand UO_1304 (O_1304,N_14984,N_14900);
nor UO_1305 (O_1305,N_14988,N_14916);
xor UO_1306 (O_1306,N_14902,N_14875);
nand UO_1307 (O_1307,N_14946,N_14918);
nor UO_1308 (O_1308,N_14925,N_14983);
nor UO_1309 (O_1309,N_14919,N_14973);
or UO_1310 (O_1310,N_14954,N_14904);
nand UO_1311 (O_1311,N_14937,N_14911);
nand UO_1312 (O_1312,N_14956,N_14933);
nor UO_1313 (O_1313,N_14936,N_14913);
nor UO_1314 (O_1314,N_14982,N_14928);
nor UO_1315 (O_1315,N_14966,N_14920);
or UO_1316 (O_1316,N_14970,N_14886);
and UO_1317 (O_1317,N_14928,N_14955);
nor UO_1318 (O_1318,N_14969,N_14950);
or UO_1319 (O_1319,N_14968,N_14881);
or UO_1320 (O_1320,N_14910,N_14913);
nor UO_1321 (O_1321,N_14949,N_14979);
nand UO_1322 (O_1322,N_14898,N_14877);
nor UO_1323 (O_1323,N_14915,N_14890);
nor UO_1324 (O_1324,N_14917,N_14961);
nand UO_1325 (O_1325,N_14917,N_14941);
nor UO_1326 (O_1326,N_14923,N_14984);
nor UO_1327 (O_1327,N_14988,N_14966);
nand UO_1328 (O_1328,N_14930,N_14937);
and UO_1329 (O_1329,N_14897,N_14945);
or UO_1330 (O_1330,N_14967,N_14990);
and UO_1331 (O_1331,N_14973,N_14975);
and UO_1332 (O_1332,N_14948,N_14956);
nor UO_1333 (O_1333,N_14971,N_14909);
and UO_1334 (O_1334,N_14976,N_14978);
nor UO_1335 (O_1335,N_14877,N_14954);
nor UO_1336 (O_1336,N_14895,N_14912);
nand UO_1337 (O_1337,N_14990,N_14949);
and UO_1338 (O_1338,N_14979,N_14888);
nor UO_1339 (O_1339,N_14945,N_14977);
nor UO_1340 (O_1340,N_14883,N_14940);
xnor UO_1341 (O_1341,N_14875,N_14999);
or UO_1342 (O_1342,N_14935,N_14885);
nand UO_1343 (O_1343,N_14889,N_14925);
and UO_1344 (O_1344,N_14950,N_14926);
and UO_1345 (O_1345,N_14955,N_14882);
or UO_1346 (O_1346,N_14965,N_14911);
nand UO_1347 (O_1347,N_14938,N_14998);
nand UO_1348 (O_1348,N_14953,N_14892);
or UO_1349 (O_1349,N_14995,N_14921);
and UO_1350 (O_1350,N_14929,N_14936);
nor UO_1351 (O_1351,N_14994,N_14987);
and UO_1352 (O_1352,N_14932,N_14985);
or UO_1353 (O_1353,N_14896,N_14981);
and UO_1354 (O_1354,N_14893,N_14948);
nor UO_1355 (O_1355,N_14922,N_14961);
or UO_1356 (O_1356,N_14893,N_14947);
nor UO_1357 (O_1357,N_14938,N_14933);
and UO_1358 (O_1358,N_14978,N_14887);
or UO_1359 (O_1359,N_14879,N_14933);
nand UO_1360 (O_1360,N_14999,N_14954);
and UO_1361 (O_1361,N_14897,N_14960);
xor UO_1362 (O_1362,N_14961,N_14911);
and UO_1363 (O_1363,N_14894,N_14909);
nand UO_1364 (O_1364,N_14885,N_14928);
or UO_1365 (O_1365,N_14949,N_14877);
and UO_1366 (O_1366,N_14970,N_14960);
nand UO_1367 (O_1367,N_14941,N_14987);
or UO_1368 (O_1368,N_14905,N_14971);
nand UO_1369 (O_1369,N_14922,N_14921);
or UO_1370 (O_1370,N_14904,N_14899);
or UO_1371 (O_1371,N_14947,N_14983);
or UO_1372 (O_1372,N_14917,N_14958);
xnor UO_1373 (O_1373,N_14988,N_14923);
or UO_1374 (O_1374,N_14894,N_14893);
and UO_1375 (O_1375,N_14889,N_14992);
nor UO_1376 (O_1376,N_14932,N_14890);
nor UO_1377 (O_1377,N_14893,N_14935);
xnor UO_1378 (O_1378,N_14976,N_14928);
nand UO_1379 (O_1379,N_14934,N_14897);
nor UO_1380 (O_1380,N_14939,N_14915);
xor UO_1381 (O_1381,N_14992,N_14883);
xor UO_1382 (O_1382,N_14993,N_14913);
nand UO_1383 (O_1383,N_14961,N_14972);
and UO_1384 (O_1384,N_14892,N_14956);
nor UO_1385 (O_1385,N_14973,N_14961);
nand UO_1386 (O_1386,N_14880,N_14879);
or UO_1387 (O_1387,N_14930,N_14901);
nor UO_1388 (O_1388,N_14931,N_14958);
nand UO_1389 (O_1389,N_14970,N_14953);
and UO_1390 (O_1390,N_14993,N_14978);
nand UO_1391 (O_1391,N_14983,N_14930);
xor UO_1392 (O_1392,N_14879,N_14985);
and UO_1393 (O_1393,N_14980,N_14916);
nand UO_1394 (O_1394,N_14876,N_14912);
or UO_1395 (O_1395,N_14987,N_14891);
nand UO_1396 (O_1396,N_14919,N_14979);
nand UO_1397 (O_1397,N_14969,N_14990);
nor UO_1398 (O_1398,N_14901,N_14899);
nor UO_1399 (O_1399,N_14995,N_14897);
or UO_1400 (O_1400,N_14991,N_14875);
and UO_1401 (O_1401,N_14937,N_14902);
and UO_1402 (O_1402,N_14969,N_14933);
or UO_1403 (O_1403,N_14931,N_14898);
xor UO_1404 (O_1404,N_14947,N_14905);
nand UO_1405 (O_1405,N_14998,N_14980);
and UO_1406 (O_1406,N_14952,N_14913);
xor UO_1407 (O_1407,N_14966,N_14967);
or UO_1408 (O_1408,N_14917,N_14881);
nand UO_1409 (O_1409,N_14925,N_14921);
or UO_1410 (O_1410,N_14887,N_14980);
and UO_1411 (O_1411,N_14977,N_14939);
xnor UO_1412 (O_1412,N_14923,N_14983);
or UO_1413 (O_1413,N_14943,N_14949);
nand UO_1414 (O_1414,N_14926,N_14917);
nor UO_1415 (O_1415,N_14990,N_14908);
nor UO_1416 (O_1416,N_14981,N_14880);
and UO_1417 (O_1417,N_14949,N_14930);
or UO_1418 (O_1418,N_14908,N_14980);
and UO_1419 (O_1419,N_14932,N_14945);
and UO_1420 (O_1420,N_14961,N_14960);
nor UO_1421 (O_1421,N_14879,N_14911);
nor UO_1422 (O_1422,N_14931,N_14981);
nand UO_1423 (O_1423,N_14909,N_14882);
nor UO_1424 (O_1424,N_14989,N_14973);
and UO_1425 (O_1425,N_14905,N_14882);
xnor UO_1426 (O_1426,N_14900,N_14979);
or UO_1427 (O_1427,N_14961,N_14946);
nor UO_1428 (O_1428,N_14977,N_14887);
xnor UO_1429 (O_1429,N_14944,N_14993);
and UO_1430 (O_1430,N_14944,N_14992);
nor UO_1431 (O_1431,N_14889,N_14967);
nand UO_1432 (O_1432,N_14882,N_14928);
and UO_1433 (O_1433,N_14890,N_14928);
or UO_1434 (O_1434,N_14897,N_14899);
or UO_1435 (O_1435,N_14998,N_14892);
or UO_1436 (O_1436,N_14989,N_14968);
or UO_1437 (O_1437,N_14875,N_14888);
and UO_1438 (O_1438,N_14898,N_14961);
nand UO_1439 (O_1439,N_14891,N_14982);
nand UO_1440 (O_1440,N_14934,N_14905);
or UO_1441 (O_1441,N_14998,N_14953);
nor UO_1442 (O_1442,N_14875,N_14925);
nor UO_1443 (O_1443,N_14907,N_14893);
xnor UO_1444 (O_1444,N_14948,N_14906);
or UO_1445 (O_1445,N_14955,N_14969);
nor UO_1446 (O_1446,N_14903,N_14918);
nor UO_1447 (O_1447,N_14977,N_14927);
nand UO_1448 (O_1448,N_14950,N_14997);
xor UO_1449 (O_1449,N_14971,N_14934);
nor UO_1450 (O_1450,N_14960,N_14991);
or UO_1451 (O_1451,N_14923,N_14931);
nand UO_1452 (O_1452,N_14969,N_14945);
nand UO_1453 (O_1453,N_14954,N_14876);
or UO_1454 (O_1454,N_14953,N_14914);
or UO_1455 (O_1455,N_14944,N_14884);
xnor UO_1456 (O_1456,N_14971,N_14996);
and UO_1457 (O_1457,N_14965,N_14933);
nor UO_1458 (O_1458,N_14925,N_14917);
nor UO_1459 (O_1459,N_14952,N_14909);
nor UO_1460 (O_1460,N_14915,N_14980);
nor UO_1461 (O_1461,N_14922,N_14893);
and UO_1462 (O_1462,N_14979,N_14908);
nor UO_1463 (O_1463,N_14927,N_14988);
nand UO_1464 (O_1464,N_14989,N_14978);
nor UO_1465 (O_1465,N_14895,N_14992);
nand UO_1466 (O_1466,N_14910,N_14935);
nor UO_1467 (O_1467,N_14976,N_14966);
and UO_1468 (O_1468,N_14937,N_14892);
or UO_1469 (O_1469,N_14969,N_14985);
or UO_1470 (O_1470,N_14949,N_14925);
and UO_1471 (O_1471,N_14983,N_14895);
nor UO_1472 (O_1472,N_14951,N_14946);
nor UO_1473 (O_1473,N_14984,N_14961);
nor UO_1474 (O_1474,N_14880,N_14990);
nand UO_1475 (O_1475,N_14987,N_14960);
nand UO_1476 (O_1476,N_14875,N_14953);
or UO_1477 (O_1477,N_14894,N_14953);
and UO_1478 (O_1478,N_14986,N_14920);
or UO_1479 (O_1479,N_14908,N_14942);
or UO_1480 (O_1480,N_14946,N_14940);
or UO_1481 (O_1481,N_14892,N_14913);
and UO_1482 (O_1482,N_14943,N_14913);
nor UO_1483 (O_1483,N_14993,N_14937);
or UO_1484 (O_1484,N_14914,N_14918);
nand UO_1485 (O_1485,N_14980,N_14902);
or UO_1486 (O_1486,N_14971,N_14973);
xor UO_1487 (O_1487,N_14883,N_14905);
or UO_1488 (O_1488,N_14984,N_14901);
nor UO_1489 (O_1489,N_14986,N_14962);
or UO_1490 (O_1490,N_14972,N_14990);
nand UO_1491 (O_1491,N_14963,N_14947);
xnor UO_1492 (O_1492,N_14952,N_14955);
nor UO_1493 (O_1493,N_14927,N_14990);
and UO_1494 (O_1494,N_14972,N_14889);
or UO_1495 (O_1495,N_14927,N_14956);
nor UO_1496 (O_1496,N_14905,N_14880);
and UO_1497 (O_1497,N_14995,N_14881);
and UO_1498 (O_1498,N_14940,N_14933);
nor UO_1499 (O_1499,N_14928,N_14902);
or UO_1500 (O_1500,N_14913,N_14918);
nand UO_1501 (O_1501,N_14996,N_14972);
nor UO_1502 (O_1502,N_14954,N_14975);
and UO_1503 (O_1503,N_14955,N_14891);
nand UO_1504 (O_1504,N_14912,N_14875);
nand UO_1505 (O_1505,N_14959,N_14893);
nor UO_1506 (O_1506,N_14907,N_14900);
or UO_1507 (O_1507,N_14953,N_14883);
nand UO_1508 (O_1508,N_14890,N_14989);
nor UO_1509 (O_1509,N_14890,N_14935);
nor UO_1510 (O_1510,N_14949,N_14957);
or UO_1511 (O_1511,N_14936,N_14972);
nand UO_1512 (O_1512,N_14961,N_14936);
xnor UO_1513 (O_1513,N_14891,N_14976);
or UO_1514 (O_1514,N_14904,N_14978);
nand UO_1515 (O_1515,N_14973,N_14952);
or UO_1516 (O_1516,N_14990,N_14907);
nand UO_1517 (O_1517,N_14958,N_14920);
nand UO_1518 (O_1518,N_14900,N_14910);
nor UO_1519 (O_1519,N_14915,N_14902);
nor UO_1520 (O_1520,N_14973,N_14991);
nand UO_1521 (O_1521,N_14916,N_14979);
or UO_1522 (O_1522,N_14985,N_14970);
or UO_1523 (O_1523,N_14937,N_14910);
and UO_1524 (O_1524,N_14932,N_14959);
nand UO_1525 (O_1525,N_14964,N_14998);
nand UO_1526 (O_1526,N_14904,N_14991);
nand UO_1527 (O_1527,N_14895,N_14997);
and UO_1528 (O_1528,N_14987,N_14908);
nand UO_1529 (O_1529,N_14899,N_14951);
xor UO_1530 (O_1530,N_14941,N_14933);
xor UO_1531 (O_1531,N_14892,N_14983);
and UO_1532 (O_1532,N_14887,N_14920);
and UO_1533 (O_1533,N_14881,N_14963);
and UO_1534 (O_1534,N_14968,N_14946);
and UO_1535 (O_1535,N_14899,N_14993);
nand UO_1536 (O_1536,N_14969,N_14952);
or UO_1537 (O_1537,N_14929,N_14975);
xnor UO_1538 (O_1538,N_14891,N_14909);
and UO_1539 (O_1539,N_14889,N_14895);
nor UO_1540 (O_1540,N_14932,N_14995);
and UO_1541 (O_1541,N_14969,N_14918);
and UO_1542 (O_1542,N_14908,N_14988);
nand UO_1543 (O_1543,N_14931,N_14988);
or UO_1544 (O_1544,N_14881,N_14927);
nor UO_1545 (O_1545,N_14931,N_14967);
nand UO_1546 (O_1546,N_14933,N_14880);
and UO_1547 (O_1547,N_14880,N_14989);
nor UO_1548 (O_1548,N_14944,N_14977);
nand UO_1549 (O_1549,N_14978,N_14928);
xor UO_1550 (O_1550,N_14920,N_14978);
nand UO_1551 (O_1551,N_14943,N_14964);
and UO_1552 (O_1552,N_14977,N_14947);
or UO_1553 (O_1553,N_14904,N_14886);
and UO_1554 (O_1554,N_14942,N_14961);
or UO_1555 (O_1555,N_14900,N_14973);
and UO_1556 (O_1556,N_14972,N_14875);
nand UO_1557 (O_1557,N_14906,N_14892);
or UO_1558 (O_1558,N_14965,N_14946);
xor UO_1559 (O_1559,N_14902,N_14990);
xor UO_1560 (O_1560,N_14893,N_14996);
xnor UO_1561 (O_1561,N_14921,N_14894);
xnor UO_1562 (O_1562,N_14915,N_14985);
xor UO_1563 (O_1563,N_14937,N_14990);
or UO_1564 (O_1564,N_14892,N_14885);
nand UO_1565 (O_1565,N_14982,N_14998);
or UO_1566 (O_1566,N_14994,N_14982);
or UO_1567 (O_1567,N_14896,N_14918);
nor UO_1568 (O_1568,N_14930,N_14927);
and UO_1569 (O_1569,N_14989,N_14905);
nand UO_1570 (O_1570,N_14998,N_14976);
and UO_1571 (O_1571,N_14942,N_14966);
nor UO_1572 (O_1572,N_14879,N_14970);
xor UO_1573 (O_1573,N_14974,N_14965);
nand UO_1574 (O_1574,N_14908,N_14915);
xor UO_1575 (O_1575,N_14981,N_14932);
nand UO_1576 (O_1576,N_14910,N_14957);
nor UO_1577 (O_1577,N_14926,N_14902);
nand UO_1578 (O_1578,N_14989,N_14930);
or UO_1579 (O_1579,N_14890,N_14889);
nor UO_1580 (O_1580,N_14992,N_14946);
xor UO_1581 (O_1581,N_14916,N_14985);
nand UO_1582 (O_1582,N_14882,N_14912);
nand UO_1583 (O_1583,N_14968,N_14973);
and UO_1584 (O_1584,N_14924,N_14911);
nand UO_1585 (O_1585,N_14990,N_14899);
and UO_1586 (O_1586,N_14930,N_14913);
nand UO_1587 (O_1587,N_14915,N_14941);
or UO_1588 (O_1588,N_14917,N_14904);
nand UO_1589 (O_1589,N_14966,N_14929);
nand UO_1590 (O_1590,N_14978,N_14895);
nand UO_1591 (O_1591,N_14930,N_14994);
or UO_1592 (O_1592,N_14963,N_14886);
and UO_1593 (O_1593,N_14881,N_14921);
nand UO_1594 (O_1594,N_14959,N_14973);
or UO_1595 (O_1595,N_14993,N_14906);
nor UO_1596 (O_1596,N_14887,N_14891);
or UO_1597 (O_1597,N_14994,N_14995);
nor UO_1598 (O_1598,N_14972,N_14973);
nand UO_1599 (O_1599,N_14887,N_14893);
and UO_1600 (O_1600,N_14954,N_14970);
nor UO_1601 (O_1601,N_14971,N_14894);
and UO_1602 (O_1602,N_14978,N_14953);
nand UO_1603 (O_1603,N_14919,N_14969);
and UO_1604 (O_1604,N_14964,N_14933);
nor UO_1605 (O_1605,N_14926,N_14954);
xnor UO_1606 (O_1606,N_14975,N_14966);
and UO_1607 (O_1607,N_14970,N_14875);
nand UO_1608 (O_1608,N_14965,N_14922);
xor UO_1609 (O_1609,N_14879,N_14940);
or UO_1610 (O_1610,N_14964,N_14913);
nand UO_1611 (O_1611,N_14990,N_14909);
or UO_1612 (O_1612,N_14923,N_14977);
nand UO_1613 (O_1613,N_14994,N_14919);
or UO_1614 (O_1614,N_14999,N_14930);
nor UO_1615 (O_1615,N_14890,N_14942);
nand UO_1616 (O_1616,N_14999,N_14876);
nand UO_1617 (O_1617,N_14930,N_14991);
or UO_1618 (O_1618,N_14978,N_14926);
nand UO_1619 (O_1619,N_14877,N_14922);
or UO_1620 (O_1620,N_14978,N_14960);
nand UO_1621 (O_1621,N_14908,N_14955);
and UO_1622 (O_1622,N_14964,N_14993);
nand UO_1623 (O_1623,N_14989,N_14929);
or UO_1624 (O_1624,N_14892,N_14923);
and UO_1625 (O_1625,N_14944,N_14921);
nand UO_1626 (O_1626,N_14996,N_14876);
nand UO_1627 (O_1627,N_14917,N_14976);
nand UO_1628 (O_1628,N_14929,N_14896);
nand UO_1629 (O_1629,N_14983,N_14890);
or UO_1630 (O_1630,N_14923,N_14934);
and UO_1631 (O_1631,N_14984,N_14978);
nor UO_1632 (O_1632,N_14939,N_14877);
nor UO_1633 (O_1633,N_14931,N_14891);
or UO_1634 (O_1634,N_14939,N_14990);
nor UO_1635 (O_1635,N_14890,N_14900);
nand UO_1636 (O_1636,N_14963,N_14884);
and UO_1637 (O_1637,N_14892,N_14899);
nand UO_1638 (O_1638,N_14919,N_14954);
nand UO_1639 (O_1639,N_14967,N_14895);
nor UO_1640 (O_1640,N_14890,N_14985);
or UO_1641 (O_1641,N_14932,N_14969);
nand UO_1642 (O_1642,N_14922,N_14911);
xor UO_1643 (O_1643,N_14910,N_14967);
or UO_1644 (O_1644,N_14962,N_14934);
and UO_1645 (O_1645,N_14906,N_14914);
or UO_1646 (O_1646,N_14984,N_14906);
nor UO_1647 (O_1647,N_14980,N_14989);
and UO_1648 (O_1648,N_14907,N_14923);
and UO_1649 (O_1649,N_14990,N_14998);
or UO_1650 (O_1650,N_14909,N_14914);
and UO_1651 (O_1651,N_14939,N_14889);
and UO_1652 (O_1652,N_14969,N_14968);
or UO_1653 (O_1653,N_14981,N_14913);
xor UO_1654 (O_1654,N_14891,N_14971);
and UO_1655 (O_1655,N_14911,N_14975);
and UO_1656 (O_1656,N_14958,N_14980);
nor UO_1657 (O_1657,N_14955,N_14983);
and UO_1658 (O_1658,N_14938,N_14984);
or UO_1659 (O_1659,N_14914,N_14983);
xor UO_1660 (O_1660,N_14971,N_14875);
nand UO_1661 (O_1661,N_14944,N_14889);
and UO_1662 (O_1662,N_14977,N_14952);
nand UO_1663 (O_1663,N_14946,N_14903);
and UO_1664 (O_1664,N_14898,N_14882);
and UO_1665 (O_1665,N_14934,N_14949);
and UO_1666 (O_1666,N_14929,N_14926);
or UO_1667 (O_1667,N_14895,N_14891);
nand UO_1668 (O_1668,N_14920,N_14989);
or UO_1669 (O_1669,N_14938,N_14972);
or UO_1670 (O_1670,N_14926,N_14969);
nand UO_1671 (O_1671,N_14988,N_14946);
nand UO_1672 (O_1672,N_14938,N_14912);
and UO_1673 (O_1673,N_14894,N_14875);
xor UO_1674 (O_1674,N_14946,N_14880);
and UO_1675 (O_1675,N_14966,N_14981);
and UO_1676 (O_1676,N_14941,N_14898);
or UO_1677 (O_1677,N_14960,N_14952);
and UO_1678 (O_1678,N_14988,N_14917);
xor UO_1679 (O_1679,N_14914,N_14885);
nand UO_1680 (O_1680,N_14954,N_14964);
nor UO_1681 (O_1681,N_14927,N_14909);
nand UO_1682 (O_1682,N_14972,N_14979);
xor UO_1683 (O_1683,N_14888,N_14935);
and UO_1684 (O_1684,N_14972,N_14885);
and UO_1685 (O_1685,N_14911,N_14916);
or UO_1686 (O_1686,N_14882,N_14946);
and UO_1687 (O_1687,N_14958,N_14875);
and UO_1688 (O_1688,N_14925,N_14989);
nand UO_1689 (O_1689,N_14944,N_14972);
nand UO_1690 (O_1690,N_14901,N_14947);
nand UO_1691 (O_1691,N_14968,N_14934);
or UO_1692 (O_1692,N_14916,N_14951);
and UO_1693 (O_1693,N_14925,N_14919);
nand UO_1694 (O_1694,N_14875,N_14955);
nand UO_1695 (O_1695,N_14911,N_14934);
and UO_1696 (O_1696,N_14960,N_14955);
and UO_1697 (O_1697,N_14939,N_14923);
xor UO_1698 (O_1698,N_14972,N_14879);
xnor UO_1699 (O_1699,N_14967,N_14997);
nand UO_1700 (O_1700,N_14978,N_14946);
nor UO_1701 (O_1701,N_14883,N_14981);
nand UO_1702 (O_1702,N_14996,N_14919);
nand UO_1703 (O_1703,N_14971,N_14965);
or UO_1704 (O_1704,N_14999,N_14964);
or UO_1705 (O_1705,N_14939,N_14891);
nand UO_1706 (O_1706,N_14928,N_14892);
nand UO_1707 (O_1707,N_14979,N_14911);
xor UO_1708 (O_1708,N_14903,N_14993);
nor UO_1709 (O_1709,N_14892,N_14893);
and UO_1710 (O_1710,N_14905,N_14889);
xnor UO_1711 (O_1711,N_14892,N_14985);
or UO_1712 (O_1712,N_14950,N_14933);
and UO_1713 (O_1713,N_14965,N_14929);
and UO_1714 (O_1714,N_14967,N_14896);
or UO_1715 (O_1715,N_14955,N_14991);
or UO_1716 (O_1716,N_14896,N_14965);
and UO_1717 (O_1717,N_14992,N_14897);
nand UO_1718 (O_1718,N_14987,N_14903);
and UO_1719 (O_1719,N_14925,N_14997);
and UO_1720 (O_1720,N_14892,N_14896);
nand UO_1721 (O_1721,N_14974,N_14884);
nor UO_1722 (O_1722,N_14904,N_14939);
nand UO_1723 (O_1723,N_14919,N_14934);
nor UO_1724 (O_1724,N_14892,N_14951);
and UO_1725 (O_1725,N_14887,N_14899);
xor UO_1726 (O_1726,N_14899,N_14875);
and UO_1727 (O_1727,N_14957,N_14966);
or UO_1728 (O_1728,N_14884,N_14942);
nor UO_1729 (O_1729,N_14888,N_14994);
or UO_1730 (O_1730,N_14930,N_14880);
nand UO_1731 (O_1731,N_14928,N_14941);
nand UO_1732 (O_1732,N_14916,N_14882);
nor UO_1733 (O_1733,N_14897,N_14883);
or UO_1734 (O_1734,N_14888,N_14894);
nand UO_1735 (O_1735,N_14894,N_14959);
nor UO_1736 (O_1736,N_14987,N_14917);
or UO_1737 (O_1737,N_14917,N_14891);
nor UO_1738 (O_1738,N_14926,N_14907);
nor UO_1739 (O_1739,N_14985,N_14886);
or UO_1740 (O_1740,N_14919,N_14951);
xor UO_1741 (O_1741,N_14971,N_14945);
nor UO_1742 (O_1742,N_14952,N_14905);
or UO_1743 (O_1743,N_14979,N_14885);
nor UO_1744 (O_1744,N_14970,N_14917);
or UO_1745 (O_1745,N_14995,N_14935);
and UO_1746 (O_1746,N_14978,N_14885);
or UO_1747 (O_1747,N_14992,N_14927);
nor UO_1748 (O_1748,N_14949,N_14940);
or UO_1749 (O_1749,N_14934,N_14985);
nor UO_1750 (O_1750,N_14927,N_14940);
and UO_1751 (O_1751,N_14974,N_14978);
nor UO_1752 (O_1752,N_14925,N_14966);
nor UO_1753 (O_1753,N_14891,N_14897);
or UO_1754 (O_1754,N_14946,N_14937);
nand UO_1755 (O_1755,N_14932,N_14991);
and UO_1756 (O_1756,N_14888,N_14928);
nand UO_1757 (O_1757,N_14878,N_14997);
nor UO_1758 (O_1758,N_14940,N_14963);
nor UO_1759 (O_1759,N_14906,N_14884);
or UO_1760 (O_1760,N_14889,N_14923);
and UO_1761 (O_1761,N_14899,N_14964);
nor UO_1762 (O_1762,N_14941,N_14963);
xnor UO_1763 (O_1763,N_14928,N_14936);
or UO_1764 (O_1764,N_14955,N_14899);
nor UO_1765 (O_1765,N_14911,N_14983);
and UO_1766 (O_1766,N_14995,N_14891);
xnor UO_1767 (O_1767,N_14904,N_14976);
nand UO_1768 (O_1768,N_14875,N_14974);
or UO_1769 (O_1769,N_14957,N_14968);
nand UO_1770 (O_1770,N_14975,N_14996);
nand UO_1771 (O_1771,N_14897,N_14914);
or UO_1772 (O_1772,N_14973,N_14946);
or UO_1773 (O_1773,N_14945,N_14893);
xor UO_1774 (O_1774,N_14982,N_14926);
or UO_1775 (O_1775,N_14914,N_14900);
nor UO_1776 (O_1776,N_14956,N_14920);
or UO_1777 (O_1777,N_14881,N_14948);
and UO_1778 (O_1778,N_14887,N_14924);
and UO_1779 (O_1779,N_14991,N_14944);
xnor UO_1780 (O_1780,N_14989,N_14875);
nand UO_1781 (O_1781,N_14958,N_14985);
or UO_1782 (O_1782,N_14877,N_14895);
nand UO_1783 (O_1783,N_14886,N_14888);
or UO_1784 (O_1784,N_14994,N_14898);
xor UO_1785 (O_1785,N_14993,N_14926);
xor UO_1786 (O_1786,N_14936,N_14947);
nand UO_1787 (O_1787,N_14890,N_14967);
nand UO_1788 (O_1788,N_14978,N_14942);
and UO_1789 (O_1789,N_14888,N_14972);
xor UO_1790 (O_1790,N_14961,N_14892);
nand UO_1791 (O_1791,N_14957,N_14993);
and UO_1792 (O_1792,N_14990,N_14938);
xnor UO_1793 (O_1793,N_14893,N_14882);
or UO_1794 (O_1794,N_14943,N_14961);
or UO_1795 (O_1795,N_14887,N_14935);
nor UO_1796 (O_1796,N_14920,N_14922);
nand UO_1797 (O_1797,N_14883,N_14935);
nand UO_1798 (O_1798,N_14926,N_14972);
and UO_1799 (O_1799,N_14936,N_14986);
nand UO_1800 (O_1800,N_14897,N_14921);
and UO_1801 (O_1801,N_14998,N_14917);
nand UO_1802 (O_1802,N_14930,N_14941);
or UO_1803 (O_1803,N_14923,N_14999);
nand UO_1804 (O_1804,N_14958,N_14924);
nand UO_1805 (O_1805,N_14989,N_14995);
and UO_1806 (O_1806,N_14921,N_14891);
xnor UO_1807 (O_1807,N_14951,N_14934);
nor UO_1808 (O_1808,N_14936,N_14949);
and UO_1809 (O_1809,N_14945,N_14948);
nor UO_1810 (O_1810,N_14982,N_14877);
or UO_1811 (O_1811,N_14988,N_14992);
or UO_1812 (O_1812,N_14880,N_14941);
and UO_1813 (O_1813,N_14902,N_14941);
and UO_1814 (O_1814,N_14926,N_14977);
or UO_1815 (O_1815,N_14876,N_14896);
nor UO_1816 (O_1816,N_14903,N_14894);
nor UO_1817 (O_1817,N_14955,N_14887);
and UO_1818 (O_1818,N_14959,N_14931);
and UO_1819 (O_1819,N_14953,N_14896);
xnor UO_1820 (O_1820,N_14942,N_14923);
nor UO_1821 (O_1821,N_14997,N_14917);
nor UO_1822 (O_1822,N_14889,N_14876);
or UO_1823 (O_1823,N_14927,N_14889);
nand UO_1824 (O_1824,N_14958,N_14912);
or UO_1825 (O_1825,N_14875,N_14897);
or UO_1826 (O_1826,N_14916,N_14913);
nor UO_1827 (O_1827,N_14976,N_14979);
nor UO_1828 (O_1828,N_14969,N_14897);
nor UO_1829 (O_1829,N_14893,N_14953);
nor UO_1830 (O_1830,N_14986,N_14960);
nand UO_1831 (O_1831,N_14909,N_14934);
nand UO_1832 (O_1832,N_14962,N_14927);
nand UO_1833 (O_1833,N_14967,N_14941);
or UO_1834 (O_1834,N_14924,N_14951);
xnor UO_1835 (O_1835,N_14966,N_14908);
nand UO_1836 (O_1836,N_14958,N_14969);
or UO_1837 (O_1837,N_14992,N_14904);
nor UO_1838 (O_1838,N_14921,N_14955);
xor UO_1839 (O_1839,N_14891,N_14954);
and UO_1840 (O_1840,N_14947,N_14966);
nand UO_1841 (O_1841,N_14914,N_14982);
or UO_1842 (O_1842,N_14978,N_14918);
nor UO_1843 (O_1843,N_14883,N_14982);
or UO_1844 (O_1844,N_14954,N_14956);
and UO_1845 (O_1845,N_14885,N_14920);
nand UO_1846 (O_1846,N_14958,N_14945);
nand UO_1847 (O_1847,N_14993,N_14984);
xor UO_1848 (O_1848,N_14965,N_14882);
and UO_1849 (O_1849,N_14909,N_14964);
nand UO_1850 (O_1850,N_14988,N_14942);
nor UO_1851 (O_1851,N_14979,N_14906);
xnor UO_1852 (O_1852,N_14936,N_14996);
and UO_1853 (O_1853,N_14922,N_14967);
and UO_1854 (O_1854,N_14898,N_14880);
and UO_1855 (O_1855,N_14928,N_14914);
and UO_1856 (O_1856,N_14883,N_14970);
or UO_1857 (O_1857,N_14919,N_14906);
or UO_1858 (O_1858,N_14941,N_14916);
or UO_1859 (O_1859,N_14880,N_14995);
nand UO_1860 (O_1860,N_14984,N_14952);
xnor UO_1861 (O_1861,N_14904,N_14884);
nor UO_1862 (O_1862,N_14888,N_14924);
xnor UO_1863 (O_1863,N_14997,N_14961);
nor UO_1864 (O_1864,N_14987,N_14928);
or UO_1865 (O_1865,N_14890,N_14978);
nor UO_1866 (O_1866,N_14910,N_14933);
nor UO_1867 (O_1867,N_14975,N_14921);
and UO_1868 (O_1868,N_14952,N_14900);
and UO_1869 (O_1869,N_14905,N_14987);
xor UO_1870 (O_1870,N_14920,N_14925);
or UO_1871 (O_1871,N_14891,N_14953);
nand UO_1872 (O_1872,N_14888,N_14990);
nor UO_1873 (O_1873,N_14894,N_14877);
or UO_1874 (O_1874,N_14960,N_14998);
nand UO_1875 (O_1875,N_14936,N_14993);
nor UO_1876 (O_1876,N_14965,N_14897);
or UO_1877 (O_1877,N_14900,N_14878);
or UO_1878 (O_1878,N_14918,N_14884);
and UO_1879 (O_1879,N_14878,N_14916);
and UO_1880 (O_1880,N_14900,N_14978);
or UO_1881 (O_1881,N_14943,N_14997);
and UO_1882 (O_1882,N_14883,N_14927);
nor UO_1883 (O_1883,N_14912,N_14939);
or UO_1884 (O_1884,N_14938,N_14877);
xor UO_1885 (O_1885,N_14922,N_14970);
or UO_1886 (O_1886,N_14905,N_14996);
nand UO_1887 (O_1887,N_14938,N_14964);
or UO_1888 (O_1888,N_14917,N_14982);
nand UO_1889 (O_1889,N_14993,N_14988);
nor UO_1890 (O_1890,N_14947,N_14981);
nand UO_1891 (O_1891,N_14882,N_14949);
and UO_1892 (O_1892,N_14940,N_14938);
nand UO_1893 (O_1893,N_14926,N_14892);
or UO_1894 (O_1894,N_14929,N_14945);
and UO_1895 (O_1895,N_14889,N_14983);
nand UO_1896 (O_1896,N_14903,N_14916);
nor UO_1897 (O_1897,N_14924,N_14905);
nor UO_1898 (O_1898,N_14978,N_14997);
or UO_1899 (O_1899,N_14964,N_14994);
or UO_1900 (O_1900,N_14952,N_14894);
and UO_1901 (O_1901,N_14953,N_14926);
and UO_1902 (O_1902,N_14895,N_14909);
or UO_1903 (O_1903,N_14912,N_14985);
and UO_1904 (O_1904,N_14886,N_14890);
or UO_1905 (O_1905,N_14997,N_14891);
nor UO_1906 (O_1906,N_14999,N_14888);
nor UO_1907 (O_1907,N_14927,N_14949);
nor UO_1908 (O_1908,N_14928,N_14875);
or UO_1909 (O_1909,N_14995,N_14962);
xor UO_1910 (O_1910,N_14965,N_14936);
and UO_1911 (O_1911,N_14912,N_14941);
nand UO_1912 (O_1912,N_14899,N_14992);
and UO_1913 (O_1913,N_14882,N_14993);
nand UO_1914 (O_1914,N_14993,N_14950);
and UO_1915 (O_1915,N_14969,N_14974);
nand UO_1916 (O_1916,N_14923,N_14970);
nand UO_1917 (O_1917,N_14955,N_14911);
nand UO_1918 (O_1918,N_14976,N_14950);
nor UO_1919 (O_1919,N_14953,N_14904);
or UO_1920 (O_1920,N_14935,N_14915);
and UO_1921 (O_1921,N_14897,N_14902);
or UO_1922 (O_1922,N_14898,N_14995);
nor UO_1923 (O_1923,N_14976,N_14940);
and UO_1924 (O_1924,N_14899,N_14886);
or UO_1925 (O_1925,N_14891,N_14974);
or UO_1926 (O_1926,N_14961,N_14945);
and UO_1927 (O_1927,N_14907,N_14976);
nor UO_1928 (O_1928,N_14889,N_14986);
nand UO_1929 (O_1929,N_14875,N_14968);
or UO_1930 (O_1930,N_14982,N_14937);
nor UO_1931 (O_1931,N_14942,N_14919);
or UO_1932 (O_1932,N_14955,N_14933);
or UO_1933 (O_1933,N_14964,N_14995);
or UO_1934 (O_1934,N_14901,N_14961);
nor UO_1935 (O_1935,N_14974,N_14953);
nand UO_1936 (O_1936,N_14940,N_14912);
nand UO_1937 (O_1937,N_14941,N_14996);
and UO_1938 (O_1938,N_14876,N_14951);
nand UO_1939 (O_1939,N_14946,N_14878);
nor UO_1940 (O_1940,N_14910,N_14931);
or UO_1941 (O_1941,N_14938,N_14949);
xnor UO_1942 (O_1942,N_14951,N_14940);
or UO_1943 (O_1943,N_14894,N_14885);
xor UO_1944 (O_1944,N_14879,N_14965);
or UO_1945 (O_1945,N_14904,N_14984);
nor UO_1946 (O_1946,N_14978,N_14981);
nand UO_1947 (O_1947,N_14984,N_14965);
nand UO_1948 (O_1948,N_14930,N_14884);
nand UO_1949 (O_1949,N_14900,N_14919);
and UO_1950 (O_1950,N_14983,N_14943);
nand UO_1951 (O_1951,N_14947,N_14988);
nor UO_1952 (O_1952,N_14887,N_14948);
nand UO_1953 (O_1953,N_14936,N_14958);
nor UO_1954 (O_1954,N_14922,N_14899);
nand UO_1955 (O_1955,N_14878,N_14981);
nand UO_1956 (O_1956,N_14993,N_14907);
nand UO_1957 (O_1957,N_14886,N_14880);
or UO_1958 (O_1958,N_14992,N_14887);
xor UO_1959 (O_1959,N_14951,N_14913);
xnor UO_1960 (O_1960,N_14878,N_14896);
or UO_1961 (O_1961,N_14899,N_14966);
and UO_1962 (O_1962,N_14885,N_14969);
xor UO_1963 (O_1963,N_14915,N_14945);
xor UO_1964 (O_1964,N_14936,N_14882);
or UO_1965 (O_1965,N_14956,N_14916);
nor UO_1966 (O_1966,N_14950,N_14988);
xnor UO_1967 (O_1967,N_14937,N_14924);
and UO_1968 (O_1968,N_14948,N_14900);
nor UO_1969 (O_1969,N_14934,N_14875);
and UO_1970 (O_1970,N_14984,N_14879);
or UO_1971 (O_1971,N_14976,N_14995);
nand UO_1972 (O_1972,N_14881,N_14986);
nor UO_1973 (O_1973,N_14957,N_14956);
and UO_1974 (O_1974,N_14988,N_14877);
xnor UO_1975 (O_1975,N_14896,N_14936);
and UO_1976 (O_1976,N_14962,N_14875);
and UO_1977 (O_1977,N_14983,N_14981);
and UO_1978 (O_1978,N_14941,N_14959);
xor UO_1979 (O_1979,N_14912,N_14896);
nand UO_1980 (O_1980,N_14895,N_14919);
nor UO_1981 (O_1981,N_14997,N_14907);
nor UO_1982 (O_1982,N_14940,N_14982);
or UO_1983 (O_1983,N_14981,N_14906);
and UO_1984 (O_1984,N_14914,N_14908);
or UO_1985 (O_1985,N_14975,N_14961);
nor UO_1986 (O_1986,N_14950,N_14980);
or UO_1987 (O_1987,N_14908,N_14899);
and UO_1988 (O_1988,N_14963,N_14944);
xnor UO_1989 (O_1989,N_14966,N_14928);
nand UO_1990 (O_1990,N_14876,N_14962);
and UO_1991 (O_1991,N_14920,N_14896);
xor UO_1992 (O_1992,N_14930,N_14969);
nand UO_1993 (O_1993,N_14934,N_14958);
or UO_1994 (O_1994,N_14948,N_14925);
nor UO_1995 (O_1995,N_14875,N_14930);
or UO_1996 (O_1996,N_14995,N_14882);
and UO_1997 (O_1997,N_14958,N_14944);
nor UO_1998 (O_1998,N_14914,N_14950);
or UO_1999 (O_1999,N_14924,N_14980);
endmodule