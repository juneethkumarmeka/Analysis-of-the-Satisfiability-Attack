module basic_2000_20000_2500_10_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
or U0 (N_0,In_701,In_531);
nand U1 (N_1,In_112,In_1040);
nor U2 (N_2,In_987,In_1785);
or U3 (N_3,In_1774,In_1397);
nand U4 (N_4,In_629,In_1739);
nand U5 (N_5,In_1208,In_1884);
nand U6 (N_6,In_1944,In_1680);
or U7 (N_7,In_1351,In_756);
nor U8 (N_8,In_1897,In_265);
and U9 (N_9,In_214,In_951);
or U10 (N_10,In_475,In_247);
and U11 (N_11,In_1698,In_971);
or U12 (N_12,In_1487,In_1558);
or U13 (N_13,In_896,In_70);
nand U14 (N_14,In_774,In_542);
or U15 (N_15,In_727,In_988);
or U16 (N_16,In_697,In_1050);
and U17 (N_17,In_1297,In_1909);
and U18 (N_18,In_857,In_627);
and U19 (N_19,In_1098,In_464);
or U20 (N_20,In_577,In_1631);
nor U21 (N_21,In_362,In_428);
xor U22 (N_22,In_337,In_1824);
nor U23 (N_23,In_92,In_1654);
nand U24 (N_24,In_132,In_1950);
or U25 (N_25,In_1356,In_405);
xnor U26 (N_26,In_1580,In_1380);
and U27 (N_27,In_1541,In_384);
and U28 (N_28,In_39,In_1783);
nor U29 (N_29,In_729,In_830);
and U30 (N_30,In_947,In_1355);
nand U31 (N_31,In_888,In_928);
nor U32 (N_32,In_239,In_670);
or U33 (N_33,In_770,In_549);
and U34 (N_34,In_559,In_1434);
and U35 (N_35,In_849,In_166);
nor U36 (N_36,In_554,In_259);
and U37 (N_37,In_1693,In_938);
or U38 (N_38,In_1623,In_939);
nor U39 (N_39,In_1057,In_19);
xnor U40 (N_40,In_1894,In_930);
or U41 (N_41,In_1927,In_927);
xor U42 (N_42,In_1460,In_103);
nand U43 (N_43,In_110,In_906);
or U44 (N_44,In_1972,In_444);
nor U45 (N_45,In_759,In_412);
nand U46 (N_46,In_71,In_1074);
or U47 (N_47,In_1923,In_710);
nand U48 (N_48,In_1552,In_1864);
and U49 (N_49,In_173,In_413);
nor U50 (N_50,In_1300,In_1462);
nor U51 (N_51,In_1047,In_1327);
and U52 (N_52,In_1402,In_536);
nand U53 (N_53,In_1362,In_1499);
nand U54 (N_54,In_735,In_1117);
or U55 (N_55,In_1649,In_1592);
xnor U56 (N_56,In_739,In_530);
and U57 (N_57,In_42,In_284);
nand U58 (N_58,In_98,In_1214);
nor U59 (N_59,In_937,In_297);
xor U60 (N_60,In_1034,In_1875);
nand U61 (N_61,In_685,In_824);
and U62 (N_62,In_1557,In_1828);
nand U63 (N_63,In_661,In_1478);
nor U64 (N_64,In_1985,In_1603);
nand U65 (N_65,In_1448,In_203);
nand U66 (N_66,In_1643,In_365);
nor U67 (N_67,In_74,In_418);
nand U68 (N_68,In_105,In_1538);
nor U69 (N_69,In_354,In_1190);
xnor U70 (N_70,In_803,In_177);
or U71 (N_71,In_163,In_963);
or U72 (N_72,In_510,In_898);
nand U73 (N_73,In_1615,In_145);
or U74 (N_74,In_473,In_1852);
nand U75 (N_75,In_1674,In_1641);
or U76 (N_76,In_711,In_1629);
or U77 (N_77,In_1962,In_424);
and U78 (N_78,In_1498,In_47);
and U79 (N_79,In_76,In_872);
nor U80 (N_80,In_737,In_1539);
nor U81 (N_81,In_1319,In_1818);
or U82 (N_82,In_644,In_728);
or U83 (N_83,In_677,In_231);
nand U84 (N_84,In_814,In_144);
or U85 (N_85,In_257,In_1400);
nand U86 (N_86,In_488,In_180);
or U87 (N_87,In_1118,In_1743);
and U88 (N_88,In_168,In_507);
xnor U89 (N_89,In_1726,In_1350);
nor U90 (N_90,In_966,In_286);
or U91 (N_91,In_1266,In_1062);
or U92 (N_92,In_1999,In_1806);
nand U93 (N_93,In_1577,In_876);
and U94 (N_94,In_537,In_1090);
and U95 (N_95,In_1429,In_1720);
nand U96 (N_96,In_34,In_1604);
and U97 (N_97,In_512,In_1312);
or U98 (N_98,In_1826,In_1468);
nor U99 (N_99,In_659,In_1282);
and U100 (N_100,In_1287,In_371);
xnor U101 (N_101,In_1292,In_1598);
and U102 (N_102,In_376,In_218);
nand U103 (N_103,In_1871,In_969);
nor U104 (N_104,In_94,In_1229);
nor U105 (N_105,In_826,In_1017);
or U106 (N_106,In_120,In_639);
or U107 (N_107,In_448,In_1669);
or U108 (N_108,In_1167,In_1484);
and U109 (N_109,In_1914,In_280);
or U110 (N_110,In_1180,In_1861);
or U111 (N_111,In_911,In_1549);
xor U112 (N_112,In_82,In_916);
nand U113 (N_113,In_887,In_264);
nand U114 (N_114,In_1919,In_1157);
nand U115 (N_115,In_1134,In_658);
or U116 (N_116,In_1658,In_1796);
nor U117 (N_117,In_1801,In_1366);
nand U118 (N_118,In_1307,In_1224);
nor U119 (N_119,In_442,In_812);
nand U120 (N_120,In_845,In_890);
or U121 (N_121,In_1381,In_1389);
or U122 (N_122,In_1045,In_210);
nand U123 (N_123,In_1501,In_419);
and U124 (N_124,In_1430,In_1947);
nand U125 (N_125,In_246,In_1590);
nor U126 (N_126,In_1955,In_1236);
xor U127 (N_127,In_614,In_1372);
nand U128 (N_128,In_1281,In_1694);
nor U129 (N_129,In_625,In_792);
nor U130 (N_130,In_744,In_605);
or U131 (N_131,In_1020,In_1417);
nor U132 (N_132,In_1465,In_1857);
xor U133 (N_133,In_806,In_611);
nor U134 (N_134,In_1958,In_244);
or U135 (N_135,In_46,In_738);
and U136 (N_136,In_400,In_63);
and U137 (N_137,In_583,In_717);
nand U138 (N_138,In_1326,In_616);
nand U139 (N_139,In_1403,In_2);
nand U140 (N_140,In_278,In_1104);
nand U141 (N_141,In_275,In_55);
and U142 (N_142,In_313,In_1252);
nor U143 (N_143,In_1918,In_692);
and U144 (N_144,In_1187,In_1833);
nand U145 (N_145,In_1636,In_471);
and U146 (N_146,In_856,In_690);
and U147 (N_147,In_267,In_955);
or U148 (N_148,In_351,In_1264);
nand U149 (N_149,In_260,In_1761);
xor U150 (N_150,In_1168,In_1870);
nand U151 (N_151,In_1701,In_1271);
or U152 (N_152,In_1343,In_199);
xor U153 (N_153,In_408,In_702);
and U154 (N_154,In_1088,In_1511);
nor U155 (N_155,In_249,In_272);
or U156 (N_156,In_1655,In_1908);
nand U157 (N_157,In_1111,In_1866);
or U158 (N_158,In_946,In_1925);
or U159 (N_159,In_1110,In_1943);
and U160 (N_160,In_1702,In_1899);
or U161 (N_161,In_957,In_188);
xor U162 (N_162,In_613,In_569);
or U163 (N_163,In_1470,In_1325);
or U164 (N_164,In_716,In_491);
nor U165 (N_165,In_848,In_1677);
nor U166 (N_166,In_967,In_1814);
nor U167 (N_167,In_1469,In_1975);
nor U168 (N_168,In_1492,In_1442);
and U169 (N_169,In_1485,In_1787);
and U170 (N_170,In_1862,In_283);
nor U171 (N_171,In_327,In_1068);
nand U172 (N_172,In_1177,In_1627);
nor U173 (N_173,In_101,In_1522);
and U174 (N_174,In_708,In_1778);
or U175 (N_175,In_385,In_1995);
and U176 (N_176,In_1059,In_331);
xor U177 (N_177,In_1471,In_1757);
and U178 (N_178,In_1817,In_321);
or U179 (N_179,In_1219,In_1392);
nor U180 (N_180,In_722,In_808);
and U181 (N_181,In_1346,In_943);
or U182 (N_182,In_1363,In_1353);
nand U183 (N_183,In_1736,In_1574);
nand U184 (N_184,In_54,In_1732);
and U185 (N_185,In_1745,In_1974);
nor U186 (N_186,In_560,In_1707);
nor U187 (N_187,In_567,In_383);
nor U188 (N_188,In_1513,In_842);
xnor U189 (N_189,In_1012,In_1039);
and U190 (N_190,In_1846,In_509);
nand U191 (N_191,In_623,In_1291);
and U192 (N_192,In_1255,In_858);
and U193 (N_193,In_109,In_1008);
nand U194 (N_194,In_31,In_1415);
nand U195 (N_195,In_1225,In_575);
nand U196 (N_196,In_960,In_870);
or U197 (N_197,In_1929,In_1609);
or U198 (N_198,In_950,In_1051);
and U199 (N_199,In_343,In_771);
nand U200 (N_200,In_1044,In_146);
nor U201 (N_201,In_1205,In_1476);
or U202 (N_202,In_1223,In_1011);
nand U203 (N_203,In_1613,In_1210);
nor U204 (N_204,In_1595,In_1107);
nand U205 (N_205,In_1547,In_1788);
or U206 (N_206,In_1024,In_402);
nor U207 (N_207,In_223,In_26);
or U208 (N_208,In_1128,In_529);
and U209 (N_209,In_454,In_1411);
xor U210 (N_210,In_443,In_116);
or U211 (N_211,In_1737,In_778);
and U212 (N_212,In_433,In_436);
nor U213 (N_213,In_1527,In_1903);
and U214 (N_214,In_130,In_645);
and U215 (N_215,In_520,In_1338);
nor U216 (N_216,In_1466,In_1583);
nand U217 (N_217,In_1530,In_1029);
and U218 (N_218,In_1032,In_336);
nand U219 (N_219,In_310,In_1644);
nand U220 (N_220,In_682,In_62);
xor U221 (N_221,In_694,In_204);
nor U222 (N_222,In_1808,In_964);
nor U223 (N_223,In_1932,In_1069);
or U224 (N_224,In_827,In_1477);
nor U225 (N_225,In_1676,In_724);
and U226 (N_226,In_1184,In_1917);
nor U227 (N_227,In_435,In_638);
nor U228 (N_228,In_407,In_820);
or U229 (N_229,In_393,In_1653);
nand U230 (N_230,In_1868,In_1869);
nor U231 (N_231,In_411,In_1172);
and U232 (N_232,In_1775,In_36);
and U233 (N_233,In_1838,In_871);
and U234 (N_234,In_1670,In_292);
or U235 (N_235,In_463,In_1865);
nor U236 (N_236,In_736,In_882);
or U237 (N_237,In_115,In_60);
and U238 (N_238,In_1145,In_1594);
xnor U239 (N_239,In_620,In_348);
and U240 (N_240,In_1367,In_1815);
xnor U241 (N_241,In_482,In_674);
or U242 (N_242,In_1130,In_483);
nand U243 (N_243,In_1451,In_176);
or U244 (N_244,In_1673,In_501);
or U245 (N_245,In_1555,In_1352);
or U246 (N_246,In_1197,In_404);
nand U247 (N_247,In_1892,In_1162);
nor U248 (N_248,In_929,In_821);
nor U249 (N_249,In_1769,In_1435);
nand U250 (N_250,In_832,In_1393);
and U251 (N_251,In_519,In_652);
nor U252 (N_252,In_16,In_32);
or U253 (N_253,In_1333,In_22);
nor U254 (N_254,In_459,In_768);
nor U255 (N_255,In_1990,In_1457);
nor U256 (N_256,In_953,In_1794);
nand U257 (N_257,In_1863,In_485);
nand U258 (N_258,In_804,In_77);
nor U259 (N_259,In_1922,In_734);
xnor U260 (N_260,In_797,In_308);
nor U261 (N_261,In_1375,In_841);
or U262 (N_262,In_1821,In_619);
nand U263 (N_263,In_1964,In_1751);
nor U264 (N_264,In_1533,In_815);
or U265 (N_265,In_174,In_135);
xor U266 (N_266,In_401,In_344);
and U267 (N_267,In_170,In_1898);
and U268 (N_268,In_477,In_1217);
xor U269 (N_269,In_1009,In_1165);
or U270 (N_270,In_1405,In_783);
and U271 (N_271,In_158,In_1792);
and U272 (N_272,In_1315,In_968);
or U273 (N_273,In_1708,In_339);
and U274 (N_274,In_587,In_245);
nor U275 (N_275,In_9,In_865);
nor U276 (N_276,In_279,In_87);
nor U277 (N_277,In_1073,In_1108);
and U278 (N_278,In_923,In_965);
xnor U279 (N_279,In_1048,In_1685);
or U280 (N_280,In_905,In_1311);
and U281 (N_281,In_1554,In_1756);
and U282 (N_282,In_506,In_1961);
nand U283 (N_283,In_1683,In_1733);
nor U284 (N_284,In_982,In_599);
and U285 (N_285,In_1013,In_1119);
and U286 (N_286,In_489,In_117);
and U287 (N_287,In_1939,In_1399);
and U288 (N_288,In_184,In_863);
or U289 (N_289,In_102,In_1998);
nor U290 (N_290,In_23,In_139);
and U291 (N_291,In_822,In_1759);
xnor U292 (N_292,In_977,In_538);
xor U293 (N_293,In_1610,In_1404);
nor U294 (N_294,In_791,In_1856);
nand U295 (N_295,In_131,In_192);
nand U296 (N_296,In_1773,In_455);
nor U297 (N_297,In_367,In_1886);
nand U298 (N_298,In_779,In_684);
nor U299 (N_299,In_466,In_975);
nor U300 (N_300,In_1719,In_979);
nand U301 (N_301,In_1005,In_1585);
and U302 (N_302,In_521,In_582);
or U303 (N_303,In_976,In_162);
or U304 (N_304,In_1387,In_228);
xor U305 (N_305,In_607,In_72);
nand U306 (N_306,In_1934,In_1959);
nor U307 (N_307,In_1647,In_360);
nor U308 (N_308,In_949,In_1444);
and U309 (N_309,In_1486,In_978);
and U310 (N_310,In_256,In_972);
nor U311 (N_311,In_113,In_1729);
nand U312 (N_312,In_478,In_1094);
or U313 (N_313,In_1900,In_755);
xor U314 (N_314,In_837,In_450);
or U315 (N_315,In_1341,In_1406);
or U316 (N_316,In_688,In_589);
xnor U317 (N_317,In_894,In_10);
and U318 (N_318,In_1529,In_1369);
nand U319 (N_319,In_998,In_1867);
nor U320 (N_320,In_1370,In_1176);
and U321 (N_321,In_762,In_1679);
nor U322 (N_322,In_631,In_1945);
nand U323 (N_323,In_1063,In_370);
or U324 (N_324,In_44,In_726);
and U325 (N_325,In_1046,In_1309);
and U326 (N_326,In_458,In_334);
nand U327 (N_327,In_504,In_1018);
or U328 (N_328,In_1087,In_942);
nand U329 (N_329,In_838,In_1154);
or U330 (N_330,In_1690,In_1185);
or U331 (N_331,In_1378,In_142);
nor U332 (N_332,In_1780,In_1593);
or U333 (N_333,In_1606,In_1278);
and U334 (N_334,In_1192,In_43);
and U335 (N_335,In_919,In_271);
nand U336 (N_336,In_99,In_1666);
or U337 (N_337,In_1078,In_1445);
nor U338 (N_338,In_1859,In_1933);
and U339 (N_339,In_991,In_1388);
nor U340 (N_340,In_307,In_1504);
or U341 (N_341,In_1576,In_1618);
and U342 (N_342,In_219,In_1956);
or U343 (N_343,In_816,In_864);
nand U344 (N_344,In_196,In_1668);
and U345 (N_345,In_1456,In_1556);
nor U346 (N_346,In_390,In_95);
or U347 (N_347,In_1239,In_1042);
and U348 (N_348,In_1201,In_1936);
or U349 (N_349,In_1268,In_1722);
and U350 (N_350,In_1957,In_1251);
nand U351 (N_351,In_349,In_441);
xnor U352 (N_352,In_83,In_1749);
nand U353 (N_353,In_819,In_997);
nand U354 (N_354,In_628,In_200);
or U355 (N_355,In_1842,In_303);
xor U356 (N_356,In_372,In_1630);
and U357 (N_357,In_730,In_273);
or U358 (N_358,In_1500,In_1037);
nor U359 (N_359,In_1276,In_472);
nor U360 (N_360,In_341,In_1439);
nand U361 (N_361,In_593,In_741);
xor U362 (N_362,In_785,In_1077);
nor U363 (N_363,In_789,In_193);
and U364 (N_364,In_1688,In_1028);
and U365 (N_365,In_563,In_1202);
nor U366 (N_366,In_1124,In_657);
nor U367 (N_367,In_1542,In_689);
nor U368 (N_368,In_1888,In_282);
nand U369 (N_369,In_1575,In_1571);
xor U370 (N_370,In_884,In_853);
xor U371 (N_371,In_794,In_1441);
or U372 (N_372,In_1713,In_1438);
nor U373 (N_373,In_835,In_434);
or U374 (N_374,In_1376,In_1133);
and U375 (N_375,In_1663,In_1083);
nand U376 (N_376,In_319,In_1335);
nand U377 (N_377,In_746,In_836);
xnor U378 (N_378,In_1030,In_1310);
xor U379 (N_379,In_1298,In_201);
and U380 (N_380,In_1318,In_300);
nor U381 (N_381,In_1426,In_1682);
or U382 (N_382,In_50,In_294);
nor U383 (N_383,In_1601,In_749);
nor U384 (N_384,In_585,In_931);
nand U385 (N_385,In_432,In_1772);
xnor U386 (N_386,In_883,In_576);
and U387 (N_387,In_1832,In_1259);
and U388 (N_388,In_517,In_781);
xnor U389 (N_389,In_213,In_899);
xnor U390 (N_390,In_106,In_346);
xor U391 (N_391,In_1109,In_750);
or U392 (N_392,In_484,In_1758);
xor U393 (N_393,In_137,In_1716);
and U394 (N_394,In_637,In_233);
xnor U395 (N_395,In_1710,In_846);
or U396 (N_396,In_250,In_129);
and U397 (N_397,In_93,In_765);
nor U398 (N_398,In_956,In_1887);
nor U399 (N_399,In_1851,In_801);
xor U400 (N_400,In_1004,In_1126);
nand U401 (N_401,In_309,In_361);
nor U402 (N_402,In_190,In_40);
nor U403 (N_403,In_533,In_45);
and U404 (N_404,In_1093,In_1967);
nand U405 (N_405,In_745,In_391);
or U406 (N_406,In_1215,In_468);
or U407 (N_407,In_232,In_1510);
and U408 (N_408,In_123,In_119);
or U409 (N_409,In_1283,In_1033);
nor U410 (N_410,In_1681,In_1473);
and U411 (N_411,In_1616,In_641);
xnor U412 (N_412,In_945,In_211);
xor U413 (N_413,In_328,In_1531);
nand U414 (N_414,In_406,In_209);
and U415 (N_415,In_457,In_378);
or U416 (N_416,In_1728,In_954);
or U417 (N_417,In_752,In_1843);
and U418 (N_418,In_229,In_290);
nor U419 (N_419,In_438,In_1599);
xnor U420 (N_420,In_557,In_1019);
or U421 (N_421,In_1305,In_1368);
nand U422 (N_422,In_1247,In_470);
nand U423 (N_423,In_1891,In_1452);
and U424 (N_424,In_1328,In_1304);
or U425 (N_425,In_1901,In_1570);
or U426 (N_426,In_1408,In_151);
or U427 (N_427,In_396,In_1453);
or U428 (N_428,In_782,In_1991);
xor U429 (N_429,In_487,In_1873);
nand U430 (N_430,In_527,In_1786);
nand U431 (N_431,In_1014,In_875);
nand U432 (N_432,In_635,In_989);
or U433 (N_433,In_636,In_523);
nand U434 (N_434,In_1482,In_1881);
nand U435 (N_435,In_451,In_1149);
and U436 (N_436,In_1596,In_1672);
or U437 (N_437,In_175,In_1260);
nor U438 (N_438,In_414,In_1686);
xor U439 (N_439,In_1520,In_134);
xnor U440 (N_440,In_602,In_695);
and U441 (N_441,In_61,In_540);
and U442 (N_442,In_1249,In_1874);
nor U443 (N_443,In_1007,In_1582);
nand U444 (N_444,In_1855,In_1802);
and U445 (N_445,In_1213,In_426);
nand U446 (N_446,In_1755,In_573);
or U447 (N_447,In_1112,In_1407);
nand U448 (N_448,In_1611,In_1921);
or U449 (N_449,In_1491,In_1203);
nand U450 (N_450,In_1220,In_1099);
xor U451 (N_451,In_1459,In_1173);
nor U452 (N_452,In_1543,In_20);
nor U453 (N_453,In_254,In_1479);
nand U454 (N_454,In_1617,In_1398);
nor U455 (N_455,In_78,In_240);
nand U456 (N_456,In_1602,In_230);
and U457 (N_457,In_1420,In_633);
nand U458 (N_458,In_1067,In_1614);
or U459 (N_459,In_1000,In_1242);
or U460 (N_460,In_543,In_649);
xnor U461 (N_461,In_1289,In_1170);
xor U462 (N_462,In_525,In_221);
and U463 (N_463,In_235,In_1928);
nor U464 (N_464,In_1505,In_80);
or U465 (N_465,In_1506,In_225);
or U466 (N_466,In_14,In_860);
and U467 (N_467,In_1391,In_111);
and U468 (N_468,In_1810,In_298);
or U469 (N_469,In_1515,In_609);
nor U470 (N_470,In_114,In_1935);
nor U471 (N_471,In_497,In_669);
xnor U472 (N_472,In_1896,In_1140);
nor U473 (N_473,In_364,In_25);
and U474 (N_474,In_1537,In_1290);
or U475 (N_475,In_1799,In_1508);
nor U476 (N_476,In_306,In_1526);
nand U477 (N_477,In_1997,In_171);
or U478 (N_478,In_161,In_1082);
nand U479 (N_479,In_676,In_1514);
and U480 (N_480,In_1054,In_1132);
nand U481 (N_481,In_843,In_1830);
nand U482 (N_482,In_403,In_1348);
and U483 (N_483,In_719,In_1700);
xnor U484 (N_484,In_1178,In_1518);
nor U485 (N_485,In_1804,In_1730);
nand U486 (N_486,In_809,In_921);
or U487 (N_487,In_597,In_1241);
nor U488 (N_488,In_1839,In_253);
nor U489 (N_489,In_48,In_227);
nand U490 (N_490,In_828,In_382);
nand U491 (N_491,In_667,In_1916);
or U492 (N_492,In_1951,In_675);
or U493 (N_493,In_1924,In_224);
or U494 (N_494,In_248,In_970);
xnor U495 (N_495,In_1568,In_160);
nor U496 (N_496,In_88,In_236);
nor U497 (N_497,In_1231,In_1904);
and U498 (N_498,In_1373,In_355);
nand U499 (N_499,In_1639,In_1805);
nand U500 (N_500,In_1640,In_1910);
nor U501 (N_501,In_1461,In_1136);
nor U502 (N_502,In_1360,In_601);
nor U503 (N_503,In_1645,In_1760);
and U504 (N_504,In_1969,In_1147);
or U505 (N_505,In_1137,In_1579);
nand U506 (N_506,In_1589,In_1450);
and U507 (N_507,In_1129,In_1727);
nor U508 (N_508,In_37,In_748);
or U509 (N_509,In_1841,In_1978);
and U510 (N_510,In_1102,In_1827);
and U511 (N_511,In_167,In_1718);
and U512 (N_512,In_1809,In_347);
nand U513 (N_513,In_1714,In_1416);
and U514 (N_514,In_1764,In_1212);
or U515 (N_515,In_269,In_1175);
nand U516 (N_516,In_461,In_775);
or U517 (N_517,In_1207,In_1424);
and U518 (N_518,In_798,In_1243);
and U519 (N_519,In_1056,In_1877);
and U520 (N_520,In_1931,In_672);
or U521 (N_521,In_1971,In_24);
nand U522 (N_522,In_1121,In_934);
or U523 (N_523,In_366,In_564);
nand U524 (N_524,In_1277,In_430);
nand U525 (N_525,In_263,In_12);
nor U526 (N_526,In_1572,In_544);
and U527 (N_527,In_800,In_266);
nand U528 (N_528,In_1777,In_7);
nor U529 (N_529,In_1221,In_1535);
xnor U530 (N_530,In_1027,In_1100);
nand U531 (N_531,In_1540,In_1354);
and U532 (N_532,In_1748,In_445);
or U533 (N_533,In_855,In_479);
nand U534 (N_534,In_663,In_154);
xor U535 (N_535,In_255,In_1497);
and U536 (N_536,In_1633,In_1994);
xnor U537 (N_537,In_387,In_1106);
or U538 (N_538,In_617,In_693);
nor U539 (N_539,In_914,In_1060);
and U540 (N_540,In_386,In_301);
nor U541 (N_541,In_1902,In_541);
nor U542 (N_542,In_881,In_1553);
and U543 (N_543,In_84,In_571);
or U544 (N_544,In_1371,In_1905);
nand U545 (N_545,In_1807,In_85);
and U546 (N_546,In_1031,In_653);
or U547 (N_547,In_141,In_121);
nor U548 (N_548,In_1652,In_302);
nand U549 (N_549,In_1996,In_1963);
nand U550 (N_550,In_1306,In_895);
and U551 (N_551,In_1089,In_1308);
or U552 (N_552,In_1564,In_1822);
nor U553 (N_553,In_133,In_18);
nand U554 (N_554,In_1689,In_6);
and U555 (N_555,In_1324,In_152);
xor U556 (N_556,In_1503,In_183);
xnor U557 (N_557,In_1767,In_565);
nand U558 (N_558,In_1819,In_1263);
and U559 (N_559,In_920,In_1320);
and U560 (N_560,In_494,In_714);
nor U561 (N_561,In_1753,In_1228);
or U562 (N_562,In_1699,In_67);
nor U563 (N_563,In_1637,In_159);
and U564 (N_564,In_547,In_417);
nand U565 (N_565,In_1752,In_1626);
xor U566 (N_566,In_1848,In_195);
nand U567 (N_567,In_904,In_1101);
and U568 (N_568,In_1322,In_1628);
and U569 (N_569,In_948,In_469);
and U570 (N_570,In_369,In_1695);
and U571 (N_571,In_900,In_902);
or U572 (N_572,In_1041,In_994);
or U573 (N_573,In_935,In_11);
or U574 (N_574,In_1742,In_1938);
and U575 (N_575,In_493,In_1559);
nor U576 (N_576,In_480,In_699);
and U577 (N_577,In_5,In_108);
and U578 (N_578,In_1664,In_1567);
and U579 (N_579,In_909,In_1196);
and U580 (N_580,In_1703,In_1684);
and U581 (N_581,In_1660,In_1091);
and U582 (N_582,In_985,In_182);
nand U583 (N_583,In_118,In_1545);
nor U584 (N_584,In_1746,In_462);
xnor U585 (N_585,In_1776,In_581);
nand U586 (N_586,In_1238,In_551);
nand U587 (N_587,In_1097,In_1174);
nand U588 (N_588,In_1002,In_1548);
and U589 (N_589,In_912,In_186);
xor U590 (N_590,In_795,In_524);
nor U591 (N_591,In_723,In_1992);
or U592 (N_592,In_1015,In_793);
nor U593 (N_593,In_1127,In_1948);
and U594 (N_594,In_908,In_1075);
and U595 (N_595,In_320,In_165);
and U596 (N_596,In_1584,In_3);
and U597 (N_597,In_304,In_591);
nand U598 (N_598,In_817,In_503);
nand U599 (N_599,In_1296,In_1454);
nor U600 (N_600,In_1563,In_1973);
or U601 (N_601,In_1474,In_1519);
and U602 (N_602,In_381,In_194);
xnor U603 (N_603,In_1779,In_878);
or U604 (N_604,In_1854,In_1987);
or U605 (N_605,In_505,In_35);
xnor U606 (N_606,In_868,In_594);
and U607 (N_607,In_936,In_604);
and U608 (N_608,In_38,In_1770);
nor U609 (N_609,In_1467,In_1141);
xnor U610 (N_610,In_992,In_570);
nor U611 (N_611,In_299,In_315);
nand U612 (N_612,In_352,In_270);
nand U613 (N_613,In_1161,In_1364);
and U614 (N_614,In_786,In_1560);
nor U615 (N_615,In_511,In_237);
nand U616 (N_616,In_73,In_1744);
or U617 (N_617,In_353,In_1820);
and U618 (N_618,In_1206,In_1735);
and U619 (N_619,In_558,In_243);
or U620 (N_620,In_712,In_831);
nor U621 (N_621,In_1412,In_1302);
nand U622 (N_622,In_397,In_1550);
nand U623 (N_623,In_1960,In_1432);
nand U624 (N_624,In_335,In_1494);
and U625 (N_625,In_97,In_664);
or U626 (N_626,In_1493,In_1706);
and U627 (N_627,In_207,In_1464);
or U628 (N_628,In_995,In_1591);
and U629 (N_629,In_643,In_1544);
and U630 (N_630,In_1386,In_1285);
and U631 (N_631,In_422,In_1656);
nand U632 (N_632,In_1665,In_743);
and U633 (N_633,In_874,In_754);
nor U634 (N_634,In_958,In_1650);
nor U635 (N_635,In_706,In_332);
or U636 (N_636,In_1692,In_656);
or U637 (N_637,In_1427,In_854);
or U638 (N_638,In_4,In_1913);
or U639 (N_639,In_30,In_1233);
nor U640 (N_640,In_640,In_788);
nor U641 (N_641,In_1988,In_1872);
nor U642 (N_642,In_1731,In_285);
or U643 (N_643,In_586,In_217);
nor U644 (N_644,In_686,In_1395);
nor U645 (N_645,In_681,In_647);
nor U646 (N_646,In_1984,In_65);
xor U647 (N_647,In_1638,In_1085);
and U648 (N_648,In_1625,In_15);
and U649 (N_649,In_1359,In_1115);
or U650 (N_650,In_1198,In_873);
or U651 (N_651,In_514,In_1261);
nor U652 (N_652,In_1534,In_446);
xnor U653 (N_653,In_867,In_1835);
and U654 (N_654,In_1659,In_1125);
xnor U655 (N_655,In_1344,In_703);
nand U656 (N_656,In_705,In_305);
and U657 (N_657,In_17,In_410);
and U658 (N_658,In_1120,In_598);
xnor U659 (N_659,In_1222,In_1347);
or U660 (N_660,In_421,In_877);
nand U661 (N_661,In_1768,In_709);
nor U662 (N_662,In_191,In_409);
nand U663 (N_663,In_1103,In_1937);
and U664 (N_664,In_449,In_548);
nand U665 (N_665,In_632,In_276);
and U666 (N_666,In_1182,In_700);
nor U667 (N_667,In_220,In_453);
or U668 (N_668,In_1723,In_148);
nor U669 (N_669,In_1691,In_289);
and U670 (N_670,In_89,In_147);
nor U671 (N_671,In_545,In_1342);
nor U672 (N_672,In_818,In_492);
and U673 (N_673,In_359,In_1840);
xnor U674 (N_674,In_1704,In_1321);
nand U675 (N_675,In_880,In_1160);
nor U676 (N_676,In_1845,In_216);
and U677 (N_677,In_1349,In_725);
nor U678 (N_678,In_1619,In_379);
or U679 (N_679,In_1717,In_772);
or U680 (N_680,In_721,In_1662);
xor U681 (N_681,In_910,In_790);
nor U682 (N_682,In_1878,In_1235);
or U683 (N_683,In_606,In_1949);
and U684 (N_684,In_1385,In_747);
or U685 (N_685,In_1295,In_1816);
and U686 (N_686,In_1850,In_1358);
and U687 (N_687,In_357,In_28);
or U688 (N_688,In_1293,In_1171);
or U689 (N_689,In_1357,In_740);
or U690 (N_690,In_392,In_1152);
and U691 (N_691,In_1023,In_1483);
or U692 (N_692,In_1377,In_1025);
or U693 (N_693,In_1741,In_859);
nor U694 (N_694,In_388,In_1186);
or U695 (N_695,In_1784,In_1284);
nand U696 (N_696,In_1472,In_1163);
nor U697 (N_697,In_751,In_715);
or U698 (N_698,In_1158,In_1270);
or U699 (N_699,In_802,In_13);
or U700 (N_700,In_897,In_1144);
nor U701 (N_701,In_1265,In_1218);
nor U702 (N_702,In_777,In_1495);
or U703 (N_703,In_322,In_918);
and U704 (N_704,In_107,In_839);
nand U705 (N_705,In_1605,In_654);
nor U706 (N_706,In_1734,In_1329);
xnor U707 (N_707,In_1058,In_981);
or U708 (N_708,In_1254,In_993);
and U709 (N_709,In_1648,In_1715);
nor U710 (N_710,In_1080,In_1431);
xor U711 (N_711,In_1642,In_476);
and U712 (N_712,In_1954,In_329);
or U713 (N_713,In_1622,In_1907);
and U714 (N_714,In_465,In_1725);
or U715 (N_715,In_1092,In_1191);
and U716 (N_716,In_1551,In_780);
or U717 (N_717,In_1789,In_1114);
or U718 (N_718,In_358,In_917);
xnor U719 (N_719,In_518,In_1523);
and U720 (N_720,In_691,In_1860);
or U721 (N_721,In_1301,In_1740);
xor U722 (N_722,In_1952,In_49);
nand U723 (N_723,In_508,In_330);
xor U724 (N_724,In_1879,In_399);
nor U725 (N_725,In_481,In_1546);
nor U726 (N_726,In_608,In_1885);
nor U727 (N_727,In_1274,In_546);
nand U728 (N_728,In_1334,In_287);
nand U729 (N_729,In_1064,In_687);
nand U730 (N_730,In_91,In_1288);
nor U731 (N_731,In_1941,In_460);
nand U732 (N_732,In_986,In_138);
xnor U733 (N_733,In_377,In_274);
nand U734 (N_734,In_668,In_251);
nand U735 (N_735,In_1061,In_179);
nor U736 (N_736,In_1148,In_630);
and U737 (N_737,In_961,In_596);
nor U738 (N_738,In_1488,In_1314);
nor U739 (N_739,In_1079,In_1428);
or U740 (N_740,In_1597,In_610);
and U741 (N_741,In_1750,In_27);
nor U742 (N_742,In_1390,In_733);
and U743 (N_743,In_1425,In_155);
xor U744 (N_744,In_143,In_1463);
or U745 (N_745,In_915,In_1588);
or U746 (N_746,In_974,In_1394);
xor U747 (N_747,In_941,In_1621);
nor U748 (N_748,In_368,In_983);
nand U749 (N_749,In_539,In_1795);
nor U750 (N_750,In_1612,In_773);
and U751 (N_751,In_1339,In_1687);
or U752 (N_752,In_502,In_1382);
nand U753 (N_753,In_1248,In_1035);
nand U754 (N_754,In_1829,In_1711);
nand U755 (N_755,In_1065,In_1766);
xnor U756 (N_756,In_590,In_1607);
or U757 (N_757,In_1262,In_1237);
nor U758 (N_758,In_398,In_1724);
xor U759 (N_759,In_526,In_415);
or U760 (N_760,In_1374,In_893);
and U761 (N_761,In_1986,In_704);
or U762 (N_762,In_932,In_833);
nor U763 (N_763,In_683,In_1496);
and U764 (N_764,In_238,In_241);
or U765 (N_765,In_58,In_496);
and U766 (N_766,In_1244,In_423);
nor U767 (N_767,In_732,In_1);
nand U768 (N_768,In_634,In_825);
nand U769 (N_769,In_317,In_1313);
xnor U770 (N_770,In_1516,In_164);
or U771 (N_771,In_456,In_1490);
and U772 (N_772,In_153,In_281);
and U773 (N_773,In_933,In_1116);
nand U774 (N_774,In_1524,In_420);
and U775 (N_775,In_104,In_764);
nand U776 (N_776,In_650,In_1299);
nor U777 (N_777,In_149,In_1413);
or U778 (N_778,In_125,In_1797);
xor U779 (N_779,In_980,In_796);
or U780 (N_780,In_618,In_1250);
nor U781 (N_781,In_622,In_262);
or U782 (N_782,In_886,In_1798);
or U783 (N_783,In_1781,In_840);
nor U784 (N_784,In_474,In_1883);
nand U785 (N_785,In_178,In_1273);
and U786 (N_786,In_532,In_498);
or U787 (N_787,In_592,In_1423);
or U788 (N_788,In_731,In_1143);
nand U789 (N_789,In_718,In_373);
nor U790 (N_790,In_1858,In_124);
nand U791 (N_791,In_522,In_150);
nand U792 (N_792,In_984,In_81);
nand U793 (N_793,In_844,In_1847);
and U794 (N_794,In_1038,In_1076);
nand U795 (N_795,In_1849,In_753);
and U796 (N_796,In_342,In_64);
and U797 (N_797,In_1257,In_1246);
and U798 (N_798,In_1072,In_568);
nand U799 (N_799,In_891,In_431);
nor U800 (N_800,In_1661,In_1139);
and U801 (N_801,In_33,In_1361);
and U802 (N_802,In_452,In_1036);
nor U803 (N_803,In_555,In_326);
nor U804 (N_804,In_258,In_1624);
xnor U805 (N_805,In_996,In_1525);
or U806 (N_806,In_41,In_1517);
or U807 (N_807,In_1436,In_427);
nand U808 (N_808,In_1365,In_56);
or U809 (N_809,In_680,In_562);
nand U810 (N_810,In_1586,In_1006);
or U811 (N_811,In_1812,In_1021);
nor U812 (N_812,In_642,In_1245);
or U813 (N_813,In_600,In_86);
nor U814 (N_814,In_1294,In_338);
or U815 (N_815,In_1230,In_1976);
nor U816 (N_816,In_1437,In_579);
nand U817 (N_817,In_850,In_75);
and U818 (N_818,In_96,In_1081);
xnor U819 (N_819,In_1876,In_678);
nor U820 (N_820,In_1317,In_1447);
nor U821 (N_821,In_1286,In_651);
and U822 (N_822,In_1489,In_198);
or U823 (N_823,In_1016,In_467);
nor U824 (N_824,In_208,In_1316);
nand U825 (N_825,In_1323,In_1193);
xor U826 (N_826,In_1480,In_1823);
nor U827 (N_827,In_1890,In_1953);
nor U828 (N_828,In_1738,In_1512);
nor U829 (N_829,In_813,In_776);
and U830 (N_830,In_671,In_769);
or U831 (N_831,In_1793,In_1421);
or U832 (N_832,In_439,In_1181);
and U833 (N_833,In_758,In_862);
and U834 (N_834,In_973,In_1410);
and U835 (N_835,In_513,In_1942);
nor U836 (N_836,In_1071,In_126);
nand U837 (N_837,In_1893,In_940);
nor U838 (N_838,In_1179,In_1790);
and U839 (N_839,In_1940,In_805);
xnor U840 (N_840,In_1123,In_1414);
nor U841 (N_841,In_8,In_1536);
or U842 (N_842,In_1565,In_1825);
nand U843 (N_843,In_1146,In_1449);
nor U844 (N_844,In_52,In_1001);
and U845 (N_845,In_1791,In_293);
and U846 (N_846,In_277,In_1880);
and U847 (N_847,In_799,In_140);
or U848 (N_848,In_892,In_1747);
and U849 (N_849,In_316,In_1209);
or U850 (N_850,In_447,In_1211);
and U851 (N_851,In_1697,In_440);
nand U852 (N_852,In_1131,In_312);
nand U853 (N_853,In_1573,In_528);
or U854 (N_854,In_851,In_1267);
nor U855 (N_855,In_1979,In_100);
nor U856 (N_856,In_1253,In_1443);
nor U857 (N_857,In_847,In_1561);
xor U858 (N_858,In_1240,In_534);
nor U859 (N_859,In_234,In_553);
xor U860 (N_860,In_1678,In_156);
nor U861 (N_861,In_852,In_1303);
and U862 (N_862,In_787,In_1234);
or U863 (N_863,In_1419,In_172);
nand U864 (N_864,In_1113,In_1084);
or U865 (N_865,In_1600,In_869);
xor U866 (N_866,In_1022,In_655);
or U867 (N_867,In_1782,In_552);
nand U868 (N_868,In_885,In_807);
xor U869 (N_869,In_1159,In_696);
or U870 (N_870,In_1155,In_1345);
and U871 (N_871,In_1834,In_962);
and U872 (N_872,In_615,In_1153);
nand U873 (N_873,In_1532,In_889);
and U874 (N_874,In_572,In_136);
nand U875 (N_875,In_296,In_202);
nor U876 (N_876,In_580,In_242);
and U877 (N_877,In_1275,In_53);
and U878 (N_878,In_901,In_1970);
xor U879 (N_879,In_425,In_1667);
nor U880 (N_880,In_1010,In_1138);
nand U881 (N_881,In_222,In_1280);
nand U882 (N_882,In_866,In_1330);
and U883 (N_883,In_1151,In_323);
nor U884 (N_884,In_1232,In_646);
nand U885 (N_885,In_1164,In_500);
nand U886 (N_886,In_333,In_157);
nor U887 (N_887,In_1566,In_1977);
nand U888 (N_888,In_1980,In_345);
nor U889 (N_889,In_57,In_1502);
and U890 (N_890,In_291,In_128);
and U891 (N_891,In_1446,In_226);
nand U892 (N_892,In_1227,In_1721);
nand U893 (N_893,In_490,In_999);
or U894 (N_894,In_288,In_1657);
nor U895 (N_895,In_584,In_1216);
or U896 (N_896,In_51,In_679);
nand U897 (N_897,In_624,In_1528);
nand U898 (N_898,In_1632,In_698);
xor U899 (N_899,In_1142,In_21);
or U900 (N_900,In_1383,In_811);
nor U901 (N_901,In_0,In_395);
or U902 (N_902,In_922,In_1475);
or U903 (N_903,In_29,In_861);
xnor U904 (N_904,In_595,In_1053);
nand U905 (N_905,In_1269,In_1831);
xor U906 (N_906,In_766,In_1169);
xor U907 (N_907,In_516,In_1981);
or U908 (N_908,In_1150,In_1578);
or U909 (N_909,In_90,In_1095);
nor U910 (N_910,In_1509,In_1562);
nand U911 (N_911,In_363,In_1912);
xor U912 (N_912,In_1811,In_1003);
nor U913 (N_913,In_1844,In_1920);
nand U914 (N_914,In_1384,In_1418);
or U915 (N_915,In_375,In_181);
nor U916 (N_916,In_784,In_1122);
nand U917 (N_917,In_205,In_665);
nand U918 (N_918,In_1635,In_1521);
or U919 (N_919,In_1340,In_1837);
xor U920 (N_920,In_197,In_1455);
or U921 (N_921,In_187,In_1026);
xor U922 (N_922,In_1675,In_325);
and U923 (N_923,In_1272,In_834);
or U924 (N_924,In_1765,In_1055);
nor U925 (N_925,In_763,In_1396);
xor U926 (N_926,In_1993,In_416);
or U927 (N_927,In_1966,In_713);
nand U928 (N_928,In_268,In_1096);
nor U929 (N_929,In_925,In_588);
nand U930 (N_930,In_1587,In_380);
or U931 (N_931,In_1634,In_79);
nand U932 (N_932,In_1895,In_1889);
and U933 (N_933,In_189,In_913);
xor U934 (N_934,In_1800,In_1043);
or U935 (N_935,In_1705,In_311);
or U936 (N_936,In_1946,In_495);
and U937 (N_937,In_1926,In_389);
xor U938 (N_938,In_903,In_1762);
nand U939 (N_939,In_1337,In_621);
nand U940 (N_940,In_1696,In_1651);
nand U941 (N_941,In_1422,In_1379);
and U942 (N_942,In_879,In_394);
nand U943 (N_943,In_535,In_1401);
or U944 (N_944,In_1803,In_1279);
nor U945 (N_945,In_1195,In_1204);
or U946 (N_946,In_1433,In_612);
or U947 (N_947,In_1194,In_429);
and U948 (N_948,In_561,In_1982);
or U949 (N_949,In_318,In_1989);
and U950 (N_950,In_1853,In_1569);
nor U951 (N_951,In_486,In_1965);
and U952 (N_952,In_760,In_1332);
and U953 (N_953,In_1166,In_1771);
xor U954 (N_954,In_1507,In_1189);
and U955 (N_955,In_1066,In_1156);
and U956 (N_956,In_1712,In_660);
nor U957 (N_957,In_314,In_122);
and U958 (N_958,In_907,In_515);
nor U959 (N_959,In_1709,In_673);
or U960 (N_960,In_574,In_1409);
nor U961 (N_961,In_212,In_1258);
or U962 (N_962,In_1763,In_1049);
and U963 (N_963,In_185,In_550);
nand U964 (N_964,In_924,In_662);
or U965 (N_965,In_1671,In_1911);
nand U966 (N_966,In_1983,In_707);
nor U967 (N_967,In_59,In_1200);
or U968 (N_968,In_1070,In_68);
nand U969 (N_969,In_374,In_1813);
nor U970 (N_970,In_1968,In_1458);
nand U971 (N_971,In_1331,In_1256);
nor U972 (N_972,In_810,In_990);
nor U973 (N_973,In_206,In_1915);
nand U974 (N_974,In_1336,In_1608);
or U975 (N_975,In_1581,In_829);
nand U976 (N_976,In_757,In_1052);
nor U977 (N_977,In_1105,In_626);
and U978 (N_978,In_1135,In_295);
and U979 (N_979,In_261,In_1183);
nor U980 (N_980,In_69,In_356);
or U981 (N_981,In_1440,In_340);
nor U982 (N_982,In_252,In_566);
or U983 (N_983,In_1199,In_169);
nor U984 (N_984,In_578,In_1836);
or U985 (N_985,In_823,In_1226);
nor U986 (N_986,In_437,In_666);
nand U987 (N_987,In_1086,In_66);
nor U988 (N_988,In_603,In_1930);
nor U989 (N_989,In_1646,In_1754);
nand U990 (N_990,In_324,In_926);
or U991 (N_991,In_944,In_1620);
and U992 (N_992,In_499,In_1882);
and U993 (N_993,In_215,In_720);
nor U994 (N_994,In_959,In_1906);
nand U995 (N_995,In_1481,In_127);
or U996 (N_996,In_761,In_648);
or U997 (N_997,In_1188,In_742);
nor U998 (N_998,In_556,In_952);
and U999 (N_999,In_767,In_350);
and U1000 (N_1000,In_1768,In_890);
nor U1001 (N_1001,In_1825,In_476);
nor U1002 (N_1002,In_1269,In_1176);
nor U1003 (N_1003,In_1051,In_618);
and U1004 (N_1004,In_900,In_136);
nor U1005 (N_1005,In_889,In_553);
and U1006 (N_1006,In_846,In_986);
or U1007 (N_1007,In_1897,In_636);
or U1008 (N_1008,In_349,In_1736);
and U1009 (N_1009,In_134,In_246);
and U1010 (N_1010,In_1943,In_626);
or U1011 (N_1011,In_1154,In_1170);
nand U1012 (N_1012,In_721,In_1365);
and U1013 (N_1013,In_1714,In_137);
xor U1014 (N_1014,In_728,In_1670);
and U1015 (N_1015,In_190,In_522);
nor U1016 (N_1016,In_833,In_829);
nand U1017 (N_1017,In_1605,In_210);
xnor U1018 (N_1018,In_568,In_757);
nand U1019 (N_1019,In_1860,In_630);
or U1020 (N_1020,In_1795,In_1619);
or U1021 (N_1021,In_1200,In_1371);
and U1022 (N_1022,In_1488,In_1793);
xnor U1023 (N_1023,In_304,In_275);
or U1024 (N_1024,In_1018,In_86);
nor U1025 (N_1025,In_49,In_1749);
or U1026 (N_1026,In_1675,In_188);
and U1027 (N_1027,In_584,In_212);
or U1028 (N_1028,In_1447,In_560);
nand U1029 (N_1029,In_1718,In_1662);
or U1030 (N_1030,In_779,In_1710);
nor U1031 (N_1031,In_10,In_1523);
nand U1032 (N_1032,In_801,In_445);
nor U1033 (N_1033,In_189,In_564);
nor U1034 (N_1034,In_1883,In_1925);
and U1035 (N_1035,In_1975,In_1753);
nor U1036 (N_1036,In_1137,In_1974);
nand U1037 (N_1037,In_1483,In_1642);
nor U1038 (N_1038,In_1310,In_1017);
and U1039 (N_1039,In_1362,In_1322);
xnor U1040 (N_1040,In_621,In_1476);
and U1041 (N_1041,In_1182,In_547);
or U1042 (N_1042,In_1170,In_399);
nor U1043 (N_1043,In_185,In_817);
xor U1044 (N_1044,In_256,In_1932);
or U1045 (N_1045,In_1353,In_1195);
nor U1046 (N_1046,In_377,In_703);
nand U1047 (N_1047,In_1745,In_1794);
nand U1048 (N_1048,In_814,In_294);
or U1049 (N_1049,In_1686,In_1771);
nand U1050 (N_1050,In_818,In_68);
or U1051 (N_1051,In_1693,In_1648);
nor U1052 (N_1052,In_1786,In_1090);
or U1053 (N_1053,In_1056,In_252);
and U1054 (N_1054,In_1876,In_1797);
or U1055 (N_1055,In_394,In_318);
nor U1056 (N_1056,In_1824,In_1881);
and U1057 (N_1057,In_457,In_1183);
and U1058 (N_1058,In_1243,In_1186);
or U1059 (N_1059,In_1590,In_856);
or U1060 (N_1060,In_839,In_1867);
nand U1061 (N_1061,In_711,In_179);
or U1062 (N_1062,In_504,In_1387);
nor U1063 (N_1063,In_363,In_986);
and U1064 (N_1064,In_763,In_124);
nand U1065 (N_1065,In_1851,In_637);
nor U1066 (N_1066,In_356,In_1442);
nand U1067 (N_1067,In_229,In_1457);
and U1068 (N_1068,In_1783,In_786);
or U1069 (N_1069,In_334,In_317);
or U1070 (N_1070,In_810,In_113);
and U1071 (N_1071,In_1621,In_600);
and U1072 (N_1072,In_318,In_1691);
or U1073 (N_1073,In_444,In_732);
nand U1074 (N_1074,In_62,In_1517);
nand U1075 (N_1075,In_986,In_1643);
nor U1076 (N_1076,In_107,In_294);
xnor U1077 (N_1077,In_946,In_929);
nand U1078 (N_1078,In_383,In_1458);
and U1079 (N_1079,In_1471,In_1588);
or U1080 (N_1080,In_222,In_1160);
and U1081 (N_1081,In_1204,In_1848);
or U1082 (N_1082,In_388,In_361);
and U1083 (N_1083,In_483,In_1011);
and U1084 (N_1084,In_125,In_1755);
and U1085 (N_1085,In_1456,In_685);
nor U1086 (N_1086,In_1060,In_1388);
nor U1087 (N_1087,In_1843,In_160);
xnor U1088 (N_1088,In_704,In_888);
or U1089 (N_1089,In_1525,In_1615);
nand U1090 (N_1090,In_855,In_645);
nor U1091 (N_1091,In_380,In_1189);
or U1092 (N_1092,In_1607,In_370);
nand U1093 (N_1093,In_615,In_601);
and U1094 (N_1094,In_1498,In_1828);
xor U1095 (N_1095,In_102,In_1701);
nand U1096 (N_1096,In_135,In_1304);
xor U1097 (N_1097,In_249,In_61);
or U1098 (N_1098,In_247,In_639);
nand U1099 (N_1099,In_388,In_1150);
and U1100 (N_1100,In_85,In_657);
nand U1101 (N_1101,In_114,In_741);
nor U1102 (N_1102,In_295,In_493);
nand U1103 (N_1103,In_1706,In_1500);
or U1104 (N_1104,In_911,In_135);
nand U1105 (N_1105,In_792,In_600);
nand U1106 (N_1106,In_345,In_1953);
nor U1107 (N_1107,In_942,In_776);
nand U1108 (N_1108,In_125,In_1764);
or U1109 (N_1109,In_608,In_868);
xor U1110 (N_1110,In_1081,In_1790);
xnor U1111 (N_1111,In_131,In_1798);
and U1112 (N_1112,In_835,In_1350);
nor U1113 (N_1113,In_116,In_1006);
and U1114 (N_1114,In_1876,In_924);
or U1115 (N_1115,In_1379,In_496);
and U1116 (N_1116,In_896,In_1790);
or U1117 (N_1117,In_796,In_27);
nor U1118 (N_1118,In_16,In_95);
nand U1119 (N_1119,In_1755,In_1842);
or U1120 (N_1120,In_1918,In_655);
or U1121 (N_1121,In_1765,In_724);
and U1122 (N_1122,In_944,In_210);
and U1123 (N_1123,In_781,In_1962);
and U1124 (N_1124,In_918,In_1901);
or U1125 (N_1125,In_1405,In_1852);
nand U1126 (N_1126,In_1723,In_161);
nand U1127 (N_1127,In_1045,In_1209);
and U1128 (N_1128,In_1684,In_1017);
nand U1129 (N_1129,In_1240,In_1662);
and U1130 (N_1130,In_1528,In_315);
nand U1131 (N_1131,In_1310,In_1534);
and U1132 (N_1132,In_1616,In_1490);
xor U1133 (N_1133,In_1795,In_808);
nand U1134 (N_1134,In_1192,In_1684);
nand U1135 (N_1135,In_547,In_427);
or U1136 (N_1136,In_1916,In_649);
or U1137 (N_1137,In_1067,In_443);
or U1138 (N_1138,In_140,In_1777);
nor U1139 (N_1139,In_847,In_1681);
or U1140 (N_1140,In_1058,In_1745);
nor U1141 (N_1141,In_639,In_1347);
or U1142 (N_1142,In_738,In_219);
nand U1143 (N_1143,In_1655,In_1446);
nor U1144 (N_1144,In_1775,In_435);
nand U1145 (N_1145,In_1560,In_1791);
nand U1146 (N_1146,In_1449,In_1750);
nor U1147 (N_1147,In_1105,In_1682);
and U1148 (N_1148,In_778,In_113);
or U1149 (N_1149,In_649,In_974);
or U1150 (N_1150,In_990,In_714);
or U1151 (N_1151,In_611,In_423);
and U1152 (N_1152,In_733,In_1512);
nand U1153 (N_1153,In_1765,In_1588);
nor U1154 (N_1154,In_277,In_1644);
nand U1155 (N_1155,In_536,In_1388);
or U1156 (N_1156,In_13,In_702);
or U1157 (N_1157,In_430,In_1471);
or U1158 (N_1158,In_1499,In_1428);
and U1159 (N_1159,In_791,In_637);
or U1160 (N_1160,In_502,In_167);
or U1161 (N_1161,In_860,In_279);
xnor U1162 (N_1162,In_1257,In_302);
or U1163 (N_1163,In_411,In_629);
or U1164 (N_1164,In_184,In_1414);
nand U1165 (N_1165,In_1040,In_647);
nor U1166 (N_1166,In_141,In_1629);
nand U1167 (N_1167,In_1559,In_1971);
nand U1168 (N_1168,In_272,In_1854);
and U1169 (N_1169,In_530,In_698);
or U1170 (N_1170,In_383,In_1022);
nand U1171 (N_1171,In_1262,In_448);
nor U1172 (N_1172,In_573,In_56);
nor U1173 (N_1173,In_1520,In_591);
nor U1174 (N_1174,In_502,In_1883);
or U1175 (N_1175,In_764,In_554);
nor U1176 (N_1176,In_1808,In_39);
nor U1177 (N_1177,In_179,In_1502);
nor U1178 (N_1178,In_998,In_1131);
nand U1179 (N_1179,In_968,In_385);
or U1180 (N_1180,In_344,In_1005);
nor U1181 (N_1181,In_161,In_584);
and U1182 (N_1182,In_1608,In_1408);
nand U1183 (N_1183,In_1466,In_326);
xnor U1184 (N_1184,In_108,In_1604);
or U1185 (N_1185,In_574,In_194);
and U1186 (N_1186,In_35,In_294);
and U1187 (N_1187,In_202,In_1764);
nand U1188 (N_1188,In_1251,In_1829);
nor U1189 (N_1189,In_1453,In_1285);
and U1190 (N_1190,In_1830,In_212);
and U1191 (N_1191,In_1553,In_459);
nand U1192 (N_1192,In_1647,In_1386);
nor U1193 (N_1193,In_1039,In_952);
nor U1194 (N_1194,In_1073,In_1003);
nor U1195 (N_1195,In_1957,In_1250);
nor U1196 (N_1196,In_1894,In_962);
nor U1197 (N_1197,In_1357,In_632);
nand U1198 (N_1198,In_1570,In_1530);
nor U1199 (N_1199,In_800,In_1990);
or U1200 (N_1200,In_563,In_0);
or U1201 (N_1201,In_808,In_423);
nand U1202 (N_1202,In_1976,In_1103);
nor U1203 (N_1203,In_524,In_683);
nand U1204 (N_1204,In_756,In_1585);
nor U1205 (N_1205,In_936,In_1880);
nor U1206 (N_1206,In_1654,In_1747);
nand U1207 (N_1207,In_992,In_215);
or U1208 (N_1208,In_848,In_136);
xnor U1209 (N_1209,In_1966,In_1768);
xor U1210 (N_1210,In_685,In_1744);
nand U1211 (N_1211,In_1785,In_1404);
nand U1212 (N_1212,In_564,In_1961);
xor U1213 (N_1213,In_788,In_665);
nand U1214 (N_1214,In_141,In_1104);
xnor U1215 (N_1215,In_882,In_1196);
or U1216 (N_1216,In_617,In_1490);
nor U1217 (N_1217,In_998,In_1361);
or U1218 (N_1218,In_1669,In_504);
nor U1219 (N_1219,In_1749,In_1135);
or U1220 (N_1220,In_2,In_1169);
xor U1221 (N_1221,In_1399,In_117);
or U1222 (N_1222,In_615,In_1952);
nand U1223 (N_1223,In_1555,In_131);
nor U1224 (N_1224,In_1983,In_1303);
or U1225 (N_1225,In_400,In_1514);
nor U1226 (N_1226,In_375,In_1463);
or U1227 (N_1227,In_440,In_567);
nand U1228 (N_1228,In_1960,In_1273);
nand U1229 (N_1229,In_439,In_235);
nand U1230 (N_1230,In_592,In_1897);
nand U1231 (N_1231,In_1666,In_277);
nor U1232 (N_1232,In_387,In_930);
xor U1233 (N_1233,In_1752,In_1201);
nand U1234 (N_1234,In_1169,In_283);
or U1235 (N_1235,In_1107,In_576);
and U1236 (N_1236,In_568,In_1280);
or U1237 (N_1237,In_1330,In_1237);
nand U1238 (N_1238,In_30,In_1124);
nor U1239 (N_1239,In_1606,In_113);
nor U1240 (N_1240,In_847,In_1478);
nand U1241 (N_1241,In_1614,In_346);
and U1242 (N_1242,In_1824,In_1591);
or U1243 (N_1243,In_1037,In_1149);
or U1244 (N_1244,In_1380,In_357);
nand U1245 (N_1245,In_1459,In_1844);
or U1246 (N_1246,In_1713,In_1587);
nor U1247 (N_1247,In_1603,In_943);
nand U1248 (N_1248,In_711,In_1582);
nand U1249 (N_1249,In_1877,In_1392);
nand U1250 (N_1250,In_455,In_148);
or U1251 (N_1251,In_1440,In_462);
xor U1252 (N_1252,In_1097,In_1535);
nand U1253 (N_1253,In_1359,In_676);
nor U1254 (N_1254,In_487,In_182);
and U1255 (N_1255,In_1417,In_1485);
nor U1256 (N_1256,In_1769,In_1045);
nand U1257 (N_1257,In_1125,In_1328);
or U1258 (N_1258,In_1788,In_1475);
nor U1259 (N_1259,In_1200,In_1881);
and U1260 (N_1260,In_1557,In_958);
and U1261 (N_1261,In_1151,In_1311);
xor U1262 (N_1262,In_1227,In_739);
or U1263 (N_1263,In_1293,In_195);
xor U1264 (N_1264,In_703,In_1554);
and U1265 (N_1265,In_1095,In_426);
nor U1266 (N_1266,In_1797,In_1346);
and U1267 (N_1267,In_1712,In_650);
and U1268 (N_1268,In_1015,In_1978);
nor U1269 (N_1269,In_1449,In_265);
nor U1270 (N_1270,In_1866,In_1917);
nand U1271 (N_1271,In_701,In_32);
nand U1272 (N_1272,In_710,In_95);
nor U1273 (N_1273,In_1250,In_572);
and U1274 (N_1274,In_713,In_1726);
nor U1275 (N_1275,In_661,In_234);
nand U1276 (N_1276,In_1419,In_1969);
or U1277 (N_1277,In_1093,In_1724);
and U1278 (N_1278,In_1109,In_734);
xnor U1279 (N_1279,In_332,In_1689);
nand U1280 (N_1280,In_1315,In_1624);
xor U1281 (N_1281,In_403,In_427);
nand U1282 (N_1282,In_935,In_496);
nand U1283 (N_1283,In_189,In_1484);
and U1284 (N_1284,In_1566,In_1932);
or U1285 (N_1285,In_1006,In_1633);
nand U1286 (N_1286,In_1483,In_867);
or U1287 (N_1287,In_1338,In_868);
nand U1288 (N_1288,In_202,In_593);
nor U1289 (N_1289,In_680,In_125);
or U1290 (N_1290,In_320,In_1086);
nor U1291 (N_1291,In_138,In_1370);
nand U1292 (N_1292,In_343,In_394);
and U1293 (N_1293,In_920,In_1821);
nor U1294 (N_1294,In_1295,In_517);
nor U1295 (N_1295,In_1792,In_1450);
nor U1296 (N_1296,In_216,In_399);
xor U1297 (N_1297,In_1556,In_145);
and U1298 (N_1298,In_1037,In_1561);
nand U1299 (N_1299,In_599,In_1417);
or U1300 (N_1300,In_1645,In_1041);
or U1301 (N_1301,In_1866,In_1842);
nand U1302 (N_1302,In_894,In_107);
nand U1303 (N_1303,In_630,In_811);
nand U1304 (N_1304,In_1050,In_657);
and U1305 (N_1305,In_9,In_813);
and U1306 (N_1306,In_354,In_985);
xor U1307 (N_1307,In_562,In_1186);
nand U1308 (N_1308,In_1553,In_1238);
and U1309 (N_1309,In_166,In_216);
or U1310 (N_1310,In_1796,In_1632);
nor U1311 (N_1311,In_1887,In_614);
xnor U1312 (N_1312,In_1849,In_1375);
nand U1313 (N_1313,In_472,In_412);
and U1314 (N_1314,In_388,In_73);
and U1315 (N_1315,In_598,In_237);
or U1316 (N_1316,In_1864,In_704);
and U1317 (N_1317,In_141,In_396);
xnor U1318 (N_1318,In_421,In_1214);
nor U1319 (N_1319,In_1176,In_1797);
and U1320 (N_1320,In_457,In_500);
nor U1321 (N_1321,In_365,In_116);
nand U1322 (N_1322,In_716,In_1410);
or U1323 (N_1323,In_805,In_1870);
or U1324 (N_1324,In_1575,In_457);
and U1325 (N_1325,In_250,In_914);
nand U1326 (N_1326,In_255,In_974);
nor U1327 (N_1327,In_1313,In_522);
and U1328 (N_1328,In_1789,In_1101);
or U1329 (N_1329,In_1594,In_1288);
and U1330 (N_1330,In_1699,In_1890);
or U1331 (N_1331,In_595,In_577);
nand U1332 (N_1332,In_643,In_1792);
xor U1333 (N_1333,In_1539,In_240);
nand U1334 (N_1334,In_56,In_1464);
or U1335 (N_1335,In_176,In_1793);
and U1336 (N_1336,In_1324,In_1158);
or U1337 (N_1337,In_117,In_302);
nor U1338 (N_1338,In_1997,In_305);
nor U1339 (N_1339,In_826,In_500);
nand U1340 (N_1340,In_591,In_1866);
and U1341 (N_1341,In_39,In_1319);
and U1342 (N_1342,In_1228,In_773);
or U1343 (N_1343,In_867,In_1074);
or U1344 (N_1344,In_1512,In_737);
nor U1345 (N_1345,In_621,In_1754);
and U1346 (N_1346,In_1958,In_1530);
nand U1347 (N_1347,In_1276,In_1358);
nand U1348 (N_1348,In_1537,In_1010);
or U1349 (N_1349,In_617,In_1871);
or U1350 (N_1350,In_1537,In_1446);
nand U1351 (N_1351,In_743,In_1279);
nor U1352 (N_1352,In_1715,In_699);
nor U1353 (N_1353,In_1617,In_348);
or U1354 (N_1354,In_1144,In_1065);
and U1355 (N_1355,In_1447,In_1318);
and U1356 (N_1356,In_1515,In_761);
nand U1357 (N_1357,In_1541,In_729);
and U1358 (N_1358,In_745,In_1811);
or U1359 (N_1359,In_661,In_898);
or U1360 (N_1360,In_969,In_1030);
xnor U1361 (N_1361,In_645,In_1464);
nor U1362 (N_1362,In_1223,In_166);
nand U1363 (N_1363,In_353,In_529);
or U1364 (N_1364,In_1128,In_287);
and U1365 (N_1365,In_187,In_331);
nor U1366 (N_1366,In_1816,In_1598);
nand U1367 (N_1367,In_1244,In_1209);
or U1368 (N_1368,In_1181,In_1945);
or U1369 (N_1369,In_883,In_1785);
and U1370 (N_1370,In_541,In_1077);
xor U1371 (N_1371,In_1178,In_257);
nor U1372 (N_1372,In_1710,In_100);
nand U1373 (N_1373,In_1642,In_1872);
and U1374 (N_1374,In_900,In_925);
and U1375 (N_1375,In_976,In_324);
or U1376 (N_1376,In_112,In_553);
nor U1377 (N_1377,In_57,In_453);
xnor U1378 (N_1378,In_658,In_1601);
and U1379 (N_1379,In_1591,In_1779);
or U1380 (N_1380,In_1901,In_1221);
nor U1381 (N_1381,In_620,In_1924);
or U1382 (N_1382,In_530,In_1289);
nor U1383 (N_1383,In_1269,In_961);
xor U1384 (N_1384,In_929,In_1154);
or U1385 (N_1385,In_846,In_1224);
xor U1386 (N_1386,In_1233,In_238);
nor U1387 (N_1387,In_1820,In_253);
xnor U1388 (N_1388,In_112,In_1775);
and U1389 (N_1389,In_1469,In_1250);
nor U1390 (N_1390,In_1985,In_110);
or U1391 (N_1391,In_802,In_1379);
xnor U1392 (N_1392,In_1491,In_272);
or U1393 (N_1393,In_831,In_1011);
nor U1394 (N_1394,In_124,In_1167);
or U1395 (N_1395,In_1179,In_306);
nand U1396 (N_1396,In_1204,In_600);
nor U1397 (N_1397,In_158,In_1644);
xor U1398 (N_1398,In_1244,In_458);
nand U1399 (N_1399,In_801,In_797);
nand U1400 (N_1400,In_589,In_1059);
nor U1401 (N_1401,In_1663,In_360);
xor U1402 (N_1402,In_606,In_219);
or U1403 (N_1403,In_612,In_294);
nor U1404 (N_1404,In_63,In_1494);
and U1405 (N_1405,In_405,In_620);
nor U1406 (N_1406,In_723,In_1667);
nor U1407 (N_1407,In_1584,In_1948);
and U1408 (N_1408,In_201,In_277);
and U1409 (N_1409,In_486,In_238);
and U1410 (N_1410,In_132,In_271);
or U1411 (N_1411,In_100,In_909);
nand U1412 (N_1412,In_137,In_882);
nor U1413 (N_1413,In_181,In_536);
xor U1414 (N_1414,In_1093,In_448);
nor U1415 (N_1415,In_145,In_1509);
nor U1416 (N_1416,In_752,In_304);
and U1417 (N_1417,In_399,In_1295);
nand U1418 (N_1418,In_1924,In_1264);
and U1419 (N_1419,In_671,In_131);
xnor U1420 (N_1420,In_1457,In_896);
or U1421 (N_1421,In_315,In_455);
or U1422 (N_1422,In_1275,In_1215);
and U1423 (N_1423,In_394,In_1665);
nor U1424 (N_1424,In_607,In_1733);
nand U1425 (N_1425,In_1182,In_1191);
xnor U1426 (N_1426,In_1410,In_1918);
xor U1427 (N_1427,In_1158,In_657);
and U1428 (N_1428,In_834,In_1531);
nor U1429 (N_1429,In_1643,In_357);
and U1430 (N_1430,In_624,In_1189);
nand U1431 (N_1431,In_1996,In_1285);
nor U1432 (N_1432,In_1413,In_239);
nor U1433 (N_1433,In_979,In_1414);
xnor U1434 (N_1434,In_619,In_1602);
and U1435 (N_1435,In_1424,In_1182);
or U1436 (N_1436,In_1712,In_918);
or U1437 (N_1437,In_769,In_1463);
and U1438 (N_1438,In_1141,In_87);
nor U1439 (N_1439,In_1520,In_1910);
nand U1440 (N_1440,In_937,In_1862);
nor U1441 (N_1441,In_758,In_1148);
and U1442 (N_1442,In_448,In_140);
or U1443 (N_1443,In_12,In_1039);
nor U1444 (N_1444,In_869,In_44);
nand U1445 (N_1445,In_536,In_1526);
and U1446 (N_1446,In_1760,In_1615);
nand U1447 (N_1447,In_1553,In_502);
and U1448 (N_1448,In_623,In_41);
xnor U1449 (N_1449,In_1972,In_661);
nor U1450 (N_1450,In_854,In_259);
nor U1451 (N_1451,In_1671,In_304);
nor U1452 (N_1452,In_1895,In_1253);
nor U1453 (N_1453,In_1905,In_899);
nand U1454 (N_1454,In_188,In_757);
or U1455 (N_1455,In_1594,In_613);
and U1456 (N_1456,In_704,In_1276);
nor U1457 (N_1457,In_1173,In_837);
or U1458 (N_1458,In_1694,In_1279);
xor U1459 (N_1459,In_1333,In_1983);
or U1460 (N_1460,In_478,In_267);
nand U1461 (N_1461,In_1882,In_1484);
nor U1462 (N_1462,In_243,In_1363);
xor U1463 (N_1463,In_1469,In_120);
xnor U1464 (N_1464,In_1720,In_1547);
xor U1465 (N_1465,In_1280,In_469);
xor U1466 (N_1466,In_271,In_18);
nand U1467 (N_1467,In_71,In_958);
or U1468 (N_1468,In_252,In_856);
and U1469 (N_1469,In_1242,In_916);
nand U1470 (N_1470,In_1275,In_975);
nand U1471 (N_1471,In_531,In_127);
nand U1472 (N_1472,In_1048,In_1178);
xor U1473 (N_1473,In_1656,In_1734);
nor U1474 (N_1474,In_527,In_79);
and U1475 (N_1475,In_1656,In_506);
nand U1476 (N_1476,In_1865,In_432);
and U1477 (N_1477,In_184,In_1879);
xnor U1478 (N_1478,In_315,In_1781);
and U1479 (N_1479,In_399,In_1439);
or U1480 (N_1480,In_1367,In_676);
nor U1481 (N_1481,In_285,In_714);
nor U1482 (N_1482,In_575,In_1853);
nand U1483 (N_1483,In_315,In_1019);
nor U1484 (N_1484,In_309,In_1648);
or U1485 (N_1485,In_226,In_348);
xor U1486 (N_1486,In_548,In_1073);
or U1487 (N_1487,In_416,In_935);
and U1488 (N_1488,In_419,In_1932);
nand U1489 (N_1489,In_1,In_35);
xor U1490 (N_1490,In_1895,In_1722);
nand U1491 (N_1491,In_420,In_106);
or U1492 (N_1492,In_1025,In_728);
nor U1493 (N_1493,In_244,In_883);
nand U1494 (N_1494,In_268,In_109);
xor U1495 (N_1495,In_1718,In_214);
nor U1496 (N_1496,In_305,In_309);
nand U1497 (N_1497,In_1054,In_1559);
or U1498 (N_1498,In_1534,In_340);
nand U1499 (N_1499,In_491,In_1176);
nand U1500 (N_1500,In_520,In_39);
or U1501 (N_1501,In_81,In_1430);
or U1502 (N_1502,In_964,In_773);
xor U1503 (N_1503,In_491,In_178);
xor U1504 (N_1504,In_1070,In_1392);
or U1505 (N_1505,In_656,In_478);
nand U1506 (N_1506,In_536,In_1734);
or U1507 (N_1507,In_1547,In_1171);
and U1508 (N_1508,In_900,In_398);
or U1509 (N_1509,In_287,In_250);
nand U1510 (N_1510,In_1364,In_451);
and U1511 (N_1511,In_597,In_920);
and U1512 (N_1512,In_1671,In_881);
nand U1513 (N_1513,In_553,In_1824);
or U1514 (N_1514,In_1695,In_1162);
nor U1515 (N_1515,In_525,In_248);
xnor U1516 (N_1516,In_1930,In_665);
nor U1517 (N_1517,In_1612,In_84);
nor U1518 (N_1518,In_150,In_1354);
xnor U1519 (N_1519,In_402,In_332);
nand U1520 (N_1520,In_278,In_1412);
nor U1521 (N_1521,In_1305,In_1405);
nor U1522 (N_1522,In_1478,In_334);
and U1523 (N_1523,In_758,In_839);
nand U1524 (N_1524,In_436,In_718);
xnor U1525 (N_1525,In_438,In_1673);
nand U1526 (N_1526,In_537,In_1045);
or U1527 (N_1527,In_1486,In_1673);
nand U1528 (N_1528,In_533,In_1834);
xor U1529 (N_1529,In_904,In_1307);
or U1530 (N_1530,In_1087,In_1377);
or U1531 (N_1531,In_1433,In_182);
or U1532 (N_1532,In_1453,In_632);
and U1533 (N_1533,In_392,In_908);
nor U1534 (N_1534,In_734,In_85);
and U1535 (N_1535,In_892,In_730);
nand U1536 (N_1536,In_492,In_1015);
nand U1537 (N_1537,In_272,In_980);
and U1538 (N_1538,In_1079,In_258);
nor U1539 (N_1539,In_1760,In_1548);
and U1540 (N_1540,In_1733,In_1647);
nor U1541 (N_1541,In_1434,In_282);
nand U1542 (N_1542,In_1811,In_548);
nor U1543 (N_1543,In_1843,In_138);
or U1544 (N_1544,In_1535,In_313);
nand U1545 (N_1545,In_956,In_171);
xnor U1546 (N_1546,In_104,In_1236);
and U1547 (N_1547,In_1135,In_1241);
and U1548 (N_1548,In_147,In_55);
xnor U1549 (N_1549,In_1561,In_1199);
nor U1550 (N_1550,In_749,In_1649);
and U1551 (N_1551,In_1652,In_1118);
nor U1552 (N_1552,In_40,In_648);
and U1553 (N_1553,In_363,In_928);
or U1554 (N_1554,In_1574,In_1129);
nand U1555 (N_1555,In_1547,In_1411);
or U1556 (N_1556,In_1471,In_1380);
xor U1557 (N_1557,In_1188,In_760);
or U1558 (N_1558,In_1650,In_1150);
or U1559 (N_1559,In_1370,In_1485);
and U1560 (N_1560,In_1439,In_273);
and U1561 (N_1561,In_742,In_1647);
nand U1562 (N_1562,In_1914,In_761);
and U1563 (N_1563,In_1642,In_76);
nor U1564 (N_1564,In_1545,In_243);
and U1565 (N_1565,In_246,In_151);
xnor U1566 (N_1566,In_502,In_742);
or U1567 (N_1567,In_525,In_910);
xor U1568 (N_1568,In_1236,In_363);
or U1569 (N_1569,In_607,In_992);
nor U1570 (N_1570,In_961,In_236);
nand U1571 (N_1571,In_216,In_576);
or U1572 (N_1572,In_1374,In_1941);
nor U1573 (N_1573,In_1340,In_832);
and U1574 (N_1574,In_43,In_1549);
or U1575 (N_1575,In_1105,In_285);
nor U1576 (N_1576,In_1070,In_1318);
nor U1577 (N_1577,In_1419,In_1175);
or U1578 (N_1578,In_1897,In_1584);
xnor U1579 (N_1579,In_1340,In_1103);
xnor U1580 (N_1580,In_1821,In_1385);
nand U1581 (N_1581,In_550,In_120);
nor U1582 (N_1582,In_1910,In_868);
and U1583 (N_1583,In_120,In_1197);
or U1584 (N_1584,In_1691,In_1653);
or U1585 (N_1585,In_11,In_524);
nand U1586 (N_1586,In_872,In_805);
nor U1587 (N_1587,In_1909,In_603);
nor U1588 (N_1588,In_1590,In_1807);
nor U1589 (N_1589,In_1801,In_1133);
nor U1590 (N_1590,In_202,In_222);
or U1591 (N_1591,In_487,In_1525);
nand U1592 (N_1592,In_1650,In_1375);
and U1593 (N_1593,In_454,In_1872);
or U1594 (N_1594,In_1169,In_913);
nor U1595 (N_1595,In_1741,In_1583);
or U1596 (N_1596,In_263,In_24);
nand U1597 (N_1597,In_182,In_279);
nor U1598 (N_1598,In_1164,In_1240);
xor U1599 (N_1599,In_100,In_872);
or U1600 (N_1600,In_545,In_1749);
nor U1601 (N_1601,In_1273,In_1001);
or U1602 (N_1602,In_1339,In_1371);
nand U1603 (N_1603,In_708,In_973);
nor U1604 (N_1604,In_1963,In_1169);
or U1605 (N_1605,In_384,In_1004);
and U1606 (N_1606,In_1988,In_865);
and U1607 (N_1607,In_1695,In_1501);
nand U1608 (N_1608,In_735,In_1370);
xnor U1609 (N_1609,In_894,In_973);
xor U1610 (N_1610,In_910,In_1883);
or U1611 (N_1611,In_142,In_151);
nand U1612 (N_1612,In_1253,In_355);
or U1613 (N_1613,In_1513,In_410);
nor U1614 (N_1614,In_24,In_1584);
nor U1615 (N_1615,In_1264,In_1129);
or U1616 (N_1616,In_643,In_462);
nand U1617 (N_1617,In_784,In_214);
and U1618 (N_1618,In_1857,In_1028);
or U1619 (N_1619,In_1989,In_134);
or U1620 (N_1620,In_831,In_956);
and U1621 (N_1621,In_388,In_40);
or U1622 (N_1622,In_1886,In_463);
or U1623 (N_1623,In_49,In_1385);
and U1624 (N_1624,In_842,In_1016);
nand U1625 (N_1625,In_1225,In_104);
and U1626 (N_1626,In_1280,In_46);
or U1627 (N_1627,In_1193,In_223);
and U1628 (N_1628,In_1536,In_1173);
and U1629 (N_1629,In_1752,In_1123);
nor U1630 (N_1630,In_1547,In_1322);
or U1631 (N_1631,In_1025,In_396);
or U1632 (N_1632,In_255,In_1735);
or U1633 (N_1633,In_513,In_1049);
xnor U1634 (N_1634,In_308,In_745);
or U1635 (N_1635,In_1231,In_155);
nor U1636 (N_1636,In_1139,In_610);
or U1637 (N_1637,In_623,In_393);
nor U1638 (N_1638,In_840,In_1818);
nor U1639 (N_1639,In_605,In_1631);
or U1640 (N_1640,In_1619,In_1094);
nor U1641 (N_1641,In_676,In_930);
nor U1642 (N_1642,In_1783,In_271);
nand U1643 (N_1643,In_40,In_709);
xnor U1644 (N_1644,In_562,In_1520);
xnor U1645 (N_1645,In_1899,In_979);
nor U1646 (N_1646,In_314,In_1069);
and U1647 (N_1647,In_355,In_132);
and U1648 (N_1648,In_549,In_1200);
or U1649 (N_1649,In_226,In_279);
xor U1650 (N_1650,In_1540,In_16);
nor U1651 (N_1651,In_1607,In_846);
xnor U1652 (N_1652,In_1326,In_1075);
nor U1653 (N_1653,In_1183,In_1649);
and U1654 (N_1654,In_103,In_175);
nand U1655 (N_1655,In_323,In_457);
nor U1656 (N_1656,In_616,In_375);
nand U1657 (N_1657,In_1291,In_1069);
nor U1658 (N_1658,In_670,In_1691);
nand U1659 (N_1659,In_549,In_837);
xor U1660 (N_1660,In_1641,In_513);
or U1661 (N_1661,In_912,In_1292);
or U1662 (N_1662,In_815,In_54);
nand U1663 (N_1663,In_1566,In_519);
nand U1664 (N_1664,In_1456,In_1418);
and U1665 (N_1665,In_748,In_1224);
nand U1666 (N_1666,In_691,In_791);
xnor U1667 (N_1667,In_1408,In_739);
nand U1668 (N_1668,In_277,In_1546);
and U1669 (N_1669,In_1774,In_1917);
xnor U1670 (N_1670,In_659,In_339);
and U1671 (N_1671,In_1644,In_1715);
nand U1672 (N_1672,In_932,In_37);
or U1673 (N_1673,In_715,In_1867);
and U1674 (N_1674,In_302,In_160);
nor U1675 (N_1675,In_1485,In_1847);
and U1676 (N_1676,In_1009,In_1543);
nand U1677 (N_1677,In_483,In_1426);
or U1678 (N_1678,In_1678,In_1898);
xor U1679 (N_1679,In_1323,In_1895);
nor U1680 (N_1680,In_145,In_1487);
or U1681 (N_1681,In_726,In_141);
or U1682 (N_1682,In_1261,In_303);
and U1683 (N_1683,In_1444,In_1736);
nor U1684 (N_1684,In_1011,In_254);
or U1685 (N_1685,In_1797,In_1949);
nor U1686 (N_1686,In_1852,In_843);
nand U1687 (N_1687,In_24,In_652);
nand U1688 (N_1688,In_1433,In_675);
or U1689 (N_1689,In_1924,In_589);
nor U1690 (N_1690,In_1942,In_1074);
or U1691 (N_1691,In_404,In_1542);
nand U1692 (N_1692,In_315,In_409);
nand U1693 (N_1693,In_1058,In_673);
and U1694 (N_1694,In_17,In_876);
nand U1695 (N_1695,In_105,In_1737);
nand U1696 (N_1696,In_90,In_1053);
and U1697 (N_1697,In_1516,In_306);
nand U1698 (N_1698,In_1805,In_503);
nor U1699 (N_1699,In_82,In_994);
nor U1700 (N_1700,In_1465,In_1926);
and U1701 (N_1701,In_5,In_1231);
and U1702 (N_1702,In_1790,In_808);
or U1703 (N_1703,In_364,In_181);
and U1704 (N_1704,In_876,In_1781);
nor U1705 (N_1705,In_809,In_499);
and U1706 (N_1706,In_537,In_1694);
or U1707 (N_1707,In_392,In_240);
nor U1708 (N_1708,In_125,In_1870);
and U1709 (N_1709,In_1564,In_1660);
nand U1710 (N_1710,In_183,In_1189);
or U1711 (N_1711,In_763,In_1920);
nand U1712 (N_1712,In_1279,In_1035);
nor U1713 (N_1713,In_1542,In_403);
or U1714 (N_1714,In_1865,In_312);
xnor U1715 (N_1715,In_1679,In_613);
nor U1716 (N_1716,In_617,In_369);
and U1717 (N_1717,In_342,In_1530);
nor U1718 (N_1718,In_1396,In_935);
nand U1719 (N_1719,In_1562,In_891);
nand U1720 (N_1720,In_296,In_845);
and U1721 (N_1721,In_1774,In_1231);
or U1722 (N_1722,In_1680,In_1638);
nand U1723 (N_1723,In_905,In_852);
or U1724 (N_1724,In_1847,In_638);
nor U1725 (N_1725,In_142,In_1720);
nor U1726 (N_1726,In_945,In_1140);
and U1727 (N_1727,In_299,In_596);
or U1728 (N_1728,In_1724,In_1023);
nand U1729 (N_1729,In_1368,In_1379);
nor U1730 (N_1730,In_414,In_1562);
or U1731 (N_1731,In_691,In_425);
nand U1732 (N_1732,In_1174,In_1905);
nand U1733 (N_1733,In_509,In_325);
and U1734 (N_1734,In_1751,In_273);
nor U1735 (N_1735,In_30,In_1617);
xor U1736 (N_1736,In_494,In_368);
xnor U1737 (N_1737,In_1574,In_202);
nor U1738 (N_1738,In_1506,In_898);
nand U1739 (N_1739,In_560,In_1199);
or U1740 (N_1740,In_512,In_1161);
and U1741 (N_1741,In_994,In_1393);
or U1742 (N_1742,In_1874,In_1229);
xnor U1743 (N_1743,In_435,In_768);
or U1744 (N_1744,In_1853,In_1273);
and U1745 (N_1745,In_243,In_858);
nand U1746 (N_1746,In_258,In_626);
nand U1747 (N_1747,In_1305,In_473);
or U1748 (N_1748,In_1515,In_1886);
xnor U1749 (N_1749,In_12,In_1757);
nand U1750 (N_1750,In_735,In_1727);
or U1751 (N_1751,In_438,In_1108);
or U1752 (N_1752,In_1885,In_312);
nor U1753 (N_1753,In_201,In_17);
xor U1754 (N_1754,In_487,In_414);
nor U1755 (N_1755,In_1597,In_1091);
nand U1756 (N_1756,In_1499,In_375);
nand U1757 (N_1757,In_166,In_463);
and U1758 (N_1758,In_1463,In_1479);
or U1759 (N_1759,In_563,In_914);
xor U1760 (N_1760,In_1272,In_1713);
and U1761 (N_1761,In_1155,In_311);
and U1762 (N_1762,In_1901,In_1076);
nor U1763 (N_1763,In_929,In_542);
nor U1764 (N_1764,In_1742,In_1139);
or U1765 (N_1765,In_1207,In_1002);
and U1766 (N_1766,In_1979,In_1849);
nand U1767 (N_1767,In_1886,In_491);
nand U1768 (N_1768,In_1079,In_351);
nor U1769 (N_1769,In_1686,In_210);
or U1770 (N_1770,In_1147,In_334);
nand U1771 (N_1771,In_1726,In_407);
or U1772 (N_1772,In_593,In_1864);
nand U1773 (N_1773,In_971,In_1034);
and U1774 (N_1774,In_914,In_202);
nor U1775 (N_1775,In_397,In_175);
or U1776 (N_1776,In_435,In_1976);
and U1777 (N_1777,In_1589,In_848);
or U1778 (N_1778,In_1059,In_176);
nand U1779 (N_1779,In_340,In_1699);
and U1780 (N_1780,In_639,In_92);
nand U1781 (N_1781,In_128,In_1493);
xor U1782 (N_1782,In_1330,In_1251);
and U1783 (N_1783,In_1825,In_221);
nor U1784 (N_1784,In_1643,In_1271);
nand U1785 (N_1785,In_1064,In_442);
nand U1786 (N_1786,In_632,In_1171);
or U1787 (N_1787,In_1246,In_582);
and U1788 (N_1788,In_1821,In_1459);
and U1789 (N_1789,In_1878,In_472);
nor U1790 (N_1790,In_1678,In_1653);
or U1791 (N_1791,In_1714,In_1493);
and U1792 (N_1792,In_691,In_396);
nand U1793 (N_1793,In_1715,In_1651);
nand U1794 (N_1794,In_97,In_1559);
and U1795 (N_1795,In_1061,In_1358);
nor U1796 (N_1796,In_874,In_626);
nor U1797 (N_1797,In_1210,In_338);
nand U1798 (N_1798,In_729,In_1931);
or U1799 (N_1799,In_1062,In_877);
and U1800 (N_1800,In_391,In_953);
and U1801 (N_1801,In_1590,In_1583);
nand U1802 (N_1802,In_1869,In_1806);
or U1803 (N_1803,In_681,In_1096);
nand U1804 (N_1804,In_1442,In_182);
nor U1805 (N_1805,In_107,In_630);
or U1806 (N_1806,In_1507,In_688);
or U1807 (N_1807,In_1511,In_1924);
nand U1808 (N_1808,In_714,In_1003);
or U1809 (N_1809,In_796,In_1647);
or U1810 (N_1810,In_1650,In_1157);
nand U1811 (N_1811,In_1771,In_974);
nor U1812 (N_1812,In_1363,In_1987);
or U1813 (N_1813,In_89,In_862);
nand U1814 (N_1814,In_589,In_1087);
nand U1815 (N_1815,In_1214,In_175);
or U1816 (N_1816,In_578,In_1598);
or U1817 (N_1817,In_1603,In_1071);
and U1818 (N_1818,In_80,In_984);
nor U1819 (N_1819,In_853,In_303);
nor U1820 (N_1820,In_1630,In_1459);
nand U1821 (N_1821,In_1489,In_1146);
and U1822 (N_1822,In_154,In_1618);
nand U1823 (N_1823,In_427,In_1168);
nor U1824 (N_1824,In_980,In_1311);
nand U1825 (N_1825,In_1972,In_1725);
xnor U1826 (N_1826,In_350,In_975);
nor U1827 (N_1827,In_1143,In_405);
and U1828 (N_1828,In_1349,In_748);
nand U1829 (N_1829,In_565,In_821);
or U1830 (N_1830,In_1277,In_99);
nor U1831 (N_1831,In_134,In_458);
or U1832 (N_1832,In_526,In_1658);
and U1833 (N_1833,In_599,In_1716);
or U1834 (N_1834,In_10,In_1207);
nand U1835 (N_1835,In_456,In_1105);
or U1836 (N_1836,In_10,In_181);
nor U1837 (N_1837,In_383,In_315);
and U1838 (N_1838,In_1299,In_1696);
and U1839 (N_1839,In_527,In_927);
and U1840 (N_1840,In_869,In_1374);
nor U1841 (N_1841,In_408,In_1384);
or U1842 (N_1842,In_1251,In_1123);
or U1843 (N_1843,In_691,In_304);
nand U1844 (N_1844,In_1076,In_1669);
xnor U1845 (N_1845,In_515,In_1234);
or U1846 (N_1846,In_1391,In_1785);
nor U1847 (N_1847,In_1394,In_536);
and U1848 (N_1848,In_377,In_1480);
nand U1849 (N_1849,In_479,In_1340);
xnor U1850 (N_1850,In_248,In_878);
or U1851 (N_1851,In_829,In_1148);
and U1852 (N_1852,In_724,In_128);
nand U1853 (N_1853,In_1220,In_1501);
or U1854 (N_1854,In_1137,In_645);
or U1855 (N_1855,In_858,In_1719);
or U1856 (N_1856,In_118,In_568);
or U1857 (N_1857,In_325,In_1874);
and U1858 (N_1858,In_484,In_203);
and U1859 (N_1859,In_342,In_1404);
nor U1860 (N_1860,In_483,In_930);
xnor U1861 (N_1861,In_1975,In_449);
and U1862 (N_1862,In_1891,In_1812);
or U1863 (N_1863,In_1118,In_1245);
nand U1864 (N_1864,In_873,In_692);
or U1865 (N_1865,In_1714,In_1730);
or U1866 (N_1866,In_663,In_1306);
nor U1867 (N_1867,In_1897,In_1135);
nand U1868 (N_1868,In_1718,In_112);
nor U1869 (N_1869,In_1998,In_1902);
or U1870 (N_1870,In_334,In_1283);
or U1871 (N_1871,In_564,In_1101);
and U1872 (N_1872,In_1056,In_1809);
nor U1873 (N_1873,In_1084,In_787);
or U1874 (N_1874,In_1103,In_822);
nor U1875 (N_1875,In_824,In_247);
or U1876 (N_1876,In_440,In_727);
and U1877 (N_1877,In_23,In_492);
or U1878 (N_1878,In_595,In_394);
and U1879 (N_1879,In_1951,In_1838);
nand U1880 (N_1880,In_912,In_537);
nand U1881 (N_1881,In_810,In_1440);
and U1882 (N_1882,In_1386,In_809);
nor U1883 (N_1883,In_1281,In_1693);
and U1884 (N_1884,In_584,In_457);
nor U1885 (N_1885,In_229,In_1435);
or U1886 (N_1886,In_1627,In_1823);
nor U1887 (N_1887,In_1371,In_733);
and U1888 (N_1888,In_766,In_1396);
xor U1889 (N_1889,In_490,In_921);
nor U1890 (N_1890,In_1287,In_1926);
nand U1891 (N_1891,In_1084,In_1457);
or U1892 (N_1892,In_99,In_1358);
nor U1893 (N_1893,In_1880,In_798);
or U1894 (N_1894,In_1215,In_1620);
nand U1895 (N_1895,In_1889,In_1039);
nand U1896 (N_1896,In_1221,In_1678);
nor U1897 (N_1897,In_1462,In_486);
nor U1898 (N_1898,In_839,In_789);
or U1899 (N_1899,In_281,In_1560);
or U1900 (N_1900,In_498,In_1110);
nand U1901 (N_1901,In_538,In_1223);
xor U1902 (N_1902,In_1909,In_7);
nand U1903 (N_1903,In_1348,In_163);
xor U1904 (N_1904,In_41,In_1465);
nor U1905 (N_1905,In_1715,In_118);
nor U1906 (N_1906,In_1823,In_981);
nand U1907 (N_1907,In_682,In_976);
xor U1908 (N_1908,In_23,In_510);
xnor U1909 (N_1909,In_1461,In_517);
or U1910 (N_1910,In_715,In_1367);
or U1911 (N_1911,In_629,In_603);
xor U1912 (N_1912,In_1266,In_1305);
and U1913 (N_1913,In_60,In_259);
or U1914 (N_1914,In_957,In_1948);
or U1915 (N_1915,In_785,In_1065);
nor U1916 (N_1916,In_1512,In_1671);
nand U1917 (N_1917,In_1341,In_327);
nor U1918 (N_1918,In_1840,In_110);
nor U1919 (N_1919,In_1220,In_1116);
or U1920 (N_1920,In_552,In_1244);
xor U1921 (N_1921,In_155,In_488);
nand U1922 (N_1922,In_703,In_312);
and U1923 (N_1923,In_1212,In_681);
and U1924 (N_1924,In_1829,In_1741);
and U1925 (N_1925,In_1452,In_327);
nor U1926 (N_1926,In_1608,In_994);
or U1927 (N_1927,In_1717,In_1404);
nand U1928 (N_1928,In_1976,In_1315);
nand U1929 (N_1929,In_1443,In_1681);
xor U1930 (N_1930,In_420,In_256);
nand U1931 (N_1931,In_1354,In_1273);
and U1932 (N_1932,In_1451,In_182);
and U1933 (N_1933,In_1464,In_1604);
xor U1934 (N_1934,In_1675,In_1780);
or U1935 (N_1935,In_1641,In_162);
nand U1936 (N_1936,In_1129,In_885);
and U1937 (N_1937,In_1404,In_331);
nor U1938 (N_1938,In_1168,In_968);
nor U1939 (N_1939,In_42,In_469);
or U1940 (N_1940,In_902,In_901);
nand U1941 (N_1941,In_413,In_246);
nor U1942 (N_1942,In_857,In_616);
or U1943 (N_1943,In_1529,In_1712);
nand U1944 (N_1944,In_1834,In_1621);
and U1945 (N_1945,In_173,In_330);
nor U1946 (N_1946,In_266,In_752);
nand U1947 (N_1947,In_1728,In_150);
or U1948 (N_1948,In_1334,In_1016);
or U1949 (N_1949,In_229,In_1285);
nand U1950 (N_1950,In_788,In_948);
nor U1951 (N_1951,In_752,In_1852);
nor U1952 (N_1952,In_1406,In_1);
or U1953 (N_1953,In_926,In_898);
or U1954 (N_1954,In_670,In_141);
xnor U1955 (N_1955,In_421,In_420);
nand U1956 (N_1956,In_377,In_950);
nand U1957 (N_1957,In_186,In_1674);
nand U1958 (N_1958,In_1371,In_1820);
nor U1959 (N_1959,In_1973,In_1171);
nand U1960 (N_1960,In_1805,In_235);
nand U1961 (N_1961,In_1652,In_528);
nor U1962 (N_1962,In_1891,In_533);
and U1963 (N_1963,In_1652,In_1937);
nand U1964 (N_1964,In_1616,In_478);
nor U1965 (N_1965,In_473,In_315);
nor U1966 (N_1966,In_964,In_20);
nor U1967 (N_1967,In_519,In_1400);
or U1968 (N_1968,In_1825,In_985);
and U1969 (N_1969,In_639,In_1205);
xnor U1970 (N_1970,In_1404,In_81);
nor U1971 (N_1971,In_1072,In_367);
nand U1972 (N_1972,In_406,In_1952);
nand U1973 (N_1973,In_1925,In_1019);
nand U1974 (N_1974,In_401,In_1283);
nand U1975 (N_1975,In_509,In_482);
nand U1976 (N_1976,In_1989,In_409);
and U1977 (N_1977,In_619,In_312);
nor U1978 (N_1978,In_1989,In_924);
and U1979 (N_1979,In_1097,In_1624);
nand U1980 (N_1980,In_1719,In_1661);
nor U1981 (N_1981,In_21,In_1138);
and U1982 (N_1982,In_871,In_610);
nor U1983 (N_1983,In_1150,In_188);
nand U1984 (N_1984,In_609,In_1772);
or U1985 (N_1985,In_1721,In_607);
nand U1986 (N_1986,In_1539,In_988);
nand U1987 (N_1987,In_905,In_1146);
nor U1988 (N_1988,In_1696,In_1720);
nand U1989 (N_1989,In_1379,In_1607);
xor U1990 (N_1990,In_1194,In_1042);
or U1991 (N_1991,In_71,In_938);
nand U1992 (N_1992,In_306,In_686);
nor U1993 (N_1993,In_37,In_1132);
or U1994 (N_1994,In_1650,In_195);
xnor U1995 (N_1995,In_1638,In_1232);
nor U1996 (N_1996,In_490,In_410);
and U1997 (N_1997,In_1251,In_1443);
nand U1998 (N_1998,In_1552,In_1187);
nor U1999 (N_1999,In_1253,In_1561);
or U2000 (N_2000,N_1970,N_671);
xnor U2001 (N_2001,N_1798,N_320);
nor U2002 (N_2002,N_1492,N_697);
nor U2003 (N_2003,N_1513,N_1483);
nand U2004 (N_2004,N_741,N_1831);
nor U2005 (N_2005,N_1774,N_102);
nor U2006 (N_2006,N_1652,N_1853);
nor U2007 (N_2007,N_1539,N_263);
nand U2008 (N_2008,N_986,N_381);
nor U2009 (N_2009,N_719,N_1886);
and U2010 (N_2010,N_894,N_258);
or U2011 (N_2011,N_1478,N_1);
xnor U2012 (N_2012,N_1087,N_1382);
or U2013 (N_2013,N_662,N_1915);
nor U2014 (N_2014,N_1583,N_397);
and U2015 (N_2015,N_1769,N_1272);
or U2016 (N_2016,N_956,N_871);
and U2017 (N_2017,N_490,N_253);
nor U2018 (N_2018,N_1653,N_961);
nor U2019 (N_2019,N_836,N_1895);
nor U2020 (N_2020,N_541,N_335);
xor U2021 (N_2021,N_1878,N_647);
nand U2022 (N_2022,N_302,N_1207);
and U2023 (N_2023,N_740,N_1787);
and U2024 (N_2024,N_1059,N_181);
or U2025 (N_2025,N_771,N_805);
and U2026 (N_2026,N_944,N_699);
nand U2027 (N_2027,N_1258,N_1727);
and U2028 (N_2028,N_1912,N_999);
and U2029 (N_2029,N_1824,N_724);
nor U2030 (N_2030,N_638,N_1393);
nor U2031 (N_2031,N_1942,N_1362);
nor U2032 (N_2032,N_1342,N_1778);
or U2033 (N_2033,N_868,N_1014);
and U2034 (N_2034,N_1407,N_1902);
and U2035 (N_2035,N_779,N_704);
nand U2036 (N_2036,N_1782,N_1255);
and U2037 (N_2037,N_1189,N_369);
xor U2038 (N_2038,N_1366,N_218);
nand U2039 (N_2039,N_217,N_818);
or U2040 (N_2040,N_1877,N_631);
or U2041 (N_2041,N_529,N_1808);
and U2042 (N_2042,N_664,N_1031);
or U2043 (N_2043,N_1452,N_1855);
nor U2044 (N_2044,N_861,N_295);
or U2045 (N_2045,N_633,N_1399);
and U2046 (N_2046,N_445,N_355);
nor U2047 (N_2047,N_920,N_1385);
nand U2048 (N_2048,N_1094,N_794);
nor U2049 (N_2049,N_789,N_1328);
and U2050 (N_2050,N_1771,N_1038);
nand U2051 (N_2051,N_185,N_336);
xnor U2052 (N_2052,N_1370,N_333);
or U2053 (N_2053,N_1130,N_389);
nor U2054 (N_2054,N_402,N_860);
xnor U2055 (N_2055,N_799,N_1923);
or U2056 (N_2056,N_1047,N_547);
nand U2057 (N_2057,N_509,N_500);
nor U2058 (N_2058,N_700,N_757);
nor U2059 (N_2059,N_776,N_1078);
nor U2060 (N_2060,N_1100,N_1269);
or U2061 (N_2061,N_1657,N_1933);
and U2062 (N_2062,N_1516,N_1065);
or U2063 (N_2063,N_682,N_1694);
nor U2064 (N_2064,N_13,N_446);
and U2065 (N_2065,N_1643,N_1437);
xor U2066 (N_2066,N_1298,N_208);
nor U2067 (N_2067,N_843,N_1637);
nand U2068 (N_2068,N_1137,N_658);
nand U2069 (N_2069,N_508,N_167);
and U2070 (N_2070,N_562,N_374);
nor U2071 (N_2071,N_331,N_1281);
or U2072 (N_2072,N_934,N_450);
nand U2073 (N_2073,N_1879,N_505);
or U2074 (N_2074,N_617,N_1979);
xor U2075 (N_2075,N_9,N_1511);
and U2076 (N_2076,N_54,N_1268);
nor U2077 (N_2077,N_1115,N_750);
nand U2078 (N_2078,N_1347,N_1501);
or U2079 (N_2079,N_813,N_1585);
nand U2080 (N_2080,N_216,N_1360);
or U2081 (N_2081,N_322,N_1019);
and U2082 (N_2082,N_1406,N_241);
and U2083 (N_2083,N_274,N_1558);
nand U2084 (N_2084,N_150,N_1940);
and U2085 (N_2085,N_1498,N_201);
or U2086 (N_2086,N_1614,N_1791);
and U2087 (N_2087,N_619,N_1166);
nor U2088 (N_2088,N_1678,N_1935);
nand U2089 (N_2089,N_391,N_1252);
nand U2090 (N_2090,N_316,N_162);
and U2091 (N_2091,N_175,N_679);
nand U2092 (N_2092,N_823,N_1487);
nor U2093 (N_2093,N_1634,N_556);
and U2094 (N_2094,N_1043,N_339);
and U2095 (N_2095,N_769,N_1075);
and U2096 (N_2096,N_387,N_904);
or U2097 (N_2097,N_1423,N_1571);
nor U2098 (N_2098,N_869,N_748);
xnor U2099 (N_2099,N_808,N_730);
and U2100 (N_2100,N_1962,N_1985);
and U2101 (N_2101,N_20,N_1835);
and U2102 (N_2102,N_1891,N_1419);
nor U2103 (N_2103,N_686,N_407);
or U2104 (N_2104,N_1421,N_1842);
xor U2105 (N_2105,N_73,N_580);
and U2106 (N_2106,N_801,N_34);
or U2107 (N_2107,N_1832,N_978);
nand U2108 (N_2108,N_1686,N_1106);
and U2109 (N_2109,N_453,N_756);
nor U2110 (N_2110,N_845,N_1804);
and U2111 (N_2111,N_1174,N_648);
nand U2112 (N_2112,N_635,N_802);
nor U2113 (N_2113,N_1265,N_1864);
nand U2114 (N_2114,N_585,N_370);
nor U2115 (N_2115,N_486,N_503);
xor U2116 (N_2116,N_388,N_1064);
or U2117 (N_2117,N_1379,N_36);
and U2118 (N_2118,N_1856,N_1779);
nor U2119 (N_2119,N_554,N_202);
and U2120 (N_2120,N_1958,N_1651);
or U2121 (N_2121,N_1742,N_1756);
nand U2122 (N_2122,N_1537,N_1629);
or U2123 (N_2123,N_672,N_159);
xnor U2124 (N_2124,N_520,N_222);
nand U2125 (N_2125,N_1044,N_713);
and U2126 (N_2126,N_1147,N_1807);
nand U2127 (N_2127,N_390,N_565);
nor U2128 (N_2128,N_607,N_1336);
nor U2129 (N_2129,N_401,N_543);
nand U2130 (N_2130,N_1949,N_1275);
nand U2131 (N_2131,N_1981,N_305);
and U2132 (N_2132,N_1202,N_523);
nand U2133 (N_2133,N_936,N_219);
nor U2134 (N_2134,N_1928,N_1077);
nand U2135 (N_2135,N_15,N_441);
xnor U2136 (N_2136,N_363,N_1323);
xor U2137 (N_2137,N_1232,N_1697);
or U2138 (N_2138,N_21,N_172);
nand U2139 (N_2139,N_1613,N_259);
nand U2140 (N_2140,N_179,N_1600);
nor U2141 (N_2141,N_1718,N_1440);
or U2142 (N_2142,N_791,N_1861);
and U2143 (N_2143,N_513,N_1123);
and U2144 (N_2144,N_1103,N_328);
or U2145 (N_2145,N_685,N_1310);
nand U2146 (N_2146,N_761,N_1001);
and U2147 (N_2147,N_116,N_449);
xor U2148 (N_2148,N_1209,N_1688);
or U2149 (N_2149,N_883,N_1527);
nor U2150 (N_2150,N_459,N_1308);
or U2151 (N_2151,N_1294,N_1518);
and U2152 (N_2152,N_35,N_1659);
nand U2153 (N_2153,N_1248,N_516);
and U2154 (N_2154,N_1346,N_1811);
or U2155 (N_2155,N_1568,N_136);
nand U2156 (N_2156,N_127,N_693);
xor U2157 (N_2157,N_429,N_260);
or U2158 (N_2158,N_135,N_729);
and U2159 (N_2159,N_651,N_1520);
nor U2160 (N_2160,N_885,N_551);
or U2161 (N_2161,N_1226,N_718);
or U2162 (N_2162,N_1561,N_1021);
nor U2163 (N_2163,N_767,N_1000);
xnor U2164 (N_2164,N_1907,N_963);
nor U2165 (N_2165,N_315,N_366);
nor U2166 (N_2166,N_1675,N_1416);
xnor U2167 (N_2167,N_1656,N_660);
xnor U2168 (N_2168,N_224,N_1556);
or U2169 (N_2169,N_0,N_1219);
or U2170 (N_2170,N_1996,N_1412);
nand U2171 (N_2171,N_1816,N_683);
nand U2172 (N_2172,N_68,N_134);
nor U2173 (N_2173,N_1277,N_1957);
nand U2174 (N_2174,N_1716,N_1300);
nor U2175 (N_2175,N_471,N_566);
and U2176 (N_2176,N_1056,N_1489);
and U2177 (N_2177,N_27,N_1647);
nor U2178 (N_2178,N_1626,N_692);
xnor U2179 (N_2179,N_884,N_1352);
nor U2180 (N_2180,N_210,N_787);
nor U2181 (N_2181,N_810,N_1107);
or U2182 (N_2182,N_1480,N_117);
nand U2183 (N_2183,N_1309,N_456);
nand U2184 (N_2184,N_1707,N_178);
or U2185 (N_2185,N_866,N_1794);
or U2186 (N_2186,N_1839,N_1569);
and U2187 (N_2187,N_182,N_1708);
nor U2188 (N_2188,N_723,N_1488);
nor U2189 (N_2189,N_442,N_993);
nand U2190 (N_2190,N_480,N_273);
xnor U2191 (N_2191,N_1129,N_564);
and U2192 (N_2192,N_1591,N_952);
nand U2193 (N_2193,N_168,N_1610);
nand U2194 (N_2194,N_1617,N_6);
nor U2195 (N_2195,N_1753,N_928);
nand U2196 (N_2196,N_408,N_1757);
or U2197 (N_2197,N_561,N_935);
xnor U2198 (N_2198,N_1010,N_838);
nor U2199 (N_2199,N_979,N_354);
and U2200 (N_2200,N_1737,N_673);
nor U2201 (N_2201,N_254,N_1947);
and U2202 (N_2202,N_737,N_1011);
nor U2203 (N_2203,N_527,N_1818);
and U2204 (N_2204,N_1354,N_1540);
and U2205 (N_2205,N_1292,N_983);
nor U2206 (N_2206,N_57,N_1074);
and U2207 (N_2207,N_1994,N_1897);
or U2208 (N_2208,N_745,N_37);
nand U2209 (N_2209,N_1266,N_312);
nand U2210 (N_2210,N_307,N_1376);
nand U2211 (N_2211,N_634,N_833);
and U2212 (N_2212,N_1836,N_1155);
and U2213 (N_2213,N_1584,N_1847);
and U2214 (N_2214,N_1948,N_92);
and U2215 (N_2215,N_1420,N_1433);
xor U2216 (N_2216,N_623,N_1734);
or U2217 (N_2217,N_998,N_1852);
or U2218 (N_2218,N_847,N_1747);
nand U2219 (N_2219,N_66,N_444);
or U2220 (N_2220,N_461,N_1187);
or U2221 (N_2221,N_1208,N_1592);
or U2222 (N_2222,N_969,N_1894);
nor U2223 (N_2223,N_828,N_874);
nand U2224 (N_2224,N_1857,N_1534);
and U2225 (N_2225,N_398,N_1544);
nand U2226 (N_2226,N_613,N_359);
and U2227 (N_2227,N_494,N_3);
and U2228 (N_2228,N_1595,N_1099);
xor U2229 (N_2229,N_716,N_394);
or U2230 (N_2230,N_596,N_760);
nand U2231 (N_2231,N_755,N_863);
nand U2232 (N_2232,N_925,N_984);
and U2233 (N_2233,N_625,N_1033);
nor U2234 (N_2234,N_1998,N_1112);
or U2235 (N_2235,N_985,N_849);
or U2236 (N_2236,N_688,N_1820);
and U2237 (N_2237,N_876,N_109);
nor U2238 (N_2238,N_1601,N_1350);
nand U2239 (N_2239,N_824,N_668);
nand U2240 (N_2240,N_75,N_327);
and U2241 (N_2241,N_226,N_1497);
nand U2242 (N_2242,N_1163,N_110);
nor U2243 (N_2243,N_129,N_85);
or U2244 (N_2244,N_678,N_393);
nand U2245 (N_2245,N_1706,N_180);
and U2246 (N_2246,N_1215,N_1250);
nand U2247 (N_2247,N_1648,N_610);
and U2248 (N_2248,N_1542,N_1562);
nand U2249 (N_2249,N_1506,N_722);
nand U2250 (N_2250,N_283,N_1224);
xnor U2251 (N_2251,N_157,N_448);
nor U2252 (N_2252,N_161,N_1759);
nor U2253 (N_2253,N_1809,N_186);
nor U2254 (N_2254,N_1453,N_152);
nor U2255 (N_2255,N_267,N_1263);
and U2256 (N_2256,N_1934,N_144);
nand U2257 (N_2257,N_1826,N_415);
xnor U2258 (N_2258,N_1335,N_131);
or U2259 (N_2259,N_962,N_1479);
nor U2260 (N_2260,N_783,N_280);
or U2261 (N_2261,N_1784,N_870);
or U2262 (N_2262,N_1810,N_227);
nand U2263 (N_2263,N_1216,N_1611);
nor U2264 (N_2264,N_1240,N_1743);
nand U2265 (N_2265,N_346,N_1276);
nor U2266 (N_2266,N_1619,N_559);
and U2267 (N_2267,N_506,N_1472);
nand U2268 (N_2268,N_878,N_544);
or U2269 (N_2269,N_468,N_463);
or U2270 (N_2270,N_923,N_593);
nor U2271 (N_2271,N_1914,N_968);
or U2272 (N_2272,N_392,N_1531);
and U2273 (N_2273,N_570,N_1750);
and U2274 (N_2274,N_209,N_451);
nor U2275 (N_2275,N_1008,N_665);
xnor U2276 (N_2276,N_1004,N_344);
nand U2277 (N_2277,N_1312,N_482);
nor U2278 (N_2278,N_362,N_534);
and U2279 (N_2279,N_1025,N_497);
nand U2280 (N_2280,N_951,N_947);
nand U2281 (N_2281,N_921,N_620);
xor U2282 (N_2282,N_1374,N_793);
nand U2283 (N_2283,N_194,N_912);
nand U2284 (N_2284,N_1548,N_1293);
xor U2285 (N_2285,N_1358,N_83);
xnor U2286 (N_2286,N_1367,N_1766);
nand U2287 (N_2287,N_933,N_1500);
and U2288 (N_2288,N_1510,N_980);
and U2289 (N_2289,N_1712,N_128);
nand U2290 (N_2290,N_959,N_841);
or U2291 (N_2291,N_204,N_1523);
nand U2292 (N_2292,N_481,N_1408);
nand U2293 (N_2293,N_1745,N_1381);
or U2294 (N_2294,N_257,N_918);
nor U2295 (N_2295,N_177,N_1638);
nand U2296 (N_2296,N_1621,N_1049);
nand U2297 (N_2297,N_1135,N_1917);
nor U2298 (N_2298,N_1509,N_153);
nand U2299 (N_2299,N_858,N_264);
nand U2300 (N_2300,N_515,N_1671);
or U2301 (N_2301,N_424,N_187);
nor U2302 (N_2302,N_1926,N_1649);
nor U2303 (N_2303,N_1175,N_1340);
nor U2304 (N_2304,N_914,N_77);
nor U2305 (N_2305,N_349,N_1426);
or U2306 (N_2306,N_304,N_709);
nor U2307 (N_2307,N_342,N_1582);
and U2308 (N_2308,N_1451,N_1222);
xnor U2309 (N_2309,N_1233,N_785);
nor U2310 (N_2310,N_1655,N_1220);
and U2311 (N_2311,N_1993,N_16);
nor U2312 (N_2312,N_1355,N_1375);
or U2313 (N_2313,N_1041,N_1630);
nand U2314 (N_2314,N_1577,N_1356);
nand U2315 (N_2315,N_364,N_1118);
and U2316 (N_2316,N_111,N_299);
xnor U2317 (N_2317,N_32,N_735);
nor U2318 (N_2318,N_1140,N_372);
and U2319 (N_2319,N_288,N_560);
nor U2320 (N_2320,N_974,N_926);
nand U2321 (N_2321,N_212,N_1225);
and U2322 (N_2322,N_1640,N_1758);
and U2323 (N_2323,N_875,N_707);
and U2324 (N_2324,N_1136,N_1625);
and U2325 (N_2325,N_742,N_1641);
nor U2326 (N_2326,N_290,N_680);
nand U2327 (N_2327,N_1093,N_151);
nand U2328 (N_2328,N_1526,N_296);
or U2329 (N_2329,N_1674,N_97);
and U2330 (N_2330,N_1170,N_1361);
or U2331 (N_2331,N_1680,N_1596);
or U2332 (N_2332,N_1262,N_303);
or U2333 (N_2333,N_525,N_71);
or U2334 (N_2334,N_28,N_950);
nand U2335 (N_2335,N_902,N_281);
nor U2336 (N_2336,N_1463,N_1830);
and U2337 (N_2337,N_286,N_604);
nand U2338 (N_2338,N_916,N_52);
nand U2339 (N_2339,N_348,N_1673);
and U2340 (N_2340,N_1654,N_887);
or U2341 (N_2341,N_426,N_436);
nor U2342 (N_2342,N_1153,N_1618);
nor U2343 (N_2343,N_119,N_826);
nand U2344 (N_2344,N_294,N_337);
nand U2345 (N_2345,N_1590,N_140);
nand U2346 (N_2346,N_1627,N_404);
and U2347 (N_2347,N_1146,N_22);
nand U2348 (N_2348,N_1055,N_1210);
xor U2349 (N_2349,N_816,N_1241);
nand U2350 (N_2350,N_375,N_550);
and U2351 (N_2351,N_1959,N_1924);
nand U2352 (N_2352,N_1700,N_1096);
and U2353 (N_2353,N_569,N_646);
nand U2354 (N_2354,N_1436,N_1402);
and U2355 (N_2355,N_1642,N_1698);
and U2356 (N_2356,N_368,N_365);
nand U2357 (N_2357,N_1971,N_937);
and U2358 (N_2358,N_1007,N_614);
nand U2359 (N_2359,N_641,N_203);
and U2360 (N_2360,N_1036,N_669);
or U2361 (N_2361,N_1338,N_1254);
nand U2362 (N_2362,N_615,N_676);
xnor U2363 (N_2363,N_1635,N_958);
or U2364 (N_2364,N_1978,N_1395);
or U2365 (N_2365,N_1111,N_1490);
nand U2366 (N_2366,N_1271,N_976);
nor U2367 (N_2367,N_1494,N_236);
or U2368 (N_2368,N_1325,N_1951);
or U2369 (N_2369,N_231,N_235);
xnor U2370 (N_2370,N_1102,N_1316);
or U2371 (N_2371,N_195,N_276);
nor U2372 (N_2372,N_432,N_1587);
or U2373 (N_2373,N_1303,N_84);
and U2374 (N_2374,N_1953,N_160);
nor U2375 (N_2375,N_311,N_220);
xor U2376 (N_2376,N_1391,N_1445);
nor U2377 (N_2377,N_141,N_1679);
nand U2378 (N_2378,N_910,N_1259);
and U2379 (N_2379,N_1054,N_1073);
and U2380 (N_2380,N_1218,N_705);
nand U2381 (N_2381,N_422,N_606);
or U2382 (N_2382,N_385,N_1564);
and U2383 (N_2383,N_1066,N_689);
nor U2384 (N_2384,N_1780,N_1372);
xor U2385 (N_2385,N_848,N_1862);
and U2386 (N_2386,N_865,N_1411);
or U2387 (N_2387,N_1841,N_329);
xor U2388 (N_2388,N_531,N_940);
or U2389 (N_2389,N_1896,N_684);
nand U2390 (N_2390,N_1670,N_746);
nand U2391 (N_2391,N_649,N_1594);
nor U2392 (N_2392,N_1318,N_39);
or U2393 (N_2393,N_1068,N_1464);
and U2394 (N_2394,N_764,N_1339);
or U2395 (N_2395,N_214,N_650);
nor U2396 (N_2396,N_1305,N_1507);
nor U2397 (N_2397,N_1612,N_50);
or U2398 (N_2398,N_1650,N_1260);
and U2399 (N_2399,N_576,N_710);
nor U2400 (N_2400,N_1976,N_1770);
and U2401 (N_2401,N_588,N_842);
or U2402 (N_2402,N_1052,N_270);
and U2403 (N_2403,N_492,N_1499);
and U2404 (N_2404,N_272,N_621);
or U2405 (N_2405,N_1828,N_200);
nand U2406 (N_2406,N_1138,N_1282);
nor U2407 (N_2407,N_1434,N_1213);
or U2408 (N_2408,N_578,N_1201);
nand U2409 (N_2409,N_1918,N_498);
nor U2410 (N_2410,N_1105,N_269);
and U2411 (N_2411,N_907,N_855);
and U2412 (N_2412,N_192,N_743);
xor U2413 (N_2413,N_64,N_1620);
nand U2414 (N_2414,N_1684,N_1161);
or U2415 (N_2415,N_230,N_1301);
or U2416 (N_2416,N_1709,N_1663);
nor U2417 (N_2417,N_188,N_1449);
nand U2418 (N_2418,N_1945,N_1660);
xor U2419 (N_2419,N_815,N_1883);
nand U2420 (N_2420,N_1899,N_949);
nor U2421 (N_2421,N_1992,N_1027);
and U2422 (N_2422,N_653,N_1113);
and U2423 (N_2423,N_674,N_759);
and U2424 (N_2424,N_618,N_1289);
and U2425 (N_2425,N_1133,N_1231);
nor U2426 (N_2426,N_145,N_1450);
nand U2427 (N_2427,N_63,N_1943);
nand U2428 (N_2428,N_1687,N_1045);
nor U2429 (N_2429,N_1868,N_681);
and U2430 (N_2430,N_104,N_1214);
or U2431 (N_2431,N_1837,N_118);
nor U2432 (N_2432,N_469,N_788);
nor U2433 (N_2433,N_1669,N_491);
nand U2434 (N_2434,N_1740,N_1768);
and U2435 (N_2435,N_1703,N_470);
nand U2436 (N_2436,N_1227,N_384);
nand U2437 (N_2437,N_1030,N_26);
nand U2438 (N_2438,N_675,N_412);
xnor U2439 (N_2439,N_1249,N_1125);
nand U2440 (N_2440,N_53,N_814);
or U2441 (N_2441,N_571,N_514);
nor U2442 (N_2442,N_1037,N_540);
and U2443 (N_2443,N_155,N_827);
nor U2444 (N_2444,N_1124,N_1405);
nor U2445 (N_2445,N_1457,N_822);
or U2446 (N_2446,N_234,N_1559);
or U2447 (N_2447,N_919,N_1997);
nor U2448 (N_2448,N_1198,N_1013);
nor U2449 (N_2449,N_247,N_542);
nand U2450 (N_2450,N_663,N_211);
nand U2451 (N_2451,N_975,N_1704);
or U2452 (N_2452,N_443,N_1474);
or U2453 (N_2453,N_95,N_1946);
and U2454 (N_2454,N_1205,N_1845);
nand U2455 (N_2455,N_1906,N_1570);
or U2456 (N_2456,N_425,N_1024);
and U2457 (N_2457,N_1206,N_1128);
nand U2458 (N_2458,N_582,N_460);
and U2459 (N_2459,N_784,N_1018);
and U2460 (N_2460,N_1473,N_1536);
nor U2461 (N_2461,N_239,N_1117);
or U2462 (N_2462,N_1023,N_1788);
nand U2463 (N_2463,N_712,N_1022);
and U2464 (N_2464,N_1481,N_163);
nor U2465 (N_2465,N_1546,N_879);
or U2466 (N_2466,N_1257,N_846);
or U2467 (N_2467,N_1397,N_1101);
and U2468 (N_2468,N_319,N_583);
or U2469 (N_2469,N_70,N_1566);
or U2470 (N_2470,N_1005,N_1741);
or U2471 (N_2471,N_1141,N_350);
nor U2472 (N_2472,N_45,N_721);
nor U2473 (N_2473,N_261,N_584);
nor U2474 (N_2474,N_1177,N_1496);
nand U2475 (N_2475,N_806,N_1203);
and U2476 (N_2476,N_1961,N_428);
xnor U2477 (N_2477,N_774,N_626);
or U2478 (N_2478,N_862,N_1916);
nand U2479 (N_2479,N_1284,N_994);
and U2480 (N_2480,N_1805,N_120);
or U2481 (N_2481,N_1563,N_40);
nor U2482 (N_2482,N_995,N_1003);
or U2483 (N_2483,N_244,N_1459);
or U2484 (N_2484,N_334,N_1705);
nand U2485 (N_2485,N_532,N_1547);
and U2486 (N_2486,N_361,N_1330);
xnor U2487 (N_2487,N_440,N_781);
or U2488 (N_2488,N_1607,N_1608);
nand U2489 (N_2489,N_243,N_1796);
nor U2490 (N_2490,N_1793,N_942);
xor U2491 (N_2491,N_1748,N_1821);
xnor U2492 (N_2492,N_640,N_1495);
nand U2493 (N_2493,N_1975,N_82);
xnor U2494 (N_2494,N_600,N_1387);
nor U2495 (N_2495,N_1152,N_587);
nand U2496 (N_2496,N_1968,N_1172);
and U2497 (N_2497,N_1280,N_1580);
or U2498 (N_2498,N_1383,N_245);
and U2499 (N_2499,N_466,N_535);
nand U2500 (N_2500,N_352,N_478);
nor U2501 (N_2501,N_1299,N_317);
nor U2502 (N_2502,N_690,N_1990);
nand U2503 (N_2503,N_237,N_1925);
nand U2504 (N_2504,N_1485,N_931);
nand U2505 (N_2505,N_301,N_1327);
nand U2506 (N_2506,N_67,N_572);
and U2507 (N_2507,N_347,N_1145);
nor U2508 (N_2508,N_637,N_1089);
or U2509 (N_2509,N_467,N_58);
nor U2510 (N_2510,N_2,N_1977);
nand U2511 (N_2511,N_1192,N_732);
nand U2512 (N_2512,N_1528,N_1825);
and U2513 (N_2513,N_898,N_176);
nand U2514 (N_2514,N_396,N_1149);
and U2515 (N_2515,N_1173,N_1866);
xnor U2516 (N_2516,N_1430,N_1631);
nand U2517 (N_2517,N_96,N_1854);
or U2518 (N_2518,N_1197,N_106);
or U2519 (N_2519,N_88,N_1726);
and U2520 (N_2520,N_538,N_1927);
nor U2521 (N_2521,N_125,N_44);
nand U2522 (N_2522,N_33,N_1448);
nor U2523 (N_2523,N_10,N_321);
nand U2524 (N_2524,N_1076,N_377);
or U2525 (N_2525,N_1091,N_376);
and U2526 (N_2526,N_233,N_1319);
nand U2527 (N_2527,N_1932,N_56);
nand U2528 (N_2528,N_313,N_1984);
or U2529 (N_2529,N_1930,N_91);
nand U2530 (N_2530,N_1936,N_291);
nand U2531 (N_2531,N_1428,N_232);
or U2532 (N_2532,N_1369,N_825);
and U2533 (N_2533,N_1567,N_338);
and U2534 (N_2534,N_652,N_1639);
or U2535 (N_2535,N_1238,N_691);
and U2536 (N_2536,N_1560,N_1988);
or U2537 (N_2537,N_807,N_798);
or U2538 (N_2538,N_1822,N_539);
and U2539 (N_2539,N_292,N_196);
nor U2540 (N_2540,N_1234,N_124);
and U2541 (N_2541,N_72,N_1632);
or U2542 (N_2542,N_715,N_1458);
or U2543 (N_2543,N_1042,N_727);
nand U2544 (N_2544,N_821,N_1179);
nor U2545 (N_2545,N_929,N_1009);
nor U2546 (N_2546,N_782,N_1151);
and U2547 (N_2547,N_1800,N_1781);
or U2548 (N_2548,N_1521,N_1603);
nand U2549 (N_2549,N_1986,N_1083);
and U2550 (N_2550,N_358,N_419);
nor U2551 (N_2551,N_55,N_835);
and U2552 (N_2552,N_832,N_545);
xnor U2553 (N_2553,N_1142,N_1874);
or U2554 (N_2554,N_438,N_1143);
or U2555 (N_2555,N_1229,N_1939);
nand U2556 (N_2556,N_656,N_1763);
or U2557 (N_2557,N_105,N_1505);
or U2558 (N_2558,N_1415,N_714);
xnor U2559 (N_2559,N_889,N_1017);
or U2560 (N_2560,N_1169,N_1760);
xnor U2561 (N_2561,N_1156,N_1191);
or U2562 (N_2562,N_972,N_927);
and U2563 (N_2563,N_455,N_1159);
or U2564 (N_2564,N_1114,N_504);
or U2565 (N_2565,N_1554,N_932);
or U2566 (N_2566,N_1493,N_1221);
or U2567 (N_2567,N_479,N_753);
or U2568 (N_2568,N_1337,N_476);
nor U2569 (N_2569,N_1815,N_24);
xor U2570 (N_2570,N_409,N_1693);
and U2571 (N_2571,N_758,N_659);
nor U2572 (N_2572,N_1817,N_711);
xor U2573 (N_2573,N_190,N_251);
and U2574 (N_2574,N_747,N_1296);
nand U2575 (N_2575,N_1164,N_1482);
xor U2576 (N_2576,N_1863,N_103);
or U2577 (N_2577,N_250,N_1551);
nor U2578 (N_2578,N_1267,N_953);
and U2579 (N_2579,N_49,N_852);
nor U2580 (N_2580,N_12,N_1178);
or U2581 (N_2581,N_122,N_1195);
nor U2582 (N_2582,N_1904,N_1287);
nor U2583 (N_2583,N_1126,N_123);
or U2584 (N_2584,N_725,N_558);
or U2585 (N_2585,N_341,N_1456);
nor U2586 (N_2586,N_255,N_734);
nand U2587 (N_2587,N_1110,N_1767);
nand U2588 (N_2588,N_901,N_1389);
nor U2589 (N_2589,N_1586,N_1719);
nor U2590 (N_2590,N_489,N_1404);
nand U2591 (N_2591,N_437,N_840);
or U2592 (N_2592,N_1460,N_1295);
xnor U2593 (N_2593,N_1477,N_1876);
nor U2594 (N_2594,N_744,N_1286);
or U2595 (N_2595,N_1194,N_353);
or U2596 (N_2596,N_1116,N_23);
or U2597 (N_2597,N_1438,N_1353);
or U2598 (N_2598,N_502,N_457);
or U2599 (N_2599,N_69,N_1755);
nand U2600 (N_2600,N_1690,N_1729);
nor U2601 (N_2601,N_1732,N_1199);
xor U2602 (N_2602,N_1792,N_1695);
or U2603 (N_2603,N_1028,N_603);
nor U2604 (N_2604,N_853,N_46);
or U2605 (N_2605,N_549,N_1502);
and U2606 (N_2606,N_1237,N_1080);
nor U2607 (N_2607,N_521,N_636);
and U2608 (N_2608,N_248,N_223);
nor U2609 (N_2609,N_616,N_643);
or U2610 (N_2610,N_1401,N_395);
or U2611 (N_2611,N_599,N_553);
and U2612 (N_2612,N_1893,N_14);
nor U2613 (N_2613,N_30,N_1331);
nand U2614 (N_2614,N_59,N_1162);
and U2615 (N_2615,N_948,N_1530);
nor U2616 (N_2616,N_971,N_60);
and U2617 (N_2617,N_1941,N_447);
nor U2618 (N_2618,N_1390,N_780);
and U2619 (N_2619,N_1851,N_1341);
nand U2620 (N_2620,N_1503,N_65);
nor U2621 (N_2621,N_1873,N_1557);
nand U2622 (N_2622,N_487,N_400);
nor U2623 (N_2623,N_38,N_1814);
nor U2624 (N_2624,N_265,N_1119);
or U2625 (N_2625,N_133,N_1762);
nor U2626 (N_2626,N_1761,N_1752);
and U2627 (N_2627,N_41,N_1960);
or U2628 (N_2628,N_1403,N_568);
nand U2629 (N_2629,N_1409,N_61);
nor U2630 (N_2630,N_752,N_1579);
nand U2631 (N_2631,N_17,N_922);
nor U2632 (N_2632,N_1400,N_454);
or U2633 (N_2633,N_1256,N_488);
or U2634 (N_2634,N_536,N_215);
and U2635 (N_2635,N_1035,N_622);
nand U2636 (N_2636,N_589,N_360);
xnor U2637 (N_2637,N_5,N_1730);
and U2638 (N_2638,N_1120,N_462);
and U2639 (N_2639,N_1398,N_930);
and U2640 (N_2640,N_666,N_114);
nor U2641 (N_2641,N_738,N_483);
or U2642 (N_2642,N_1311,N_1302);
nor U2643 (N_2643,N_1865,N_495);
xnor U2644 (N_2644,N_148,N_262);
xnor U2645 (N_2645,N_472,N_1965);
or U2646 (N_2646,N_1046,N_1604);
or U2647 (N_2647,N_1565,N_1744);
and U2648 (N_2648,N_1871,N_1533);
or U2649 (N_2649,N_1462,N_48);
nand U2650 (N_2650,N_1728,N_1593);
or U2651 (N_2651,N_537,N_1016);
nand U2652 (N_2652,N_913,N_7);
nand U2653 (N_2653,N_1026,N_51);
nand U2654 (N_2654,N_1860,N_899);
nor U2655 (N_2655,N_1622,N_1581);
nor U2656 (N_2656,N_991,N_886);
or U2657 (N_2657,N_1278,N_1364);
xor U2658 (N_2658,N_477,N_1314);
and U2659 (N_2659,N_1966,N_4);
nand U2660 (N_2660,N_590,N_1633);
xnor U2661 (N_2661,N_1081,N_1733);
nand U2662 (N_2662,N_698,N_511);
and U2663 (N_2663,N_1307,N_1980);
or U2664 (N_2664,N_1273,N_25);
nor U2665 (N_2665,N_581,N_228);
nor U2666 (N_2666,N_800,N_1783);
nand U2667 (N_2667,N_1908,N_1410);
nor U2668 (N_2668,N_1185,N_1849);
nor U2669 (N_2669,N_1995,N_642);
or U2670 (N_2670,N_864,N_905);
and U2671 (N_2671,N_1713,N_1384);
nor U2672 (N_2672,N_687,N_1425);
nand U2673 (N_2673,N_1722,N_786);
or U2674 (N_2674,N_1439,N_1589);
and U2675 (N_2675,N_1060,N_795);
xnor U2676 (N_2676,N_277,N_1486);
and U2677 (N_2677,N_733,N_739);
nor U2678 (N_2678,N_1550,N_112);
or U2679 (N_2679,N_225,N_891);
and U2680 (N_2680,N_183,N_1944);
nor U2681 (N_2681,N_938,N_829);
or U2682 (N_2682,N_796,N_897);
and U2683 (N_2683,N_1880,N_1834);
or U2684 (N_2684,N_1132,N_323);
nor U2685 (N_2685,N_708,N_1875);
nor U2686 (N_2686,N_1545,N_1846);
nor U2687 (N_2687,N_867,N_1989);
xnor U2688 (N_2688,N_1061,N_1461);
or U2689 (N_2689,N_1098,N_1085);
or U2690 (N_2690,N_1454,N_1084);
nor U2691 (N_2691,N_1020,N_895);
xor U2692 (N_2692,N_977,N_1204);
and U2693 (N_2693,N_1819,N_1666);
xor U2694 (N_2694,N_430,N_507);
and U2695 (N_2695,N_577,N_1188);
and U2696 (N_2696,N_1168,N_1662);
and U2697 (N_2697,N_702,N_667);
nor U2698 (N_2698,N_1881,N_598);
and U2699 (N_2699,N_1380,N_1212);
nor U2700 (N_2700,N_1676,N_1514);
and U2701 (N_2701,N_414,N_252);
and U2702 (N_2702,N_1973,N_1285);
nand U2703 (N_2703,N_728,N_249);
xor U2704 (N_2704,N_143,N_1731);
and U2705 (N_2705,N_174,N_1910);
and U2706 (N_2706,N_941,N_81);
xnor U2707 (N_2707,N_1736,N_1435);
or U2708 (N_2708,N_1573,N_844);
and U2709 (N_2709,N_1963,N_1051);
nor U2710 (N_2710,N_915,N_271);
nand U2711 (N_2711,N_512,N_79);
and U2712 (N_2712,N_1812,N_1371);
nor U2713 (N_2713,N_1795,N_475);
or U2714 (N_2714,N_293,N_594);
or U2715 (N_2715,N_1711,N_1572);
or U2716 (N_2716,N_213,N_1739);
xor U2717 (N_2717,N_306,N_147);
nor U2718 (N_2718,N_115,N_1326);
nor U2719 (N_2719,N_1343,N_199);
and U2720 (N_2720,N_900,N_189);
xor U2721 (N_2721,N_1628,N_1870);
or U2722 (N_2722,N_62,N_1664);
xor U2723 (N_2723,N_592,N_906);
xnor U2724 (N_2724,N_609,N_778);
nand U2725 (N_2725,N_1476,N_1522);
or U2726 (N_2726,N_101,N_1901);
xnor U2727 (N_2727,N_1443,N_1150);
and U2728 (N_2728,N_790,N_1377);
xor U2729 (N_2729,N_1725,N_146);
and U2730 (N_2730,N_946,N_1180);
nor U2731 (N_2731,N_42,N_435);
nor U2732 (N_2732,N_1181,N_1806);
nand U2733 (N_2733,N_1685,N_1900);
nand U2734 (N_2734,N_158,N_138);
nand U2735 (N_2735,N_1144,N_812);
nand U2736 (N_2736,N_1491,N_282);
xnor U2737 (N_2737,N_1840,N_1444);
nor U2738 (N_2738,N_526,N_1598);
nand U2739 (N_2739,N_1576,N_1691);
and U2740 (N_2740,N_1131,N_318);
and U2741 (N_2741,N_166,N_1006);
nor U2742 (N_2742,N_100,N_1315);
xor U2743 (N_2743,N_957,N_1710);
nand U2744 (N_2744,N_1313,N_238);
nor U2745 (N_2745,N_1665,N_1394);
xor U2746 (N_2746,N_205,N_1789);
or U2747 (N_2747,N_591,N_207);
and U2748 (N_2748,N_413,N_1247);
nor U2749 (N_2749,N_1040,N_881);
and U2750 (N_2750,N_1898,N_1348);
xnor U2751 (N_2751,N_1843,N_1378);
nand U2752 (N_2752,N_47,N_1261);
or U2753 (N_2753,N_1274,N_1599);
nor U2754 (N_2754,N_696,N_1414);
xor U2755 (N_2755,N_1974,N_657);
nor U2756 (N_2756,N_1801,N_1972);
nand U2757 (N_2757,N_1699,N_1386);
nand U2758 (N_2758,N_1190,N_1967);
or U2759 (N_2759,N_221,N_1441);
or U2760 (N_2760,N_420,N_1121);
or U2761 (N_2761,N_1606,N_1334);
or U2762 (N_2762,N_98,N_229);
nor U2763 (N_2763,N_1646,N_522);
or U2764 (N_2764,N_960,N_820);
and U2765 (N_2765,N_309,N_164);
xnor U2766 (N_2766,N_1890,N_608);
nor U2767 (N_2767,N_421,N_416);
or U2768 (N_2768,N_279,N_1034);
or U2769 (N_2769,N_380,N_1701);
xor U2770 (N_2770,N_519,N_1658);
and U2771 (N_2771,N_1552,N_1413);
nor U2772 (N_2772,N_169,N_1242);
nor U2773 (N_2773,N_1359,N_546);
xnor U2774 (N_2774,N_763,N_268);
nor U2775 (N_2775,N_510,N_1848);
nand U2776 (N_2776,N_330,N_629);
and U2777 (N_2777,N_1243,N_1465);
nand U2778 (N_2778,N_831,N_1029);
nor U2779 (N_2779,N_126,N_29);
nor U2780 (N_2780,N_345,N_139);
nand U2781 (N_2781,N_121,N_893);
or U2782 (N_2782,N_406,N_242);
nor U2783 (N_2783,N_1239,N_1471);
and U2784 (N_2784,N_197,N_908);
nor U2785 (N_2785,N_314,N_275);
xor U2786 (N_2786,N_1786,N_78);
xnor U2787 (N_2787,N_1681,N_1365);
and U2788 (N_2788,N_1983,N_854);
nor U2789 (N_2789,N_1602,N_1160);
xnor U2790 (N_2790,N_992,N_1291);
and U2791 (N_2791,N_1182,N_811);
nor U2792 (N_2792,N_1667,N_367);
or U2793 (N_2793,N_1193,N_1931);
nor U2794 (N_2794,N_1538,N_108);
nand U2795 (N_2795,N_772,N_357);
nand U2796 (N_2796,N_1644,N_198);
nand U2797 (N_2797,N_1270,N_1363);
nor U2798 (N_2798,N_452,N_1070);
xnor U2799 (N_2799,N_1575,N_206);
or U2800 (N_2800,N_611,N_1723);
nor U2801 (N_2801,N_1517,N_837);
or U2802 (N_2802,N_1519,N_191);
and U2803 (N_2803,N_1134,N_1885);
and U2804 (N_2804,N_1991,N_954);
and U2805 (N_2805,N_499,N_1859);
or U2806 (N_2806,N_1223,N_877);
and U2807 (N_2807,N_880,N_1797);
xor U2808 (N_2808,N_1455,N_1623);
and U2809 (N_2809,N_1468,N_966);
xor U2810 (N_2810,N_340,N_1597);
and U2811 (N_2811,N_1803,N_1373);
or U2812 (N_2812,N_911,N_563);
xor U2813 (N_2813,N_284,N_982);
nand U2814 (N_2814,N_624,N_1154);
and U2815 (N_2815,N_1749,N_1504);
or U2816 (N_2816,N_809,N_256);
xnor U2817 (N_2817,N_1344,N_903);
or U2818 (N_2818,N_173,N_1541);
or U2819 (N_2819,N_382,N_851);
and U2820 (N_2820,N_1772,N_1512);
and U2821 (N_2821,N_300,N_967);
and U2822 (N_2822,N_1888,N_1071);
and U2823 (N_2823,N_1555,N_1802);
and U2824 (N_2824,N_403,N_1324);
nor U2825 (N_2825,N_80,N_1682);
or U2826 (N_2826,N_1715,N_973);
nand U2827 (N_2827,N_632,N_1850);
and U2828 (N_2828,N_1069,N_433);
or U2829 (N_2829,N_1167,N_766);
and U2830 (N_2830,N_246,N_132);
nand U2831 (N_2831,N_1889,N_726);
nor U2832 (N_2832,N_107,N_76);
nor U2833 (N_2833,N_1909,N_1724);
nand U2834 (N_2834,N_325,N_990);
nor U2835 (N_2835,N_1090,N_1431);
and U2836 (N_2836,N_892,N_1905);
and U2837 (N_2837,N_1790,N_1283);
nor U2838 (N_2838,N_1251,N_1092);
and U2839 (N_2839,N_19,N_89);
or U2840 (N_2840,N_1470,N_1689);
and U2841 (N_2841,N_997,N_1515);
and U2842 (N_2842,N_285,N_765);
and U2843 (N_2843,N_524,N_298);
and U2844 (N_2844,N_1012,N_156);
nand U2845 (N_2845,N_736,N_1062);
or U2846 (N_2846,N_1735,N_1432);
and U2847 (N_2847,N_373,N_981);
nor U2848 (N_2848,N_310,N_628);
or U2849 (N_2849,N_493,N_1345);
and U2850 (N_2850,N_184,N_278);
nand U2851 (N_2851,N_701,N_1264);
nor U2852 (N_2852,N_165,N_1467);
xor U2853 (N_2853,N_1320,N_1543);
and U2854 (N_2854,N_427,N_1838);
and U2855 (N_2855,N_775,N_1388);
xnor U2856 (N_2856,N_830,N_1304);
xnor U2857 (N_2857,N_458,N_1982);
and U2858 (N_2858,N_1253,N_1196);
or U2859 (N_2859,N_1892,N_1721);
or U2860 (N_2860,N_574,N_1176);
nand U2861 (N_2861,N_1184,N_555);
and U2862 (N_2862,N_943,N_1692);
nand U2863 (N_2863,N_856,N_1524);
nand U2864 (N_2864,N_1082,N_1245);
nor U2865 (N_2865,N_1535,N_1754);
and U2866 (N_2866,N_1158,N_1244);
nor U2867 (N_2867,N_1764,N_1329);
nand U2868 (N_2868,N_1702,N_955);
and U2869 (N_2869,N_1938,N_1636);
or U2870 (N_2870,N_1952,N_431);
nor U2871 (N_2871,N_1058,N_1050);
and U2872 (N_2872,N_803,N_1418);
nand U2873 (N_2873,N_1833,N_872);
xor U2874 (N_2874,N_706,N_1148);
and U2875 (N_2875,N_87,N_797);
or U2876 (N_2876,N_804,N_1235);
or U2877 (N_2877,N_439,N_1858);
or U2878 (N_2878,N_266,N_1053);
nor U2879 (N_2879,N_1279,N_882);
and U2880 (N_2880,N_43,N_31);
nor U2881 (N_2881,N_703,N_754);
xnor U2882 (N_2882,N_1911,N_612);
nand U2883 (N_2883,N_11,N_93);
nor U2884 (N_2884,N_1532,N_644);
nor U2885 (N_2885,N_1429,N_888);
or U2886 (N_2886,N_1922,N_289);
and U2887 (N_2887,N_405,N_1211);
or U2888 (N_2888,N_1086,N_773);
nand U2889 (N_2889,N_1777,N_1236);
nor U2890 (N_2890,N_170,N_1827);
or U2891 (N_2891,N_1882,N_1157);
xor U2892 (N_2892,N_630,N_485);
and U2893 (N_2893,N_762,N_149);
nor U2894 (N_2894,N_1048,N_1139);
or U2895 (N_2895,N_1368,N_474);
or U2896 (N_2896,N_694,N_1127);
or U2897 (N_2897,N_1351,N_1508);
or U2898 (N_2898,N_595,N_351);
and U2899 (N_2899,N_418,N_324);
and U2900 (N_2900,N_939,N_518);
and U2901 (N_2901,N_1773,N_792);
and U2902 (N_2902,N_586,N_1549);
and U2903 (N_2903,N_1392,N_193);
nand U2904 (N_2904,N_297,N_501);
nor U2905 (N_2905,N_1751,N_859);
xor U2906 (N_2906,N_1165,N_1466);
and U2907 (N_2907,N_965,N_18);
xor U2908 (N_2908,N_1869,N_417);
nand U2909 (N_2909,N_670,N_1624);
xor U2910 (N_2910,N_1717,N_770);
or U2911 (N_2911,N_86,N_1937);
nand U2912 (N_2912,N_1872,N_1306);
nand U2913 (N_2913,N_113,N_1903);
nor U2914 (N_2914,N_1574,N_1661);
or U2915 (N_2915,N_602,N_240);
nand U2916 (N_2916,N_410,N_1427);
or U2917 (N_2917,N_1823,N_1714);
nand U2918 (N_2918,N_1955,N_1672);
or U2919 (N_2919,N_1884,N_379);
or U2920 (N_2920,N_1921,N_1525);
or U2921 (N_2921,N_326,N_1447);
nand U2922 (N_2922,N_1609,N_1738);
and U2923 (N_2923,N_1104,N_1929);
nand U2924 (N_2924,N_917,N_1079);
nor U2925 (N_2925,N_496,N_970);
nor U2926 (N_2926,N_1095,N_1217);
nor U2927 (N_2927,N_749,N_90);
xor U2928 (N_2928,N_896,N_378);
nor U2929 (N_2929,N_1039,N_1776);
and U2930 (N_2930,N_371,N_1668);
nand U2931 (N_2931,N_695,N_533);
nand U2932 (N_2932,N_528,N_1317);
and U2933 (N_2933,N_1015,N_575);
nor U2934 (N_2934,N_751,N_768);
xnor U2935 (N_2935,N_873,N_857);
nand U2936 (N_2936,N_987,N_356);
and U2937 (N_2937,N_1964,N_343);
nor U2938 (N_2938,N_1183,N_655);
nor U2939 (N_2939,N_1067,N_1063);
xor U2940 (N_2940,N_557,N_1200);
xnor U2941 (N_2941,N_945,N_1785);
or U2942 (N_2942,N_484,N_464);
nand U2943 (N_2943,N_654,N_530);
nand U2944 (N_2944,N_1956,N_1696);
xnor U2945 (N_2945,N_1605,N_777);
or U2946 (N_2946,N_1775,N_567);
and U2947 (N_2947,N_383,N_1288);
nor U2948 (N_2948,N_1424,N_850);
or U2949 (N_2949,N_1002,N_731);
nand U2950 (N_2950,N_661,N_1969);
and U2951 (N_2951,N_1122,N_1171);
or U2952 (N_2952,N_605,N_1920);
and U2953 (N_2953,N_1615,N_1765);
and U2954 (N_2954,N_1097,N_154);
nand U2955 (N_2955,N_1332,N_130);
or U2956 (N_2956,N_411,N_1186);
or U2957 (N_2957,N_1333,N_423);
xor U2958 (N_2958,N_137,N_717);
and U2959 (N_2959,N_332,N_1290);
or U2960 (N_2960,N_839,N_1829);
or U2961 (N_2961,N_964,N_720);
nor U2962 (N_2962,N_74,N_1057);
and U2963 (N_2963,N_1954,N_386);
or U2964 (N_2964,N_1867,N_1645);
or U2965 (N_2965,N_1357,N_1588);
or U2966 (N_2966,N_1475,N_171);
nor U2967 (N_2967,N_399,N_1396);
or U2968 (N_2968,N_1799,N_517);
xor U2969 (N_2969,N_1616,N_1887);
or U2970 (N_2970,N_1442,N_473);
nor U2971 (N_2971,N_573,N_1230);
or U2972 (N_2972,N_597,N_1297);
nor U2973 (N_2973,N_1813,N_1422);
or U2974 (N_2974,N_1746,N_988);
nor U2975 (N_2975,N_1109,N_1228);
and U2976 (N_2976,N_1484,N_579);
and U2977 (N_2977,N_1469,N_677);
nor U2978 (N_2978,N_1999,N_890);
nand U2979 (N_2979,N_8,N_142);
and U2980 (N_2980,N_1417,N_1950);
or U2981 (N_2981,N_1987,N_1446);
nand U2982 (N_2982,N_1322,N_1321);
or U2983 (N_2983,N_627,N_1553);
nor U2984 (N_2984,N_1578,N_1246);
nor U2985 (N_2985,N_1677,N_645);
and U2986 (N_2986,N_287,N_434);
and U2987 (N_2987,N_99,N_817);
and U2988 (N_2988,N_1720,N_1919);
and U2989 (N_2989,N_465,N_1349);
nand U2990 (N_2990,N_308,N_1529);
and U2991 (N_2991,N_1108,N_1088);
or U2992 (N_2992,N_834,N_1072);
nor U2993 (N_2993,N_1032,N_819);
and U2994 (N_2994,N_548,N_94);
and U2995 (N_2995,N_639,N_989);
nor U2996 (N_2996,N_601,N_1683);
nand U2997 (N_2997,N_552,N_909);
nor U2998 (N_2998,N_924,N_1913);
and U2999 (N_2999,N_1844,N_996);
and U3000 (N_3000,N_1536,N_515);
or U3001 (N_3001,N_15,N_681);
xnor U3002 (N_3002,N_406,N_1269);
and U3003 (N_3003,N_3,N_1625);
or U3004 (N_3004,N_1865,N_1066);
and U3005 (N_3005,N_86,N_623);
nand U3006 (N_3006,N_604,N_619);
nor U3007 (N_3007,N_1937,N_618);
nor U3008 (N_3008,N_438,N_69);
and U3009 (N_3009,N_494,N_37);
nand U3010 (N_3010,N_328,N_125);
nand U3011 (N_3011,N_771,N_838);
nor U3012 (N_3012,N_912,N_1568);
xor U3013 (N_3013,N_1395,N_1324);
nand U3014 (N_3014,N_723,N_1519);
or U3015 (N_3015,N_1217,N_1809);
and U3016 (N_3016,N_1963,N_1465);
xnor U3017 (N_3017,N_1771,N_1374);
nand U3018 (N_3018,N_800,N_838);
or U3019 (N_3019,N_962,N_1841);
or U3020 (N_3020,N_342,N_1204);
or U3021 (N_3021,N_55,N_1447);
nand U3022 (N_3022,N_1567,N_578);
nand U3023 (N_3023,N_1581,N_1346);
xor U3024 (N_3024,N_287,N_116);
or U3025 (N_3025,N_1797,N_358);
nand U3026 (N_3026,N_225,N_1265);
or U3027 (N_3027,N_1894,N_1282);
nor U3028 (N_3028,N_1468,N_285);
nand U3029 (N_3029,N_1738,N_1036);
xnor U3030 (N_3030,N_1071,N_748);
nand U3031 (N_3031,N_1709,N_147);
or U3032 (N_3032,N_1158,N_38);
xnor U3033 (N_3033,N_1388,N_32);
nor U3034 (N_3034,N_1835,N_1870);
nand U3035 (N_3035,N_757,N_904);
or U3036 (N_3036,N_670,N_1528);
nand U3037 (N_3037,N_749,N_1158);
or U3038 (N_3038,N_81,N_89);
nand U3039 (N_3039,N_1539,N_1418);
nand U3040 (N_3040,N_42,N_1980);
nor U3041 (N_3041,N_38,N_1419);
nor U3042 (N_3042,N_1504,N_1869);
nor U3043 (N_3043,N_865,N_1791);
xor U3044 (N_3044,N_1893,N_224);
nor U3045 (N_3045,N_833,N_132);
nand U3046 (N_3046,N_567,N_1722);
or U3047 (N_3047,N_1849,N_1948);
and U3048 (N_3048,N_1824,N_998);
xor U3049 (N_3049,N_635,N_1715);
and U3050 (N_3050,N_1303,N_212);
and U3051 (N_3051,N_405,N_1715);
nand U3052 (N_3052,N_180,N_905);
nor U3053 (N_3053,N_341,N_234);
nor U3054 (N_3054,N_1018,N_1511);
and U3055 (N_3055,N_98,N_1730);
and U3056 (N_3056,N_610,N_1228);
or U3057 (N_3057,N_1573,N_1738);
nor U3058 (N_3058,N_617,N_831);
xnor U3059 (N_3059,N_869,N_1498);
and U3060 (N_3060,N_213,N_846);
nor U3061 (N_3061,N_333,N_1949);
nand U3062 (N_3062,N_1344,N_0);
nor U3063 (N_3063,N_1354,N_604);
xnor U3064 (N_3064,N_1335,N_1617);
nor U3065 (N_3065,N_213,N_1471);
nand U3066 (N_3066,N_1857,N_704);
and U3067 (N_3067,N_343,N_1131);
and U3068 (N_3068,N_369,N_1768);
nor U3069 (N_3069,N_706,N_483);
and U3070 (N_3070,N_1600,N_335);
or U3071 (N_3071,N_577,N_1886);
and U3072 (N_3072,N_1012,N_57);
nor U3073 (N_3073,N_814,N_264);
and U3074 (N_3074,N_1795,N_394);
nand U3075 (N_3075,N_1167,N_491);
nand U3076 (N_3076,N_1651,N_1244);
or U3077 (N_3077,N_164,N_486);
nor U3078 (N_3078,N_1779,N_654);
and U3079 (N_3079,N_1920,N_783);
or U3080 (N_3080,N_1652,N_1830);
nand U3081 (N_3081,N_1432,N_1430);
and U3082 (N_3082,N_653,N_30);
nand U3083 (N_3083,N_1688,N_570);
and U3084 (N_3084,N_528,N_688);
nand U3085 (N_3085,N_687,N_1694);
nor U3086 (N_3086,N_1209,N_1354);
xor U3087 (N_3087,N_1851,N_418);
nand U3088 (N_3088,N_156,N_1912);
nand U3089 (N_3089,N_86,N_445);
nor U3090 (N_3090,N_1663,N_1209);
and U3091 (N_3091,N_1136,N_355);
nor U3092 (N_3092,N_766,N_43);
nand U3093 (N_3093,N_544,N_1445);
and U3094 (N_3094,N_497,N_70);
nor U3095 (N_3095,N_756,N_1463);
and U3096 (N_3096,N_1749,N_1613);
or U3097 (N_3097,N_1570,N_1142);
and U3098 (N_3098,N_159,N_331);
nand U3099 (N_3099,N_1108,N_1464);
xor U3100 (N_3100,N_801,N_790);
and U3101 (N_3101,N_461,N_1102);
and U3102 (N_3102,N_763,N_1044);
or U3103 (N_3103,N_1994,N_1690);
nor U3104 (N_3104,N_318,N_1358);
nand U3105 (N_3105,N_877,N_1257);
nor U3106 (N_3106,N_1575,N_859);
nor U3107 (N_3107,N_401,N_482);
or U3108 (N_3108,N_287,N_647);
or U3109 (N_3109,N_1784,N_1054);
or U3110 (N_3110,N_1124,N_1266);
and U3111 (N_3111,N_341,N_1799);
or U3112 (N_3112,N_1036,N_1717);
and U3113 (N_3113,N_1667,N_308);
and U3114 (N_3114,N_1154,N_943);
nand U3115 (N_3115,N_899,N_369);
or U3116 (N_3116,N_1043,N_1656);
nor U3117 (N_3117,N_1310,N_1557);
and U3118 (N_3118,N_1906,N_1185);
nand U3119 (N_3119,N_1732,N_1262);
xnor U3120 (N_3120,N_1862,N_368);
nand U3121 (N_3121,N_1244,N_321);
nor U3122 (N_3122,N_678,N_1910);
or U3123 (N_3123,N_1798,N_1152);
nand U3124 (N_3124,N_111,N_605);
nand U3125 (N_3125,N_1229,N_215);
nor U3126 (N_3126,N_1649,N_1276);
and U3127 (N_3127,N_999,N_864);
and U3128 (N_3128,N_455,N_1112);
nand U3129 (N_3129,N_1317,N_140);
or U3130 (N_3130,N_645,N_437);
and U3131 (N_3131,N_143,N_1932);
xor U3132 (N_3132,N_1207,N_329);
xnor U3133 (N_3133,N_6,N_912);
xor U3134 (N_3134,N_1716,N_180);
nand U3135 (N_3135,N_212,N_1807);
and U3136 (N_3136,N_575,N_1951);
nor U3137 (N_3137,N_907,N_637);
and U3138 (N_3138,N_884,N_1555);
and U3139 (N_3139,N_399,N_1640);
or U3140 (N_3140,N_228,N_1606);
nand U3141 (N_3141,N_392,N_790);
nand U3142 (N_3142,N_1639,N_159);
nand U3143 (N_3143,N_1461,N_890);
xnor U3144 (N_3144,N_365,N_1974);
nor U3145 (N_3145,N_763,N_959);
nor U3146 (N_3146,N_1016,N_1702);
and U3147 (N_3147,N_953,N_240);
nand U3148 (N_3148,N_390,N_1334);
xor U3149 (N_3149,N_1029,N_845);
or U3150 (N_3150,N_483,N_933);
or U3151 (N_3151,N_1510,N_906);
xnor U3152 (N_3152,N_1603,N_1573);
and U3153 (N_3153,N_699,N_1908);
nor U3154 (N_3154,N_690,N_1634);
nor U3155 (N_3155,N_1410,N_594);
nor U3156 (N_3156,N_1079,N_0);
nor U3157 (N_3157,N_369,N_1052);
and U3158 (N_3158,N_645,N_1466);
xor U3159 (N_3159,N_5,N_37);
and U3160 (N_3160,N_382,N_1794);
nand U3161 (N_3161,N_1922,N_804);
and U3162 (N_3162,N_1225,N_902);
and U3163 (N_3163,N_1358,N_397);
or U3164 (N_3164,N_378,N_818);
nand U3165 (N_3165,N_419,N_1435);
xor U3166 (N_3166,N_1085,N_1120);
nor U3167 (N_3167,N_1414,N_449);
xor U3168 (N_3168,N_145,N_159);
xnor U3169 (N_3169,N_1255,N_1548);
and U3170 (N_3170,N_1371,N_201);
and U3171 (N_3171,N_1975,N_1743);
xor U3172 (N_3172,N_608,N_1336);
nand U3173 (N_3173,N_366,N_1400);
xnor U3174 (N_3174,N_1934,N_1609);
xnor U3175 (N_3175,N_748,N_1264);
or U3176 (N_3176,N_1968,N_825);
xnor U3177 (N_3177,N_218,N_1813);
nand U3178 (N_3178,N_1572,N_1692);
or U3179 (N_3179,N_1790,N_250);
nand U3180 (N_3180,N_277,N_1259);
or U3181 (N_3181,N_302,N_31);
and U3182 (N_3182,N_1188,N_735);
or U3183 (N_3183,N_1159,N_1971);
nand U3184 (N_3184,N_1192,N_1840);
and U3185 (N_3185,N_765,N_588);
and U3186 (N_3186,N_955,N_811);
xnor U3187 (N_3187,N_797,N_1724);
or U3188 (N_3188,N_314,N_536);
and U3189 (N_3189,N_1303,N_945);
or U3190 (N_3190,N_77,N_736);
or U3191 (N_3191,N_864,N_21);
nand U3192 (N_3192,N_537,N_102);
or U3193 (N_3193,N_750,N_1651);
and U3194 (N_3194,N_1997,N_760);
and U3195 (N_3195,N_1794,N_355);
and U3196 (N_3196,N_907,N_1117);
nand U3197 (N_3197,N_1809,N_924);
nand U3198 (N_3198,N_1974,N_1218);
nor U3199 (N_3199,N_835,N_668);
or U3200 (N_3200,N_283,N_1672);
and U3201 (N_3201,N_1213,N_217);
and U3202 (N_3202,N_742,N_247);
and U3203 (N_3203,N_454,N_576);
nor U3204 (N_3204,N_1043,N_549);
nor U3205 (N_3205,N_609,N_918);
or U3206 (N_3206,N_1451,N_20);
or U3207 (N_3207,N_1634,N_1385);
nor U3208 (N_3208,N_1225,N_1633);
or U3209 (N_3209,N_1817,N_1134);
nor U3210 (N_3210,N_399,N_957);
nor U3211 (N_3211,N_616,N_1658);
and U3212 (N_3212,N_1251,N_387);
nand U3213 (N_3213,N_273,N_1494);
and U3214 (N_3214,N_459,N_402);
and U3215 (N_3215,N_13,N_5);
nor U3216 (N_3216,N_82,N_1014);
nor U3217 (N_3217,N_1100,N_323);
and U3218 (N_3218,N_907,N_142);
and U3219 (N_3219,N_1186,N_263);
nand U3220 (N_3220,N_1379,N_514);
nand U3221 (N_3221,N_1120,N_797);
or U3222 (N_3222,N_622,N_1067);
nand U3223 (N_3223,N_632,N_1933);
nor U3224 (N_3224,N_343,N_915);
xor U3225 (N_3225,N_1522,N_1121);
and U3226 (N_3226,N_1211,N_885);
nand U3227 (N_3227,N_473,N_392);
and U3228 (N_3228,N_981,N_1349);
nand U3229 (N_3229,N_989,N_1003);
or U3230 (N_3230,N_616,N_1412);
nand U3231 (N_3231,N_315,N_665);
and U3232 (N_3232,N_398,N_716);
nand U3233 (N_3233,N_557,N_1607);
or U3234 (N_3234,N_1916,N_1763);
nand U3235 (N_3235,N_979,N_769);
and U3236 (N_3236,N_830,N_639);
or U3237 (N_3237,N_959,N_1058);
and U3238 (N_3238,N_1844,N_1805);
and U3239 (N_3239,N_1373,N_247);
and U3240 (N_3240,N_1846,N_1135);
nand U3241 (N_3241,N_702,N_301);
nor U3242 (N_3242,N_1203,N_1558);
nand U3243 (N_3243,N_565,N_412);
nor U3244 (N_3244,N_1827,N_915);
nor U3245 (N_3245,N_1533,N_1109);
nand U3246 (N_3246,N_721,N_594);
and U3247 (N_3247,N_102,N_1501);
or U3248 (N_3248,N_879,N_1696);
nand U3249 (N_3249,N_1448,N_541);
nor U3250 (N_3250,N_0,N_704);
and U3251 (N_3251,N_1662,N_974);
or U3252 (N_3252,N_5,N_1767);
nand U3253 (N_3253,N_1133,N_1405);
nor U3254 (N_3254,N_1894,N_70);
nand U3255 (N_3255,N_1648,N_493);
and U3256 (N_3256,N_278,N_1202);
nor U3257 (N_3257,N_310,N_1440);
nand U3258 (N_3258,N_749,N_624);
xnor U3259 (N_3259,N_506,N_795);
nor U3260 (N_3260,N_1676,N_112);
nand U3261 (N_3261,N_1127,N_558);
nand U3262 (N_3262,N_1966,N_202);
and U3263 (N_3263,N_268,N_848);
or U3264 (N_3264,N_1539,N_449);
nor U3265 (N_3265,N_1961,N_867);
nand U3266 (N_3266,N_1170,N_1237);
and U3267 (N_3267,N_231,N_1922);
nor U3268 (N_3268,N_1159,N_833);
or U3269 (N_3269,N_19,N_486);
nand U3270 (N_3270,N_140,N_950);
and U3271 (N_3271,N_80,N_1094);
or U3272 (N_3272,N_1589,N_1248);
and U3273 (N_3273,N_1279,N_1953);
xor U3274 (N_3274,N_936,N_789);
and U3275 (N_3275,N_1357,N_615);
and U3276 (N_3276,N_126,N_544);
xnor U3277 (N_3277,N_1396,N_1435);
xnor U3278 (N_3278,N_535,N_1431);
nor U3279 (N_3279,N_1188,N_1424);
nor U3280 (N_3280,N_639,N_1345);
or U3281 (N_3281,N_1909,N_1598);
nor U3282 (N_3282,N_1285,N_810);
or U3283 (N_3283,N_1097,N_1169);
or U3284 (N_3284,N_1132,N_865);
or U3285 (N_3285,N_499,N_1201);
nor U3286 (N_3286,N_1829,N_1329);
xnor U3287 (N_3287,N_80,N_1949);
and U3288 (N_3288,N_1701,N_54);
and U3289 (N_3289,N_611,N_633);
and U3290 (N_3290,N_630,N_1359);
nand U3291 (N_3291,N_918,N_814);
or U3292 (N_3292,N_905,N_574);
and U3293 (N_3293,N_789,N_613);
and U3294 (N_3294,N_637,N_1555);
xor U3295 (N_3295,N_578,N_18);
xor U3296 (N_3296,N_751,N_1810);
and U3297 (N_3297,N_1460,N_309);
nand U3298 (N_3298,N_1501,N_638);
or U3299 (N_3299,N_943,N_484);
or U3300 (N_3300,N_639,N_1168);
nand U3301 (N_3301,N_1595,N_1434);
nor U3302 (N_3302,N_1109,N_482);
or U3303 (N_3303,N_999,N_1355);
or U3304 (N_3304,N_400,N_1624);
or U3305 (N_3305,N_42,N_883);
or U3306 (N_3306,N_1065,N_1926);
nand U3307 (N_3307,N_90,N_294);
nor U3308 (N_3308,N_818,N_1165);
nor U3309 (N_3309,N_1292,N_810);
nand U3310 (N_3310,N_1939,N_1227);
or U3311 (N_3311,N_652,N_1047);
nor U3312 (N_3312,N_1933,N_848);
or U3313 (N_3313,N_896,N_805);
xor U3314 (N_3314,N_1647,N_585);
nor U3315 (N_3315,N_679,N_1562);
or U3316 (N_3316,N_1078,N_1563);
or U3317 (N_3317,N_322,N_1588);
and U3318 (N_3318,N_1776,N_1830);
nand U3319 (N_3319,N_146,N_24);
nand U3320 (N_3320,N_1014,N_246);
and U3321 (N_3321,N_95,N_377);
nand U3322 (N_3322,N_1053,N_790);
or U3323 (N_3323,N_259,N_1922);
and U3324 (N_3324,N_211,N_111);
and U3325 (N_3325,N_1559,N_1466);
and U3326 (N_3326,N_1271,N_645);
or U3327 (N_3327,N_1138,N_747);
and U3328 (N_3328,N_1773,N_484);
nand U3329 (N_3329,N_519,N_1766);
and U3330 (N_3330,N_1708,N_1502);
xor U3331 (N_3331,N_1943,N_861);
or U3332 (N_3332,N_416,N_886);
nor U3333 (N_3333,N_553,N_1965);
nand U3334 (N_3334,N_671,N_1755);
or U3335 (N_3335,N_1005,N_832);
xor U3336 (N_3336,N_583,N_1436);
or U3337 (N_3337,N_75,N_1526);
nor U3338 (N_3338,N_1606,N_1104);
nand U3339 (N_3339,N_1584,N_932);
and U3340 (N_3340,N_1288,N_222);
and U3341 (N_3341,N_1765,N_1269);
xnor U3342 (N_3342,N_1905,N_271);
nor U3343 (N_3343,N_1840,N_1049);
and U3344 (N_3344,N_809,N_858);
or U3345 (N_3345,N_108,N_802);
and U3346 (N_3346,N_1744,N_759);
nand U3347 (N_3347,N_1874,N_272);
or U3348 (N_3348,N_631,N_131);
and U3349 (N_3349,N_1646,N_505);
and U3350 (N_3350,N_1620,N_1114);
xor U3351 (N_3351,N_1904,N_583);
nor U3352 (N_3352,N_491,N_1697);
nand U3353 (N_3353,N_1772,N_902);
xnor U3354 (N_3354,N_1561,N_767);
xnor U3355 (N_3355,N_1510,N_1369);
or U3356 (N_3356,N_310,N_586);
and U3357 (N_3357,N_619,N_753);
and U3358 (N_3358,N_1442,N_724);
or U3359 (N_3359,N_833,N_1281);
nand U3360 (N_3360,N_1223,N_562);
nand U3361 (N_3361,N_399,N_650);
and U3362 (N_3362,N_1418,N_1579);
nor U3363 (N_3363,N_1106,N_1938);
or U3364 (N_3364,N_215,N_765);
nor U3365 (N_3365,N_518,N_914);
and U3366 (N_3366,N_167,N_719);
and U3367 (N_3367,N_1257,N_1577);
nor U3368 (N_3368,N_517,N_819);
and U3369 (N_3369,N_444,N_1020);
or U3370 (N_3370,N_884,N_628);
and U3371 (N_3371,N_612,N_251);
nor U3372 (N_3372,N_1162,N_263);
or U3373 (N_3373,N_1350,N_617);
or U3374 (N_3374,N_627,N_1617);
and U3375 (N_3375,N_732,N_474);
or U3376 (N_3376,N_1069,N_1382);
nor U3377 (N_3377,N_1191,N_1136);
nor U3378 (N_3378,N_1850,N_70);
and U3379 (N_3379,N_1271,N_88);
or U3380 (N_3380,N_1712,N_1120);
xnor U3381 (N_3381,N_1070,N_1939);
nand U3382 (N_3382,N_312,N_625);
nand U3383 (N_3383,N_1420,N_1704);
nor U3384 (N_3384,N_1428,N_717);
or U3385 (N_3385,N_436,N_6);
xnor U3386 (N_3386,N_879,N_153);
nand U3387 (N_3387,N_1318,N_1248);
and U3388 (N_3388,N_1315,N_216);
nand U3389 (N_3389,N_856,N_216);
xnor U3390 (N_3390,N_654,N_4);
nand U3391 (N_3391,N_1966,N_997);
or U3392 (N_3392,N_884,N_968);
xor U3393 (N_3393,N_1857,N_1273);
or U3394 (N_3394,N_962,N_1602);
xor U3395 (N_3395,N_529,N_1456);
nor U3396 (N_3396,N_647,N_1907);
nand U3397 (N_3397,N_963,N_68);
and U3398 (N_3398,N_821,N_533);
nand U3399 (N_3399,N_181,N_478);
or U3400 (N_3400,N_1962,N_316);
nor U3401 (N_3401,N_1123,N_772);
or U3402 (N_3402,N_1676,N_436);
nor U3403 (N_3403,N_127,N_1450);
and U3404 (N_3404,N_1160,N_1647);
nand U3405 (N_3405,N_1939,N_1464);
and U3406 (N_3406,N_852,N_1008);
nor U3407 (N_3407,N_1367,N_1596);
and U3408 (N_3408,N_1251,N_1599);
or U3409 (N_3409,N_1514,N_761);
and U3410 (N_3410,N_952,N_631);
xnor U3411 (N_3411,N_485,N_1645);
xor U3412 (N_3412,N_1377,N_478);
nand U3413 (N_3413,N_359,N_1369);
or U3414 (N_3414,N_619,N_613);
nand U3415 (N_3415,N_1396,N_124);
and U3416 (N_3416,N_1053,N_732);
nor U3417 (N_3417,N_1860,N_1924);
xnor U3418 (N_3418,N_1059,N_356);
xnor U3419 (N_3419,N_1003,N_1421);
nor U3420 (N_3420,N_869,N_35);
nand U3421 (N_3421,N_990,N_1712);
nor U3422 (N_3422,N_1893,N_1125);
nor U3423 (N_3423,N_1042,N_1206);
nand U3424 (N_3424,N_211,N_1965);
and U3425 (N_3425,N_437,N_1175);
nand U3426 (N_3426,N_1249,N_1317);
nor U3427 (N_3427,N_77,N_1333);
nor U3428 (N_3428,N_1494,N_912);
nor U3429 (N_3429,N_1979,N_1681);
nor U3430 (N_3430,N_1241,N_509);
nand U3431 (N_3431,N_1159,N_1021);
and U3432 (N_3432,N_1962,N_1067);
nor U3433 (N_3433,N_1699,N_290);
or U3434 (N_3434,N_786,N_1541);
or U3435 (N_3435,N_1744,N_254);
nand U3436 (N_3436,N_535,N_319);
xor U3437 (N_3437,N_398,N_6);
nand U3438 (N_3438,N_574,N_620);
nor U3439 (N_3439,N_120,N_1487);
nand U3440 (N_3440,N_1148,N_1222);
nand U3441 (N_3441,N_988,N_299);
or U3442 (N_3442,N_366,N_1700);
or U3443 (N_3443,N_1090,N_1925);
nand U3444 (N_3444,N_305,N_441);
nand U3445 (N_3445,N_578,N_1041);
or U3446 (N_3446,N_1626,N_805);
nand U3447 (N_3447,N_517,N_151);
nand U3448 (N_3448,N_118,N_721);
and U3449 (N_3449,N_1854,N_653);
or U3450 (N_3450,N_1152,N_1819);
nor U3451 (N_3451,N_810,N_1887);
or U3452 (N_3452,N_1553,N_1154);
nand U3453 (N_3453,N_1719,N_186);
xor U3454 (N_3454,N_1920,N_526);
or U3455 (N_3455,N_1704,N_1599);
nor U3456 (N_3456,N_1537,N_1417);
or U3457 (N_3457,N_1334,N_1550);
nor U3458 (N_3458,N_1044,N_1131);
and U3459 (N_3459,N_900,N_1794);
nand U3460 (N_3460,N_1391,N_1116);
or U3461 (N_3461,N_176,N_141);
nand U3462 (N_3462,N_511,N_1574);
nand U3463 (N_3463,N_1487,N_338);
or U3464 (N_3464,N_1794,N_1453);
or U3465 (N_3465,N_597,N_1574);
and U3466 (N_3466,N_1636,N_1726);
nand U3467 (N_3467,N_185,N_8);
and U3468 (N_3468,N_1487,N_1932);
nor U3469 (N_3469,N_77,N_574);
nor U3470 (N_3470,N_1888,N_1531);
nand U3471 (N_3471,N_1745,N_812);
xor U3472 (N_3472,N_352,N_1959);
or U3473 (N_3473,N_365,N_1118);
nand U3474 (N_3474,N_940,N_1520);
or U3475 (N_3475,N_754,N_1832);
or U3476 (N_3476,N_756,N_1987);
xor U3477 (N_3477,N_385,N_1820);
and U3478 (N_3478,N_296,N_1466);
or U3479 (N_3479,N_248,N_1992);
nand U3480 (N_3480,N_782,N_407);
nand U3481 (N_3481,N_257,N_1515);
nand U3482 (N_3482,N_497,N_1972);
nor U3483 (N_3483,N_662,N_1648);
xor U3484 (N_3484,N_697,N_803);
and U3485 (N_3485,N_824,N_209);
xnor U3486 (N_3486,N_357,N_1665);
xor U3487 (N_3487,N_231,N_1628);
and U3488 (N_3488,N_706,N_1332);
and U3489 (N_3489,N_1944,N_940);
nor U3490 (N_3490,N_1081,N_171);
and U3491 (N_3491,N_718,N_1619);
and U3492 (N_3492,N_125,N_1195);
nand U3493 (N_3493,N_1734,N_1052);
or U3494 (N_3494,N_435,N_1598);
or U3495 (N_3495,N_1024,N_202);
xnor U3496 (N_3496,N_774,N_954);
nor U3497 (N_3497,N_1667,N_1827);
nor U3498 (N_3498,N_799,N_350);
nand U3499 (N_3499,N_883,N_1383);
nor U3500 (N_3500,N_1878,N_1287);
or U3501 (N_3501,N_1998,N_267);
or U3502 (N_3502,N_1849,N_78);
and U3503 (N_3503,N_657,N_1462);
and U3504 (N_3504,N_490,N_896);
and U3505 (N_3505,N_1696,N_481);
xnor U3506 (N_3506,N_1375,N_233);
or U3507 (N_3507,N_175,N_1208);
nand U3508 (N_3508,N_920,N_1846);
or U3509 (N_3509,N_1484,N_284);
nand U3510 (N_3510,N_961,N_552);
and U3511 (N_3511,N_1306,N_221);
and U3512 (N_3512,N_1598,N_1281);
and U3513 (N_3513,N_1720,N_711);
nand U3514 (N_3514,N_1638,N_1987);
nor U3515 (N_3515,N_1048,N_1574);
nor U3516 (N_3516,N_545,N_1807);
xor U3517 (N_3517,N_974,N_900);
and U3518 (N_3518,N_1238,N_862);
and U3519 (N_3519,N_1148,N_82);
and U3520 (N_3520,N_610,N_295);
nor U3521 (N_3521,N_554,N_1450);
and U3522 (N_3522,N_1032,N_1754);
or U3523 (N_3523,N_782,N_1096);
and U3524 (N_3524,N_1110,N_1737);
nor U3525 (N_3525,N_1199,N_344);
xor U3526 (N_3526,N_1394,N_377);
or U3527 (N_3527,N_1319,N_1306);
nor U3528 (N_3528,N_123,N_1937);
nand U3529 (N_3529,N_703,N_136);
xnor U3530 (N_3530,N_87,N_389);
nand U3531 (N_3531,N_1154,N_585);
and U3532 (N_3532,N_116,N_83);
and U3533 (N_3533,N_662,N_1834);
xnor U3534 (N_3534,N_337,N_353);
and U3535 (N_3535,N_1436,N_1755);
and U3536 (N_3536,N_123,N_1572);
nor U3537 (N_3537,N_1731,N_317);
and U3538 (N_3538,N_1375,N_1996);
or U3539 (N_3539,N_484,N_314);
or U3540 (N_3540,N_1650,N_1293);
nor U3541 (N_3541,N_1849,N_1488);
or U3542 (N_3542,N_192,N_1786);
and U3543 (N_3543,N_1841,N_33);
and U3544 (N_3544,N_276,N_615);
or U3545 (N_3545,N_857,N_368);
nor U3546 (N_3546,N_1030,N_1351);
nor U3547 (N_3547,N_1930,N_1585);
nand U3548 (N_3548,N_793,N_421);
or U3549 (N_3549,N_931,N_80);
or U3550 (N_3550,N_1692,N_1482);
and U3551 (N_3551,N_478,N_272);
and U3552 (N_3552,N_1906,N_1854);
nand U3553 (N_3553,N_1243,N_233);
xor U3554 (N_3554,N_1113,N_1171);
or U3555 (N_3555,N_243,N_45);
or U3556 (N_3556,N_649,N_1237);
or U3557 (N_3557,N_1334,N_710);
nand U3558 (N_3558,N_768,N_417);
nor U3559 (N_3559,N_187,N_65);
and U3560 (N_3560,N_1476,N_1841);
or U3561 (N_3561,N_283,N_1119);
and U3562 (N_3562,N_204,N_1987);
nor U3563 (N_3563,N_1834,N_1660);
and U3564 (N_3564,N_811,N_1622);
xnor U3565 (N_3565,N_922,N_1555);
and U3566 (N_3566,N_852,N_643);
or U3567 (N_3567,N_1946,N_441);
xnor U3568 (N_3568,N_928,N_764);
nand U3569 (N_3569,N_1647,N_855);
xnor U3570 (N_3570,N_534,N_1554);
xor U3571 (N_3571,N_785,N_687);
or U3572 (N_3572,N_939,N_629);
and U3573 (N_3573,N_1072,N_519);
and U3574 (N_3574,N_317,N_1428);
and U3575 (N_3575,N_448,N_1016);
nand U3576 (N_3576,N_850,N_96);
xor U3577 (N_3577,N_738,N_1724);
nand U3578 (N_3578,N_967,N_1797);
and U3579 (N_3579,N_722,N_283);
and U3580 (N_3580,N_1451,N_1577);
nor U3581 (N_3581,N_419,N_509);
nor U3582 (N_3582,N_739,N_1414);
and U3583 (N_3583,N_1209,N_199);
nand U3584 (N_3584,N_1628,N_1061);
and U3585 (N_3585,N_1836,N_1096);
and U3586 (N_3586,N_731,N_678);
nor U3587 (N_3587,N_283,N_1379);
xor U3588 (N_3588,N_1329,N_1992);
or U3589 (N_3589,N_1837,N_1290);
and U3590 (N_3590,N_561,N_1351);
nor U3591 (N_3591,N_466,N_1486);
or U3592 (N_3592,N_943,N_998);
nor U3593 (N_3593,N_237,N_1425);
and U3594 (N_3594,N_1470,N_260);
and U3595 (N_3595,N_1356,N_1054);
nor U3596 (N_3596,N_1763,N_515);
nor U3597 (N_3597,N_1018,N_34);
nand U3598 (N_3598,N_508,N_1550);
xor U3599 (N_3599,N_675,N_764);
nor U3600 (N_3600,N_824,N_1285);
nor U3601 (N_3601,N_1559,N_811);
nand U3602 (N_3602,N_1343,N_102);
or U3603 (N_3603,N_947,N_703);
nor U3604 (N_3604,N_59,N_1402);
xnor U3605 (N_3605,N_1629,N_1497);
nand U3606 (N_3606,N_751,N_1843);
nand U3607 (N_3607,N_858,N_324);
and U3608 (N_3608,N_1589,N_1066);
nor U3609 (N_3609,N_74,N_1930);
or U3610 (N_3610,N_1974,N_1270);
and U3611 (N_3611,N_640,N_370);
and U3612 (N_3612,N_1836,N_122);
nand U3613 (N_3613,N_82,N_334);
or U3614 (N_3614,N_393,N_1268);
or U3615 (N_3615,N_1892,N_1275);
and U3616 (N_3616,N_758,N_751);
and U3617 (N_3617,N_1541,N_700);
nand U3618 (N_3618,N_1191,N_1006);
nor U3619 (N_3619,N_1333,N_1578);
nand U3620 (N_3620,N_243,N_1733);
nand U3621 (N_3621,N_54,N_1637);
nand U3622 (N_3622,N_1052,N_1265);
or U3623 (N_3623,N_1267,N_1447);
nand U3624 (N_3624,N_62,N_1212);
nor U3625 (N_3625,N_1618,N_1384);
xor U3626 (N_3626,N_888,N_51);
nor U3627 (N_3627,N_1352,N_1928);
nand U3628 (N_3628,N_1308,N_1763);
nand U3629 (N_3629,N_1782,N_1795);
nor U3630 (N_3630,N_1478,N_1443);
nand U3631 (N_3631,N_1817,N_485);
or U3632 (N_3632,N_1058,N_1136);
nor U3633 (N_3633,N_1680,N_1512);
nor U3634 (N_3634,N_150,N_1630);
or U3635 (N_3635,N_297,N_1096);
or U3636 (N_3636,N_1389,N_906);
xnor U3637 (N_3637,N_1122,N_1962);
nor U3638 (N_3638,N_1388,N_299);
and U3639 (N_3639,N_1541,N_345);
and U3640 (N_3640,N_954,N_496);
and U3641 (N_3641,N_1339,N_978);
and U3642 (N_3642,N_1534,N_1612);
or U3643 (N_3643,N_972,N_768);
or U3644 (N_3644,N_1167,N_729);
and U3645 (N_3645,N_19,N_279);
xor U3646 (N_3646,N_1242,N_1487);
and U3647 (N_3647,N_1724,N_779);
or U3648 (N_3648,N_859,N_1501);
and U3649 (N_3649,N_1180,N_1277);
and U3650 (N_3650,N_467,N_513);
and U3651 (N_3651,N_1837,N_235);
nand U3652 (N_3652,N_544,N_241);
xnor U3653 (N_3653,N_1030,N_272);
and U3654 (N_3654,N_1836,N_1797);
and U3655 (N_3655,N_1461,N_1849);
nor U3656 (N_3656,N_1215,N_1810);
xor U3657 (N_3657,N_1513,N_1371);
nor U3658 (N_3658,N_129,N_1847);
or U3659 (N_3659,N_1934,N_650);
nand U3660 (N_3660,N_1732,N_337);
or U3661 (N_3661,N_1377,N_635);
nand U3662 (N_3662,N_1775,N_1478);
and U3663 (N_3663,N_855,N_634);
nand U3664 (N_3664,N_1087,N_1483);
and U3665 (N_3665,N_1013,N_650);
or U3666 (N_3666,N_365,N_1864);
or U3667 (N_3667,N_410,N_1835);
and U3668 (N_3668,N_1313,N_32);
nor U3669 (N_3669,N_398,N_720);
xor U3670 (N_3670,N_204,N_974);
or U3671 (N_3671,N_1492,N_1062);
or U3672 (N_3672,N_516,N_506);
nand U3673 (N_3673,N_529,N_375);
and U3674 (N_3674,N_1147,N_1542);
nand U3675 (N_3675,N_1778,N_768);
xnor U3676 (N_3676,N_1678,N_999);
or U3677 (N_3677,N_809,N_1721);
nand U3678 (N_3678,N_1692,N_1045);
nor U3679 (N_3679,N_977,N_1859);
and U3680 (N_3680,N_897,N_453);
or U3681 (N_3681,N_380,N_1237);
nand U3682 (N_3682,N_1301,N_17);
or U3683 (N_3683,N_1957,N_284);
or U3684 (N_3684,N_1462,N_1103);
and U3685 (N_3685,N_1290,N_1790);
nor U3686 (N_3686,N_1860,N_1513);
nand U3687 (N_3687,N_41,N_210);
nand U3688 (N_3688,N_1269,N_1510);
and U3689 (N_3689,N_1997,N_1049);
and U3690 (N_3690,N_1258,N_1897);
nor U3691 (N_3691,N_640,N_1936);
nor U3692 (N_3692,N_1253,N_261);
and U3693 (N_3693,N_1633,N_57);
xor U3694 (N_3694,N_719,N_266);
and U3695 (N_3695,N_1804,N_417);
or U3696 (N_3696,N_452,N_1242);
or U3697 (N_3697,N_658,N_858);
or U3698 (N_3698,N_839,N_1810);
or U3699 (N_3699,N_1663,N_1118);
nor U3700 (N_3700,N_465,N_375);
xnor U3701 (N_3701,N_783,N_558);
xor U3702 (N_3702,N_366,N_1191);
and U3703 (N_3703,N_644,N_276);
and U3704 (N_3704,N_1910,N_814);
or U3705 (N_3705,N_234,N_30);
nand U3706 (N_3706,N_129,N_1554);
or U3707 (N_3707,N_919,N_799);
nand U3708 (N_3708,N_266,N_731);
nor U3709 (N_3709,N_1127,N_481);
nor U3710 (N_3710,N_380,N_1076);
nand U3711 (N_3711,N_557,N_871);
nand U3712 (N_3712,N_845,N_1929);
and U3713 (N_3713,N_1872,N_1921);
nor U3714 (N_3714,N_118,N_241);
or U3715 (N_3715,N_1463,N_1603);
and U3716 (N_3716,N_1054,N_55);
xor U3717 (N_3717,N_303,N_1914);
nor U3718 (N_3718,N_907,N_1725);
nand U3719 (N_3719,N_503,N_1147);
nand U3720 (N_3720,N_1475,N_21);
xor U3721 (N_3721,N_220,N_1507);
or U3722 (N_3722,N_1703,N_1419);
xor U3723 (N_3723,N_977,N_476);
nand U3724 (N_3724,N_1691,N_488);
and U3725 (N_3725,N_139,N_143);
nor U3726 (N_3726,N_609,N_691);
or U3727 (N_3727,N_1921,N_188);
nor U3728 (N_3728,N_1955,N_1903);
or U3729 (N_3729,N_1300,N_711);
and U3730 (N_3730,N_564,N_654);
and U3731 (N_3731,N_1716,N_529);
and U3732 (N_3732,N_1970,N_615);
or U3733 (N_3733,N_195,N_190);
or U3734 (N_3734,N_995,N_1568);
nor U3735 (N_3735,N_561,N_566);
nand U3736 (N_3736,N_1209,N_759);
or U3737 (N_3737,N_1963,N_893);
xor U3738 (N_3738,N_1644,N_1206);
or U3739 (N_3739,N_1768,N_1759);
nand U3740 (N_3740,N_1399,N_879);
and U3741 (N_3741,N_989,N_773);
and U3742 (N_3742,N_883,N_67);
nor U3743 (N_3743,N_1313,N_1049);
nor U3744 (N_3744,N_1052,N_220);
or U3745 (N_3745,N_1614,N_189);
and U3746 (N_3746,N_1901,N_1273);
nand U3747 (N_3747,N_1417,N_1637);
and U3748 (N_3748,N_905,N_662);
and U3749 (N_3749,N_1545,N_901);
xnor U3750 (N_3750,N_681,N_805);
nor U3751 (N_3751,N_1068,N_1493);
and U3752 (N_3752,N_1146,N_1672);
nand U3753 (N_3753,N_575,N_177);
xnor U3754 (N_3754,N_748,N_239);
or U3755 (N_3755,N_236,N_188);
nand U3756 (N_3756,N_1004,N_1347);
and U3757 (N_3757,N_1631,N_1470);
nand U3758 (N_3758,N_1986,N_958);
xor U3759 (N_3759,N_1242,N_16);
or U3760 (N_3760,N_919,N_1424);
nand U3761 (N_3761,N_1816,N_1222);
and U3762 (N_3762,N_403,N_125);
nor U3763 (N_3763,N_1598,N_1406);
xor U3764 (N_3764,N_1523,N_1613);
and U3765 (N_3765,N_1122,N_919);
and U3766 (N_3766,N_1779,N_1223);
xnor U3767 (N_3767,N_734,N_319);
and U3768 (N_3768,N_444,N_1662);
or U3769 (N_3769,N_539,N_1748);
nand U3770 (N_3770,N_822,N_872);
nand U3771 (N_3771,N_1526,N_683);
or U3772 (N_3772,N_1138,N_114);
nand U3773 (N_3773,N_458,N_1641);
nand U3774 (N_3774,N_1356,N_389);
or U3775 (N_3775,N_1885,N_1108);
nor U3776 (N_3776,N_1008,N_81);
xor U3777 (N_3777,N_362,N_1019);
xnor U3778 (N_3778,N_1846,N_1836);
and U3779 (N_3779,N_149,N_312);
or U3780 (N_3780,N_83,N_1790);
and U3781 (N_3781,N_1581,N_1459);
xor U3782 (N_3782,N_1767,N_1108);
nor U3783 (N_3783,N_1459,N_56);
nand U3784 (N_3784,N_887,N_32);
nor U3785 (N_3785,N_1226,N_1442);
nor U3786 (N_3786,N_753,N_1217);
nor U3787 (N_3787,N_1160,N_1507);
nand U3788 (N_3788,N_1742,N_470);
or U3789 (N_3789,N_414,N_473);
or U3790 (N_3790,N_1275,N_257);
nor U3791 (N_3791,N_1824,N_1169);
nor U3792 (N_3792,N_1221,N_1045);
nor U3793 (N_3793,N_1102,N_469);
or U3794 (N_3794,N_1355,N_912);
nand U3795 (N_3795,N_1204,N_930);
and U3796 (N_3796,N_508,N_1784);
nor U3797 (N_3797,N_1985,N_1170);
nand U3798 (N_3798,N_1271,N_651);
nor U3799 (N_3799,N_1858,N_144);
or U3800 (N_3800,N_0,N_1922);
nand U3801 (N_3801,N_1697,N_1940);
nor U3802 (N_3802,N_1407,N_346);
nor U3803 (N_3803,N_1325,N_1753);
nand U3804 (N_3804,N_1652,N_379);
and U3805 (N_3805,N_524,N_320);
nor U3806 (N_3806,N_5,N_237);
and U3807 (N_3807,N_240,N_1022);
and U3808 (N_3808,N_1276,N_908);
xor U3809 (N_3809,N_491,N_880);
nand U3810 (N_3810,N_869,N_1480);
nor U3811 (N_3811,N_1376,N_955);
and U3812 (N_3812,N_1641,N_333);
xnor U3813 (N_3813,N_1306,N_495);
or U3814 (N_3814,N_299,N_400);
and U3815 (N_3815,N_1487,N_1578);
and U3816 (N_3816,N_565,N_17);
nand U3817 (N_3817,N_488,N_1993);
or U3818 (N_3818,N_1168,N_17);
xor U3819 (N_3819,N_170,N_910);
and U3820 (N_3820,N_832,N_116);
and U3821 (N_3821,N_60,N_1399);
nand U3822 (N_3822,N_1579,N_277);
xor U3823 (N_3823,N_1684,N_1941);
nand U3824 (N_3824,N_1834,N_247);
and U3825 (N_3825,N_1460,N_555);
nor U3826 (N_3826,N_35,N_569);
and U3827 (N_3827,N_1685,N_259);
or U3828 (N_3828,N_449,N_1286);
xor U3829 (N_3829,N_1947,N_212);
or U3830 (N_3830,N_498,N_1429);
and U3831 (N_3831,N_976,N_1658);
and U3832 (N_3832,N_1389,N_927);
and U3833 (N_3833,N_1060,N_1839);
or U3834 (N_3834,N_447,N_1370);
and U3835 (N_3835,N_664,N_1673);
nand U3836 (N_3836,N_1668,N_242);
nor U3837 (N_3837,N_1448,N_714);
nor U3838 (N_3838,N_1771,N_1667);
and U3839 (N_3839,N_1165,N_1112);
xnor U3840 (N_3840,N_263,N_1693);
or U3841 (N_3841,N_1081,N_1351);
and U3842 (N_3842,N_1621,N_1602);
and U3843 (N_3843,N_1941,N_995);
nor U3844 (N_3844,N_632,N_64);
or U3845 (N_3845,N_322,N_586);
xnor U3846 (N_3846,N_553,N_1558);
nand U3847 (N_3847,N_256,N_597);
nor U3848 (N_3848,N_1332,N_83);
nand U3849 (N_3849,N_1292,N_976);
nand U3850 (N_3850,N_1843,N_367);
nor U3851 (N_3851,N_1642,N_688);
nor U3852 (N_3852,N_1139,N_910);
nor U3853 (N_3853,N_36,N_1123);
nor U3854 (N_3854,N_1663,N_21);
or U3855 (N_3855,N_1483,N_1577);
and U3856 (N_3856,N_505,N_789);
or U3857 (N_3857,N_1157,N_1745);
nor U3858 (N_3858,N_1024,N_440);
and U3859 (N_3859,N_323,N_1733);
and U3860 (N_3860,N_1786,N_993);
or U3861 (N_3861,N_1025,N_1836);
xor U3862 (N_3862,N_1556,N_416);
nor U3863 (N_3863,N_1579,N_592);
xor U3864 (N_3864,N_1487,N_1485);
nor U3865 (N_3865,N_218,N_1033);
nand U3866 (N_3866,N_302,N_893);
and U3867 (N_3867,N_640,N_942);
nand U3868 (N_3868,N_1119,N_1919);
nor U3869 (N_3869,N_821,N_1225);
or U3870 (N_3870,N_633,N_169);
and U3871 (N_3871,N_1033,N_1612);
nor U3872 (N_3872,N_1167,N_735);
nor U3873 (N_3873,N_982,N_1513);
nand U3874 (N_3874,N_1815,N_682);
nand U3875 (N_3875,N_899,N_1863);
and U3876 (N_3876,N_1369,N_1392);
xor U3877 (N_3877,N_1499,N_157);
nand U3878 (N_3878,N_1975,N_1578);
nor U3879 (N_3879,N_1154,N_784);
nand U3880 (N_3880,N_653,N_1303);
or U3881 (N_3881,N_990,N_1825);
nor U3882 (N_3882,N_662,N_1606);
xnor U3883 (N_3883,N_1678,N_1037);
nand U3884 (N_3884,N_1952,N_298);
nor U3885 (N_3885,N_1728,N_1150);
or U3886 (N_3886,N_1623,N_1501);
nor U3887 (N_3887,N_1631,N_1657);
nand U3888 (N_3888,N_1157,N_672);
nand U3889 (N_3889,N_1596,N_1998);
nand U3890 (N_3890,N_1255,N_730);
xnor U3891 (N_3891,N_1779,N_1320);
nor U3892 (N_3892,N_127,N_681);
or U3893 (N_3893,N_1591,N_180);
and U3894 (N_3894,N_941,N_1178);
and U3895 (N_3895,N_1000,N_728);
nand U3896 (N_3896,N_1429,N_204);
and U3897 (N_3897,N_1855,N_1954);
nor U3898 (N_3898,N_1216,N_1342);
nor U3899 (N_3899,N_1071,N_1801);
and U3900 (N_3900,N_1520,N_439);
nor U3901 (N_3901,N_331,N_1248);
nor U3902 (N_3902,N_278,N_1653);
nor U3903 (N_3903,N_1025,N_163);
nand U3904 (N_3904,N_280,N_398);
and U3905 (N_3905,N_1373,N_1949);
and U3906 (N_3906,N_151,N_212);
nand U3907 (N_3907,N_1100,N_758);
xnor U3908 (N_3908,N_215,N_527);
and U3909 (N_3909,N_1074,N_371);
nand U3910 (N_3910,N_1734,N_942);
nor U3911 (N_3911,N_386,N_1930);
nand U3912 (N_3912,N_1117,N_1828);
or U3913 (N_3913,N_1272,N_1408);
nor U3914 (N_3914,N_392,N_763);
or U3915 (N_3915,N_1502,N_461);
nor U3916 (N_3916,N_594,N_895);
and U3917 (N_3917,N_939,N_756);
and U3918 (N_3918,N_1662,N_1152);
and U3919 (N_3919,N_477,N_986);
or U3920 (N_3920,N_194,N_852);
xor U3921 (N_3921,N_1053,N_1345);
and U3922 (N_3922,N_1570,N_309);
nand U3923 (N_3923,N_1699,N_763);
xnor U3924 (N_3924,N_433,N_583);
nand U3925 (N_3925,N_1734,N_224);
and U3926 (N_3926,N_1171,N_1275);
nand U3927 (N_3927,N_997,N_722);
nor U3928 (N_3928,N_151,N_1163);
nand U3929 (N_3929,N_290,N_322);
or U3930 (N_3930,N_1420,N_1310);
nor U3931 (N_3931,N_1249,N_1513);
or U3932 (N_3932,N_1245,N_30);
nor U3933 (N_3933,N_1927,N_840);
and U3934 (N_3934,N_170,N_316);
nand U3935 (N_3935,N_1731,N_1106);
and U3936 (N_3936,N_173,N_695);
nand U3937 (N_3937,N_1817,N_231);
nor U3938 (N_3938,N_828,N_867);
nor U3939 (N_3939,N_649,N_1156);
or U3940 (N_3940,N_1663,N_534);
nand U3941 (N_3941,N_1874,N_66);
nor U3942 (N_3942,N_1432,N_764);
nor U3943 (N_3943,N_1783,N_1684);
xnor U3944 (N_3944,N_737,N_920);
or U3945 (N_3945,N_946,N_1699);
nor U3946 (N_3946,N_906,N_531);
nor U3947 (N_3947,N_48,N_350);
and U3948 (N_3948,N_654,N_265);
xnor U3949 (N_3949,N_4,N_1829);
nor U3950 (N_3950,N_1305,N_1378);
nand U3951 (N_3951,N_795,N_1143);
nand U3952 (N_3952,N_154,N_1566);
or U3953 (N_3953,N_693,N_1208);
nor U3954 (N_3954,N_1507,N_1008);
nand U3955 (N_3955,N_481,N_1974);
xnor U3956 (N_3956,N_155,N_747);
or U3957 (N_3957,N_1688,N_1744);
nor U3958 (N_3958,N_1790,N_1386);
and U3959 (N_3959,N_1381,N_863);
and U3960 (N_3960,N_352,N_836);
nor U3961 (N_3961,N_1002,N_415);
or U3962 (N_3962,N_517,N_364);
or U3963 (N_3963,N_1576,N_107);
or U3964 (N_3964,N_1501,N_443);
nand U3965 (N_3965,N_2,N_1420);
xor U3966 (N_3966,N_1083,N_1515);
nand U3967 (N_3967,N_337,N_721);
nand U3968 (N_3968,N_1727,N_733);
and U3969 (N_3969,N_1176,N_795);
and U3970 (N_3970,N_276,N_396);
xnor U3971 (N_3971,N_1564,N_683);
or U3972 (N_3972,N_671,N_122);
nand U3973 (N_3973,N_245,N_539);
and U3974 (N_3974,N_105,N_634);
or U3975 (N_3975,N_1399,N_509);
and U3976 (N_3976,N_1321,N_227);
or U3977 (N_3977,N_1138,N_354);
nand U3978 (N_3978,N_1664,N_1412);
nor U3979 (N_3979,N_1893,N_937);
and U3980 (N_3980,N_1851,N_1697);
and U3981 (N_3981,N_574,N_694);
or U3982 (N_3982,N_1836,N_816);
nand U3983 (N_3983,N_227,N_1091);
nand U3984 (N_3984,N_465,N_338);
nand U3985 (N_3985,N_1499,N_108);
nand U3986 (N_3986,N_75,N_879);
nor U3987 (N_3987,N_1288,N_1581);
nand U3988 (N_3988,N_1590,N_775);
xnor U3989 (N_3989,N_549,N_191);
nor U3990 (N_3990,N_1382,N_523);
or U3991 (N_3991,N_696,N_30);
or U3992 (N_3992,N_778,N_57);
or U3993 (N_3993,N_182,N_115);
nand U3994 (N_3994,N_1105,N_1622);
nand U3995 (N_3995,N_1630,N_315);
or U3996 (N_3996,N_500,N_535);
nor U3997 (N_3997,N_671,N_922);
or U3998 (N_3998,N_377,N_1524);
or U3999 (N_3999,N_1501,N_325);
nor U4000 (N_4000,N_3283,N_3875);
and U4001 (N_4001,N_2960,N_2852);
xnor U4002 (N_4002,N_2439,N_3656);
nor U4003 (N_4003,N_3608,N_2004);
and U4004 (N_4004,N_3105,N_2118);
or U4005 (N_4005,N_3449,N_2443);
nor U4006 (N_4006,N_3243,N_3421);
nor U4007 (N_4007,N_3998,N_3521);
nor U4008 (N_4008,N_2766,N_3987);
nor U4009 (N_4009,N_2088,N_2661);
or U4010 (N_4010,N_2208,N_3353);
xnor U4011 (N_4011,N_3821,N_3325);
or U4012 (N_4012,N_2281,N_3742);
nor U4013 (N_4013,N_3358,N_2069);
and U4014 (N_4014,N_3642,N_2093);
or U4015 (N_4015,N_2372,N_2235);
xnor U4016 (N_4016,N_3307,N_2655);
xor U4017 (N_4017,N_2258,N_3462);
xnor U4018 (N_4018,N_3944,N_3126);
or U4019 (N_4019,N_3936,N_2108);
nor U4020 (N_4020,N_2212,N_3756);
nand U4021 (N_4021,N_3092,N_3037);
nand U4022 (N_4022,N_3593,N_2283);
nand U4023 (N_4023,N_2177,N_2652);
and U4024 (N_4024,N_2651,N_2286);
nand U4025 (N_4025,N_3945,N_2775);
or U4026 (N_4026,N_2566,N_2006);
or U4027 (N_4027,N_3925,N_3946);
nor U4028 (N_4028,N_3724,N_3226);
nand U4029 (N_4029,N_2115,N_3577);
nand U4030 (N_4030,N_3197,N_3695);
and U4031 (N_4031,N_2047,N_3453);
or U4032 (N_4032,N_3108,N_2748);
nor U4033 (N_4033,N_2071,N_2070);
or U4034 (N_4034,N_3069,N_2995);
nand U4035 (N_4035,N_2389,N_3511);
nand U4036 (N_4036,N_3788,N_2242);
or U4037 (N_4037,N_3324,N_3061);
nor U4038 (N_4038,N_3908,N_2180);
nor U4039 (N_4039,N_2739,N_3240);
nor U4040 (N_4040,N_2464,N_2928);
nor U4041 (N_4041,N_3560,N_2440);
nor U4042 (N_4042,N_2476,N_3774);
or U4043 (N_4043,N_3904,N_2428);
or U4044 (N_4044,N_2862,N_2947);
nand U4045 (N_4045,N_2777,N_3464);
or U4046 (N_4046,N_2379,N_2012);
and U4047 (N_4047,N_3293,N_2229);
and U4048 (N_4048,N_2854,N_2020);
nor U4049 (N_4049,N_2581,N_2972);
or U4050 (N_4050,N_2203,N_3305);
nand U4051 (N_4051,N_2137,N_3991);
or U4052 (N_4052,N_2030,N_2847);
or U4053 (N_4053,N_3550,N_3207);
xnor U4054 (N_4054,N_2261,N_3984);
xor U4055 (N_4055,N_2446,N_3344);
xor U4056 (N_4056,N_2523,N_2551);
nand U4057 (N_4057,N_2561,N_2684);
nor U4058 (N_4058,N_3536,N_3627);
or U4059 (N_4059,N_2239,N_3191);
xnor U4060 (N_4060,N_3159,N_3481);
or U4061 (N_4061,N_2291,N_3466);
and U4062 (N_4062,N_2448,N_2410);
nand U4063 (N_4063,N_3186,N_3120);
and U4064 (N_4064,N_3757,N_3165);
nor U4065 (N_4065,N_3856,N_2654);
or U4066 (N_4066,N_3204,N_3628);
or U4067 (N_4067,N_2259,N_3026);
nand U4068 (N_4068,N_3149,N_3429);
nand U4069 (N_4069,N_3030,N_3490);
nor U4070 (N_4070,N_2250,N_2631);
xnor U4071 (N_4071,N_3672,N_2934);
nor U4072 (N_4072,N_2290,N_2043);
or U4073 (N_4073,N_3712,N_2929);
and U4074 (N_4074,N_3430,N_3309);
and U4075 (N_4075,N_3488,N_2569);
and U4076 (N_4076,N_2393,N_2185);
and U4077 (N_4077,N_2016,N_2577);
and U4078 (N_4078,N_3110,N_2114);
or U4079 (N_4079,N_2041,N_3295);
xnor U4080 (N_4080,N_3340,N_3096);
nor U4081 (N_4081,N_2754,N_3112);
nand U4082 (N_4082,N_3826,N_2207);
nand U4083 (N_4083,N_3799,N_2697);
and U4084 (N_4084,N_2518,N_3732);
xor U4085 (N_4085,N_3103,N_3715);
or U4086 (N_4086,N_3828,N_2075);
xor U4087 (N_4087,N_2447,N_3257);
nand U4088 (N_4088,N_3919,N_3836);
nand U4089 (N_4089,N_3569,N_2142);
or U4090 (N_4090,N_2001,N_2026);
xnor U4091 (N_4091,N_2877,N_3993);
nor U4092 (N_4092,N_3179,N_3044);
or U4093 (N_4093,N_3900,N_2462);
or U4094 (N_4094,N_2723,N_2365);
or U4095 (N_4095,N_3534,N_3510);
nor U4096 (N_4096,N_3762,N_2730);
nand U4097 (N_4097,N_2780,N_3468);
or U4098 (N_4098,N_2420,N_2715);
or U4099 (N_4099,N_3530,N_3520);
nor U4100 (N_4100,N_2138,N_2818);
and U4101 (N_4101,N_2712,N_3576);
and U4102 (N_4102,N_2935,N_2418);
and U4103 (N_4103,N_2441,N_3248);
xor U4104 (N_4104,N_3002,N_3291);
or U4105 (N_4105,N_3880,N_3425);
nor U4106 (N_4106,N_3956,N_3053);
nor U4107 (N_4107,N_3411,N_3010);
xnor U4108 (N_4108,N_2366,N_3460);
and U4109 (N_4109,N_2473,N_3995);
and U4110 (N_4110,N_2053,N_3189);
and U4111 (N_4111,N_3977,N_3845);
or U4112 (N_4112,N_3773,N_3540);
nand U4113 (N_4113,N_3161,N_3516);
nor U4114 (N_4114,N_2845,N_3583);
or U4115 (N_4115,N_3461,N_3673);
nand U4116 (N_4116,N_2155,N_2857);
or U4117 (N_4117,N_3615,N_2424);
nor U4118 (N_4118,N_2284,N_3194);
nand U4119 (N_4119,N_2753,N_3048);
and U4120 (N_4120,N_3643,N_3780);
and U4121 (N_4121,N_2668,N_3062);
nand U4122 (N_4122,N_3391,N_2160);
nand U4123 (N_4123,N_3087,N_2653);
and U4124 (N_4124,N_3630,N_3999);
nor U4125 (N_4125,N_2762,N_2450);
nand U4126 (N_4126,N_3174,N_2222);
nand U4127 (N_4127,N_2343,N_2918);
nor U4128 (N_4128,N_3227,N_2367);
nor U4129 (N_4129,N_2179,N_3035);
nand U4130 (N_4130,N_3491,N_3851);
and U4131 (N_4131,N_2451,N_3806);
or U4132 (N_4132,N_3365,N_3965);
and U4133 (N_4133,N_2205,N_2911);
or U4134 (N_4134,N_2033,N_2336);
xnor U4135 (N_4135,N_2216,N_2621);
or U4136 (N_4136,N_2681,N_2732);
or U4137 (N_4137,N_3199,N_2036);
nand U4138 (N_4138,N_3524,N_2781);
nand U4139 (N_4139,N_3299,N_3041);
and U4140 (N_4140,N_3146,N_3758);
nand U4141 (N_4141,N_2545,N_3704);
nand U4142 (N_4142,N_3888,N_2072);
nand U4143 (N_4143,N_2568,N_2397);
xor U4144 (N_4144,N_2804,N_2570);
or U4145 (N_4145,N_3924,N_3273);
and U4146 (N_4146,N_3156,N_3417);
nor U4147 (N_4147,N_3316,N_2198);
nor U4148 (N_4148,N_2884,N_3013);
nor U4149 (N_4149,N_3388,N_3371);
or U4150 (N_4150,N_3022,N_3487);
and U4151 (N_4151,N_3731,N_2442);
or U4152 (N_4152,N_2629,N_3889);
xor U4153 (N_4153,N_2988,N_3746);
nor U4154 (N_4154,N_2735,N_3675);
xor U4155 (N_4155,N_2294,N_2802);
nor U4156 (N_4156,N_3831,N_3260);
nand U4157 (N_4157,N_3117,N_3394);
xnor U4158 (N_4158,N_3119,N_3431);
or U4159 (N_4159,N_2392,N_3896);
nor U4160 (N_4160,N_3726,N_3887);
or U4161 (N_4161,N_2484,N_3741);
and U4162 (N_4162,N_2694,N_3616);
or U4163 (N_4163,N_3548,N_3378);
xnor U4164 (N_4164,N_3346,N_3021);
nand U4165 (N_4165,N_3162,N_2806);
nand U4166 (N_4166,N_2508,N_3674);
nand U4167 (N_4167,N_2676,N_2463);
xnor U4168 (N_4168,N_3469,N_2076);
nor U4169 (N_4169,N_2002,N_3983);
and U4170 (N_4170,N_3533,N_2387);
or U4171 (N_4171,N_3529,N_3747);
nand U4172 (N_4172,N_3444,N_3658);
nand U4173 (N_4173,N_2201,N_2940);
nand U4174 (N_4174,N_2337,N_2872);
or U4175 (N_4175,N_2547,N_2202);
nand U4176 (N_4176,N_2639,N_2117);
and U4177 (N_4177,N_2840,N_3566);
and U4178 (N_4178,N_2050,N_2223);
nand U4179 (N_4179,N_3404,N_3218);
or U4180 (N_4180,N_3640,N_3122);
and U4181 (N_4181,N_2221,N_2713);
and U4182 (N_4182,N_3585,N_3646);
or U4183 (N_4183,N_2412,N_3623);
nor U4184 (N_4184,N_2782,N_2326);
nand U4185 (N_4185,N_3793,N_2526);
and U4186 (N_4186,N_2161,N_3660);
nor U4187 (N_4187,N_2186,N_2495);
nor U4188 (N_4188,N_3125,N_2218);
and U4189 (N_4189,N_3150,N_2328);
or U4190 (N_4190,N_2738,N_2452);
nand U4191 (N_4191,N_2437,N_3805);
nand U4192 (N_4192,N_3023,N_2747);
or U4193 (N_4193,N_3154,N_3538);
nand U4194 (N_4194,N_3800,N_2822);
or U4195 (N_4195,N_2896,N_2571);
nand U4196 (N_4196,N_3937,N_3663);
nand U4197 (N_4197,N_3060,N_2292);
nand U4198 (N_4198,N_3228,N_3361);
or U4199 (N_4199,N_3933,N_2932);
nor U4200 (N_4200,N_3101,N_3072);
nor U4201 (N_4201,N_2612,N_3236);
or U4202 (N_4202,N_3867,N_3434);
nand U4203 (N_4203,N_3779,N_3068);
nor U4204 (N_4204,N_3824,N_3230);
nor U4205 (N_4205,N_2910,N_3745);
nor U4206 (N_4206,N_3959,N_3819);
or U4207 (N_4207,N_3850,N_3258);
nor U4208 (N_4208,N_2238,N_2345);
nor U4209 (N_4209,N_2482,N_3990);
and U4210 (N_4210,N_2882,N_2425);
and U4211 (N_4211,N_3523,N_2725);
nor U4212 (N_4212,N_2321,N_2266);
nor U4213 (N_4213,N_2987,N_2111);
and U4214 (N_4214,N_2426,N_2542);
or U4215 (N_4215,N_3211,N_3437);
nor U4216 (N_4216,N_2469,N_2206);
nand U4217 (N_4217,N_3234,N_3853);
nor U4218 (N_4218,N_3222,N_3383);
or U4219 (N_4219,N_3213,N_2962);
nand U4220 (N_4220,N_2106,N_3225);
xor U4221 (N_4221,N_2512,N_2151);
and U4222 (N_4222,N_2431,N_3129);
and U4223 (N_4223,N_2623,N_2788);
nor U4224 (N_4224,N_2973,N_2092);
nor U4225 (N_4225,N_3954,N_3907);
nor U4226 (N_4226,N_2900,N_3329);
nor U4227 (N_4227,N_2130,N_3484);
and U4228 (N_4228,N_3242,N_3501);
and U4229 (N_4229,N_2383,N_3892);
nand U4230 (N_4230,N_3972,N_2538);
nor U4231 (N_4231,N_2491,N_2786);
and U4232 (N_4232,N_2699,N_2922);
nor U4233 (N_4233,N_2164,N_2855);
nand U4234 (N_4234,N_2646,N_3849);
or U4235 (N_4235,N_2253,N_3514);
and U4236 (N_4236,N_2187,N_3190);
and U4237 (N_4237,N_2722,N_3337);
or U4238 (N_4238,N_3463,N_3333);
nand U4239 (N_4239,N_3679,N_3609);
nand U4240 (N_4240,N_3351,N_3564);
nor U4241 (N_4241,N_3852,N_3091);
or U4242 (N_4242,N_3376,N_2307);
nor U4243 (N_4243,N_2673,N_2376);
and U4244 (N_4244,N_2023,N_2596);
nand U4245 (N_4245,N_3178,N_2524);
xor U4246 (N_4246,N_2773,N_2658);
xnor U4247 (N_4247,N_2247,N_2056);
nor U4248 (N_4248,N_2578,N_2487);
nor U4249 (N_4249,N_2841,N_3281);
nand U4250 (N_4250,N_2790,N_2772);
xor U4251 (N_4251,N_2955,N_2992);
nor U4252 (N_4252,N_2468,N_2087);
or U4253 (N_4253,N_2683,N_2795);
xnor U4254 (N_4254,N_3176,N_3531);
nand U4255 (N_4255,N_3350,N_3102);
or U4256 (N_4256,N_3345,N_2957);
xor U4257 (N_4257,N_3767,N_3251);
nand U4258 (N_4258,N_3175,N_3541);
and U4259 (N_4259,N_2249,N_3360);
nor U4260 (N_4260,N_2996,N_2246);
nor U4261 (N_4261,N_2488,N_2306);
and U4262 (N_4262,N_2776,N_3668);
and U4263 (N_4263,N_2920,N_2527);
nor U4264 (N_4264,N_3539,N_3625);
and U4265 (N_4265,N_3277,N_2403);
nor U4266 (N_4266,N_2685,N_3571);
or U4267 (N_4267,N_2436,N_2904);
xnor U4268 (N_4268,N_3310,N_2613);
or U4269 (N_4269,N_3144,N_3844);
or U4270 (N_4270,N_2836,N_3137);
nand U4271 (N_4271,N_2969,N_2324);
or U4272 (N_4272,N_3607,N_3064);
nor U4273 (N_4273,N_2583,N_3389);
nor U4274 (N_4274,N_3155,N_2793);
nor U4275 (N_4275,N_3858,N_2391);
nor U4276 (N_4276,N_2984,N_3184);
or U4277 (N_4277,N_2099,N_3777);
or U4278 (N_4278,N_3147,N_2849);
xnor U4279 (N_4279,N_3294,N_2686);
nand U4280 (N_4280,N_2312,N_2770);
or U4281 (N_4281,N_3339,N_2815);
and U4282 (N_4282,N_3470,N_2758);
nand U4283 (N_4283,N_2273,N_3879);
nand U4284 (N_4284,N_2693,N_2368);
nand U4285 (N_4285,N_2913,N_3089);
or U4286 (N_4286,N_2122,N_3635);
or U4287 (N_4287,N_2774,N_3677);
nor U4288 (N_4288,N_2975,N_3133);
and U4289 (N_4289,N_2251,N_3413);
nand U4290 (N_4290,N_2347,N_3323);
and U4291 (N_4291,N_2921,N_2267);
and U4292 (N_4292,N_2690,N_3574);
and U4293 (N_4293,N_3676,N_2978);
nor U4294 (N_4294,N_2131,N_2977);
and U4295 (N_4295,N_3503,N_3870);
nor U4296 (N_4296,N_3986,N_3580);
nor U4297 (N_4297,N_2744,N_3405);
and U4298 (N_4298,N_3220,N_2217);
or U4299 (N_4299,N_3597,N_3423);
nand U4300 (N_4300,N_2190,N_2586);
nor U4301 (N_4301,N_2799,N_2214);
nor U4302 (N_4302,N_3620,N_3698);
and U4303 (N_4303,N_2554,N_2846);
or U4304 (N_4304,N_2671,N_2572);
or U4305 (N_4305,N_3868,N_2666);
or U4306 (N_4306,N_2152,N_2467);
or U4307 (N_4307,N_2188,N_2810);
or U4308 (N_4308,N_3771,N_2537);
nor U4309 (N_4309,N_2502,N_2765);
nand U4310 (N_4310,N_3153,N_3930);
and U4311 (N_4311,N_3884,N_3474);
nand U4312 (N_4312,N_2172,N_2669);
nor U4313 (N_4313,N_2851,N_3359);
nand U4314 (N_4314,N_2165,N_2119);
nor U4315 (N_4315,N_2121,N_3835);
and U4316 (N_4316,N_2670,N_2278);
or U4317 (N_4317,N_2060,N_2084);
nand U4318 (N_4318,N_3736,N_3205);
or U4319 (N_4319,N_3974,N_3653);
and U4320 (N_4320,N_2887,N_3210);
xnor U4321 (N_4321,N_2796,N_2374);
and U4322 (N_4322,N_3238,N_2194);
nand U4323 (N_4323,N_2734,N_2067);
and U4324 (N_4324,N_2506,N_2298);
and U4325 (N_4325,N_3586,N_3526);
or U4326 (N_4326,N_2279,N_3543);
and U4327 (N_4327,N_3500,N_2309);
nor U4328 (N_4328,N_2416,N_3038);
nor U4329 (N_4329,N_2381,N_3871);
and U4330 (N_4330,N_3231,N_2147);
xor U4331 (N_4331,N_3019,N_2127);
or U4332 (N_4332,N_3822,N_2938);
nor U4333 (N_4333,N_3381,N_3705);
nor U4334 (N_4334,N_2677,N_2285);
nor U4335 (N_4335,N_3246,N_2909);
or U4336 (N_4336,N_3951,N_2102);
and U4337 (N_4337,N_3497,N_3393);
nand U4338 (N_4338,N_3832,N_2891);
and U4339 (N_4339,N_2834,N_3400);
nor U4340 (N_4340,N_3588,N_3978);
nand U4341 (N_4341,N_2630,N_2498);
nor U4342 (N_4342,N_2963,N_2870);
nor U4343 (N_4343,N_2522,N_2716);
nor U4344 (N_4344,N_3776,N_3233);
or U4345 (N_4345,N_3182,N_2024);
nand U4346 (N_4346,N_2879,N_3941);
or U4347 (N_4347,N_2602,N_2875);
nand U4348 (N_4348,N_3567,N_2401);
and U4349 (N_4349,N_2892,N_2028);
or U4350 (N_4350,N_2032,N_2740);
and U4351 (N_4351,N_2532,N_2329);
or U4352 (N_4352,N_3012,N_2791);
and U4353 (N_4353,N_2477,N_2149);
nand U4354 (N_4354,N_3882,N_3076);
xor U4355 (N_4355,N_2953,N_3031);
and U4356 (N_4356,N_3684,N_3634);
nor U4357 (N_4357,N_3442,N_3054);
nor U4358 (N_4358,N_2595,N_3599);
or U4359 (N_4359,N_3901,N_2080);
and U4360 (N_4360,N_3740,N_3432);
and U4361 (N_4361,N_3886,N_3052);
nor U4362 (N_4362,N_3005,N_3838);
nor U4363 (N_4363,N_2556,N_2660);
nor U4364 (N_4364,N_2183,N_2338);
nor U4365 (N_4365,N_2480,N_2785);
and U4366 (N_4366,N_3717,N_3390);
or U4367 (N_4367,N_2479,N_3621);
and U4368 (N_4368,N_3572,N_2702);
xnor U4369 (N_4369,N_3934,N_3931);
or U4370 (N_4370,N_2618,N_2270);
nand U4371 (N_4371,N_3438,N_2609);
or U4372 (N_4372,N_3697,N_3810);
or U4373 (N_4373,N_3558,N_3809);
nor U4374 (N_4374,N_2301,N_3232);
and U4375 (N_4375,N_2701,N_2966);
or U4376 (N_4376,N_2755,N_3169);
nor U4377 (N_4377,N_2807,N_2869);
nor U4378 (N_4378,N_3168,N_3467);
and U4379 (N_4379,N_3426,N_3334);
nand U4380 (N_4380,N_2726,N_2148);
or U4381 (N_4381,N_3483,N_2800);
nand U4382 (N_4382,N_2634,N_3532);
nand U4383 (N_4383,N_3632,N_2489);
or U4384 (N_4384,N_2504,N_3727);
nor U4385 (N_4385,N_2994,N_3976);
and U4386 (N_4386,N_3703,N_2109);
nand U4387 (N_4387,N_2413,N_2297);
nor U4388 (N_4388,N_3575,N_3947);
or U4389 (N_4389,N_2159,N_3926);
and U4390 (N_4390,N_3290,N_2768);
or U4391 (N_4391,N_3024,N_2145);
nand U4392 (N_4392,N_2674,N_2287);
nor U4393 (N_4393,N_3172,N_2895);
or U4394 (N_4394,N_3286,N_2456);
nand U4395 (N_4395,N_2228,N_3229);
or U4396 (N_4396,N_3357,N_3256);
xnor U4397 (N_4397,N_3505,N_2430);
nor U4398 (N_4398,N_3367,N_3303);
and U4399 (N_4399,N_2961,N_2444);
or U4400 (N_4400,N_3605,N_2268);
or U4401 (N_4401,N_3363,N_2980);
and U4402 (N_4402,N_3591,N_3496);
xnor U4403 (N_4403,N_3298,N_2333);
nand U4404 (N_4404,N_2303,N_3499);
nor U4405 (N_4405,N_2949,N_2230);
nor U4406 (N_4406,N_3802,N_2906);
xnor U4407 (N_4407,N_3691,N_2588);
nor U4408 (N_4408,N_3099,N_3781);
xnor U4409 (N_4409,N_3410,N_3269);
nor U4410 (N_4410,N_2013,N_2354);
xor U4411 (N_4411,N_3042,N_2927);
or U4412 (N_4412,N_3565,N_3265);
nand U4413 (N_4413,N_3473,N_2601);
and U4414 (N_4414,N_3897,N_2954);
nor U4415 (N_4415,N_2589,N_3107);
and U4416 (N_4416,N_3266,N_2763);
xor U4417 (N_4417,N_3763,N_2521);
and U4418 (N_4418,N_2626,N_2003);
xor U4419 (N_4419,N_3783,N_2915);
or U4420 (N_4420,N_3519,N_3927);
and U4421 (N_4421,N_3314,N_3166);
or U4422 (N_4422,N_3247,N_3160);
nor U4423 (N_4423,N_3895,N_3513);
nand U4424 (N_4424,N_3195,N_3083);
xor U4425 (N_4425,N_2617,N_2649);
and U4426 (N_4426,N_3713,N_2096);
nand U4427 (N_4427,N_3098,N_3113);
and U4428 (N_4428,N_3903,N_2457);
or U4429 (N_4429,N_2582,N_2181);
and U4430 (N_4430,N_2931,N_2888);
nor U4431 (N_4431,N_3614,N_2411);
nor U4432 (N_4432,N_2304,N_2946);
xnor U4433 (N_4433,N_2089,N_3167);
and U4434 (N_4434,N_3949,N_3447);
nor U4435 (N_4435,N_2505,N_2339);
xor U4436 (N_4436,N_3797,N_2591);
xnor U4437 (N_4437,N_2704,N_3796);
nand U4438 (N_4438,N_3036,N_3855);
or U4439 (N_4439,N_3553,N_2274);
xor U4440 (N_4440,N_3507,N_3770);
or U4441 (N_4441,N_3744,N_2046);
or U4442 (N_4442,N_2959,N_3111);
xnor U4443 (N_4443,N_2794,N_3482);
and U4444 (N_4444,N_2375,N_2128);
and U4445 (N_4445,N_3457,N_3080);
and U4446 (N_4446,N_2272,N_2672);
and U4447 (N_4447,N_3839,N_3029);
or U4448 (N_4448,N_3948,N_3960);
and U4449 (N_4449,N_3163,N_2429);
nor U4450 (N_4450,N_2700,N_2536);
and U4451 (N_4451,N_2453,N_2843);
nand U4452 (N_4452,N_2398,N_3138);
and U4453 (N_4453,N_2562,N_3016);
nand U4454 (N_4454,N_3775,N_3073);
xor U4455 (N_4455,N_3912,N_2507);
and U4456 (N_4456,N_3047,N_2607);
nor U4457 (N_4457,N_3581,N_2741);
nor U4458 (N_4458,N_2717,N_2531);
and U4459 (N_4459,N_2637,N_3477);
nand U4460 (N_4460,N_3396,N_2245);
xor U4461 (N_4461,N_3552,N_2399);
nor U4462 (N_4462,N_3848,N_3040);
nand U4463 (N_4463,N_3046,N_2720);
nor U4464 (N_4464,N_3475,N_3015);
nor U4465 (N_4465,N_3790,N_3428);
nand U4466 (N_4466,N_2627,N_3081);
nor U4467 (N_4467,N_2757,N_2133);
nand U4468 (N_4468,N_3170,N_3950);
nand U4469 (N_4469,N_2395,N_3890);
nor U4470 (N_4470,N_3215,N_3600);
and U4471 (N_4471,N_3644,N_2317);
or U4472 (N_4472,N_2867,N_2539);
or U4473 (N_4473,N_3097,N_3768);
or U4474 (N_4474,N_2824,N_2255);
or U4475 (N_4475,N_2318,N_2850);
and U4476 (N_4476,N_3455,N_3711);
nor U4477 (N_4477,N_2974,N_3789);
and U4478 (N_4478,N_2787,N_2210);
or U4479 (N_4479,N_2344,N_2129);
nand U4480 (N_4480,N_3865,N_2600);
xnor U4481 (N_4481,N_3559,N_2211);
or U4482 (N_4482,N_2737,N_3459);
or U4483 (N_4483,N_2055,N_3465);
and U4484 (N_4484,N_2865,N_3356);
and U4485 (N_4485,N_2943,N_3568);
or U4486 (N_4486,N_3725,N_3734);
and U4487 (N_4487,N_3506,N_3878);
nor U4488 (N_4488,N_3001,N_3384);
and U4489 (N_4489,N_2976,N_3288);
xor U4490 (N_4490,N_3368,N_2811);
and U4491 (N_4491,N_3480,N_2587);
and U4492 (N_4492,N_3239,N_3893);
nor U4493 (N_4493,N_3331,N_3084);
xnor U4494 (N_4494,N_3573,N_2608);
nand U4495 (N_4495,N_3018,N_2598);
nand U4496 (N_4496,N_3859,N_2624);
and U4497 (N_4497,N_2769,N_3885);
nor U4498 (N_4498,N_2908,N_2530);
or U4499 (N_4499,N_3847,N_3648);
or U4500 (N_4500,N_2146,N_3834);
or U4501 (N_4501,N_2100,N_3249);
or U4502 (N_4502,N_2341,N_2018);
nand U4503 (N_4503,N_2174,N_2615);
nor U4504 (N_4504,N_2760,N_2349);
and U4505 (N_4505,N_2893,N_2474);
or U4506 (N_4506,N_3151,N_2058);
nor U4507 (N_4507,N_3275,N_2166);
and U4508 (N_4508,N_2842,N_3082);
nand U4509 (N_4509,N_2346,N_2721);
nand U4510 (N_4510,N_3051,N_3669);
and U4511 (N_4511,N_3399,N_2240);
or U4512 (N_4512,N_3688,N_2157);
or U4513 (N_4513,N_2384,N_3905);
nor U4514 (N_4514,N_2005,N_3347);
xor U4515 (N_4515,N_2029,N_2021);
nor U4516 (N_4516,N_2856,N_2982);
or U4517 (N_4517,N_2901,N_3639);
and U4518 (N_4518,N_3039,N_3241);
or U4519 (N_4519,N_2396,N_3579);
or U4520 (N_4520,N_2490,N_2125);
nand U4521 (N_4521,N_2065,N_2358);
nor U4522 (N_4522,N_3424,N_2880);
or U4523 (N_4523,N_2073,N_3718);
nor U4524 (N_4524,N_3451,N_2853);
nand U4525 (N_4525,N_3386,N_3158);
or U4526 (N_4526,N_3284,N_3964);
or U4527 (N_4527,N_3173,N_2729);
and U4528 (N_4528,N_3985,N_3439);
and U4529 (N_4529,N_3883,N_3320);
nand U4530 (N_4530,N_3263,N_3686);
or U4531 (N_4531,N_2656,N_2034);
or U4532 (N_4532,N_3706,N_2552);
or U4533 (N_4533,N_2812,N_2141);
or U4534 (N_4534,N_2406,N_3671);
xnor U4535 (N_4535,N_3913,N_2580);
and U4536 (N_4536,N_2792,N_2647);
or U4537 (N_4537,N_3055,N_3795);
or U4538 (N_4538,N_3300,N_2478);
nor U4539 (N_4539,N_3094,N_2163);
or U4540 (N_4540,N_3751,N_3221);
and U4541 (N_4541,N_3631,N_2455);
and U4542 (N_4542,N_3709,N_2320);
nor U4543 (N_4543,N_2308,N_3784);
and U4544 (N_4544,N_3765,N_2866);
nand U4545 (N_4545,N_3065,N_2549);
xor U4546 (N_4546,N_2733,N_3833);
or U4547 (N_4547,N_2745,N_3909);
and U4548 (N_4548,N_2942,N_2832);
and U4549 (N_4549,N_2644,N_3454);
nand U4550 (N_4550,N_2956,N_2085);
and U4551 (N_4551,N_2027,N_2132);
nand U4552 (N_4552,N_3409,N_2319);
or U4553 (N_4553,N_2905,N_2593);
or U4554 (N_4554,N_2625,N_2497);
nor U4555 (N_4555,N_3610,N_3661);
and U4556 (N_4556,N_2025,N_3816);
or U4557 (N_4557,N_2643,N_2944);
and U4558 (N_4558,N_3406,N_2124);
or U4559 (N_4559,N_2232,N_2178);
nor U4560 (N_4560,N_2068,N_2361);
and U4561 (N_4561,N_3760,N_3422);
and U4562 (N_4562,N_2558,N_2574);
nand U4563 (N_4563,N_3289,N_2579);
or U4564 (N_4564,N_3274,N_2209);
nand U4565 (N_4565,N_2560,N_3025);
nand U4566 (N_4566,N_2327,N_3910);
nand U4567 (N_4567,N_2470,N_2064);
xnor U4568 (N_4568,N_2362,N_3911);
or U4569 (N_4569,N_2019,N_3450);
nor U4570 (N_4570,N_3652,N_3132);
nand U4571 (N_4571,N_3134,N_3441);
or U4572 (N_4572,N_2858,N_3446);
and U4573 (N_4573,N_3994,N_3319);
nor U4574 (N_4574,N_3659,N_2848);
or U4575 (N_4575,N_2813,N_2371);
nand U4576 (N_4576,N_2486,N_3276);
nand U4577 (N_4577,N_3928,N_2534);
xor U4578 (N_4578,N_3297,N_2861);
nand U4579 (N_4579,N_3813,N_2837);
xnor U4580 (N_4580,N_3121,N_2914);
or U4581 (N_4581,N_3443,N_3471);
and U4582 (N_4582,N_3008,N_3562);
nand U4583 (N_4583,N_3177,N_2830);
and U4584 (N_4584,N_3814,N_2585);
nor U4585 (N_4585,N_2241,N_2123);
or U4586 (N_4586,N_3478,N_3891);
nor U4587 (N_4587,N_2062,N_2311);
nor U4588 (N_4588,N_2705,N_3311);
nor U4589 (N_4589,N_2827,N_3722);
nor U4590 (N_4590,N_2323,N_3750);
nand U4591 (N_4591,N_2313,N_2260);
xnor U4592 (N_4592,N_2682,N_3335);
nand U4593 (N_4593,N_2638,N_2199);
nor U4594 (N_4594,N_3645,N_2466);
and U4595 (N_4595,N_2679,N_2271);
nor U4596 (N_4596,N_3820,N_2711);
and U4597 (N_4597,N_2353,N_2378);
nand U4598 (N_4598,N_2243,N_3369);
and U4599 (N_4599,N_3056,N_2985);
nor U4600 (N_4600,N_3380,N_2153);
nand U4601 (N_4601,N_2640,N_2828);
xor U4602 (N_4602,N_3187,N_3433);
and U4603 (N_4603,N_2264,N_2883);
xnor U4604 (N_4604,N_3354,N_2066);
and U4605 (N_4605,N_3124,N_3594);
nor U4606 (N_4606,N_3104,N_3595);
nand U4607 (N_4607,N_2965,N_3807);
and U4608 (N_4608,N_3748,N_2864);
and U4609 (N_4609,N_2759,N_3654);
nand U4610 (N_4610,N_2325,N_3071);
nand U4611 (N_4611,N_2404,N_3296);
xor U4612 (N_4612,N_2548,N_3864);
nand U4613 (N_4613,N_2269,N_2874);
nand U4614 (N_4614,N_2926,N_3254);
or U4615 (N_4615,N_2438,N_2897);
or U4616 (N_4616,N_2173,N_3382);
and U4617 (N_4617,N_3996,N_3004);
nor U4618 (N_4618,N_3650,N_3313);
nand U4619 (N_4619,N_3330,N_3665);
and U4620 (N_4620,N_3957,N_2220);
xor U4621 (N_4621,N_3407,N_2310);
and U4622 (N_4622,N_3445,N_2516);
or U4623 (N_4623,N_2993,N_2083);
xor U4624 (N_4624,N_2315,N_2225);
xnor U4625 (N_4625,N_3095,N_2805);
and U4626 (N_4626,N_2628,N_2423);
and U4627 (N_4627,N_2280,N_2917);
nand U4628 (N_4628,N_3808,N_3115);
or U4629 (N_4629,N_3148,N_3837);
nor U4630 (N_4630,N_2419,N_3321);
nand U4631 (N_4631,N_3604,N_3551);
nand U4632 (N_4632,N_3448,N_3074);
or U4633 (N_4633,N_2844,N_3504);
nand U4634 (N_4634,N_3743,N_2543);
and U4635 (N_4635,N_2081,N_2829);
and U4636 (N_4636,N_2999,N_2158);
and U4637 (N_4637,N_2696,N_2752);
or U4638 (N_4638,N_2642,N_3214);
nor U4639 (N_4639,N_2256,N_3561);
nand U4640 (N_4640,N_2881,N_2688);
nand U4641 (N_4641,N_3626,N_2465);
and U4642 (N_4642,N_3181,N_2667);
nor U4643 (N_4643,N_3458,N_3708);
nor U4644 (N_4644,N_3685,N_3612);
xnor U4645 (N_4645,N_3145,N_3922);
or U4646 (N_4646,N_3292,N_2557);
or U4647 (N_4647,N_3403,N_2098);
nand U4648 (N_4648,N_3815,N_2204);
and U4649 (N_4649,N_3690,N_2923);
or U4650 (N_4650,N_3606,N_3077);
nand U4651 (N_4651,N_3918,N_3366);
nand U4652 (N_4652,N_2360,N_2611);
and U4653 (N_4653,N_3655,N_2435);
nor U4654 (N_4654,N_3906,N_3268);
and U4655 (N_4655,N_2662,N_3079);
nor U4656 (N_4656,N_3827,N_3769);
and U4657 (N_4657,N_2051,N_2622);
or U4658 (N_4658,N_2104,N_3203);
and U4659 (N_4659,N_2641,N_2833);
and U4660 (N_4660,N_3270,N_2784);
nor U4661 (N_4661,N_3000,N_2665);
and U4662 (N_4662,N_2958,N_2449);
xnor U4663 (N_4663,N_3735,N_2535);
xnor U4664 (N_4664,N_2689,N_2196);
nor U4665 (N_4665,N_2645,N_2471);
or U4666 (N_4666,N_2370,N_3988);
or U4667 (N_4667,N_2434,N_3136);
xnor U4668 (N_4668,N_3192,N_2322);
or U4669 (N_4669,N_3613,N_3131);
or U4670 (N_4670,N_2097,N_2890);
nand U4671 (N_4671,N_3772,N_3877);
xor U4672 (N_4672,N_2878,N_3687);
and U4673 (N_4673,N_2680,N_3106);
and U4674 (N_4674,N_3578,N_3200);
nor U4675 (N_4675,N_2743,N_3201);
and U4676 (N_4676,N_3692,N_2541);
xor U4677 (N_4677,N_3970,N_2724);
nor U4678 (N_4678,N_2567,N_2778);
nand U4679 (N_4679,N_2967,N_2385);
nand U4680 (N_4680,N_2632,N_3180);
nor U4681 (N_4681,N_2779,N_2709);
or U4682 (N_4682,N_3494,N_3755);
or U4683 (N_4683,N_2135,N_3527);
and U4684 (N_4684,N_2749,N_3118);
and U4685 (N_4685,N_3932,N_3485);
nand U4686 (N_4686,N_2421,N_2902);
or U4687 (N_4687,N_3619,N_2983);
or U4688 (N_4688,N_3007,N_2952);
and U4689 (N_4689,N_2636,N_2971);
or U4690 (N_4690,N_2564,N_3915);
or U4691 (N_4691,N_3401,N_2200);
nand U4692 (N_4692,N_2606,N_2710);
nand U4693 (N_4693,N_3267,N_3395);
nand U4694 (N_4694,N_3057,N_3237);
nand U4695 (N_4695,N_2889,N_3641);
and U4696 (N_4696,N_2048,N_3415);
nor U4697 (N_4697,N_2664,N_3252);
or U4698 (N_4698,N_2819,N_3377);
or U4699 (N_4699,N_3486,N_3418);
nor U4700 (N_4700,N_2509,N_2120);
nor U4701 (N_4701,N_3728,N_3596);
nand U4702 (N_4702,N_3992,N_2458);
or U4703 (N_4703,N_3343,N_3093);
or U4704 (N_4704,N_2154,N_3235);
xnor U4705 (N_4705,N_2650,N_3963);
nor U4706 (N_4706,N_3598,N_2288);
xnor U4707 (N_4707,N_3306,N_3302);
or U4708 (N_4708,N_2356,N_2394);
nor U4709 (N_4709,N_3792,N_3823);
or U4710 (N_4710,N_2871,N_2803);
xnor U4711 (N_4711,N_2771,N_2254);
and U4712 (N_4712,N_3636,N_3899);
and U4713 (N_4713,N_3961,N_3866);
nand U4714 (N_4714,N_2414,N_3955);
and U4715 (N_4715,N_3554,N_2350);
or U4716 (N_4716,N_3312,N_3841);
or U4717 (N_4717,N_2226,N_2584);
or U4718 (N_4718,N_3301,N_2126);
or U4719 (N_4719,N_2045,N_3355);
and U4720 (N_4720,N_3271,N_2409);
and U4721 (N_4721,N_2059,N_2839);
or U4722 (N_4722,N_3375,N_2727);
nor U4723 (N_4723,N_2432,N_3971);
and U4724 (N_4724,N_2500,N_2886);
or U4725 (N_4725,N_3058,N_2373);
and U4726 (N_4726,N_3419,N_2936);
nand U4727 (N_4727,N_3157,N_2485);
nor U4728 (N_4728,N_2868,N_3436);
nor U4729 (N_4729,N_2816,N_3515);
nand U4730 (N_4730,N_2499,N_2110);
nor U4731 (N_4731,N_2090,N_2275);
nor U4732 (N_4732,N_2382,N_3707);
nand U4733 (N_4733,N_3397,N_3414);
or U4734 (N_4734,N_2826,N_3590);
or U4735 (N_4735,N_2355,N_2764);
nor U4736 (N_4736,N_2332,N_3385);
nand U4737 (N_4737,N_3262,N_3223);
and U4738 (N_4738,N_3611,N_3843);
nand U4739 (N_4739,N_3085,N_3127);
nor U4740 (N_4740,N_2797,N_2573);
and U4741 (N_4741,N_3374,N_3049);
nor U4742 (N_4742,N_3317,N_2077);
or U4743 (N_4743,N_3130,N_2427);
and U4744 (N_4744,N_2907,N_3261);
and U4745 (N_4745,N_3920,N_3253);
nor U4746 (N_4746,N_3857,N_2687);
nor U4747 (N_4747,N_3128,N_3791);
nand U4748 (N_4748,N_3716,N_3537);
nor U4749 (N_4749,N_2916,N_2657);
nor U4750 (N_4750,N_2074,N_3973);
nor U4751 (N_4751,N_3753,N_2227);
nor U4752 (N_4752,N_2691,N_2529);
or U4753 (N_4753,N_3570,N_2989);
and U4754 (N_4754,N_3332,N_3557);
or U4755 (N_4755,N_2599,N_3141);
xnor U4756 (N_4756,N_3278,N_3556);
and U4757 (N_4757,N_2038,N_2835);
nor U4758 (N_4758,N_3142,N_2620);
or U4759 (N_4759,N_2300,N_2176);
nand U4760 (N_4760,N_3328,N_3545);
nor U4761 (N_4761,N_3923,N_3617);
nor U4762 (N_4762,N_2107,N_2742);
xnor U4763 (N_4763,N_3045,N_2714);
and U4764 (N_4764,N_3370,N_2054);
nand U4765 (N_4765,N_3308,N_3416);
or U4766 (N_4766,N_3752,N_2718);
or U4767 (N_4767,N_2052,N_3589);
or U4768 (N_4768,N_3969,N_2305);
xnor U4769 (N_4769,N_2514,N_3522);
nor U4770 (N_4770,N_2219,N_3981);
nand U4771 (N_4771,N_2825,N_2454);
and U4772 (N_4772,N_3647,N_2798);
or U4773 (N_4773,N_3694,N_2417);
nand U4774 (N_4774,N_3364,N_2078);
or U4775 (N_4775,N_3185,N_3341);
nand U4776 (N_4776,N_2592,N_2789);
nand U4777 (N_4777,N_2565,N_2299);
or U4778 (N_4778,N_3967,N_3699);
and U4779 (N_4779,N_2678,N_2663);
nor U4780 (N_4780,N_2042,N_2061);
and U4781 (N_4781,N_2170,N_3412);
nand U4782 (N_4782,N_3245,N_3206);
and U4783 (N_4783,N_2501,N_2248);
and U4784 (N_4784,N_3714,N_2105);
nor U4785 (N_4785,N_2633,N_3502);
nand U4786 (N_4786,N_2302,N_3362);
or U4787 (N_4787,N_2698,N_3188);
nand U4788 (N_4788,N_2898,N_2289);
or U4789 (N_4789,N_3392,N_3662);
or U4790 (N_4790,N_2244,N_2459);
nand U4791 (N_4791,N_3535,N_3739);
or U4792 (N_4792,N_2731,N_3701);
and U4793 (N_4793,N_2175,N_3966);
or U4794 (N_4794,N_3678,N_2619);
nor U4795 (N_4795,N_3997,N_2692);
nor U4796 (N_4796,N_3067,N_3387);
nor U4797 (N_4797,N_3980,N_3420);
xnor U4798 (N_4798,N_3602,N_2388);
or U4799 (N_4799,N_2351,N_2357);
nand U4800 (N_4800,N_2340,N_3547);
and U4801 (N_4801,N_2948,N_3894);
and U4802 (N_4802,N_2924,N_3090);
or U4803 (N_4803,N_2728,N_3508);
or U4804 (N_4804,N_3782,N_3326);
or U4805 (N_4805,N_2257,N_3898);
nor U4806 (N_4806,N_3975,N_3408);
xor U4807 (N_4807,N_3398,N_3942);
and U4808 (N_4808,N_2400,N_3140);
nor U4809 (N_4809,N_3733,N_3754);
or U4810 (N_4810,N_3028,N_3618);
nand U4811 (N_4811,N_3829,N_2330);
and U4812 (N_4812,N_3009,N_2193);
xor U4813 (N_4813,N_2503,N_3721);
nand U4814 (N_4814,N_3584,N_3962);
nor U4815 (N_4815,N_3812,N_3279);
or U4816 (N_4816,N_2386,N_2991);
nor U4817 (N_4817,N_3710,N_3861);
nor U4818 (N_4818,N_3803,N_3066);
and U4819 (N_4819,N_2496,N_3059);
and U4820 (N_4820,N_2493,N_2197);
nand U4821 (N_4821,N_2334,N_3968);
or U4822 (N_4822,N_3264,N_3555);
nand U4823 (N_4823,N_3348,N_2997);
nand U4824 (N_4824,N_2746,N_2614);
or U4825 (N_4825,N_2912,N_2037);
and U4826 (N_4826,N_3033,N_3953);
and U4827 (N_4827,N_2086,N_2009);
nand U4828 (N_4828,N_2899,N_3452);
and U4829 (N_4829,N_2143,N_2873);
or U4830 (N_4830,N_2544,N_2553);
nor U4831 (N_4831,N_3702,N_3881);
nand U4832 (N_4832,N_2979,N_3622);
nor U4833 (N_4833,N_3862,N_2616);
nor U4834 (N_4834,N_2750,N_3014);
or U4835 (N_4835,N_3872,N_2236);
nor U4836 (N_4836,N_2094,N_2377);
nor U4837 (N_4837,N_3876,N_3766);
and U4838 (N_4838,N_3512,N_2014);
nand U4839 (N_4839,N_2184,N_3318);
or U4840 (N_4840,N_3842,N_3139);
and U4841 (N_4841,N_3801,N_2998);
or U4842 (N_4842,N_2095,N_3629);
xor U4843 (N_4843,N_3592,N_3342);
xor U4844 (N_4844,N_3285,N_2859);
or U4845 (N_4845,N_3003,N_2276);
and U4846 (N_4846,N_2231,N_2761);
nor U4847 (N_4847,N_3208,N_2838);
nor U4848 (N_4848,N_2894,N_2550);
or U4849 (N_4849,N_3798,N_2433);
xor U4850 (N_4850,N_2937,N_3587);
nand U4851 (N_4851,N_2144,N_2559);
nor U4852 (N_4852,N_2113,N_3649);
or U4853 (N_4853,N_3952,N_3738);
or U4854 (N_4854,N_2648,N_2407);
or U4855 (N_4855,N_3349,N_2981);
or U4856 (N_4856,N_2101,N_2555);
nor U4857 (N_4857,N_3196,N_2951);
nand U4858 (N_4858,N_3664,N_2817);
nand U4859 (N_4859,N_3929,N_2492);
nand U4860 (N_4860,N_3078,N_2930);
nor U4861 (N_4861,N_3982,N_3027);
nand U4862 (N_4862,N_3219,N_3917);
nand U4863 (N_4863,N_2597,N_3456);
or U4864 (N_4864,N_3123,N_2316);
nand U4865 (N_4865,N_2610,N_2167);
or U4866 (N_4866,N_2380,N_3050);
nor U4867 (N_4867,N_2103,N_3152);
nand U4868 (N_4868,N_3860,N_3786);
nand U4869 (N_4869,N_3440,N_3011);
or U4870 (N_4870,N_2017,N_2445);
nor U4871 (N_4871,N_3840,N_3100);
or U4872 (N_4872,N_3811,N_3785);
nor U4873 (N_4873,N_2168,N_3749);
nor U4874 (N_4874,N_3517,N_3938);
nand U4875 (N_4875,N_2265,N_2296);
nor U4876 (N_4876,N_2461,N_2191);
or U4877 (N_4877,N_3667,N_3304);
nor U4878 (N_4878,N_3109,N_2342);
nor U4879 (N_4879,N_3498,N_2405);
nand U4880 (N_4880,N_2546,N_3255);
nor U4881 (N_4881,N_3683,N_2941);
and U4882 (N_4882,N_2528,N_2314);
nand U4883 (N_4883,N_2708,N_3244);
nor U4884 (N_4884,N_3493,N_2082);
nand U4885 (N_4885,N_3914,N_3794);
nand U4886 (N_4886,N_3116,N_2821);
xnor U4887 (N_4887,N_3544,N_2252);
and U4888 (N_4888,N_2801,N_3818);
nor U4889 (N_4889,N_3689,N_3525);
or U4890 (N_4890,N_3693,N_3250);
or U4891 (N_4891,N_3681,N_2919);
nor U4892 (N_4892,N_2335,N_3830);
or U4893 (N_4893,N_3135,N_2903);
nand U4894 (N_4894,N_2939,N_2831);
or U4895 (N_4895,N_2282,N_3670);
nor U4896 (N_4896,N_3546,N_2007);
xnor U4897 (N_4897,N_2233,N_2860);
and U4898 (N_4898,N_3916,N_3217);
nor U4899 (N_4899,N_3601,N_2112);
and U4900 (N_4900,N_2422,N_3088);
and U4901 (N_4901,N_2945,N_2359);
xor U4902 (N_4902,N_3287,N_3171);
or U4903 (N_4903,N_2134,N_2162);
nand U4904 (N_4904,N_2237,N_2970);
nand U4905 (N_4905,N_2277,N_2010);
and U4906 (N_4906,N_3216,N_2820);
or U4907 (N_4907,N_3582,N_2814);
nor U4908 (N_4908,N_2364,N_3259);
or U4909 (N_4909,N_3680,N_2192);
nand U4910 (N_4910,N_3666,N_2964);
or U4911 (N_4911,N_3921,N_3472);
nor U4912 (N_4912,N_2136,N_3528);
nor U4913 (N_4913,N_2363,N_2213);
and U4914 (N_4914,N_3193,N_3327);
or U4915 (N_4915,N_2031,N_2767);
nor U4916 (N_4916,N_2295,N_3825);
and U4917 (N_4917,N_2605,N_2224);
nand U4918 (N_4918,N_2703,N_3164);
nand U4919 (N_4919,N_2520,N_3846);
or U4920 (N_4920,N_3518,N_3479);
nor U4921 (N_4921,N_2950,N_2515);
or U4922 (N_4922,N_2169,N_3902);
or U4923 (N_4923,N_2933,N_3939);
xnor U4924 (N_4924,N_2594,N_2719);
nor U4925 (N_4925,N_3759,N_2517);
and U4926 (N_4926,N_2079,N_2563);
and U4927 (N_4927,N_2139,N_3633);
and U4928 (N_4928,N_3315,N_2525);
nand U4929 (N_4929,N_2369,N_3737);
or U4930 (N_4930,N_3729,N_3202);
nor U4931 (N_4931,N_3070,N_2576);
nor U4932 (N_4932,N_2635,N_2408);
nor U4933 (N_4933,N_3280,N_2182);
or U4934 (N_4934,N_2063,N_3657);
nand U4935 (N_4935,N_2150,N_2040);
nor U4936 (N_4936,N_3272,N_3804);
or U4937 (N_4937,N_2293,N_3489);
and U4938 (N_4938,N_3402,N_2590);
and U4939 (N_4939,N_3730,N_2736);
or U4940 (N_4940,N_3020,N_3032);
xor U4941 (N_4941,N_2039,N_2783);
nand U4942 (N_4942,N_2263,N_2519);
and U4943 (N_4943,N_3979,N_3063);
and U4944 (N_4944,N_3209,N_2415);
nand U4945 (N_4945,N_2603,N_2695);
nor U4946 (N_4946,N_3006,N_3787);
nor U4947 (N_4947,N_2000,N_3682);
and U4948 (N_4948,N_3720,N_2140);
or U4949 (N_4949,N_3509,N_3958);
xor U4950 (N_4950,N_3043,N_3435);
nor U4951 (N_4951,N_2171,N_3322);
or U4952 (N_4952,N_2604,N_2540);
nor U4953 (N_4953,N_3869,N_2885);
nand U4954 (N_4954,N_2483,N_2035);
nand U4955 (N_4955,N_3492,N_3352);
and U4956 (N_4956,N_3373,N_3282);
or U4957 (N_4957,N_3075,N_2659);
xor U4958 (N_4958,N_2390,N_2348);
or U4959 (N_4959,N_2011,N_2472);
nor U4960 (N_4960,N_3017,N_2022);
and U4961 (N_4961,N_3114,N_3700);
nand U4962 (N_4962,N_2876,N_3224);
and U4963 (N_4963,N_2925,N_3336);
or U4964 (N_4964,N_3723,N_3854);
and U4965 (N_4965,N_2751,N_3563);
or U4966 (N_4966,N_3764,N_3935);
nor U4967 (N_4967,N_2481,N_2511);
nand U4968 (N_4968,N_2510,N_3542);
nor U4969 (N_4969,N_2057,N_2863);
or U4970 (N_4970,N_3143,N_2215);
nor U4971 (N_4971,N_2675,N_2575);
or U4972 (N_4972,N_2402,N_2990);
and U4973 (N_4973,N_2494,N_3719);
xor U4974 (N_4974,N_2091,N_3549);
or U4975 (N_4975,N_2475,N_3379);
nand U4976 (N_4976,N_3696,N_3761);
nand U4977 (N_4977,N_2234,N_3874);
nand U4978 (N_4978,N_2707,N_2986);
nor U4979 (N_4979,N_2808,N_2533);
nor U4980 (N_4980,N_3989,N_2809);
nand U4981 (N_4981,N_3372,N_2049);
nand U4982 (N_4982,N_3183,N_2189);
or U4983 (N_4983,N_3940,N_2116);
and U4984 (N_4984,N_3338,N_2262);
nor U4985 (N_4985,N_3863,N_2968);
nor U4986 (N_4986,N_3637,N_2352);
or U4987 (N_4987,N_2015,N_3476);
xor U4988 (N_4988,N_3212,N_3651);
or U4989 (N_4989,N_2460,N_2156);
nor U4990 (N_4990,N_3034,N_2513);
or U4991 (N_4991,N_2331,N_2008);
xnor U4992 (N_4992,N_3817,N_3943);
nand U4993 (N_4993,N_3495,N_2706);
nand U4994 (N_4994,N_3873,N_2756);
nor U4995 (N_4995,N_3198,N_2044);
and U4996 (N_4996,N_2823,N_3427);
or U4997 (N_4997,N_3603,N_3624);
and U4998 (N_4998,N_3778,N_3086);
nor U4999 (N_4999,N_3638,N_2195);
nor U5000 (N_5000,N_2638,N_3668);
and U5001 (N_5001,N_2686,N_3447);
nor U5002 (N_5002,N_2203,N_3839);
and U5003 (N_5003,N_3088,N_2759);
and U5004 (N_5004,N_2584,N_2077);
xor U5005 (N_5005,N_2863,N_2292);
and U5006 (N_5006,N_3261,N_3386);
xnor U5007 (N_5007,N_3076,N_3281);
or U5008 (N_5008,N_3685,N_3603);
or U5009 (N_5009,N_3255,N_2470);
xnor U5010 (N_5010,N_2109,N_2271);
and U5011 (N_5011,N_2708,N_3010);
nor U5012 (N_5012,N_3231,N_3154);
or U5013 (N_5013,N_3449,N_2690);
and U5014 (N_5014,N_3915,N_3760);
xnor U5015 (N_5015,N_2990,N_2567);
nand U5016 (N_5016,N_2940,N_3326);
nand U5017 (N_5017,N_2770,N_3522);
or U5018 (N_5018,N_3358,N_2984);
and U5019 (N_5019,N_2602,N_3826);
or U5020 (N_5020,N_3497,N_2718);
nand U5021 (N_5021,N_2048,N_3898);
or U5022 (N_5022,N_3305,N_2348);
nor U5023 (N_5023,N_2523,N_2989);
nand U5024 (N_5024,N_2096,N_3780);
or U5025 (N_5025,N_2123,N_3554);
xnor U5026 (N_5026,N_2527,N_3472);
nand U5027 (N_5027,N_3945,N_2459);
nand U5028 (N_5028,N_3474,N_2676);
nand U5029 (N_5029,N_3944,N_2377);
or U5030 (N_5030,N_2345,N_3533);
or U5031 (N_5031,N_3410,N_3334);
nor U5032 (N_5032,N_2130,N_2815);
nor U5033 (N_5033,N_2980,N_3440);
nand U5034 (N_5034,N_2118,N_3049);
nor U5035 (N_5035,N_3408,N_2286);
and U5036 (N_5036,N_2498,N_2908);
nand U5037 (N_5037,N_2538,N_3266);
or U5038 (N_5038,N_3797,N_3795);
and U5039 (N_5039,N_2320,N_2589);
nor U5040 (N_5040,N_3777,N_3905);
nand U5041 (N_5041,N_3596,N_2745);
or U5042 (N_5042,N_2638,N_3529);
and U5043 (N_5043,N_2160,N_2684);
nor U5044 (N_5044,N_3495,N_3745);
or U5045 (N_5045,N_2757,N_3450);
nand U5046 (N_5046,N_3325,N_2018);
xor U5047 (N_5047,N_3972,N_3273);
nor U5048 (N_5048,N_2197,N_2602);
or U5049 (N_5049,N_2975,N_2333);
nand U5050 (N_5050,N_3605,N_3836);
or U5051 (N_5051,N_2219,N_3255);
nor U5052 (N_5052,N_2955,N_2765);
nand U5053 (N_5053,N_2262,N_2561);
nor U5054 (N_5054,N_2350,N_2694);
xor U5055 (N_5055,N_3349,N_2932);
nand U5056 (N_5056,N_2334,N_2295);
or U5057 (N_5057,N_2702,N_3979);
xnor U5058 (N_5058,N_3699,N_3321);
and U5059 (N_5059,N_3966,N_2785);
nor U5060 (N_5060,N_2540,N_3000);
and U5061 (N_5061,N_3538,N_3605);
or U5062 (N_5062,N_2199,N_2823);
nor U5063 (N_5063,N_2789,N_2358);
or U5064 (N_5064,N_2646,N_2693);
and U5065 (N_5065,N_2175,N_3148);
nor U5066 (N_5066,N_2549,N_2252);
and U5067 (N_5067,N_2350,N_2334);
or U5068 (N_5068,N_2425,N_2969);
nand U5069 (N_5069,N_2002,N_3714);
or U5070 (N_5070,N_2662,N_3570);
and U5071 (N_5071,N_2023,N_2629);
nand U5072 (N_5072,N_3306,N_2265);
nand U5073 (N_5073,N_3696,N_2374);
nor U5074 (N_5074,N_2940,N_2023);
and U5075 (N_5075,N_2613,N_2368);
xnor U5076 (N_5076,N_2629,N_2597);
nor U5077 (N_5077,N_2375,N_3405);
nand U5078 (N_5078,N_2762,N_3512);
nor U5079 (N_5079,N_3560,N_2103);
or U5080 (N_5080,N_3589,N_2982);
and U5081 (N_5081,N_2816,N_3171);
nand U5082 (N_5082,N_2073,N_3975);
nor U5083 (N_5083,N_3299,N_2631);
nand U5084 (N_5084,N_3433,N_2684);
nand U5085 (N_5085,N_3553,N_3500);
or U5086 (N_5086,N_3053,N_3414);
and U5087 (N_5087,N_2858,N_2664);
and U5088 (N_5088,N_2080,N_2683);
nand U5089 (N_5089,N_2119,N_3062);
or U5090 (N_5090,N_2904,N_2102);
nand U5091 (N_5091,N_2085,N_3144);
nand U5092 (N_5092,N_2105,N_3232);
nand U5093 (N_5093,N_2836,N_2036);
nand U5094 (N_5094,N_2527,N_2302);
nand U5095 (N_5095,N_2252,N_2930);
nand U5096 (N_5096,N_3332,N_2152);
nand U5097 (N_5097,N_2969,N_2174);
nor U5098 (N_5098,N_2749,N_3388);
or U5099 (N_5099,N_2921,N_2715);
xor U5100 (N_5100,N_2067,N_2902);
nor U5101 (N_5101,N_3563,N_2710);
and U5102 (N_5102,N_3876,N_2998);
nor U5103 (N_5103,N_2705,N_2880);
or U5104 (N_5104,N_3701,N_3732);
or U5105 (N_5105,N_3543,N_3456);
nand U5106 (N_5106,N_2027,N_3441);
xnor U5107 (N_5107,N_2920,N_2724);
nand U5108 (N_5108,N_2016,N_3768);
or U5109 (N_5109,N_2226,N_2040);
nand U5110 (N_5110,N_2261,N_2611);
and U5111 (N_5111,N_2747,N_2532);
nor U5112 (N_5112,N_2457,N_3080);
nor U5113 (N_5113,N_2461,N_2001);
nor U5114 (N_5114,N_2774,N_3608);
xor U5115 (N_5115,N_2931,N_3731);
and U5116 (N_5116,N_2624,N_3165);
or U5117 (N_5117,N_3773,N_2560);
or U5118 (N_5118,N_3869,N_3750);
nor U5119 (N_5119,N_2053,N_2036);
nor U5120 (N_5120,N_2021,N_3333);
nor U5121 (N_5121,N_3816,N_2032);
or U5122 (N_5122,N_2382,N_3180);
and U5123 (N_5123,N_2732,N_3521);
or U5124 (N_5124,N_2540,N_2226);
nand U5125 (N_5125,N_2966,N_2352);
xor U5126 (N_5126,N_3768,N_3562);
nor U5127 (N_5127,N_2549,N_2687);
nor U5128 (N_5128,N_3459,N_2592);
nand U5129 (N_5129,N_2491,N_3176);
or U5130 (N_5130,N_2946,N_2704);
xor U5131 (N_5131,N_3276,N_3713);
nor U5132 (N_5132,N_3859,N_3114);
and U5133 (N_5133,N_3179,N_3607);
or U5134 (N_5134,N_3174,N_2589);
nand U5135 (N_5135,N_2363,N_3099);
and U5136 (N_5136,N_3241,N_3804);
and U5137 (N_5137,N_2528,N_2228);
nand U5138 (N_5138,N_3931,N_3457);
nor U5139 (N_5139,N_3187,N_3558);
or U5140 (N_5140,N_3751,N_2315);
and U5141 (N_5141,N_3508,N_2158);
nor U5142 (N_5142,N_3289,N_3481);
or U5143 (N_5143,N_2477,N_3201);
or U5144 (N_5144,N_2304,N_2609);
nor U5145 (N_5145,N_3252,N_2517);
or U5146 (N_5146,N_2501,N_2560);
nor U5147 (N_5147,N_3935,N_2615);
or U5148 (N_5148,N_3413,N_2244);
and U5149 (N_5149,N_2098,N_2525);
and U5150 (N_5150,N_2076,N_2307);
and U5151 (N_5151,N_3898,N_2280);
nand U5152 (N_5152,N_2859,N_3936);
or U5153 (N_5153,N_3264,N_3556);
or U5154 (N_5154,N_3224,N_2068);
nor U5155 (N_5155,N_2735,N_2704);
nand U5156 (N_5156,N_3021,N_2812);
and U5157 (N_5157,N_2307,N_2353);
or U5158 (N_5158,N_2916,N_2502);
nand U5159 (N_5159,N_2382,N_2327);
and U5160 (N_5160,N_3774,N_3724);
xnor U5161 (N_5161,N_2627,N_3314);
and U5162 (N_5162,N_2335,N_2778);
nand U5163 (N_5163,N_3818,N_3057);
nor U5164 (N_5164,N_2760,N_3884);
nor U5165 (N_5165,N_2065,N_2631);
xor U5166 (N_5166,N_3331,N_3582);
nor U5167 (N_5167,N_2239,N_2446);
and U5168 (N_5168,N_2705,N_3330);
nand U5169 (N_5169,N_2075,N_3840);
xnor U5170 (N_5170,N_2878,N_2368);
nor U5171 (N_5171,N_3891,N_2934);
or U5172 (N_5172,N_2735,N_3716);
nand U5173 (N_5173,N_2894,N_2523);
or U5174 (N_5174,N_3186,N_2376);
xor U5175 (N_5175,N_3873,N_3291);
xnor U5176 (N_5176,N_2178,N_2384);
and U5177 (N_5177,N_3876,N_3727);
and U5178 (N_5178,N_2742,N_2532);
and U5179 (N_5179,N_3341,N_2604);
or U5180 (N_5180,N_3159,N_2032);
nor U5181 (N_5181,N_3017,N_3952);
and U5182 (N_5182,N_2763,N_3910);
or U5183 (N_5183,N_2847,N_2169);
and U5184 (N_5184,N_2603,N_2381);
nand U5185 (N_5185,N_3285,N_2345);
nand U5186 (N_5186,N_2138,N_3429);
nor U5187 (N_5187,N_2424,N_3990);
or U5188 (N_5188,N_2170,N_3323);
xor U5189 (N_5189,N_2928,N_2295);
or U5190 (N_5190,N_2166,N_3239);
and U5191 (N_5191,N_3757,N_2128);
nor U5192 (N_5192,N_3808,N_2469);
and U5193 (N_5193,N_2398,N_3967);
or U5194 (N_5194,N_3643,N_3281);
nor U5195 (N_5195,N_2685,N_2635);
nand U5196 (N_5196,N_2368,N_2668);
or U5197 (N_5197,N_3933,N_2229);
xnor U5198 (N_5198,N_3638,N_3823);
or U5199 (N_5199,N_2044,N_3650);
or U5200 (N_5200,N_2615,N_2973);
xor U5201 (N_5201,N_3699,N_3734);
nor U5202 (N_5202,N_2423,N_2823);
nand U5203 (N_5203,N_2122,N_2962);
or U5204 (N_5204,N_3487,N_3096);
nand U5205 (N_5205,N_2553,N_2235);
nor U5206 (N_5206,N_3222,N_2133);
nor U5207 (N_5207,N_3777,N_2219);
and U5208 (N_5208,N_2737,N_3587);
nor U5209 (N_5209,N_3237,N_2861);
and U5210 (N_5210,N_2082,N_3227);
or U5211 (N_5211,N_2862,N_3910);
or U5212 (N_5212,N_2790,N_2389);
nor U5213 (N_5213,N_3062,N_3583);
and U5214 (N_5214,N_3382,N_2354);
nor U5215 (N_5215,N_3984,N_3281);
nor U5216 (N_5216,N_3558,N_2950);
and U5217 (N_5217,N_3750,N_3369);
nand U5218 (N_5218,N_2219,N_2882);
and U5219 (N_5219,N_3204,N_3016);
nor U5220 (N_5220,N_2075,N_3305);
or U5221 (N_5221,N_3974,N_2108);
nor U5222 (N_5222,N_3156,N_3815);
or U5223 (N_5223,N_3765,N_2234);
nor U5224 (N_5224,N_3302,N_2409);
xor U5225 (N_5225,N_3535,N_2735);
or U5226 (N_5226,N_2258,N_3414);
or U5227 (N_5227,N_2012,N_2218);
nand U5228 (N_5228,N_3192,N_3896);
and U5229 (N_5229,N_3679,N_3221);
nor U5230 (N_5230,N_2736,N_3348);
nand U5231 (N_5231,N_3058,N_3640);
nand U5232 (N_5232,N_2676,N_3840);
nand U5233 (N_5233,N_3956,N_3158);
and U5234 (N_5234,N_3384,N_3024);
nor U5235 (N_5235,N_3204,N_2691);
xor U5236 (N_5236,N_3072,N_2121);
or U5237 (N_5237,N_3403,N_3107);
or U5238 (N_5238,N_3705,N_2573);
or U5239 (N_5239,N_3635,N_3818);
nand U5240 (N_5240,N_3422,N_2136);
xor U5241 (N_5241,N_2143,N_2864);
nor U5242 (N_5242,N_2962,N_2517);
or U5243 (N_5243,N_2980,N_3751);
and U5244 (N_5244,N_2757,N_3404);
or U5245 (N_5245,N_2437,N_2969);
or U5246 (N_5246,N_2211,N_3747);
nand U5247 (N_5247,N_3185,N_3726);
xnor U5248 (N_5248,N_3531,N_2568);
and U5249 (N_5249,N_2374,N_2331);
and U5250 (N_5250,N_2441,N_3014);
nor U5251 (N_5251,N_2224,N_3550);
or U5252 (N_5252,N_3269,N_2840);
nand U5253 (N_5253,N_3390,N_2246);
nand U5254 (N_5254,N_3121,N_2910);
nor U5255 (N_5255,N_3662,N_3971);
nor U5256 (N_5256,N_2348,N_3706);
or U5257 (N_5257,N_2378,N_3771);
and U5258 (N_5258,N_3184,N_3653);
nand U5259 (N_5259,N_3500,N_2185);
nor U5260 (N_5260,N_2174,N_3869);
or U5261 (N_5261,N_2294,N_3164);
nor U5262 (N_5262,N_2981,N_3108);
or U5263 (N_5263,N_2350,N_3274);
nor U5264 (N_5264,N_3300,N_3046);
and U5265 (N_5265,N_3653,N_3941);
and U5266 (N_5266,N_3717,N_2002);
nand U5267 (N_5267,N_2732,N_3698);
nor U5268 (N_5268,N_3280,N_3438);
xnor U5269 (N_5269,N_2399,N_3839);
xnor U5270 (N_5270,N_2136,N_3892);
xnor U5271 (N_5271,N_3589,N_2275);
nor U5272 (N_5272,N_2361,N_2929);
nand U5273 (N_5273,N_2383,N_3846);
nor U5274 (N_5274,N_2839,N_3368);
nor U5275 (N_5275,N_3582,N_2622);
xor U5276 (N_5276,N_2836,N_3144);
nand U5277 (N_5277,N_3368,N_3987);
nor U5278 (N_5278,N_2001,N_2546);
xor U5279 (N_5279,N_2446,N_3356);
or U5280 (N_5280,N_3837,N_3068);
xnor U5281 (N_5281,N_3516,N_3909);
nand U5282 (N_5282,N_2980,N_3508);
and U5283 (N_5283,N_2035,N_3440);
and U5284 (N_5284,N_2933,N_2210);
nor U5285 (N_5285,N_3067,N_3469);
nand U5286 (N_5286,N_3597,N_3005);
or U5287 (N_5287,N_3955,N_3017);
or U5288 (N_5288,N_3545,N_3686);
and U5289 (N_5289,N_3119,N_3957);
or U5290 (N_5290,N_2335,N_2824);
xor U5291 (N_5291,N_2874,N_3267);
nor U5292 (N_5292,N_2368,N_2574);
nand U5293 (N_5293,N_2844,N_3435);
nor U5294 (N_5294,N_3089,N_2266);
nand U5295 (N_5295,N_3139,N_3410);
and U5296 (N_5296,N_2504,N_2216);
nand U5297 (N_5297,N_2657,N_3264);
and U5298 (N_5298,N_2150,N_2021);
nor U5299 (N_5299,N_2388,N_2324);
xor U5300 (N_5300,N_2239,N_2347);
xor U5301 (N_5301,N_3685,N_3555);
or U5302 (N_5302,N_3058,N_2972);
xor U5303 (N_5303,N_3425,N_2203);
nand U5304 (N_5304,N_2030,N_2409);
or U5305 (N_5305,N_3834,N_2711);
nor U5306 (N_5306,N_2326,N_3417);
nand U5307 (N_5307,N_3963,N_3673);
nand U5308 (N_5308,N_3605,N_2127);
xnor U5309 (N_5309,N_3939,N_2176);
nor U5310 (N_5310,N_3153,N_2154);
nor U5311 (N_5311,N_3330,N_3718);
and U5312 (N_5312,N_3904,N_3408);
and U5313 (N_5313,N_3274,N_2197);
or U5314 (N_5314,N_2244,N_2667);
and U5315 (N_5315,N_2299,N_2239);
or U5316 (N_5316,N_2463,N_3980);
and U5317 (N_5317,N_3325,N_3189);
nor U5318 (N_5318,N_2638,N_3437);
and U5319 (N_5319,N_2155,N_2351);
nand U5320 (N_5320,N_2755,N_2862);
nor U5321 (N_5321,N_3499,N_3047);
nand U5322 (N_5322,N_3553,N_3051);
and U5323 (N_5323,N_3116,N_2290);
or U5324 (N_5324,N_3298,N_2556);
nor U5325 (N_5325,N_2700,N_2753);
or U5326 (N_5326,N_3865,N_3947);
or U5327 (N_5327,N_2570,N_3346);
or U5328 (N_5328,N_2239,N_2036);
or U5329 (N_5329,N_3095,N_3908);
xnor U5330 (N_5330,N_2419,N_3271);
or U5331 (N_5331,N_3164,N_3505);
nor U5332 (N_5332,N_2128,N_2455);
xor U5333 (N_5333,N_3667,N_3766);
and U5334 (N_5334,N_2902,N_3666);
and U5335 (N_5335,N_3412,N_3279);
nand U5336 (N_5336,N_2628,N_3474);
nand U5337 (N_5337,N_2121,N_2255);
nand U5338 (N_5338,N_3613,N_2682);
nand U5339 (N_5339,N_2327,N_2636);
or U5340 (N_5340,N_3734,N_2083);
nand U5341 (N_5341,N_3492,N_2624);
and U5342 (N_5342,N_3292,N_2710);
nand U5343 (N_5343,N_3219,N_2457);
nor U5344 (N_5344,N_2573,N_3501);
nor U5345 (N_5345,N_2667,N_2003);
nand U5346 (N_5346,N_2367,N_3756);
or U5347 (N_5347,N_2874,N_3877);
or U5348 (N_5348,N_2944,N_3039);
nand U5349 (N_5349,N_2974,N_3547);
and U5350 (N_5350,N_3260,N_3193);
and U5351 (N_5351,N_3020,N_3013);
nand U5352 (N_5352,N_3789,N_3228);
or U5353 (N_5353,N_2488,N_3783);
nor U5354 (N_5354,N_2220,N_2187);
or U5355 (N_5355,N_3916,N_2263);
or U5356 (N_5356,N_2814,N_3191);
or U5357 (N_5357,N_2525,N_3240);
nor U5358 (N_5358,N_3776,N_2286);
or U5359 (N_5359,N_2097,N_3429);
nor U5360 (N_5360,N_2697,N_2287);
or U5361 (N_5361,N_2603,N_2401);
nor U5362 (N_5362,N_2489,N_2621);
nor U5363 (N_5363,N_3498,N_2858);
nand U5364 (N_5364,N_2012,N_2820);
or U5365 (N_5365,N_3857,N_2084);
and U5366 (N_5366,N_3109,N_2244);
nand U5367 (N_5367,N_2199,N_3006);
nor U5368 (N_5368,N_2920,N_3605);
nand U5369 (N_5369,N_3187,N_2112);
nand U5370 (N_5370,N_2092,N_3370);
or U5371 (N_5371,N_3507,N_2363);
or U5372 (N_5372,N_2511,N_2948);
and U5373 (N_5373,N_3754,N_3907);
xor U5374 (N_5374,N_2936,N_2652);
nand U5375 (N_5375,N_2580,N_2289);
and U5376 (N_5376,N_3410,N_3818);
nand U5377 (N_5377,N_2071,N_3951);
or U5378 (N_5378,N_2042,N_2831);
and U5379 (N_5379,N_2744,N_3832);
and U5380 (N_5380,N_2864,N_2413);
and U5381 (N_5381,N_2165,N_2536);
or U5382 (N_5382,N_3975,N_3327);
and U5383 (N_5383,N_2475,N_2008);
nor U5384 (N_5384,N_3217,N_3466);
xnor U5385 (N_5385,N_2519,N_3355);
nand U5386 (N_5386,N_3013,N_3094);
and U5387 (N_5387,N_2248,N_3572);
or U5388 (N_5388,N_3988,N_2269);
nand U5389 (N_5389,N_3525,N_2859);
nand U5390 (N_5390,N_3979,N_3231);
or U5391 (N_5391,N_2439,N_2502);
xor U5392 (N_5392,N_2136,N_2350);
and U5393 (N_5393,N_2018,N_2908);
and U5394 (N_5394,N_3423,N_2037);
nor U5395 (N_5395,N_2348,N_2110);
and U5396 (N_5396,N_3898,N_3532);
or U5397 (N_5397,N_2238,N_3339);
and U5398 (N_5398,N_3086,N_2393);
nand U5399 (N_5399,N_3185,N_2274);
nand U5400 (N_5400,N_3137,N_3753);
nand U5401 (N_5401,N_2479,N_3924);
nor U5402 (N_5402,N_3066,N_3492);
nand U5403 (N_5403,N_3573,N_2277);
nor U5404 (N_5404,N_3690,N_3674);
and U5405 (N_5405,N_2189,N_2347);
nand U5406 (N_5406,N_2250,N_3089);
or U5407 (N_5407,N_3925,N_2484);
and U5408 (N_5408,N_3043,N_2155);
xor U5409 (N_5409,N_3575,N_3390);
and U5410 (N_5410,N_2778,N_3470);
nand U5411 (N_5411,N_3779,N_2202);
and U5412 (N_5412,N_3741,N_2725);
xor U5413 (N_5413,N_3388,N_2650);
nand U5414 (N_5414,N_2932,N_3744);
xor U5415 (N_5415,N_2886,N_3527);
and U5416 (N_5416,N_3147,N_2995);
or U5417 (N_5417,N_3748,N_3595);
nor U5418 (N_5418,N_2678,N_2155);
or U5419 (N_5419,N_2660,N_2965);
nand U5420 (N_5420,N_3821,N_2881);
xnor U5421 (N_5421,N_3079,N_2942);
and U5422 (N_5422,N_3609,N_3474);
and U5423 (N_5423,N_3379,N_3356);
nand U5424 (N_5424,N_3840,N_3961);
and U5425 (N_5425,N_3586,N_2902);
or U5426 (N_5426,N_3301,N_3343);
and U5427 (N_5427,N_3456,N_3532);
and U5428 (N_5428,N_3874,N_3006);
and U5429 (N_5429,N_2257,N_3529);
nor U5430 (N_5430,N_3495,N_2482);
nand U5431 (N_5431,N_3838,N_2956);
or U5432 (N_5432,N_2359,N_2194);
or U5433 (N_5433,N_3331,N_3488);
nand U5434 (N_5434,N_3923,N_3630);
nor U5435 (N_5435,N_2793,N_2787);
or U5436 (N_5436,N_2437,N_3371);
nand U5437 (N_5437,N_3275,N_2044);
nor U5438 (N_5438,N_2841,N_2296);
and U5439 (N_5439,N_2240,N_2134);
and U5440 (N_5440,N_2809,N_3316);
and U5441 (N_5441,N_2166,N_2469);
nand U5442 (N_5442,N_3805,N_2529);
or U5443 (N_5443,N_2755,N_2233);
nand U5444 (N_5444,N_2797,N_3793);
or U5445 (N_5445,N_3921,N_2666);
or U5446 (N_5446,N_2903,N_2493);
and U5447 (N_5447,N_3072,N_2305);
nor U5448 (N_5448,N_3034,N_2613);
nor U5449 (N_5449,N_3288,N_3758);
or U5450 (N_5450,N_3271,N_3536);
nand U5451 (N_5451,N_3104,N_3261);
xnor U5452 (N_5452,N_3665,N_3176);
and U5453 (N_5453,N_3017,N_3341);
nand U5454 (N_5454,N_2680,N_3742);
nor U5455 (N_5455,N_3476,N_2104);
and U5456 (N_5456,N_3484,N_3119);
and U5457 (N_5457,N_3668,N_2541);
nand U5458 (N_5458,N_3798,N_3384);
nor U5459 (N_5459,N_3784,N_3465);
and U5460 (N_5460,N_3096,N_2615);
and U5461 (N_5461,N_3796,N_3081);
xnor U5462 (N_5462,N_2829,N_2887);
or U5463 (N_5463,N_3748,N_2825);
or U5464 (N_5464,N_2787,N_2893);
and U5465 (N_5465,N_2531,N_2571);
nor U5466 (N_5466,N_3647,N_3891);
nor U5467 (N_5467,N_2686,N_2988);
nand U5468 (N_5468,N_3027,N_2989);
and U5469 (N_5469,N_2196,N_2341);
and U5470 (N_5470,N_2207,N_3051);
nor U5471 (N_5471,N_3075,N_2352);
and U5472 (N_5472,N_2075,N_3615);
nor U5473 (N_5473,N_2554,N_3935);
nand U5474 (N_5474,N_3753,N_2867);
nor U5475 (N_5475,N_3459,N_2117);
or U5476 (N_5476,N_3184,N_2748);
nor U5477 (N_5477,N_3771,N_2286);
or U5478 (N_5478,N_2030,N_3550);
or U5479 (N_5479,N_2356,N_3656);
xnor U5480 (N_5480,N_3571,N_3509);
nand U5481 (N_5481,N_2993,N_2865);
or U5482 (N_5482,N_2798,N_2150);
xor U5483 (N_5483,N_3917,N_3471);
or U5484 (N_5484,N_3744,N_3061);
nor U5485 (N_5485,N_3470,N_3144);
or U5486 (N_5486,N_2933,N_3343);
xnor U5487 (N_5487,N_2636,N_2556);
or U5488 (N_5488,N_2551,N_2708);
and U5489 (N_5489,N_3596,N_3376);
xor U5490 (N_5490,N_2201,N_2392);
or U5491 (N_5491,N_2093,N_2347);
and U5492 (N_5492,N_2777,N_3867);
and U5493 (N_5493,N_3387,N_2921);
or U5494 (N_5494,N_3185,N_3302);
nor U5495 (N_5495,N_3064,N_3897);
nor U5496 (N_5496,N_3916,N_2616);
or U5497 (N_5497,N_2972,N_3175);
and U5498 (N_5498,N_3384,N_3372);
nor U5499 (N_5499,N_3775,N_3827);
or U5500 (N_5500,N_3773,N_3398);
xor U5501 (N_5501,N_2288,N_2810);
nand U5502 (N_5502,N_3794,N_2114);
nand U5503 (N_5503,N_2428,N_3633);
xor U5504 (N_5504,N_2209,N_2722);
or U5505 (N_5505,N_2833,N_3459);
and U5506 (N_5506,N_3065,N_3815);
or U5507 (N_5507,N_3876,N_2873);
or U5508 (N_5508,N_2948,N_3706);
or U5509 (N_5509,N_2841,N_2706);
or U5510 (N_5510,N_3120,N_2495);
nor U5511 (N_5511,N_3794,N_3193);
or U5512 (N_5512,N_3700,N_2324);
and U5513 (N_5513,N_3573,N_2289);
and U5514 (N_5514,N_2791,N_3253);
nor U5515 (N_5515,N_2983,N_2992);
nand U5516 (N_5516,N_2794,N_2757);
or U5517 (N_5517,N_3933,N_2230);
xor U5518 (N_5518,N_3349,N_3734);
and U5519 (N_5519,N_3898,N_2670);
xor U5520 (N_5520,N_2913,N_2098);
nand U5521 (N_5521,N_2528,N_3725);
or U5522 (N_5522,N_2770,N_3032);
xnor U5523 (N_5523,N_2269,N_3162);
or U5524 (N_5524,N_3200,N_2738);
nor U5525 (N_5525,N_2574,N_2510);
nor U5526 (N_5526,N_2226,N_2548);
nand U5527 (N_5527,N_3097,N_3062);
and U5528 (N_5528,N_3819,N_3522);
nand U5529 (N_5529,N_2760,N_3815);
nand U5530 (N_5530,N_3443,N_2581);
or U5531 (N_5531,N_3633,N_3440);
and U5532 (N_5532,N_2864,N_3904);
and U5533 (N_5533,N_2151,N_3524);
and U5534 (N_5534,N_3866,N_2963);
xor U5535 (N_5535,N_2043,N_3893);
xor U5536 (N_5536,N_3467,N_2779);
nand U5537 (N_5537,N_2334,N_3019);
nand U5538 (N_5538,N_2193,N_3702);
nor U5539 (N_5539,N_2274,N_3694);
nor U5540 (N_5540,N_2554,N_3850);
or U5541 (N_5541,N_3843,N_2116);
and U5542 (N_5542,N_2493,N_3048);
nor U5543 (N_5543,N_3098,N_3418);
nor U5544 (N_5544,N_2205,N_2421);
or U5545 (N_5545,N_3080,N_2202);
or U5546 (N_5546,N_2367,N_2464);
nor U5547 (N_5547,N_2937,N_2131);
or U5548 (N_5548,N_2890,N_2394);
or U5549 (N_5549,N_2306,N_3311);
and U5550 (N_5550,N_3267,N_2883);
nor U5551 (N_5551,N_2849,N_3618);
or U5552 (N_5552,N_3875,N_3569);
or U5553 (N_5553,N_2720,N_2965);
nand U5554 (N_5554,N_2650,N_2857);
or U5555 (N_5555,N_2485,N_3039);
and U5556 (N_5556,N_3289,N_2360);
nand U5557 (N_5557,N_2060,N_3563);
nand U5558 (N_5558,N_3395,N_3795);
or U5559 (N_5559,N_3431,N_2971);
or U5560 (N_5560,N_2646,N_2525);
xnor U5561 (N_5561,N_3287,N_2790);
nand U5562 (N_5562,N_3174,N_2815);
nor U5563 (N_5563,N_2503,N_3904);
or U5564 (N_5564,N_2695,N_3291);
nand U5565 (N_5565,N_3229,N_2956);
or U5566 (N_5566,N_2180,N_2390);
or U5567 (N_5567,N_2826,N_3889);
nand U5568 (N_5568,N_3790,N_2393);
nor U5569 (N_5569,N_2461,N_3039);
or U5570 (N_5570,N_2701,N_3307);
and U5571 (N_5571,N_2894,N_3758);
or U5572 (N_5572,N_2936,N_2139);
and U5573 (N_5573,N_3842,N_3946);
nand U5574 (N_5574,N_3864,N_2963);
nand U5575 (N_5575,N_3570,N_2374);
and U5576 (N_5576,N_3161,N_2862);
nor U5577 (N_5577,N_2058,N_3139);
and U5578 (N_5578,N_2006,N_2016);
nand U5579 (N_5579,N_2063,N_2159);
nand U5580 (N_5580,N_3937,N_2676);
nor U5581 (N_5581,N_3730,N_3645);
or U5582 (N_5582,N_2524,N_3778);
nor U5583 (N_5583,N_2681,N_3740);
or U5584 (N_5584,N_2764,N_3687);
and U5585 (N_5585,N_3282,N_2757);
nand U5586 (N_5586,N_2558,N_3752);
xor U5587 (N_5587,N_3398,N_3522);
nand U5588 (N_5588,N_2732,N_2705);
and U5589 (N_5589,N_2689,N_3520);
and U5590 (N_5590,N_3276,N_2153);
nor U5591 (N_5591,N_2418,N_2917);
nor U5592 (N_5592,N_3271,N_2814);
nor U5593 (N_5593,N_3023,N_3207);
or U5594 (N_5594,N_3832,N_3817);
nand U5595 (N_5595,N_2077,N_2096);
and U5596 (N_5596,N_3373,N_3729);
or U5597 (N_5597,N_2440,N_2011);
nand U5598 (N_5598,N_3315,N_3229);
nor U5599 (N_5599,N_2460,N_2649);
nand U5600 (N_5600,N_2098,N_3017);
nand U5601 (N_5601,N_3500,N_2214);
nor U5602 (N_5602,N_3473,N_3457);
or U5603 (N_5603,N_3981,N_2384);
and U5604 (N_5604,N_2680,N_2533);
and U5605 (N_5605,N_2184,N_2472);
xor U5606 (N_5606,N_3968,N_3350);
nand U5607 (N_5607,N_2557,N_2463);
and U5608 (N_5608,N_2497,N_3500);
and U5609 (N_5609,N_3744,N_3123);
nor U5610 (N_5610,N_2264,N_3527);
and U5611 (N_5611,N_2435,N_2895);
nand U5612 (N_5612,N_3608,N_3060);
nor U5613 (N_5613,N_2179,N_2932);
nand U5614 (N_5614,N_3520,N_2021);
or U5615 (N_5615,N_3286,N_3958);
nand U5616 (N_5616,N_3083,N_2942);
nor U5617 (N_5617,N_3175,N_3249);
nor U5618 (N_5618,N_3400,N_3821);
and U5619 (N_5619,N_3582,N_2689);
nand U5620 (N_5620,N_3942,N_2017);
or U5621 (N_5621,N_2696,N_3289);
or U5622 (N_5622,N_2425,N_2494);
and U5623 (N_5623,N_3286,N_3538);
and U5624 (N_5624,N_2369,N_2668);
or U5625 (N_5625,N_3981,N_3271);
nor U5626 (N_5626,N_3885,N_3587);
or U5627 (N_5627,N_3391,N_2714);
and U5628 (N_5628,N_3663,N_3674);
nand U5629 (N_5629,N_3874,N_2795);
nand U5630 (N_5630,N_3779,N_2670);
or U5631 (N_5631,N_2518,N_3285);
or U5632 (N_5632,N_3745,N_2630);
nand U5633 (N_5633,N_3483,N_3331);
nor U5634 (N_5634,N_3000,N_2468);
or U5635 (N_5635,N_2933,N_2041);
and U5636 (N_5636,N_2163,N_3842);
nor U5637 (N_5637,N_2432,N_2739);
nor U5638 (N_5638,N_3691,N_3380);
nor U5639 (N_5639,N_3208,N_2653);
and U5640 (N_5640,N_3415,N_2363);
nor U5641 (N_5641,N_2204,N_2427);
nand U5642 (N_5642,N_2603,N_3694);
or U5643 (N_5643,N_2813,N_3189);
nor U5644 (N_5644,N_3143,N_3122);
or U5645 (N_5645,N_2197,N_3681);
and U5646 (N_5646,N_2156,N_3155);
and U5647 (N_5647,N_3119,N_2982);
nor U5648 (N_5648,N_3170,N_3286);
or U5649 (N_5649,N_2711,N_2135);
nand U5650 (N_5650,N_2645,N_2635);
nand U5651 (N_5651,N_3064,N_3194);
nor U5652 (N_5652,N_3236,N_2915);
or U5653 (N_5653,N_3010,N_2666);
and U5654 (N_5654,N_3548,N_2860);
nor U5655 (N_5655,N_2379,N_2291);
or U5656 (N_5656,N_3076,N_2261);
and U5657 (N_5657,N_2693,N_3729);
nor U5658 (N_5658,N_3600,N_2706);
nor U5659 (N_5659,N_2614,N_3562);
nor U5660 (N_5660,N_2349,N_2556);
nor U5661 (N_5661,N_2049,N_3274);
nand U5662 (N_5662,N_2722,N_3483);
nand U5663 (N_5663,N_3499,N_2203);
and U5664 (N_5664,N_2453,N_2018);
xnor U5665 (N_5665,N_2605,N_3356);
nand U5666 (N_5666,N_3879,N_2627);
and U5667 (N_5667,N_2248,N_2635);
xor U5668 (N_5668,N_3700,N_3449);
and U5669 (N_5669,N_3983,N_3984);
or U5670 (N_5670,N_3141,N_3873);
nor U5671 (N_5671,N_2102,N_2729);
xor U5672 (N_5672,N_2547,N_3445);
and U5673 (N_5673,N_2972,N_3432);
and U5674 (N_5674,N_2602,N_2278);
nand U5675 (N_5675,N_2311,N_2321);
nor U5676 (N_5676,N_2726,N_3494);
xor U5677 (N_5677,N_3562,N_3346);
nor U5678 (N_5678,N_2567,N_3384);
xor U5679 (N_5679,N_2528,N_2039);
nor U5680 (N_5680,N_2635,N_3397);
nand U5681 (N_5681,N_3881,N_3298);
nand U5682 (N_5682,N_2266,N_2130);
nand U5683 (N_5683,N_2274,N_3243);
or U5684 (N_5684,N_2936,N_3797);
or U5685 (N_5685,N_2344,N_2431);
nand U5686 (N_5686,N_2775,N_2647);
or U5687 (N_5687,N_3038,N_3340);
or U5688 (N_5688,N_2468,N_2832);
nor U5689 (N_5689,N_2891,N_3190);
or U5690 (N_5690,N_3941,N_2903);
and U5691 (N_5691,N_2001,N_3353);
and U5692 (N_5692,N_2646,N_3088);
xnor U5693 (N_5693,N_3020,N_2711);
nor U5694 (N_5694,N_3936,N_3978);
nor U5695 (N_5695,N_3358,N_2027);
nand U5696 (N_5696,N_3470,N_2966);
or U5697 (N_5697,N_3183,N_2646);
nor U5698 (N_5698,N_3890,N_2012);
nand U5699 (N_5699,N_3918,N_2990);
nor U5700 (N_5700,N_3421,N_3681);
nand U5701 (N_5701,N_3737,N_3189);
and U5702 (N_5702,N_3147,N_3969);
nand U5703 (N_5703,N_3473,N_2121);
or U5704 (N_5704,N_2221,N_2407);
xor U5705 (N_5705,N_3398,N_2813);
or U5706 (N_5706,N_3521,N_3572);
nand U5707 (N_5707,N_2551,N_3968);
nand U5708 (N_5708,N_3872,N_3203);
nor U5709 (N_5709,N_3034,N_2033);
nand U5710 (N_5710,N_2407,N_3897);
nand U5711 (N_5711,N_3952,N_2831);
or U5712 (N_5712,N_3416,N_3404);
xnor U5713 (N_5713,N_3387,N_2240);
nand U5714 (N_5714,N_3671,N_2683);
nor U5715 (N_5715,N_3034,N_3039);
and U5716 (N_5716,N_3267,N_3485);
or U5717 (N_5717,N_3139,N_3641);
nand U5718 (N_5718,N_2666,N_3432);
xor U5719 (N_5719,N_3511,N_2047);
nand U5720 (N_5720,N_3529,N_2333);
xnor U5721 (N_5721,N_2437,N_3090);
nand U5722 (N_5722,N_2328,N_3085);
or U5723 (N_5723,N_2332,N_2087);
or U5724 (N_5724,N_2596,N_2537);
nor U5725 (N_5725,N_3292,N_2358);
nor U5726 (N_5726,N_3551,N_3731);
and U5727 (N_5727,N_3920,N_2848);
and U5728 (N_5728,N_2808,N_3262);
nor U5729 (N_5729,N_3032,N_3490);
and U5730 (N_5730,N_2986,N_2700);
or U5731 (N_5731,N_2762,N_3382);
nand U5732 (N_5732,N_2451,N_3755);
or U5733 (N_5733,N_2421,N_2698);
and U5734 (N_5734,N_3652,N_2654);
or U5735 (N_5735,N_2060,N_3444);
xor U5736 (N_5736,N_2638,N_2288);
nor U5737 (N_5737,N_3559,N_3740);
nor U5738 (N_5738,N_3787,N_3571);
nor U5739 (N_5739,N_3565,N_3275);
nand U5740 (N_5740,N_2444,N_3024);
and U5741 (N_5741,N_2784,N_3186);
or U5742 (N_5742,N_3868,N_2664);
or U5743 (N_5743,N_3392,N_2396);
nand U5744 (N_5744,N_2435,N_2759);
xnor U5745 (N_5745,N_3698,N_2785);
or U5746 (N_5746,N_3278,N_2025);
nand U5747 (N_5747,N_2947,N_3207);
and U5748 (N_5748,N_3213,N_2606);
or U5749 (N_5749,N_3016,N_3305);
nor U5750 (N_5750,N_2686,N_2724);
nor U5751 (N_5751,N_2672,N_2090);
nand U5752 (N_5752,N_2534,N_2023);
xor U5753 (N_5753,N_3764,N_2797);
or U5754 (N_5754,N_3677,N_2562);
nor U5755 (N_5755,N_3749,N_2511);
and U5756 (N_5756,N_3581,N_3865);
nand U5757 (N_5757,N_3018,N_2033);
nor U5758 (N_5758,N_2661,N_3225);
nor U5759 (N_5759,N_2772,N_2103);
nand U5760 (N_5760,N_3166,N_3888);
nor U5761 (N_5761,N_3094,N_2290);
and U5762 (N_5762,N_3220,N_2595);
or U5763 (N_5763,N_3907,N_2454);
or U5764 (N_5764,N_2618,N_3957);
or U5765 (N_5765,N_2952,N_3625);
nand U5766 (N_5766,N_2474,N_3476);
and U5767 (N_5767,N_2556,N_3801);
nand U5768 (N_5768,N_3220,N_2157);
nor U5769 (N_5769,N_2768,N_3020);
xor U5770 (N_5770,N_2264,N_2695);
nor U5771 (N_5771,N_3184,N_3393);
nand U5772 (N_5772,N_2406,N_2123);
xor U5773 (N_5773,N_3068,N_2639);
nand U5774 (N_5774,N_3315,N_3011);
and U5775 (N_5775,N_3027,N_3655);
xnor U5776 (N_5776,N_2562,N_2306);
or U5777 (N_5777,N_2256,N_3708);
or U5778 (N_5778,N_3733,N_2712);
or U5779 (N_5779,N_3104,N_3609);
and U5780 (N_5780,N_3475,N_2636);
or U5781 (N_5781,N_3499,N_2759);
xnor U5782 (N_5782,N_3575,N_2615);
and U5783 (N_5783,N_3958,N_3861);
nand U5784 (N_5784,N_2548,N_3342);
nand U5785 (N_5785,N_2168,N_2209);
nand U5786 (N_5786,N_3669,N_2136);
and U5787 (N_5787,N_2699,N_2429);
nor U5788 (N_5788,N_2525,N_2531);
nor U5789 (N_5789,N_3303,N_2680);
and U5790 (N_5790,N_2589,N_3197);
or U5791 (N_5791,N_3903,N_2025);
nor U5792 (N_5792,N_2357,N_2395);
nor U5793 (N_5793,N_3546,N_2139);
and U5794 (N_5794,N_2534,N_2118);
or U5795 (N_5795,N_2029,N_2533);
nor U5796 (N_5796,N_3055,N_3641);
or U5797 (N_5797,N_3727,N_3233);
or U5798 (N_5798,N_3613,N_2208);
and U5799 (N_5799,N_2028,N_3635);
or U5800 (N_5800,N_3923,N_3712);
or U5801 (N_5801,N_3062,N_2080);
xor U5802 (N_5802,N_2435,N_3904);
nand U5803 (N_5803,N_3409,N_2735);
nor U5804 (N_5804,N_3394,N_2905);
and U5805 (N_5805,N_2204,N_2297);
nand U5806 (N_5806,N_3673,N_3224);
or U5807 (N_5807,N_2534,N_3588);
or U5808 (N_5808,N_3983,N_2107);
and U5809 (N_5809,N_3489,N_2105);
nand U5810 (N_5810,N_3970,N_3648);
or U5811 (N_5811,N_2612,N_2964);
or U5812 (N_5812,N_2968,N_2586);
or U5813 (N_5813,N_3874,N_3962);
and U5814 (N_5814,N_2552,N_2604);
and U5815 (N_5815,N_3781,N_2044);
or U5816 (N_5816,N_3272,N_2026);
or U5817 (N_5817,N_3063,N_2238);
xor U5818 (N_5818,N_3378,N_2215);
or U5819 (N_5819,N_2766,N_3345);
or U5820 (N_5820,N_2707,N_3683);
or U5821 (N_5821,N_2705,N_3713);
xor U5822 (N_5822,N_3258,N_3714);
xnor U5823 (N_5823,N_2294,N_3671);
and U5824 (N_5824,N_2761,N_3180);
nand U5825 (N_5825,N_3282,N_2841);
and U5826 (N_5826,N_3874,N_3934);
or U5827 (N_5827,N_3109,N_3017);
nor U5828 (N_5828,N_3787,N_2355);
nand U5829 (N_5829,N_2369,N_2658);
or U5830 (N_5830,N_2990,N_2926);
or U5831 (N_5831,N_2834,N_2794);
or U5832 (N_5832,N_2984,N_2053);
nor U5833 (N_5833,N_2187,N_2724);
xor U5834 (N_5834,N_3813,N_3283);
or U5835 (N_5835,N_2204,N_2410);
xnor U5836 (N_5836,N_3648,N_2112);
and U5837 (N_5837,N_2754,N_3540);
and U5838 (N_5838,N_3983,N_3962);
nand U5839 (N_5839,N_3210,N_2409);
nand U5840 (N_5840,N_3536,N_2042);
nor U5841 (N_5841,N_2800,N_2561);
and U5842 (N_5842,N_3261,N_2508);
xor U5843 (N_5843,N_3343,N_3056);
nand U5844 (N_5844,N_3380,N_2223);
nor U5845 (N_5845,N_3299,N_3303);
nor U5846 (N_5846,N_2918,N_2827);
nor U5847 (N_5847,N_3908,N_3181);
or U5848 (N_5848,N_3280,N_3648);
nand U5849 (N_5849,N_3141,N_2200);
nor U5850 (N_5850,N_3136,N_2013);
and U5851 (N_5851,N_3650,N_3211);
nor U5852 (N_5852,N_3361,N_3060);
xor U5853 (N_5853,N_3132,N_3181);
xor U5854 (N_5854,N_2381,N_3349);
or U5855 (N_5855,N_3951,N_2521);
xor U5856 (N_5856,N_2147,N_3045);
nor U5857 (N_5857,N_3361,N_3270);
nand U5858 (N_5858,N_2218,N_3445);
and U5859 (N_5859,N_3669,N_2547);
nor U5860 (N_5860,N_2638,N_3902);
nor U5861 (N_5861,N_3321,N_3052);
nor U5862 (N_5862,N_2449,N_3963);
and U5863 (N_5863,N_3536,N_2675);
nand U5864 (N_5864,N_3347,N_2831);
nand U5865 (N_5865,N_3185,N_2672);
nand U5866 (N_5866,N_3040,N_3369);
and U5867 (N_5867,N_3926,N_2796);
or U5868 (N_5868,N_3452,N_3774);
or U5869 (N_5869,N_3507,N_2502);
nor U5870 (N_5870,N_3994,N_3586);
nand U5871 (N_5871,N_3696,N_2925);
and U5872 (N_5872,N_3956,N_3120);
and U5873 (N_5873,N_3528,N_2465);
nand U5874 (N_5874,N_2397,N_2371);
and U5875 (N_5875,N_2579,N_2757);
nand U5876 (N_5876,N_3844,N_2166);
and U5877 (N_5877,N_2391,N_3330);
nor U5878 (N_5878,N_3838,N_3843);
nor U5879 (N_5879,N_2669,N_2709);
nand U5880 (N_5880,N_3397,N_3270);
and U5881 (N_5881,N_3284,N_2744);
and U5882 (N_5882,N_3851,N_2209);
and U5883 (N_5883,N_2805,N_2089);
nor U5884 (N_5884,N_3737,N_3069);
or U5885 (N_5885,N_2213,N_3929);
xor U5886 (N_5886,N_3905,N_3147);
or U5887 (N_5887,N_2728,N_3355);
or U5888 (N_5888,N_3008,N_3504);
nor U5889 (N_5889,N_3192,N_3529);
or U5890 (N_5890,N_3144,N_2533);
and U5891 (N_5891,N_3578,N_3569);
and U5892 (N_5892,N_2919,N_2908);
and U5893 (N_5893,N_2111,N_2523);
or U5894 (N_5894,N_2746,N_3314);
nor U5895 (N_5895,N_2763,N_3358);
nor U5896 (N_5896,N_3775,N_2604);
nor U5897 (N_5897,N_3873,N_2701);
or U5898 (N_5898,N_2803,N_2243);
or U5899 (N_5899,N_3910,N_2712);
xnor U5900 (N_5900,N_3109,N_3812);
nand U5901 (N_5901,N_3699,N_2079);
nor U5902 (N_5902,N_2864,N_2755);
and U5903 (N_5903,N_2452,N_3852);
and U5904 (N_5904,N_2398,N_3615);
nor U5905 (N_5905,N_3533,N_2689);
nand U5906 (N_5906,N_3493,N_3412);
nand U5907 (N_5907,N_3657,N_3356);
nor U5908 (N_5908,N_2010,N_3706);
or U5909 (N_5909,N_3143,N_2816);
nor U5910 (N_5910,N_2986,N_3657);
nand U5911 (N_5911,N_2502,N_3542);
and U5912 (N_5912,N_2963,N_3519);
nor U5913 (N_5913,N_2878,N_2596);
nand U5914 (N_5914,N_2154,N_3757);
nand U5915 (N_5915,N_2578,N_2876);
or U5916 (N_5916,N_3021,N_2477);
or U5917 (N_5917,N_2162,N_2283);
nor U5918 (N_5918,N_3356,N_2896);
and U5919 (N_5919,N_2392,N_2817);
and U5920 (N_5920,N_3552,N_2730);
xnor U5921 (N_5921,N_3821,N_3585);
nor U5922 (N_5922,N_2164,N_3807);
nor U5923 (N_5923,N_3043,N_3606);
nand U5924 (N_5924,N_2200,N_3721);
or U5925 (N_5925,N_2637,N_3345);
nand U5926 (N_5926,N_3172,N_2555);
nor U5927 (N_5927,N_3543,N_2239);
or U5928 (N_5928,N_3731,N_3792);
nand U5929 (N_5929,N_3512,N_2805);
xnor U5930 (N_5930,N_3435,N_2446);
nor U5931 (N_5931,N_3099,N_3264);
and U5932 (N_5932,N_3949,N_2377);
or U5933 (N_5933,N_3064,N_3872);
nand U5934 (N_5934,N_3674,N_3398);
nand U5935 (N_5935,N_3116,N_2624);
nand U5936 (N_5936,N_3030,N_3448);
nor U5937 (N_5937,N_3271,N_3259);
xnor U5938 (N_5938,N_2804,N_2744);
or U5939 (N_5939,N_3367,N_2497);
and U5940 (N_5940,N_3548,N_3125);
and U5941 (N_5941,N_2307,N_3912);
and U5942 (N_5942,N_3205,N_2812);
nand U5943 (N_5943,N_3856,N_3583);
or U5944 (N_5944,N_3487,N_2402);
or U5945 (N_5945,N_2400,N_3026);
and U5946 (N_5946,N_3002,N_3132);
nor U5947 (N_5947,N_2762,N_2573);
and U5948 (N_5948,N_3475,N_3636);
nor U5949 (N_5949,N_2160,N_2848);
and U5950 (N_5950,N_2813,N_3580);
nand U5951 (N_5951,N_3126,N_3557);
and U5952 (N_5952,N_2762,N_2180);
and U5953 (N_5953,N_2156,N_3833);
or U5954 (N_5954,N_2081,N_2870);
and U5955 (N_5955,N_3674,N_2254);
xnor U5956 (N_5956,N_3522,N_3665);
and U5957 (N_5957,N_3625,N_2377);
nand U5958 (N_5958,N_3192,N_3473);
and U5959 (N_5959,N_2047,N_3380);
nor U5960 (N_5960,N_3214,N_2036);
or U5961 (N_5961,N_2947,N_3967);
or U5962 (N_5962,N_2307,N_3689);
and U5963 (N_5963,N_2012,N_2021);
and U5964 (N_5964,N_2612,N_2122);
or U5965 (N_5965,N_2878,N_3060);
or U5966 (N_5966,N_2462,N_2222);
and U5967 (N_5967,N_3884,N_3148);
nor U5968 (N_5968,N_2575,N_3223);
or U5969 (N_5969,N_2616,N_2968);
and U5970 (N_5970,N_2185,N_2571);
and U5971 (N_5971,N_2166,N_2413);
xnor U5972 (N_5972,N_3685,N_3194);
nor U5973 (N_5973,N_2330,N_3126);
and U5974 (N_5974,N_3383,N_3454);
xor U5975 (N_5975,N_2021,N_2219);
or U5976 (N_5976,N_2703,N_3864);
nand U5977 (N_5977,N_2305,N_2810);
nor U5978 (N_5978,N_2203,N_2910);
and U5979 (N_5979,N_2206,N_2360);
or U5980 (N_5980,N_3773,N_3718);
and U5981 (N_5981,N_2526,N_3323);
and U5982 (N_5982,N_2217,N_2404);
or U5983 (N_5983,N_2467,N_3414);
or U5984 (N_5984,N_2085,N_2543);
and U5985 (N_5985,N_2637,N_2915);
nand U5986 (N_5986,N_2014,N_2372);
or U5987 (N_5987,N_2659,N_2895);
nor U5988 (N_5988,N_2904,N_3388);
nand U5989 (N_5989,N_3174,N_3698);
or U5990 (N_5990,N_2556,N_3457);
or U5991 (N_5991,N_3786,N_2172);
nand U5992 (N_5992,N_2241,N_3620);
or U5993 (N_5993,N_2541,N_3748);
nor U5994 (N_5994,N_3860,N_2263);
nor U5995 (N_5995,N_3856,N_2337);
nand U5996 (N_5996,N_2572,N_2275);
xnor U5997 (N_5997,N_3869,N_3870);
or U5998 (N_5998,N_2047,N_3928);
nand U5999 (N_5999,N_2103,N_3537);
and U6000 (N_6000,N_4477,N_5131);
nand U6001 (N_6001,N_4705,N_5578);
nand U6002 (N_6002,N_4579,N_5859);
and U6003 (N_6003,N_4243,N_5823);
and U6004 (N_6004,N_5213,N_5776);
nor U6005 (N_6005,N_5509,N_4524);
nand U6006 (N_6006,N_5898,N_5928);
nand U6007 (N_6007,N_5821,N_5433);
nand U6008 (N_6008,N_4887,N_4924);
nor U6009 (N_6009,N_4922,N_5956);
or U6010 (N_6010,N_5865,N_5669);
and U6011 (N_6011,N_4398,N_4874);
and U6012 (N_6012,N_5701,N_4995);
and U6013 (N_6013,N_5276,N_4619);
and U6014 (N_6014,N_4960,N_5263);
nand U6015 (N_6015,N_4590,N_5251);
nor U6016 (N_6016,N_5296,N_5284);
nand U6017 (N_6017,N_5930,N_4907);
nand U6018 (N_6018,N_4656,N_4645);
nor U6019 (N_6019,N_4510,N_5222);
or U6020 (N_6020,N_5507,N_4967);
nand U6021 (N_6021,N_4839,N_4739);
nor U6022 (N_6022,N_4013,N_4559);
nor U6023 (N_6023,N_5416,N_4220);
xor U6024 (N_6024,N_4991,N_4728);
or U6025 (N_6025,N_4657,N_4555);
or U6026 (N_6026,N_5958,N_5918);
nand U6027 (N_6027,N_5711,N_5972);
xor U6028 (N_6028,N_5603,N_4878);
and U6029 (N_6029,N_4517,N_4153);
nor U6030 (N_6030,N_4148,N_4060);
nand U6031 (N_6031,N_5627,N_5818);
or U6032 (N_6032,N_4514,N_4549);
nor U6033 (N_6033,N_4344,N_4411);
nor U6034 (N_6034,N_4568,N_5656);
and U6035 (N_6035,N_5550,N_4198);
nor U6036 (N_6036,N_4968,N_5308);
nand U6037 (N_6037,N_5620,N_4055);
or U6038 (N_6038,N_5986,N_4953);
nor U6039 (N_6039,N_4276,N_5531);
xor U6040 (N_6040,N_5867,N_5607);
xnor U6041 (N_6041,N_4342,N_4004);
nor U6042 (N_6042,N_5574,N_4377);
nor U6043 (N_6043,N_5992,N_5398);
or U6044 (N_6044,N_4522,N_5408);
and U6045 (N_6045,N_4070,N_5758);
nand U6046 (N_6046,N_4025,N_4719);
and U6047 (N_6047,N_4942,N_4260);
and U6048 (N_6048,N_4600,N_5070);
and U6049 (N_6049,N_4999,N_4893);
nand U6050 (N_6050,N_4591,N_4012);
and U6051 (N_6051,N_4241,N_5193);
nand U6052 (N_6052,N_4604,N_5725);
and U6053 (N_6053,N_5185,N_4875);
or U6054 (N_6054,N_5490,N_4184);
and U6055 (N_6055,N_4867,N_5526);
xor U6056 (N_6056,N_5335,N_4601);
or U6057 (N_6057,N_5011,N_5508);
nand U6058 (N_6058,N_4786,N_5318);
nand U6059 (N_6059,N_5941,N_4468);
or U6060 (N_6060,N_5903,N_5896);
nor U6061 (N_6061,N_4981,N_5617);
or U6062 (N_6062,N_4909,N_4677);
or U6063 (N_6063,N_5741,N_5740);
nand U6064 (N_6064,N_4481,N_4159);
nor U6065 (N_6065,N_4445,N_4102);
nor U6066 (N_6066,N_4833,N_5238);
or U6067 (N_6067,N_4714,N_4262);
xnor U6068 (N_6068,N_5583,N_5947);
and U6069 (N_6069,N_4441,N_5180);
and U6070 (N_6070,N_4296,N_5715);
nor U6071 (N_6071,N_5114,N_4862);
or U6072 (N_6072,N_4743,N_4024);
or U6073 (N_6073,N_4817,N_5889);
or U6074 (N_6074,N_4501,N_5040);
or U6075 (N_6075,N_5570,N_4451);
nor U6076 (N_6076,N_4882,N_5935);
xnor U6077 (N_6077,N_5932,N_4438);
or U6078 (N_6078,N_4765,N_5985);
nand U6079 (N_6079,N_5913,N_4808);
or U6080 (N_6080,N_4941,N_4248);
nand U6081 (N_6081,N_5475,N_4630);
or U6082 (N_6082,N_4515,N_5563);
nor U6083 (N_6083,N_5236,N_4454);
xnor U6084 (N_6084,N_4574,N_5658);
nor U6085 (N_6085,N_4672,N_5220);
and U6086 (N_6086,N_4972,N_5478);
and U6087 (N_6087,N_4338,N_5053);
xnor U6088 (N_6088,N_4232,N_4927);
or U6089 (N_6089,N_4300,N_4780);
and U6090 (N_6090,N_4416,N_4382);
or U6091 (N_6091,N_4368,N_4309);
nor U6092 (N_6092,N_4230,N_4208);
or U6093 (N_6093,N_5469,N_4692);
and U6094 (N_6094,N_4312,N_4353);
nor U6095 (N_6095,N_5397,N_4422);
and U6096 (N_6096,N_5424,N_5439);
or U6097 (N_6097,N_5144,N_4035);
nor U6098 (N_6098,N_4031,N_4831);
or U6099 (N_6099,N_4150,N_5780);
nand U6100 (N_6100,N_4412,N_4879);
nand U6101 (N_6101,N_5927,N_5165);
and U6102 (N_6102,N_4162,N_5218);
nor U6103 (N_6103,N_4059,N_5227);
nor U6104 (N_6104,N_5179,N_4166);
nand U6105 (N_6105,N_4538,N_4550);
nor U6106 (N_6106,N_4583,N_5366);
and U6107 (N_6107,N_5018,N_4043);
nor U6108 (N_6108,N_4014,N_4302);
nand U6109 (N_6109,N_5266,N_4211);
nor U6110 (N_6110,N_5072,N_5784);
and U6111 (N_6111,N_5599,N_5606);
or U6112 (N_6112,N_5019,N_5571);
and U6113 (N_6113,N_5094,N_4572);
nor U6114 (N_6114,N_5733,N_5565);
xor U6115 (N_6115,N_5997,N_4023);
nand U6116 (N_6116,N_5166,N_5501);
or U6117 (N_6117,N_4897,N_4753);
or U6118 (N_6118,N_4815,N_4824);
nand U6119 (N_6119,N_4401,N_4969);
nand U6120 (N_6120,N_5737,N_5510);
nor U6121 (N_6121,N_4192,N_4744);
nor U6122 (N_6122,N_5000,N_5857);
nor U6123 (N_6123,N_5499,N_5077);
and U6124 (N_6124,N_5003,N_5175);
nor U6125 (N_6125,N_4201,N_5736);
nand U6126 (N_6126,N_4493,N_4320);
or U6127 (N_6127,N_4627,N_5204);
xor U6128 (N_6128,N_4337,N_5217);
and U6129 (N_6129,N_4877,N_4852);
or U6130 (N_6130,N_5500,N_5128);
and U6131 (N_6131,N_5703,N_4284);
or U6132 (N_6132,N_5329,N_5528);
or U6133 (N_6133,N_5641,N_5259);
xnor U6134 (N_6134,N_5436,N_5451);
or U6135 (N_6135,N_4779,N_5315);
and U6136 (N_6136,N_5517,N_4135);
or U6137 (N_6137,N_4912,N_4101);
nor U6138 (N_6138,N_4567,N_5484);
nand U6139 (N_6139,N_5624,N_5240);
or U6140 (N_6140,N_5016,N_4233);
and U6141 (N_6141,N_4492,N_4499);
nor U6142 (N_6142,N_5904,N_4247);
xnor U6143 (N_6143,N_5172,N_5730);
xnor U6144 (N_6144,N_4904,N_5893);
and U6145 (N_6145,N_5846,N_5886);
and U6146 (N_6146,N_5026,N_5468);
nand U6147 (N_6147,N_5549,N_4266);
or U6148 (N_6148,N_5769,N_4527);
and U6149 (N_6149,N_5153,N_4997);
nand U6150 (N_6150,N_4327,N_4142);
and U6151 (N_6151,N_4027,N_5540);
nand U6152 (N_6152,N_4678,N_5502);
nand U6153 (N_6153,N_5303,N_5147);
or U6154 (N_6154,N_4303,N_5618);
and U6155 (N_6155,N_5158,N_4740);
and U6156 (N_6156,N_5432,N_4446);
xnor U6157 (N_6157,N_4890,N_5581);
nor U6158 (N_6158,N_5545,N_5404);
xor U6159 (N_6159,N_5515,N_4239);
nand U6160 (N_6160,N_5243,N_4116);
nand U6161 (N_6161,N_5285,N_5321);
nor U6162 (N_6162,N_4990,N_5208);
or U6163 (N_6163,N_4206,N_5721);
xnor U6164 (N_6164,N_4378,N_4305);
nor U6165 (N_6165,N_4749,N_4461);
or U6166 (N_6166,N_4330,N_4745);
or U6167 (N_6167,N_5562,N_4397);
nor U6168 (N_6168,N_4127,N_4996);
or U6169 (N_6169,N_5024,N_4970);
nor U6170 (N_6170,N_5148,N_5134);
and U6171 (N_6171,N_5901,N_5648);
xnor U6172 (N_6172,N_5173,N_5640);
nor U6173 (N_6173,N_4222,N_4623);
and U6174 (N_6174,N_5497,N_5378);
and U6175 (N_6175,N_4103,N_4058);
and U6176 (N_6176,N_4314,N_4006);
and U6177 (N_6177,N_5911,N_4372);
nand U6178 (N_6178,N_4690,N_5386);
and U6179 (N_6179,N_5761,N_5727);
and U6180 (N_6180,N_5446,N_5105);
and U6181 (N_6181,N_5108,N_4662);
or U6182 (N_6182,N_5664,N_5281);
nand U6183 (N_6183,N_5113,N_5435);
nand U6184 (N_6184,N_4861,N_4959);
or U6185 (N_6185,N_4729,N_5852);
xnor U6186 (N_6186,N_5677,N_5504);
nor U6187 (N_6187,N_4005,N_5413);
or U6188 (N_6188,N_4008,N_5023);
nand U6189 (N_6189,N_5075,N_4435);
nand U6190 (N_6190,N_4773,N_4784);
and U6191 (N_6191,N_5773,N_5112);
or U6192 (N_6192,N_5407,N_5798);
and U6193 (N_6193,N_5010,N_4646);
or U6194 (N_6194,N_4597,N_4074);
and U6195 (N_6195,N_5048,N_5529);
or U6196 (N_6196,N_4557,N_4424);
and U6197 (N_6197,N_5051,N_5327);
and U6198 (N_6198,N_4195,N_4843);
xnor U6199 (N_6199,N_4563,N_4731);
and U6200 (N_6200,N_5316,N_4631);
nand U6201 (N_6201,N_5861,N_4383);
nor U6202 (N_6202,N_5096,N_5675);
or U6203 (N_6203,N_4225,N_5044);
xor U6204 (N_6204,N_5091,N_4180);
nor U6205 (N_6205,N_4654,N_4902);
or U6206 (N_6206,N_4380,N_4847);
and U6207 (N_6207,N_5709,N_5860);
or U6208 (N_6208,N_4310,N_4123);
or U6209 (N_6209,N_4287,N_5399);
nand U6210 (N_6210,N_4947,N_4506);
and U6211 (N_6211,N_5788,N_4850);
nor U6212 (N_6212,N_5961,N_4571);
and U6213 (N_6213,N_4291,N_4029);
nor U6214 (N_6214,N_5577,N_5965);
and U6215 (N_6215,N_4836,N_5665);
and U6216 (N_6216,N_4275,N_4525);
and U6217 (N_6217,N_4323,N_4781);
and U6218 (N_6218,N_5748,N_5001);
nand U6219 (N_6219,N_5631,N_5920);
nand U6220 (N_6220,N_4532,N_5789);
and U6221 (N_6221,N_5199,N_4444);
nand U6222 (N_6222,N_5184,N_5899);
nand U6223 (N_6223,N_4044,N_5045);
or U6224 (N_6224,N_5483,N_5155);
xnor U6225 (N_6225,N_5305,N_5628);
and U6226 (N_6226,N_5383,N_4292);
nand U6227 (N_6227,N_5560,N_5167);
nor U6228 (N_6228,N_5879,N_4431);
or U6229 (N_6229,N_4294,N_5306);
xnor U6230 (N_6230,N_4119,N_4387);
nand U6231 (N_6231,N_5356,N_4668);
xnor U6232 (N_6232,N_4581,N_5004);
nor U6233 (N_6233,N_5200,N_5568);
nor U6234 (N_6234,N_4226,N_5120);
or U6235 (N_6235,N_4139,N_4428);
and U6236 (N_6236,N_4189,N_5360);
nor U6237 (N_6237,N_5792,N_5286);
and U6238 (N_6238,N_4639,N_5696);
xor U6239 (N_6239,N_4760,N_5104);
or U6240 (N_6240,N_4965,N_5950);
or U6241 (N_6241,N_4828,N_4526);
nor U6242 (N_6242,N_5519,N_4939);
nand U6243 (N_6243,N_4174,N_4873);
nand U6244 (N_6244,N_4482,N_4702);
nor U6245 (N_6245,N_4315,N_4820);
nand U6246 (N_6246,N_4202,N_4485);
and U6247 (N_6247,N_4573,N_5659);
and U6248 (N_6248,N_5754,N_4569);
nor U6249 (N_6249,N_5385,N_4234);
or U6250 (N_6250,N_4066,N_5007);
nor U6251 (N_6251,N_4178,N_5968);
nand U6252 (N_6252,N_4010,N_5833);
nor U6253 (N_6253,N_5834,N_4280);
or U6254 (N_6254,N_5520,N_4696);
and U6255 (N_6255,N_5270,N_4437);
nor U6256 (N_6256,N_4976,N_4011);
xnor U6257 (N_6257,N_4405,N_4134);
xnor U6258 (N_6258,N_5216,N_5351);
nor U6259 (N_6259,N_4715,N_5197);
and U6260 (N_6260,N_5336,N_4084);
or U6261 (N_6261,N_4293,N_4339);
nor U6262 (N_6262,N_4210,N_4876);
nand U6263 (N_6263,N_4761,N_5869);
or U6264 (N_6264,N_4994,N_4295);
nand U6265 (N_6265,N_5422,N_4727);
and U6266 (N_6266,N_4319,N_5393);
nand U6267 (N_6267,N_5461,N_5738);
and U6268 (N_6268,N_4316,N_4754);
xor U6269 (N_6269,N_4673,N_4472);
nor U6270 (N_6270,N_4980,N_4707);
and U6271 (N_6271,N_5592,N_5731);
nor U6272 (N_6272,N_5826,N_5202);
nand U6273 (N_6273,N_4795,N_4341);
and U6274 (N_6274,N_5492,N_4722);
and U6275 (N_6275,N_4270,N_5460);
nor U6276 (N_6276,N_4486,N_4950);
or U6277 (N_6277,N_5015,N_5609);
or U6278 (N_6278,N_5625,N_4889);
or U6279 (N_6279,N_4062,N_5396);
and U6280 (N_6280,N_5729,N_4124);
nor U6281 (N_6281,N_4157,N_4973);
nor U6282 (N_6282,N_4307,N_5850);
or U6283 (N_6283,N_4512,N_4271);
or U6284 (N_6284,N_5143,N_4399);
and U6285 (N_6285,N_4089,N_4735);
nand U6286 (N_6286,N_5192,N_5099);
nand U6287 (N_6287,N_5699,N_4078);
or U6288 (N_6288,N_5829,N_5002);
xor U6289 (N_6289,N_4957,N_4214);
nor U6290 (N_6290,N_5489,N_4450);
nor U6291 (N_6291,N_4746,N_4511);
or U6292 (N_6292,N_5714,N_5931);
or U6293 (N_6293,N_5645,N_4603);
and U6294 (N_6294,N_5837,N_4496);
nor U6295 (N_6295,N_4643,N_4229);
nor U6296 (N_6296,N_4859,N_5816);
xor U6297 (N_6297,N_5800,N_5843);
and U6298 (N_6298,N_4509,N_5839);
nor U6299 (N_6299,N_4865,N_5410);
nand U6300 (N_6300,N_4164,N_4177);
xor U6301 (N_6301,N_4465,N_5635);
nor U6302 (N_6302,N_4389,N_5514);
or U6303 (N_6303,N_4548,N_5300);
and U6304 (N_6304,N_5323,N_4082);
or U6305 (N_6305,N_4594,N_4317);
and U6306 (N_6306,N_4434,N_4151);
nand U6307 (N_6307,N_4268,N_5875);
or U6308 (N_6308,N_4863,N_5226);
xor U6309 (N_6309,N_5417,N_4975);
nor U6310 (N_6310,N_4483,N_5629);
nor U6311 (N_6311,N_5479,N_5566);
and U6312 (N_6312,N_5851,N_5427);
or U6313 (N_6313,N_4608,N_5457);
and U6314 (N_6314,N_5589,N_4423);
or U6315 (N_6315,N_4580,N_4329);
nor U6316 (N_6316,N_5496,N_5473);
or U6317 (N_6317,N_4217,N_4986);
nand U6318 (N_6318,N_5052,N_4194);
or U6319 (N_6319,N_5674,N_4653);
and U6320 (N_6320,N_4279,N_4750);
nor U6321 (N_6321,N_4708,N_5041);
xor U6322 (N_6322,N_5275,N_4647);
nor U6323 (N_6323,N_4456,N_5543);
nor U6324 (N_6324,N_4365,N_4348);
and U6325 (N_6325,N_4856,N_4263);
nor U6326 (N_6326,N_5981,N_5732);
nor U6327 (N_6327,N_4562,N_4622);
and U6328 (N_6328,N_4688,N_4938);
nand U6329 (N_6329,N_4682,N_5828);
and U6330 (N_6330,N_4855,N_4609);
nor U6331 (N_6331,N_5842,N_5313);
nand U6332 (N_6332,N_4962,N_5081);
nand U6333 (N_6333,N_4872,N_5890);
nor U6334 (N_6334,N_4686,N_4885);
and U6335 (N_6335,N_4469,N_5279);
xor U6336 (N_6336,N_4350,N_4846);
or U6337 (N_6337,N_5434,N_5146);
or U6338 (N_6338,N_4738,N_4899);
xor U6339 (N_6339,N_4479,N_4057);
or U6340 (N_6340,N_5121,N_5685);
nor U6341 (N_6341,N_4473,N_4711);
xor U6342 (N_6342,N_4274,N_5066);
and U6343 (N_6343,N_4290,N_5298);
nand U6344 (N_6344,N_4063,N_5764);
xor U6345 (N_6345,N_5812,N_5666);
nor U6346 (N_6346,N_5678,N_4989);
or U6347 (N_6347,N_5778,N_4545);
xnor U6348 (N_6348,N_4179,N_4018);
or U6349 (N_6349,N_5786,N_4787);
nor U6350 (N_6350,N_5363,N_5759);
nor U6351 (N_6351,N_4611,N_4388);
nor U6352 (N_6352,N_5916,N_5722);
or U6353 (N_6353,N_4193,N_5633);
nor U6354 (N_6354,N_5459,N_5274);
nand U6355 (N_6355,N_4810,N_4851);
nand U6356 (N_6356,N_5785,N_4724);
xor U6357 (N_6357,N_5106,N_4768);
xnor U6358 (N_6358,N_5705,N_5750);
and U6359 (N_6359,N_4935,N_4625);
and U6360 (N_6360,N_5505,N_5177);
xor U6361 (N_6361,N_5814,N_5485);
xor U6362 (N_6362,N_5803,N_5389);
xnor U6363 (N_6363,N_5588,N_4649);
and U6364 (N_6364,N_5743,N_4258);
nor U6365 (N_6365,N_4118,N_5337);
and U6366 (N_6366,N_4841,N_4026);
and U6367 (N_6367,N_5720,N_4204);
or U6368 (N_6368,N_4945,N_5744);
nor U6369 (N_6369,N_5999,N_4832);
or U6370 (N_6370,N_4183,N_4440);
nand U6371 (N_6371,N_5576,N_5988);
nor U6372 (N_6372,N_4369,N_4886);
nand U6373 (N_6373,N_4447,N_5832);
or U6374 (N_6374,N_4072,N_5283);
nor U6375 (N_6375,N_5982,N_4905);
and U6376 (N_6376,N_5195,N_5320);
or U6377 (N_6377,N_5855,N_5799);
nand U6378 (N_6378,N_5116,N_4598);
or U6379 (N_6379,N_5029,N_5572);
xnor U6380 (N_6380,N_4704,N_4659);
and U6381 (N_6381,N_5353,N_4663);
or U6382 (N_6382,N_5595,N_5888);
nand U6383 (N_6383,N_5511,N_4925);
nor U6384 (N_6384,N_5256,N_5845);
nand U6385 (N_6385,N_4073,N_5174);
nor U6386 (N_6386,N_5486,N_4826);
nor U6387 (N_6387,N_4126,N_4147);
nand U6388 (N_6388,N_5157,N_4956);
nand U6389 (N_6389,N_5912,N_4149);
nand U6390 (N_6390,N_4932,N_4710);
nand U6391 (N_6391,N_4106,N_5698);
nand U6392 (N_6392,N_5753,N_5718);
nand U6393 (N_6393,N_4117,N_4409);
nand U6394 (N_6394,N_5097,N_5723);
and U6395 (N_6395,N_4895,N_4634);
xnor U6396 (N_6396,N_4910,N_5244);
nand U6397 (N_6397,N_5819,N_4536);
or U6398 (N_6398,N_5466,N_5159);
or U6399 (N_6399,N_5462,N_5414);
and U6400 (N_6400,N_5960,N_5293);
or U6401 (N_6401,N_5995,N_4671);
or U6402 (N_6402,N_4720,N_4531);
or U6403 (N_6403,N_4046,N_4079);
xnor U6404 (N_6404,N_4362,N_5013);
or U6405 (N_6405,N_5373,N_4065);
nor U6406 (N_6406,N_4616,N_5067);
nand U6407 (N_6407,N_5973,N_4652);
nor U6408 (N_6408,N_5169,N_5268);
or U6409 (N_6409,N_5838,N_4666);
nor U6410 (N_6410,N_5394,N_5584);
nand U6411 (N_6411,N_4094,N_4617);
xor U6412 (N_6412,N_5940,N_4054);
nor U6413 (N_6413,N_5951,N_5152);
nor U6414 (N_6414,N_5235,N_5171);
nand U6415 (N_6415,N_4811,N_4977);
and U6416 (N_6416,N_5591,N_5984);
nor U6417 (N_6417,N_5391,N_4791);
nand U6418 (N_6418,N_5253,N_4050);
nand U6419 (N_6419,N_5194,N_5807);
xnor U6420 (N_6420,N_5343,N_5921);
nor U6421 (N_6421,N_5371,N_5516);
nand U6422 (N_6422,N_5034,N_4758);
xor U6423 (N_6423,N_5110,N_4929);
and U6424 (N_6424,N_4186,N_4529);
or U6425 (N_6425,N_5506,N_5684);
and U6426 (N_6426,N_4769,N_5221);
nor U6427 (N_6427,N_5437,N_4086);
nor U6428 (N_6428,N_5975,N_5269);
nor U6429 (N_6429,N_5690,N_4191);
and U6430 (N_6430,N_5757,N_5512);
xor U6431 (N_6431,N_4570,N_5555);
and U6432 (N_6432,N_4576,N_4311);
nand U6433 (N_6433,N_5670,N_4931);
and U6434 (N_6434,N_5687,N_5909);
nand U6435 (N_6435,N_4528,N_5450);
xor U6436 (N_6436,N_5746,N_5206);
or U6437 (N_6437,N_4114,N_4543);
and U6438 (N_6438,N_4726,N_4488);
or U6439 (N_6439,N_4442,N_4381);
or U6440 (N_6440,N_4056,N_5442);
nand U6441 (N_6441,N_5693,N_5210);
and U6442 (N_6442,N_5418,N_5919);
nand U6443 (N_6443,N_4009,N_5022);
nand U6444 (N_6444,N_5564,N_4301);
nor U6445 (N_6445,N_5035,N_4624);
nor U6446 (N_6446,N_4170,N_5639);
nor U6447 (N_6447,N_5957,N_4099);
or U6448 (N_6448,N_4644,N_4415);
or U6449 (N_6449,N_5125,N_5074);
and U6450 (N_6450,N_4595,N_5594);
nand U6451 (N_6451,N_5060,N_4252);
and U6452 (N_6452,N_5644,N_5561);
or U6453 (N_6453,N_4407,N_4100);
nor U6454 (N_6454,N_4508,N_5247);
nor U6455 (N_6455,N_4593,N_5805);
or U6456 (N_6456,N_5554,N_5419);
nand U6457 (N_6457,N_4534,N_4667);
and U6458 (N_6458,N_4869,N_4813);
nor U6459 (N_6459,N_4694,N_4200);
xor U6460 (N_6460,N_4129,N_5662);
or U6461 (N_6461,N_5254,N_5161);
nand U6462 (N_6462,N_4703,N_5695);
nand U6463 (N_6463,N_4650,N_5043);
or U6464 (N_6464,N_5534,N_4685);
or U6465 (N_6465,N_5841,N_5370);
or U6466 (N_6466,N_4376,N_5168);
nor U6467 (N_6467,N_5728,N_4419);
and U6468 (N_6468,N_5381,N_5946);
xnor U6469 (N_6469,N_4115,N_5338);
xor U6470 (N_6470,N_5170,N_5129);
nor U6471 (N_6471,N_4108,N_4433);
nor U6472 (N_6472,N_5186,N_4830);
and U6473 (N_6473,N_4130,N_5771);
xnor U6474 (N_6474,N_4402,N_5580);
nand U6475 (N_6475,N_5073,N_5616);
and U6476 (N_6476,N_5264,N_5646);
nand U6477 (N_6477,N_4695,N_4818);
nand U6478 (N_6478,N_5802,N_5781);
and U6479 (N_6479,N_4244,N_4919);
nor U6480 (N_6480,N_4809,N_5223);
nand U6481 (N_6481,N_5282,N_4418);
nand U6482 (N_6482,N_5702,N_4098);
nor U6483 (N_6483,N_5287,N_5650);
nand U6484 (N_6484,N_5063,N_4641);
and U6485 (N_6485,N_4199,N_4107);
nor U6486 (N_6486,N_5638,N_4949);
xnor U6487 (N_6487,N_4837,N_4840);
nand U6488 (N_6488,N_4281,N_4785);
nand U6489 (N_6489,N_5140,N_5513);
nand U6490 (N_6490,N_4385,N_4757);
nand U6491 (N_6491,N_5472,N_5822);
or U6492 (N_6492,N_4687,N_4961);
nor U6493 (N_6493,N_4606,N_5942);
xnor U6494 (N_6494,N_5849,N_5990);
nand U6495 (N_6495,N_4914,N_5630);
nand U6496 (N_6496,N_4019,N_4801);
xnor U6497 (N_6497,N_4335,N_5815);
nor U6498 (N_6498,N_5765,N_4269);
or U6499 (N_6499,N_4790,N_4661);
or U6500 (N_6500,N_5605,N_4346);
nor U6501 (N_6501,N_4453,N_5069);
xnor U6502 (N_6502,N_5133,N_4664);
or U6503 (N_6503,N_5214,N_4988);
xor U6504 (N_6504,N_4881,N_4121);
xnor U6505 (N_6505,N_4097,N_4723);
or U6506 (N_6506,N_4400,N_5196);
nand U6507 (N_6507,N_4906,N_5036);
nand U6508 (N_6508,N_4037,N_4592);
or U6509 (N_6509,N_5367,N_5278);
nand U6510 (N_6510,N_4913,N_4257);
nand U6511 (N_6511,N_4427,N_5025);
and U6512 (N_6512,N_5447,N_5949);
and U6513 (N_6513,N_4172,N_5280);
or U6514 (N_6514,N_5820,N_4636);
and U6515 (N_6515,N_5556,N_4987);
and U6516 (N_6516,N_5248,N_4819);
nand U6517 (N_6517,N_5525,N_5539);
nand U6518 (N_6518,N_5405,N_4459);
or U6519 (N_6519,N_5453,N_4629);
nand U6520 (N_6520,N_4777,N_4674);
or U6521 (N_6521,N_5612,N_5831);
and U6522 (N_6522,N_4144,N_5686);
nor U6523 (N_6523,N_4575,N_4742);
nand U6524 (N_6524,N_5395,N_4911);
nor U6525 (N_6525,N_5038,N_4599);
xnor U6526 (N_6526,N_4032,N_4030);
or U6527 (N_6527,N_4755,N_5544);
or U6528 (N_6528,N_4283,N_4535);
or U6529 (N_6529,N_5953,N_4952);
xor U6530 (N_6530,N_5796,N_4051);
or U6531 (N_6531,N_4752,N_4104);
xor U6532 (N_6532,N_4940,N_5871);
nor U6533 (N_6533,N_5521,N_5980);
nor U6534 (N_6534,N_5421,N_4816);
xor U6535 (N_6535,N_5978,N_4087);
nand U6536 (N_6536,N_4137,N_4898);
nand U6537 (N_6537,N_4132,N_5079);
nor U6538 (N_6538,N_5182,N_4917);
and U6539 (N_6539,N_4783,N_4505);
nor U6540 (N_6540,N_4467,N_5465);
and U6541 (N_6541,N_5426,N_5062);
nor U6542 (N_6542,N_4552,N_5122);
or U6543 (N_6543,N_4466,N_5575);
or U6544 (N_6544,N_4848,N_4113);
nand U6545 (N_6545,N_4979,N_5585);
and U6546 (N_6546,N_5760,N_4173);
xor U6547 (N_6547,N_5058,N_5660);
nand U6548 (N_6548,N_4921,N_4937);
nor U6549 (N_6549,N_4655,N_5944);
nor U6550 (N_6550,N_5267,N_4391);
nor U6551 (N_6551,N_4168,N_4577);
nand U6552 (N_6552,N_5181,N_4806);
xnor U6553 (N_6553,N_4304,N_4282);
nand U6554 (N_6554,N_5825,N_5557);
nand U6555 (N_6555,N_5241,N_5623);
xnor U6556 (N_6556,N_5955,N_5255);
nor U6557 (N_6557,N_4523,N_5952);
and U6558 (N_6558,N_4069,N_4533);
nand U6559 (N_6559,N_5610,N_4520);
nor U6560 (N_6560,N_5601,N_5503);
or U6561 (N_6561,N_5668,N_4618);
nand U6562 (N_6562,N_5836,N_5880);
or U6563 (N_6563,N_4313,N_4197);
nor U6564 (N_6564,N_4566,N_4448);
nand U6565 (N_6565,N_5331,N_5477);
nand U6566 (N_6566,N_5290,N_5005);
xor U6567 (N_6567,N_5061,N_5021);
and U6568 (N_6568,N_4138,N_5691);
nand U6569 (N_6569,N_5963,N_4039);
or U6570 (N_6570,N_4789,N_4665);
nor U6571 (N_6571,N_4718,N_5622);
nand U6572 (N_6572,N_5891,N_4395);
nand U6573 (N_6573,N_4775,N_5726);
nand U6574 (N_6574,N_4406,N_5569);
and U6575 (N_6575,N_5787,N_5219);
or U6576 (N_6576,N_4918,N_4125);
nor U6577 (N_6577,N_4240,N_5615);
or U6578 (N_6578,N_5530,N_4021);
nor U6579 (N_6579,N_5943,N_5132);
and U6580 (N_6580,N_4414,N_4143);
nand U6581 (N_6581,N_5683,N_4546);
nand U6582 (N_6582,N_4077,N_4582);
or U6583 (N_6583,N_4396,N_4596);
xor U6584 (N_6584,N_5680,N_4308);
nor U6585 (N_6585,N_5535,N_4612);
and U6586 (N_6586,N_5127,N_5900);
nand U6587 (N_6587,N_4883,N_5136);
or U6588 (N_6588,N_4061,N_5139);
xnor U6589 (N_6589,N_4471,N_5877);
xnor U6590 (N_6590,N_4835,N_5203);
nor U6591 (N_6591,N_4954,N_4015);
and U6592 (N_6592,N_4870,N_5359);
nand U6593 (N_6593,N_4449,N_4267);
and U6594 (N_6594,N_5892,N_5375);
nand U6595 (N_6595,N_5076,N_5190);
nor U6596 (N_6596,N_4497,N_5883);
nand U6597 (N_6597,N_4521,N_5795);
nand U6598 (N_6598,N_4829,N_5304);
and U6599 (N_6599,N_4513,N_5102);
and U6600 (N_6600,N_4966,N_5917);
nand U6601 (N_6601,N_4734,N_4154);
or U6602 (N_6602,N_5739,N_4748);
nor U6603 (N_6603,N_4896,N_4489);
nand U6604 (N_6604,N_5876,N_4145);
xor U6605 (N_6605,N_5654,N_4554);
or U6606 (N_6606,N_4507,N_5467);
xnor U6607 (N_6607,N_4128,N_4626);
nor U6608 (N_6608,N_5423,N_5775);
nand U6609 (N_6609,N_4822,N_4175);
xor U6610 (N_6610,N_4171,N_5537);
or U6611 (N_6611,N_4460,N_4076);
xor U6612 (N_6612,N_5162,N_5250);
nor U6613 (N_6613,N_5587,N_5527);
and U6614 (N_6614,N_5160,N_4788);
nor U6615 (N_6615,N_5794,N_5724);
nor U6616 (N_6616,N_5452,N_5017);
xor U6617 (N_6617,N_4345,N_5872);
and U6618 (N_6618,N_4756,N_4998);
or U6619 (N_6619,N_5491,N_4880);
and U6620 (N_6620,N_5692,N_5887);
nor U6621 (N_6621,N_5130,N_4249);
or U6622 (N_6622,N_5064,N_5402);
and U6623 (N_6623,N_4476,N_4187);
nor U6624 (N_6624,N_4285,N_4227);
nand U6625 (N_6625,N_4894,N_4003);
xnor U6626 (N_6626,N_5086,N_5598);
nand U6627 (N_6627,N_4892,N_5101);
nand U6628 (N_6628,N_4948,N_5314);
and U6629 (N_6629,N_5149,N_4736);
or U6630 (N_6630,N_5292,N_5811);
nor U6631 (N_6631,N_4000,N_5649);
xor U6632 (N_6632,N_4321,N_5938);
nor U6633 (N_6633,N_5632,N_4158);
nand U6634 (N_6634,N_5707,N_5415);
nor U6635 (N_6635,N_4908,N_5350);
nor U6636 (N_6636,N_5552,N_5933);
nand U6637 (N_6637,N_5783,N_4767);
nand U6638 (N_6638,N_4455,N_4347);
or U6639 (N_6639,N_4374,N_5532);
nand U6640 (N_6640,N_4891,N_4658);
or U6641 (N_6641,N_4155,N_5456);
and U6642 (N_6642,N_4751,N_5365);
and U6643 (N_6643,N_5345,N_4943);
nor U6644 (N_6644,N_4854,N_4693);
and U6645 (N_6645,N_4484,N_4064);
nor U6646 (N_6646,N_4699,N_5334);
and U6647 (N_6647,N_4564,N_5225);
xor U6648 (N_6648,N_4993,N_5387);
nand U6649 (N_6649,N_5907,N_4558);
and U6650 (N_6650,N_4298,N_5156);
or U6651 (N_6651,N_4928,N_5969);
nor U6652 (N_6652,N_5124,N_4709);
xnor U6653 (N_6653,N_4958,N_4857);
nor U6654 (N_6654,N_5966,N_4163);
nand U6655 (N_6655,N_5117,N_4858);
and U6656 (N_6656,N_5797,N_4944);
and U6657 (N_6657,N_4605,N_4036);
or U6658 (N_6658,N_4551,N_4971);
nor U6659 (N_6659,N_4530,N_5643);
xor U6660 (N_6660,N_4498,N_4691);
and U6661 (N_6661,N_5377,N_4716);
or U6662 (N_6662,N_5260,N_4264);
nand U6663 (N_6663,N_4022,N_5976);
nor U6664 (N_6664,N_4358,N_4793);
nor U6665 (N_6665,N_5614,N_4985);
or U6666 (N_6666,N_4007,N_5481);
and U6667 (N_6667,N_4404,N_5804);
or U6668 (N_6668,N_4081,N_5294);
nand U6669 (N_6669,N_5936,N_5009);
xnor U6670 (N_6670,N_4110,N_4494);
or U6671 (N_6671,N_5354,N_4706);
nand U6672 (N_6672,N_4242,N_5634);
nor U6673 (N_6673,N_4133,N_4286);
xor U6674 (N_6674,N_5895,N_5590);
nand U6675 (N_6675,N_5374,N_4978);
and U6676 (N_6676,N_5384,N_5908);
and U6677 (N_6677,N_5454,N_4963);
and U6678 (N_6678,N_4585,N_5777);
nor U6679 (N_6679,N_5772,N_4717);
xor U6680 (N_6680,N_5376,N_4105);
nor U6681 (N_6681,N_5636,N_4464);
nor U6682 (N_6682,N_4457,N_5925);
or U6683 (N_6683,N_5390,N_4930);
and U6684 (N_6684,N_4689,N_5229);
or U6685 (N_6685,N_5245,N_5150);
nand U6686 (N_6686,N_4196,N_4721);
or U6687 (N_6687,N_5311,N_4621);
nor U6688 (N_6688,N_4152,N_5745);
or U6689 (N_6689,N_5090,N_5224);
nand U6690 (N_6690,N_5881,N_4518);
or U6691 (N_6691,N_4821,N_5118);
nand U6692 (N_6692,N_5071,N_5937);
and U6693 (N_6693,N_4933,N_4111);
xnor U6694 (N_6694,N_5325,N_5923);
and U6695 (N_6695,N_5926,N_5302);
or U6696 (N_6696,N_4246,N_5717);
and U6697 (N_6697,N_5830,N_5809);
or U6698 (N_6698,N_5027,N_5870);
and U6699 (N_6699,N_5012,N_5987);
xor U6700 (N_6700,N_4236,N_4713);
xnor U6701 (N_6701,N_5145,N_4730);
nor U6702 (N_6702,N_4425,N_5597);
nand U6703 (N_6703,N_5559,N_4700);
nand U6704 (N_6704,N_5271,N_5790);
xor U6705 (N_6705,N_4190,N_4185);
nand U6706 (N_6706,N_4430,N_4480);
nand U6707 (N_6707,N_4068,N_4357);
nand U6708 (N_6708,N_4432,N_4849);
nand U6709 (N_6709,N_5346,N_4860);
nor U6710 (N_6710,N_4737,N_5482);
or U6711 (N_6711,N_4209,N_4237);
nor U6712 (N_6712,N_4651,N_5242);
nor U6713 (N_6713,N_4868,N_4002);
nor U6714 (N_6714,N_5536,N_4181);
nand U6715 (N_6715,N_4273,N_4864);
or U6716 (N_6716,N_4470,N_5905);
nor U6717 (N_6717,N_5403,N_5824);
and U6718 (N_6718,N_5663,N_4112);
nand U6719 (N_6719,N_5835,N_5317);
or U6720 (N_6720,N_5198,N_4903);
or U6721 (N_6721,N_4040,N_5854);
and U6722 (N_6722,N_5364,N_5455);
or U6723 (N_6723,N_4642,N_4245);
nand U6724 (N_6724,N_4701,N_5866);
or U6725 (N_6725,N_5672,N_5655);
nor U6726 (N_6726,N_5032,N_5348);
nand U6727 (N_6727,N_4394,N_5964);
xnor U6728 (N_6728,N_5948,N_5910);
or U6729 (N_6729,N_5848,N_4614);
nor U6730 (N_6730,N_5369,N_5747);
xnor U6731 (N_6731,N_4725,N_5355);
xor U6732 (N_6732,N_5409,N_5289);
and U6733 (N_6733,N_4556,N_5994);
xnor U6734 (N_6734,N_4429,N_5388);
nand U6735 (N_6735,N_4299,N_5411);
or U6736 (N_6736,N_5706,N_5085);
nor U6737 (N_6737,N_5463,N_5430);
or U6738 (N_6738,N_5098,N_5084);
or U6739 (N_6739,N_5712,N_5688);
or U6740 (N_6740,N_5553,N_5401);
nor U6741 (N_6741,N_4028,N_4544);
and U6742 (N_6742,N_5600,N_4165);
or U6743 (N_6743,N_4083,N_5135);
and U6744 (N_6744,N_4578,N_5261);
nand U6745 (N_6745,N_5163,N_4771);
or U6746 (N_6746,N_5914,N_4410);
nand U6747 (N_6747,N_5347,N_4683);
and U6748 (N_6748,N_4141,N_4238);
and U6749 (N_6749,N_4503,N_4373);
and U6750 (N_6750,N_4272,N_5103);
and U6751 (N_6751,N_5400,N_4637);
xnor U6752 (N_6752,N_5586,N_5996);
nand U6753 (N_6753,N_4393,N_5762);
nor U6754 (N_6754,N_4747,N_5734);
and U6755 (N_6755,N_5428,N_5671);
nand U6756 (N_6756,N_5042,N_5897);
nor U6757 (N_6757,N_5154,N_5551);
or U6758 (N_6758,N_4602,N_4140);
and U6759 (N_6759,N_5231,N_5768);
nor U6760 (N_6760,N_5653,N_4992);
or U6761 (N_6761,N_5682,N_5495);
nand U6762 (N_6762,N_4542,N_5357);
xnor U6763 (N_6763,N_4782,N_4146);
xor U6764 (N_6764,N_4697,N_5431);
or U6765 (N_6765,N_4763,N_4539);
and U6766 (N_6766,N_5751,N_5474);
and U6767 (N_6767,N_4660,N_4045);
xnor U6768 (N_6768,N_5710,N_5252);
or U6769 (N_6769,N_4215,N_5087);
xor U6770 (N_6770,N_4020,N_4205);
and U6771 (N_6771,N_5138,N_4982);
nand U6772 (N_6772,N_4770,N_4712);
or U6773 (N_6773,N_5088,N_5989);
or U6774 (N_6774,N_5111,N_5107);
nor U6775 (N_6775,N_4049,N_4250);
nand U6776 (N_6776,N_5862,N_4436);
or U6777 (N_6777,N_4561,N_4462);
nor U6778 (N_6778,N_4920,N_4363);
nor U6779 (N_6779,N_5954,N_4136);
nand U6780 (N_6780,N_5262,N_5046);
nand U6781 (N_6781,N_5212,N_5689);
or U6782 (N_6782,N_4681,N_4254);
nor U6783 (N_6783,N_4216,N_4176);
nand U6784 (N_6784,N_4096,N_4131);
xnor U6785 (N_6785,N_4648,N_4318);
and U6786 (N_6786,N_5324,N_4804);
nor U6787 (N_6787,N_4265,N_5441);
xor U6788 (N_6788,N_5657,N_5915);
nand U6789 (N_6789,N_4328,N_5779);
or U6790 (N_6790,N_4182,N_5030);
nor U6791 (N_6791,N_5488,N_5420);
nor U6792 (N_6792,N_5602,N_5448);
nor U6793 (N_6793,N_4356,N_5100);
and U6794 (N_6794,N_5037,N_4092);
nand U6795 (N_6795,N_5299,N_5059);
and U6796 (N_6796,N_4386,N_4231);
or U6797 (N_6797,N_4502,N_4038);
xnor U6798 (N_6798,N_5847,N_5774);
or U6799 (N_6799,N_4071,N_5358);
and U6800 (N_6800,N_4915,N_4500);
nor U6801 (N_6801,N_4766,N_4814);
and U6802 (N_6802,N_4160,N_4504);
nor U6803 (N_6803,N_5538,N_5647);
nor U6804 (N_6804,N_5380,N_4088);
nor U6805 (N_6805,N_5310,N_5694);
and U6806 (N_6806,N_4838,N_4916);
nor U6807 (N_6807,N_5611,N_5755);
nand U6808 (N_6808,N_4680,N_5868);
and U6809 (N_6809,N_5246,N_4120);
and U6810 (N_6810,N_4490,N_4827);
nor U6811 (N_6811,N_4844,N_4188);
nand U6812 (N_6812,N_5593,N_5211);
nor U6813 (N_6813,N_5178,N_5681);
xnor U6814 (N_6814,N_5445,N_5049);
nand U6815 (N_6815,N_4762,N_4109);
nor U6816 (N_6816,N_5704,N_5604);
or U6817 (N_6817,N_4080,N_4733);
nor U6818 (N_6818,N_5801,N_4355);
nand U6819 (N_6819,N_4669,N_4053);
nor U6820 (N_6820,N_4475,N_4370);
or U6821 (N_6821,N_4122,N_4306);
or U6822 (N_6822,N_5793,N_5449);
and U6823 (N_6823,N_4322,N_4364);
and U6824 (N_6824,N_5970,N_5379);
nand U6825 (N_6825,N_5115,N_5230);
nand U6826 (N_6826,N_4834,N_4048);
or U6827 (N_6827,N_4458,N_4842);
or U6828 (N_6828,N_5763,N_4812);
nand U6829 (N_6829,N_4679,N_4228);
nor U6830 (N_6830,N_5808,N_5817);
nand U6831 (N_6831,N_5806,N_4845);
and U6832 (N_6832,N_4093,N_5109);
or U6833 (N_6833,N_4349,N_4219);
and U6834 (N_6834,N_4797,N_5273);
xor U6835 (N_6835,N_5006,N_5546);
nand U6836 (N_6836,N_5082,N_4277);
or U6837 (N_6837,N_5297,N_5922);
or U6838 (N_6838,N_4017,N_5362);
and U6839 (N_6839,N_5939,N_4366);
nor U6840 (N_6840,N_4776,N_5945);
nor U6841 (N_6841,N_4426,N_4901);
nand U6842 (N_6842,N_4741,N_4297);
nand U6843 (N_6843,N_5183,N_4560);
xnor U6844 (N_6844,N_5716,N_5476);
and U6845 (N_6845,N_5392,N_4420);
nand U6846 (N_6846,N_4085,N_5330);
or U6847 (N_6847,N_4798,N_5328);
nor U6848 (N_6848,N_5873,N_4221);
or U6849 (N_6849,N_4421,N_4823);
nand U6850 (N_6850,N_4326,N_4871);
nor U6851 (N_6851,N_5258,N_4615);
or U6852 (N_6852,N_4491,N_5494);
and U6853 (N_6853,N_4684,N_5301);
nor U6854 (N_6854,N_5608,N_5295);
and U6855 (N_6855,N_5429,N_5651);
nor U6856 (N_6856,N_5679,N_5498);
or U6857 (N_6857,N_4796,N_5582);
or U6858 (N_6858,N_4799,N_5288);
or U6859 (N_6859,N_5993,N_5189);
xor U6860 (N_6860,N_4588,N_4259);
nand U6861 (N_6861,N_4256,N_5307);
or U6862 (N_6862,N_4413,N_5444);
nand U6863 (N_6863,N_5188,N_5470);
or U6864 (N_6864,N_4169,N_4589);
xnor U6865 (N_6865,N_5766,N_5191);
or U6866 (N_6866,N_4212,N_4884);
or U6867 (N_6867,N_5673,N_4670);
nand U6868 (N_6868,N_5810,N_4207);
and U6869 (N_6869,N_4607,N_4774);
and U6870 (N_6870,N_4516,N_5339);
and U6871 (N_6871,N_4794,N_4034);
nand U6872 (N_6872,N_5440,N_4235);
and U6873 (N_6873,N_4336,N_5406);
nor U6874 (N_6874,N_4091,N_5558);
nand U6875 (N_6875,N_5014,N_5878);
and U6876 (N_6876,N_4635,N_4439);
nor U6877 (N_6877,N_4463,N_5319);
nor U6878 (N_6878,N_4803,N_4587);
nor U6879 (N_6879,N_5092,N_4540);
nand U6880 (N_6880,N_4371,N_5265);
and U6881 (N_6881,N_5924,N_5425);
nor U6882 (N_6882,N_4288,N_4047);
nor U6883 (N_6883,N_4900,N_5567);
nand U6884 (N_6884,N_5541,N_5232);
and U6885 (N_6885,N_4584,N_4946);
or U6886 (N_6886,N_4361,N_5322);
nor U6887 (N_6887,N_4633,N_5234);
nor U6888 (N_6888,N_5756,N_5055);
nand U6889 (N_6889,N_4095,N_4698);
and U6890 (N_6890,N_5767,N_5983);
nor U6891 (N_6891,N_5742,N_5257);
nand U6892 (N_6892,N_4379,N_5080);
xnor U6893 (N_6893,N_5464,N_4443);
nor U6894 (N_6894,N_4033,N_4161);
nand U6895 (N_6895,N_5205,N_5542);
nor U6896 (N_6896,N_4333,N_5791);
or U6897 (N_6897,N_5057,N_4923);
nor U6898 (N_6898,N_4983,N_5874);
nor U6899 (N_6899,N_5719,N_5884);
or U6900 (N_6900,N_5735,N_4974);
nand U6901 (N_6901,N_4067,N_5137);
nor U6902 (N_6902,N_5309,N_4223);
or U6903 (N_6903,N_5813,N_5054);
nand U6904 (N_6904,N_5613,N_4586);
nand U6905 (N_6905,N_5700,N_5493);
or U6906 (N_6906,N_5028,N_4261);
or U6907 (N_6907,N_5142,N_5164);
nand U6908 (N_6908,N_4792,N_5228);
nand U6909 (N_6909,N_5065,N_5083);
or U6910 (N_6910,N_4640,N_4090);
and U6911 (N_6911,N_5697,N_4936);
and U6912 (N_6912,N_5095,N_5676);
and U6913 (N_6913,N_4800,N_5524);
and U6914 (N_6914,N_5661,N_4408);
nor U6915 (N_6915,N_4732,N_4926);
or U6916 (N_6916,N_5412,N_5579);
nor U6917 (N_6917,N_4638,N_4553);
and U6918 (N_6918,N_4825,N_4541);
and U6919 (N_6919,N_5176,N_4334);
nand U6920 (N_6920,N_4417,N_5642);
or U6921 (N_6921,N_5443,N_4360);
or U6922 (N_6922,N_5342,N_4675);
nand U6923 (N_6923,N_4390,N_5885);
or U6924 (N_6924,N_4984,N_5522);
and U6925 (N_6925,N_5998,N_4213);
or U6926 (N_6926,N_5201,N_4764);
nand U6927 (N_6927,N_4772,N_5548);
or U6928 (N_6928,N_4041,N_4375);
or U6929 (N_6929,N_5233,N_5863);
nand U6930 (N_6930,N_5882,N_5047);
nand U6931 (N_6931,N_4367,N_5906);
nand U6932 (N_6932,N_5621,N_5333);
and U6933 (N_6933,N_4676,N_4167);
xor U6934 (N_6934,N_5126,N_5749);
nand U6935 (N_6935,N_5207,N_4487);
and U6936 (N_6936,N_5078,N_5856);
or U6937 (N_6937,N_5151,N_5929);
nor U6938 (N_6938,N_5341,N_5008);
and U6939 (N_6939,N_4253,N_5332);
or U6940 (N_6940,N_5056,N_4955);
or U6941 (N_6941,N_4610,N_5840);
and U6942 (N_6942,N_4519,N_5209);
or U6943 (N_6943,N_5312,N_5523);
and U6944 (N_6944,N_4156,N_5858);
nand U6945 (N_6945,N_5959,N_4474);
or U6946 (N_6946,N_4354,N_5902);
or U6947 (N_6947,N_5237,N_4001);
nor U6948 (N_6948,N_5326,N_5033);
or U6949 (N_6949,N_5977,N_5438);
nor U6950 (N_6950,N_5093,N_4403);
or U6951 (N_6951,N_4628,N_5894);
nand U6952 (N_6952,N_5187,N_5518);
or U6953 (N_6953,N_5119,N_4565);
xor U6954 (N_6954,N_4537,N_5827);
nor U6955 (N_6955,N_5547,N_5020);
or U6956 (N_6956,N_5372,N_5123);
nand U6957 (N_6957,N_5596,N_4964);
or U6958 (N_6958,N_4934,N_5573);
nor U6959 (N_6959,N_4866,N_5039);
nor U6960 (N_6960,N_4251,N_5971);
nand U6961 (N_6961,N_4218,N_5487);
and U6962 (N_6962,N_4052,N_5667);
or U6963 (N_6963,N_4325,N_5031);
or U6964 (N_6964,N_5853,N_4289);
nor U6965 (N_6965,N_5368,N_4331);
nor U6966 (N_6966,N_5967,N_4392);
nand U6967 (N_6967,N_5782,N_4203);
and U6968 (N_6968,N_5533,N_5962);
nand U6969 (N_6969,N_5272,N_5291);
nor U6970 (N_6970,N_4951,N_4807);
nand U6971 (N_6971,N_5934,N_4384);
and U6972 (N_6972,N_4853,N_5864);
or U6973 (N_6973,N_5239,N_4351);
and U6974 (N_6974,N_4343,N_5979);
nand U6975 (N_6975,N_5277,N_5626);
and U6976 (N_6976,N_5458,N_4278);
nor U6977 (N_6977,N_4613,N_4495);
xor U6978 (N_6978,N_5382,N_4547);
or U6979 (N_6979,N_4324,N_4620);
and U6980 (N_6980,N_4075,N_5713);
nand U6981 (N_6981,N_4255,N_4332);
or U6982 (N_6982,N_5637,N_4359);
and U6983 (N_6983,N_5471,N_5844);
and U6984 (N_6984,N_5340,N_5974);
or U6985 (N_6985,N_4888,N_5480);
or U6986 (N_6986,N_5361,N_5770);
nand U6987 (N_6987,N_4802,N_5991);
nand U6988 (N_6988,N_4759,N_5141);
nand U6989 (N_6989,N_4632,N_4042);
and U6990 (N_6990,N_5752,N_5349);
or U6991 (N_6991,N_5708,N_5344);
nor U6992 (N_6992,N_5050,N_5352);
nand U6993 (N_6993,N_5089,N_5068);
and U6994 (N_6994,N_5652,N_4452);
xor U6995 (N_6995,N_5215,N_4016);
or U6996 (N_6996,N_4805,N_4478);
nand U6997 (N_6997,N_4224,N_5249);
nand U6998 (N_6998,N_4778,N_4340);
and U6999 (N_6999,N_4352,N_5619);
or U7000 (N_7000,N_4899,N_5586);
nor U7001 (N_7001,N_4451,N_4396);
nor U7002 (N_7002,N_5576,N_4116);
nand U7003 (N_7003,N_5542,N_5097);
and U7004 (N_7004,N_4855,N_5983);
xor U7005 (N_7005,N_5714,N_5029);
or U7006 (N_7006,N_5933,N_5155);
and U7007 (N_7007,N_4675,N_4526);
and U7008 (N_7008,N_5825,N_5149);
nand U7009 (N_7009,N_4539,N_4964);
and U7010 (N_7010,N_4772,N_4915);
nor U7011 (N_7011,N_4960,N_4188);
nand U7012 (N_7012,N_5479,N_4500);
nor U7013 (N_7013,N_4848,N_5327);
and U7014 (N_7014,N_5438,N_4204);
nand U7015 (N_7015,N_4581,N_4456);
nor U7016 (N_7016,N_4921,N_4164);
and U7017 (N_7017,N_5884,N_4886);
and U7018 (N_7018,N_4560,N_4801);
and U7019 (N_7019,N_4857,N_5759);
xor U7020 (N_7020,N_5649,N_5767);
and U7021 (N_7021,N_4266,N_5708);
nor U7022 (N_7022,N_5754,N_4204);
xnor U7023 (N_7023,N_4825,N_5823);
xor U7024 (N_7024,N_5278,N_4478);
nand U7025 (N_7025,N_4725,N_4160);
nor U7026 (N_7026,N_4143,N_4233);
and U7027 (N_7027,N_4647,N_5388);
nor U7028 (N_7028,N_5147,N_5113);
nor U7029 (N_7029,N_5639,N_5910);
xor U7030 (N_7030,N_5480,N_4924);
and U7031 (N_7031,N_5366,N_4916);
nand U7032 (N_7032,N_4547,N_4847);
nand U7033 (N_7033,N_5840,N_5238);
xnor U7034 (N_7034,N_5315,N_5226);
or U7035 (N_7035,N_4419,N_4066);
nand U7036 (N_7036,N_4447,N_4716);
or U7037 (N_7037,N_4835,N_4291);
or U7038 (N_7038,N_4328,N_5814);
or U7039 (N_7039,N_5655,N_5813);
nand U7040 (N_7040,N_4508,N_4636);
or U7041 (N_7041,N_4536,N_4575);
or U7042 (N_7042,N_5754,N_5311);
nor U7043 (N_7043,N_5386,N_5858);
nor U7044 (N_7044,N_5924,N_5205);
or U7045 (N_7045,N_4833,N_5676);
and U7046 (N_7046,N_5507,N_5906);
and U7047 (N_7047,N_4067,N_5615);
nor U7048 (N_7048,N_4046,N_5874);
xnor U7049 (N_7049,N_5009,N_5350);
and U7050 (N_7050,N_5400,N_4066);
or U7051 (N_7051,N_5980,N_5772);
or U7052 (N_7052,N_5937,N_5000);
or U7053 (N_7053,N_4480,N_4649);
xor U7054 (N_7054,N_5410,N_5533);
nand U7055 (N_7055,N_4402,N_5388);
nand U7056 (N_7056,N_4883,N_4038);
nor U7057 (N_7057,N_5600,N_4867);
and U7058 (N_7058,N_4027,N_5805);
or U7059 (N_7059,N_5776,N_4819);
nor U7060 (N_7060,N_5522,N_4595);
xor U7061 (N_7061,N_4442,N_5693);
and U7062 (N_7062,N_4631,N_4626);
or U7063 (N_7063,N_4110,N_5628);
nor U7064 (N_7064,N_5103,N_4198);
nor U7065 (N_7065,N_4396,N_4541);
or U7066 (N_7066,N_4464,N_5955);
nor U7067 (N_7067,N_4921,N_4719);
nor U7068 (N_7068,N_4143,N_5786);
nand U7069 (N_7069,N_4856,N_5450);
nor U7070 (N_7070,N_5636,N_5904);
or U7071 (N_7071,N_5875,N_4473);
or U7072 (N_7072,N_5130,N_5511);
xor U7073 (N_7073,N_5372,N_4228);
or U7074 (N_7074,N_4113,N_4670);
or U7075 (N_7075,N_5391,N_5829);
or U7076 (N_7076,N_5820,N_4383);
or U7077 (N_7077,N_5308,N_5006);
xnor U7078 (N_7078,N_5153,N_4983);
nand U7079 (N_7079,N_4898,N_5478);
nor U7080 (N_7080,N_4595,N_5176);
and U7081 (N_7081,N_4761,N_4484);
and U7082 (N_7082,N_5057,N_5055);
nor U7083 (N_7083,N_5686,N_5459);
and U7084 (N_7084,N_5073,N_5165);
or U7085 (N_7085,N_4129,N_4466);
nor U7086 (N_7086,N_5561,N_4759);
or U7087 (N_7087,N_5775,N_5469);
or U7088 (N_7088,N_4714,N_4917);
nand U7089 (N_7089,N_5679,N_5714);
nand U7090 (N_7090,N_4637,N_5760);
nor U7091 (N_7091,N_5300,N_4135);
nand U7092 (N_7092,N_4207,N_4107);
nand U7093 (N_7093,N_4912,N_5684);
nor U7094 (N_7094,N_5233,N_5969);
nand U7095 (N_7095,N_4950,N_4193);
and U7096 (N_7096,N_4188,N_5212);
and U7097 (N_7097,N_5971,N_4169);
nand U7098 (N_7098,N_5977,N_4244);
nand U7099 (N_7099,N_4879,N_5798);
and U7100 (N_7100,N_5445,N_5991);
nor U7101 (N_7101,N_4893,N_5106);
nor U7102 (N_7102,N_4682,N_4801);
nor U7103 (N_7103,N_5278,N_4322);
and U7104 (N_7104,N_4697,N_4825);
nand U7105 (N_7105,N_4785,N_5903);
nand U7106 (N_7106,N_4074,N_4068);
or U7107 (N_7107,N_4499,N_5677);
or U7108 (N_7108,N_4273,N_5346);
nor U7109 (N_7109,N_5949,N_5636);
xnor U7110 (N_7110,N_5260,N_4807);
xor U7111 (N_7111,N_5434,N_4194);
or U7112 (N_7112,N_4810,N_4409);
and U7113 (N_7113,N_4702,N_4385);
or U7114 (N_7114,N_5404,N_5397);
or U7115 (N_7115,N_4602,N_5391);
xnor U7116 (N_7116,N_5826,N_4503);
nand U7117 (N_7117,N_5281,N_5946);
or U7118 (N_7118,N_5859,N_4726);
nor U7119 (N_7119,N_5690,N_4883);
nand U7120 (N_7120,N_4080,N_5432);
nand U7121 (N_7121,N_4304,N_5881);
nor U7122 (N_7122,N_4892,N_5507);
or U7123 (N_7123,N_5514,N_5524);
nor U7124 (N_7124,N_4402,N_5732);
and U7125 (N_7125,N_4582,N_4495);
and U7126 (N_7126,N_4524,N_4186);
nand U7127 (N_7127,N_5296,N_4410);
or U7128 (N_7128,N_5825,N_5946);
nand U7129 (N_7129,N_5009,N_5471);
nand U7130 (N_7130,N_4875,N_4923);
nand U7131 (N_7131,N_5889,N_4519);
nand U7132 (N_7132,N_5683,N_5168);
or U7133 (N_7133,N_4716,N_4407);
or U7134 (N_7134,N_5852,N_4269);
xnor U7135 (N_7135,N_5748,N_4560);
or U7136 (N_7136,N_4210,N_4115);
xnor U7137 (N_7137,N_5635,N_4484);
nor U7138 (N_7138,N_4373,N_5708);
nand U7139 (N_7139,N_4109,N_4071);
and U7140 (N_7140,N_5318,N_5271);
or U7141 (N_7141,N_4074,N_5227);
nand U7142 (N_7142,N_5692,N_4117);
and U7143 (N_7143,N_4737,N_5301);
and U7144 (N_7144,N_4630,N_5013);
nand U7145 (N_7145,N_5834,N_5289);
nor U7146 (N_7146,N_5487,N_4546);
or U7147 (N_7147,N_5348,N_4037);
and U7148 (N_7148,N_4675,N_4966);
nor U7149 (N_7149,N_4480,N_5390);
nand U7150 (N_7150,N_5551,N_5238);
nor U7151 (N_7151,N_4223,N_5283);
nand U7152 (N_7152,N_4080,N_4433);
nor U7153 (N_7153,N_4608,N_4809);
or U7154 (N_7154,N_4733,N_5627);
or U7155 (N_7155,N_5364,N_5516);
nand U7156 (N_7156,N_5775,N_4949);
or U7157 (N_7157,N_4411,N_5185);
and U7158 (N_7158,N_5464,N_5754);
or U7159 (N_7159,N_5823,N_4224);
nand U7160 (N_7160,N_5450,N_4995);
nor U7161 (N_7161,N_4284,N_4729);
and U7162 (N_7162,N_4945,N_4984);
or U7163 (N_7163,N_4590,N_5811);
nand U7164 (N_7164,N_5961,N_4745);
and U7165 (N_7165,N_4534,N_5965);
or U7166 (N_7166,N_5298,N_4193);
nor U7167 (N_7167,N_5497,N_5266);
and U7168 (N_7168,N_5349,N_5050);
and U7169 (N_7169,N_5197,N_5458);
nor U7170 (N_7170,N_4014,N_5377);
and U7171 (N_7171,N_4932,N_4844);
nor U7172 (N_7172,N_5097,N_4919);
nor U7173 (N_7173,N_4132,N_5167);
nand U7174 (N_7174,N_5226,N_4023);
nand U7175 (N_7175,N_5741,N_5661);
or U7176 (N_7176,N_4810,N_5615);
or U7177 (N_7177,N_5869,N_4393);
or U7178 (N_7178,N_5317,N_4631);
and U7179 (N_7179,N_4334,N_4571);
or U7180 (N_7180,N_5882,N_4894);
or U7181 (N_7181,N_5708,N_5162);
nand U7182 (N_7182,N_5804,N_4323);
nand U7183 (N_7183,N_5408,N_4482);
or U7184 (N_7184,N_5079,N_5609);
and U7185 (N_7185,N_5756,N_4147);
and U7186 (N_7186,N_5267,N_5251);
nand U7187 (N_7187,N_4069,N_4986);
xnor U7188 (N_7188,N_4697,N_4383);
or U7189 (N_7189,N_5716,N_5891);
nand U7190 (N_7190,N_5336,N_5545);
nor U7191 (N_7191,N_4743,N_5480);
nor U7192 (N_7192,N_5059,N_5892);
or U7193 (N_7193,N_4850,N_5409);
xor U7194 (N_7194,N_4718,N_4978);
or U7195 (N_7195,N_4411,N_4736);
nor U7196 (N_7196,N_5807,N_5155);
or U7197 (N_7197,N_5141,N_5677);
and U7198 (N_7198,N_4123,N_4621);
nand U7199 (N_7199,N_5322,N_5985);
nand U7200 (N_7200,N_5997,N_5526);
nor U7201 (N_7201,N_4211,N_4743);
nor U7202 (N_7202,N_4958,N_5417);
xor U7203 (N_7203,N_5646,N_5582);
or U7204 (N_7204,N_4366,N_5286);
or U7205 (N_7205,N_4538,N_4724);
xor U7206 (N_7206,N_5265,N_5990);
nor U7207 (N_7207,N_4790,N_4944);
nor U7208 (N_7208,N_5697,N_5594);
nand U7209 (N_7209,N_5416,N_5864);
and U7210 (N_7210,N_4922,N_5026);
nand U7211 (N_7211,N_4360,N_5642);
and U7212 (N_7212,N_4021,N_4146);
nand U7213 (N_7213,N_5268,N_4411);
nand U7214 (N_7214,N_4145,N_4733);
and U7215 (N_7215,N_5680,N_5057);
or U7216 (N_7216,N_4425,N_4139);
and U7217 (N_7217,N_4995,N_4698);
nor U7218 (N_7218,N_4223,N_4881);
nor U7219 (N_7219,N_5878,N_4162);
nand U7220 (N_7220,N_5770,N_4663);
nand U7221 (N_7221,N_5948,N_4855);
nor U7222 (N_7222,N_5309,N_5842);
nand U7223 (N_7223,N_4662,N_5810);
nor U7224 (N_7224,N_4438,N_5223);
or U7225 (N_7225,N_4660,N_4033);
nand U7226 (N_7226,N_5526,N_4539);
nand U7227 (N_7227,N_5519,N_5807);
nor U7228 (N_7228,N_5666,N_5150);
and U7229 (N_7229,N_5078,N_5764);
and U7230 (N_7230,N_4084,N_4904);
nand U7231 (N_7231,N_4443,N_4766);
nor U7232 (N_7232,N_5073,N_5898);
and U7233 (N_7233,N_5080,N_5684);
or U7234 (N_7234,N_5640,N_4591);
and U7235 (N_7235,N_4680,N_5857);
nor U7236 (N_7236,N_4807,N_5593);
nand U7237 (N_7237,N_4606,N_4125);
and U7238 (N_7238,N_5682,N_4941);
and U7239 (N_7239,N_4595,N_4759);
or U7240 (N_7240,N_5486,N_5302);
nand U7241 (N_7241,N_5551,N_5760);
nor U7242 (N_7242,N_4463,N_4267);
and U7243 (N_7243,N_5179,N_4848);
nor U7244 (N_7244,N_5688,N_5996);
or U7245 (N_7245,N_5979,N_5969);
xnor U7246 (N_7246,N_4755,N_5737);
nand U7247 (N_7247,N_4497,N_4000);
nand U7248 (N_7248,N_5698,N_4493);
xnor U7249 (N_7249,N_5705,N_4073);
nor U7250 (N_7250,N_4051,N_5851);
nand U7251 (N_7251,N_4600,N_4282);
xnor U7252 (N_7252,N_5047,N_4630);
and U7253 (N_7253,N_5205,N_5647);
and U7254 (N_7254,N_4431,N_4686);
nand U7255 (N_7255,N_5317,N_5706);
xnor U7256 (N_7256,N_5044,N_5482);
nor U7257 (N_7257,N_4801,N_5395);
nand U7258 (N_7258,N_5234,N_5840);
nor U7259 (N_7259,N_5989,N_5565);
nor U7260 (N_7260,N_4921,N_4923);
and U7261 (N_7261,N_5823,N_5947);
or U7262 (N_7262,N_5751,N_4655);
and U7263 (N_7263,N_4421,N_4731);
nor U7264 (N_7264,N_5545,N_5038);
nand U7265 (N_7265,N_4363,N_5169);
nor U7266 (N_7266,N_4509,N_4988);
and U7267 (N_7267,N_5231,N_4887);
and U7268 (N_7268,N_4013,N_4839);
and U7269 (N_7269,N_4582,N_5910);
xor U7270 (N_7270,N_5245,N_5534);
or U7271 (N_7271,N_4094,N_5913);
and U7272 (N_7272,N_4293,N_5374);
nand U7273 (N_7273,N_5177,N_5402);
and U7274 (N_7274,N_4448,N_4873);
and U7275 (N_7275,N_5167,N_5657);
or U7276 (N_7276,N_5292,N_4773);
nand U7277 (N_7277,N_5796,N_5559);
nor U7278 (N_7278,N_5366,N_5355);
nor U7279 (N_7279,N_5664,N_4643);
or U7280 (N_7280,N_4106,N_5183);
nor U7281 (N_7281,N_4094,N_4482);
nand U7282 (N_7282,N_4364,N_4615);
and U7283 (N_7283,N_5204,N_4883);
or U7284 (N_7284,N_4182,N_4878);
nor U7285 (N_7285,N_5028,N_5950);
nor U7286 (N_7286,N_5679,N_5586);
and U7287 (N_7287,N_5796,N_4020);
or U7288 (N_7288,N_5188,N_5021);
and U7289 (N_7289,N_4142,N_4208);
or U7290 (N_7290,N_4650,N_5539);
nand U7291 (N_7291,N_4188,N_5014);
nor U7292 (N_7292,N_5412,N_4049);
and U7293 (N_7293,N_5397,N_5473);
nand U7294 (N_7294,N_5075,N_5968);
or U7295 (N_7295,N_4606,N_5296);
or U7296 (N_7296,N_4101,N_4276);
nand U7297 (N_7297,N_5232,N_5244);
xor U7298 (N_7298,N_5754,N_5696);
or U7299 (N_7299,N_5729,N_5966);
nand U7300 (N_7300,N_4785,N_4161);
xor U7301 (N_7301,N_5263,N_4344);
and U7302 (N_7302,N_5441,N_5241);
nor U7303 (N_7303,N_4720,N_4248);
nor U7304 (N_7304,N_5337,N_4918);
or U7305 (N_7305,N_5585,N_4560);
nand U7306 (N_7306,N_4689,N_5269);
nand U7307 (N_7307,N_4602,N_5360);
or U7308 (N_7308,N_5097,N_5499);
nand U7309 (N_7309,N_4898,N_4171);
or U7310 (N_7310,N_5023,N_5442);
nand U7311 (N_7311,N_4730,N_4959);
nor U7312 (N_7312,N_4285,N_4163);
and U7313 (N_7313,N_4811,N_5288);
and U7314 (N_7314,N_5945,N_5006);
nor U7315 (N_7315,N_5837,N_4834);
or U7316 (N_7316,N_5643,N_4378);
nor U7317 (N_7317,N_4311,N_4468);
nand U7318 (N_7318,N_4810,N_5596);
and U7319 (N_7319,N_4034,N_5167);
and U7320 (N_7320,N_4128,N_4288);
nor U7321 (N_7321,N_5776,N_4108);
nand U7322 (N_7322,N_4932,N_5022);
nor U7323 (N_7323,N_4576,N_4146);
or U7324 (N_7324,N_4018,N_4826);
or U7325 (N_7325,N_4311,N_4865);
or U7326 (N_7326,N_4698,N_5045);
nor U7327 (N_7327,N_4071,N_5890);
nand U7328 (N_7328,N_5101,N_4393);
nand U7329 (N_7329,N_5448,N_5796);
nand U7330 (N_7330,N_5914,N_4664);
or U7331 (N_7331,N_4021,N_5404);
or U7332 (N_7332,N_5634,N_4669);
nand U7333 (N_7333,N_4743,N_4444);
xor U7334 (N_7334,N_4134,N_4422);
nand U7335 (N_7335,N_5816,N_4335);
nand U7336 (N_7336,N_4142,N_5098);
nand U7337 (N_7337,N_5890,N_4356);
or U7338 (N_7338,N_4388,N_5241);
nand U7339 (N_7339,N_4977,N_4287);
or U7340 (N_7340,N_5428,N_4739);
nand U7341 (N_7341,N_4225,N_5796);
and U7342 (N_7342,N_4446,N_4226);
and U7343 (N_7343,N_4233,N_4146);
or U7344 (N_7344,N_5826,N_4867);
and U7345 (N_7345,N_5990,N_5128);
and U7346 (N_7346,N_5468,N_4355);
nor U7347 (N_7347,N_4526,N_4073);
xor U7348 (N_7348,N_5033,N_5094);
and U7349 (N_7349,N_5382,N_4958);
nor U7350 (N_7350,N_5369,N_4105);
nor U7351 (N_7351,N_5464,N_4827);
or U7352 (N_7352,N_5412,N_5914);
or U7353 (N_7353,N_5512,N_5642);
nor U7354 (N_7354,N_5573,N_4110);
nor U7355 (N_7355,N_5565,N_4944);
or U7356 (N_7356,N_4828,N_5652);
or U7357 (N_7357,N_4770,N_4123);
xor U7358 (N_7358,N_4276,N_5751);
xnor U7359 (N_7359,N_5571,N_5727);
and U7360 (N_7360,N_5078,N_4305);
nand U7361 (N_7361,N_5574,N_4215);
xor U7362 (N_7362,N_4971,N_4314);
and U7363 (N_7363,N_5688,N_5436);
and U7364 (N_7364,N_5650,N_5994);
or U7365 (N_7365,N_5613,N_4013);
or U7366 (N_7366,N_4783,N_4021);
nand U7367 (N_7367,N_5696,N_5705);
nand U7368 (N_7368,N_5107,N_4485);
nor U7369 (N_7369,N_5818,N_5522);
xor U7370 (N_7370,N_5056,N_5600);
and U7371 (N_7371,N_4907,N_4268);
nand U7372 (N_7372,N_5304,N_5360);
nor U7373 (N_7373,N_5098,N_4196);
nor U7374 (N_7374,N_5553,N_4483);
nand U7375 (N_7375,N_4428,N_5179);
nor U7376 (N_7376,N_5794,N_4839);
or U7377 (N_7377,N_4813,N_4471);
or U7378 (N_7378,N_5643,N_5687);
or U7379 (N_7379,N_4706,N_4408);
nand U7380 (N_7380,N_5240,N_4269);
nor U7381 (N_7381,N_4585,N_5134);
or U7382 (N_7382,N_4812,N_4793);
nor U7383 (N_7383,N_5114,N_5419);
nand U7384 (N_7384,N_4777,N_4806);
nand U7385 (N_7385,N_4028,N_4922);
xor U7386 (N_7386,N_4742,N_4760);
and U7387 (N_7387,N_5779,N_5003);
xnor U7388 (N_7388,N_5586,N_4896);
xnor U7389 (N_7389,N_4778,N_4150);
or U7390 (N_7390,N_5339,N_4725);
nor U7391 (N_7391,N_4974,N_5018);
or U7392 (N_7392,N_4127,N_5820);
or U7393 (N_7393,N_5455,N_5998);
or U7394 (N_7394,N_4235,N_4194);
or U7395 (N_7395,N_5157,N_5297);
or U7396 (N_7396,N_4140,N_5545);
or U7397 (N_7397,N_5390,N_4670);
or U7398 (N_7398,N_4389,N_5967);
nor U7399 (N_7399,N_4311,N_4157);
nand U7400 (N_7400,N_4731,N_4713);
nand U7401 (N_7401,N_4382,N_5076);
or U7402 (N_7402,N_4595,N_4791);
nor U7403 (N_7403,N_5608,N_5402);
or U7404 (N_7404,N_5540,N_5062);
nand U7405 (N_7405,N_4392,N_4595);
xnor U7406 (N_7406,N_5905,N_4033);
and U7407 (N_7407,N_4444,N_5741);
nor U7408 (N_7408,N_5472,N_4475);
nand U7409 (N_7409,N_5900,N_4179);
and U7410 (N_7410,N_5529,N_5791);
nor U7411 (N_7411,N_4527,N_5661);
xor U7412 (N_7412,N_4931,N_5904);
and U7413 (N_7413,N_4171,N_4465);
nand U7414 (N_7414,N_4305,N_4096);
or U7415 (N_7415,N_4724,N_4793);
and U7416 (N_7416,N_5950,N_5250);
nor U7417 (N_7417,N_4554,N_5301);
or U7418 (N_7418,N_5615,N_5919);
nor U7419 (N_7419,N_4186,N_5250);
or U7420 (N_7420,N_5925,N_5605);
or U7421 (N_7421,N_5296,N_4504);
xor U7422 (N_7422,N_4303,N_4164);
nand U7423 (N_7423,N_4503,N_4971);
or U7424 (N_7424,N_5646,N_5428);
or U7425 (N_7425,N_4955,N_4775);
nor U7426 (N_7426,N_4686,N_5382);
nor U7427 (N_7427,N_4939,N_5250);
nand U7428 (N_7428,N_5046,N_5770);
and U7429 (N_7429,N_4414,N_4253);
or U7430 (N_7430,N_5545,N_4877);
nor U7431 (N_7431,N_5349,N_5092);
or U7432 (N_7432,N_4069,N_4177);
xnor U7433 (N_7433,N_5674,N_4501);
nand U7434 (N_7434,N_4282,N_4594);
or U7435 (N_7435,N_4494,N_5288);
and U7436 (N_7436,N_5770,N_5949);
nand U7437 (N_7437,N_5787,N_4256);
or U7438 (N_7438,N_4024,N_4060);
or U7439 (N_7439,N_5887,N_4916);
or U7440 (N_7440,N_4367,N_5058);
nor U7441 (N_7441,N_5392,N_4131);
and U7442 (N_7442,N_5177,N_4940);
or U7443 (N_7443,N_4066,N_4549);
or U7444 (N_7444,N_5498,N_5727);
or U7445 (N_7445,N_4225,N_4243);
or U7446 (N_7446,N_5696,N_4622);
nand U7447 (N_7447,N_4351,N_4071);
nand U7448 (N_7448,N_5333,N_5063);
or U7449 (N_7449,N_5469,N_4147);
xnor U7450 (N_7450,N_5393,N_5926);
nor U7451 (N_7451,N_5846,N_4173);
nand U7452 (N_7452,N_5463,N_5650);
nor U7453 (N_7453,N_4429,N_4611);
nand U7454 (N_7454,N_4515,N_4199);
xnor U7455 (N_7455,N_5830,N_4861);
nand U7456 (N_7456,N_4318,N_4442);
nor U7457 (N_7457,N_5336,N_5428);
nor U7458 (N_7458,N_4595,N_5541);
nand U7459 (N_7459,N_5694,N_5178);
nor U7460 (N_7460,N_4309,N_4393);
nand U7461 (N_7461,N_5294,N_4090);
nand U7462 (N_7462,N_5812,N_4569);
xor U7463 (N_7463,N_4731,N_4612);
and U7464 (N_7464,N_4576,N_5851);
nor U7465 (N_7465,N_4509,N_5408);
and U7466 (N_7466,N_5629,N_4882);
nand U7467 (N_7467,N_4640,N_5582);
or U7468 (N_7468,N_5981,N_5382);
and U7469 (N_7469,N_5966,N_5736);
nand U7470 (N_7470,N_4873,N_4182);
nand U7471 (N_7471,N_4970,N_5893);
and U7472 (N_7472,N_5664,N_4601);
nor U7473 (N_7473,N_4491,N_5872);
or U7474 (N_7474,N_4431,N_4152);
nand U7475 (N_7475,N_4066,N_4465);
nand U7476 (N_7476,N_5505,N_5248);
nor U7477 (N_7477,N_4268,N_5474);
and U7478 (N_7478,N_5604,N_5526);
nand U7479 (N_7479,N_4012,N_4038);
nand U7480 (N_7480,N_5793,N_4016);
nand U7481 (N_7481,N_4327,N_4416);
xor U7482 (N_7482,N_4684,N_5592);
nand U7483 (N_7483,N_5537,N_5011);
or U7484 (N_7484,N_5277,N_4349);
or U7485 (N_7485,N_4297,N_5785);
nor U7486 (N_7486,N_4531,N_5576);
nand U7487 (N_7487,N_5720,N_5553);
nand U7488 (N_7488,N_4122,N_4731);
xor U7489 (N_7489,N_5455,N_5168);
nor U7490 (N_7490,N_5905,N_4441);
nand U7491 (N_7491,N_5081,N_4542);
or U7492 (N_7492,N_5302,N_5330);
and U7493 (N_7493,N_4211,N_5906);
and U7494 (N_7494,N_5792,N_4894);
and U7495 (N_7495,N_4450,N_5478);
nand U7496 (N_7496,N_4626,N_4114);
or U7497 (N_7497,N_5715,N_5071);
nor U7498 (N_7498,N_5214,N_4148);
and U7499 (N_7499,N_4388,N_5299);
and U7500 (N_7500,N_5881,N_4879);
xnor U7501 (N_7501,N_4085,N_5109);
nand U7502 (N_7502,N_5571,N_5158);
nor U7503 (N_7503,N_5175,N_5784);
xor U7504 (N_7504,N_5860,N_4730);
nor U7505 (N_7505,N_5747,N_4856);
nor U7506 (N_7506,N_5907,N_4344);
or U7507 (N_7507,N_4574,N_5483);
and U7508 (N_7508,N_4898,N_5320);
nor U7509 (N_7509,N_5863,N_5483);
or U7510 (N_7510,N_5938,N_4857);
and U7511 (N_7511,N_5480,N_4660);
nor U7512 (N_7512,N_5986,N_5175);
and U7513 (N_7513,N_5182,N_5406);
or U7514 (N_7514,N_5412,N_5066);
or U7515 (N_7515,N_5523,N_5873);
or U7516 (N_7516,N_5531,N_5467);
nor U7517 (N_7517,N_4868,N_4493);
nand U7518 (N_7518,N_5410,N_4299);
or U7519 (N_7519,N_5945,N_4027);
or U7520 (N_7520,N_5626,N_4164);
and U7521 (N_7521,N_4637,N_5117);
nand U7522 (N_7522,N_5356,N_5951);
or U7523 (N_7523,N_4616,N_4235);
or U7524 (N_7524,N_4268,N_5454);
and U7525 (N_7525,N_4431,N_5002);
or U7526 (N_7526,N_4375,N_4213);
nor U7527 (N_7527,N_4825,N_5083);
xnor U7528 (N_7528,N_4846,N_5213);
or U7529 (N_7529,N_4161,N_5909);
and U7530 (N_7530,N_4060,N_4900);
nand U7531 (N_7531,N_5953,N_4863);
and U7532 (N_7532,N_5534,N_4416);
or U7533 (N_7533,N_4251,N_5506);
xnor U7534 (N_7534,N_4163,N_4316);
and U7535 (N_7535,N_4734,N_5674);
nand U7536 (N_7536,N_4653,N_5391);
or U7537 (N_7537,N_4779,N_4918);
nor U7538 (N_7538,N_5637,N_4022);
nor U7539 (N_7539,N_5864,N_5797);
xor U7540 (N_7540,N_4446,N_5704);
or U7541 (N_7541,N_4288,N_5614);
nand U7542 (N_7542,N_5300,N_5882);
or U7543 (N_7543,N_5261,N_4059);
or U7544 (N_7544,N_4694,N_5753);
nor U7545 (N_7545,N_4374,N_4981);
or U7546 (N_7546,N_4793,N_4388);
xor U7547 (N_7547,N_4423,N_4952);
nor U7548 (N_7548,N_5689,N_4647);
or U7549 (N_7549,N_5705,N_5368);
nand U7550 (N_7550,N_5731,N_4778);
and U7551 (N_7551,N_4754,N_5554);
or U7552 (N_7552,N_5449,N_5353);
nor U7553 (N_7553,N_4152,N_5172);
nor U7554 (N_7554,N_4508,N_5523);
nand U7555 (N_7555,N_5825,N_5812);
or U7556 (N_7556,N_5791,N_4088);
or U7557 (N_7557,N_5854,N_5102);
or U7558 (N_7558,N_5070,N_5617);
nand U7559 (N_7559,N_5142,N_5724);
and U7560 (N_7560,N_4461,N_5547);
nand U7561 (N_7561,N_5890,N_5269);
xor U7562 (N_7562,N_4541,N_5639);
nor U7563 (N_7563,N_5852,N_5836);
nand U7564 (N_7564,N_5896,N_4937);
nor U7565 (N_7565,N_5454,N_5130);
xnor U7566 (N_7566,N_5532,N_5912);
or U7567 (N_7567,N_4832,N_4368);
nand U7568 (N_7568,N_4644,N_4546);
or U7569 (N_7569,N_4514,N_4646);
nor U7570 (N_7570,N_5810,N_4263);
or U7571 (N_7571,N_5702,N_5963);
and U7572 (N_7572,N_5609,N_5921);
or U7573 (N_7573,N_4955,N_5563);
and U7574 (N_7574,N_5210,N_5240);
or U7575 (N_7575,N_5791,N_5625);
or U7576 (N_7576,N_4199,N_4814);
nand U7577 (N_7577,N_5216,N_5492);
and U7578 (N_7578,N_4728,N_4047);
nand U7579 (N_7579,N_4005,N_4575);
nand U7580 (N_7580,N_5228,N_5983);
xor U7581 (N_7581,N_4479,N_5942);
or U7582 (N_7582,N_4340,N_5282);
nand U7583 (N_7583,N_5693,N_4333);
xor U7584 (N_7584,N_5923,N_5205);
and U7585 (N_7585,N_5106,N_4511);
and U7586 (N_7586,N_4661,N_4521);
nor U7587 (N_7587,N_4349,N_4238);
nand U7588 (N_7588,N_4929,N_5100);
nor U7589 (N_7589,N_5559,N_5493);
and U7590 (N_7590,N_5315,N_4877);
nand U7591 (N_7591,N_5242,N_4783);
and U7592 (N_7592,N_4123,N_4427);
nor U7593 (N_7593,N_5052,N_4503);
nor U7594 (N_7594,N_4260,N_4446);
or U7595 (N_7595,N_4955,N_4806);
or U7596 (N_7596,N_4508,N_5585);
and U7597 (N_7597,N_4659,N_4058);
nand U7598 (N_7598,N_4713,N_4154);
and U7599 (N_7599,N_5003,N_5162);
nor U7600 (N_7600,N_4464,N_4846);
nor U7601 (N_7601,N_4412,N_5361);
xor U7602 (N_7602,N_4910,N_5459);
nor U7603 (N_7603,N_5865,N_4047);
and U7604 (N_7604,N_4201,N_4694);
nor U7605 (N_7605,N_4112,N_5432);
nor U7606 (N_7606,N_4810,N_4941);
nor U7607 (N_7607,N_5527,N_5591);
xor U7608 (N_7608,N_4314,N_4298);
and U7609 (N_7609,N_5207,N_5369);
or U7610 (N_7610,N_4350,N_5137);
nand U7611 (N_7611,N_5324,N_5275);
and U7612 (N_7612,N_4505,N_4768);
nand U7613 (N_7613,N_5857,N_5667);
and U7614 (N_7614,N_5279,N_5579);
and U7615 (N_7615,N_5433,N_5615);
nand U7616 (N_7616,N_5920,N_4524);
and U7617 (N_7617,N_4547,N_5808);
nor U7618 (N_7618,N_4799,N_4500);
and U7619 (N_7619,N_4430,N_5998);
nor U7620 (N_7620,N_4849,N_5616);
and U7621 (N_7621,N_5646,N_5072);
xor U7622 (N_7622,N_4591,N_5078);
and U7623 (N_7623,N_5564,N_4554);
nor U7624 (N_7624,N_5338,N_5849);
nor U7625 (N_7625,N_4412,N_4640);
nor U7626 (N_7626,N_4794,N_5675);
or U7627 (N_7627,N_5796,N_4421);
nor U7628 (N_7628,N_5055,N_5922);
nand U7629 (N_7629,N_4917,N_5955);
nor U7630 (N_7630,N_4647,N_4213);
nor U7631 (N_7631,N_4137,N_4971);
nand U7632 (N_7632,N_4996,N_5120);
and U7633 (N_7633,N_5497,N_5911);
nand U7634 (N_7634,N_4095,N_4220);
nand U7635 (N_7635,N_4825,N_5163);
nand U7636 (N_7636,N_4288,N_4322);
and U7637 (N_7637,N_4173,N_5504);
nand U7638 (N_7638,N_5804,N_5173);
xnor U7639 (N_7639,N_4564,N_4478);
nand U7640 (N_7640,N_5732,N_5125);
nand U7641 (N_7641,N_4004,N_5217);
xor U7642 (N_7642,N_5587,N_4239);
or U7643 (N_7643,N_4685,N_5604);
or U7644 (N_7644,N_4215,N_5891);
nand U7645 (N_7645,N_5441,N_4527);
or U7646 (N_7646,N_4211,N_4397);
or U7647 (N_7647,N_5266,N_5369);
nor U7648 (N_7648,N_5393,N_4792);
nor U7649 (N_7649,N_5537,N_5164);
nor U7650 (N_7650,N_5671,N_4800);
xnor U7651 (N_7651,N_4510,N_4702);
xor U7652 (N_7652,N_4953,N_4677);
and U7653 (N_7653,N_5465,N_5567);
nor U7654 (N_7654,N_5719,N_4907);
nor U7655 (N_7655,N_5713,N_4548);
nand U7656 (N_7656,N_5617,N_5217);
and U7657 (N_7657,N_5899,N_4067);
nor U7658 (N_7658,N_5166,N_4265);
nand U7659 (N_7659,N_5823,N_4565);
or U7660 (N_7660,N_4885,N_5255);
or U7661 (N_7661,N_5386,N_5237);
nor U7662 (N_7662,N_4873,N_5033);
and U7663 (N_7663,N_4741,N_5090);
or U7664 (N_7664,N_5406,N_5894);
or U7665 (N_7665,N_5451,N_4548);
and U7666 (N_7666,N_4103,N_4560);
xnor U7667 (N_7667,N_5805,N_5781);
and U7668 (N_7668,N_5592,N_5285);
and U7669 (N_7669,N_5338,N_4142);
nand U7670 (N_7670,N_4848,N_5756);
nand U7671 (N_7671,N_4214,N_5767);
xor U7672 (N_7672,N_4798,N_4162);
or U7673 (N_7673,N_4162,N_4680);
and U7674 (N_7674,N_4392,N_4236);
or U7675 (N_7675,N_4602,N_4295);
nand U7676 (N_7676,N_4210,N_4740);
nand U7677 (N_7677,N_5371,N_4075);
nor U7678 (N_7678,N_4739,N_5355);
nor U7679 (N_7679,N_4523,N_4532);
or U7680 (N_7680,N_4112,N_5306);
nand U7681 (N_7681,N_4606,N_5986);
nor U7682 (N_7682,N_5805,N_5489);
nor U7683 (N_7683,N_4136,N_5770);
and U7684 (N_7684,N_5139,N_4343);
nand U7685 (N_7685,N_4914,N_4810);
or U7686 (N_7686,N_5552,N_5704);
and U7687 (N_7687,N_4877,N_5625);
and U7688 (N_7688,N_5986,N_5780);
nor U7689 (N_7689,N_5933,N_5391);
xor U7690 (N_7690,N_5525,N_4728);
and U7691 (N_7691,N_5941,N_5871);
nand U7692 (N_7692,N_4496,N_4818);
nand U7693 (N_7693,N_4694,N_4409);
nor U7694 (N_7694,N_4505,N_5388);
or U7695 (N_7695,N_5559,N_4638);
or U7696 (N_7696,N_5061,N_4745);
or U7697 (N_7697,N_4155,N_4981);
and U7698 (N_7698,N_4869,N_4665);
or U7699 (N_7699,N_5612,N_5288);
nor U7700 (N_7700,N_4950,N_4482);
or U7701 (N_7701,N_4732,N_5127);
and U7702 (N_7702,N_4887,N_5483);
nor U7703 (N_7703,N_4402,N_5048);
or U7704 (N_7704,N_5982,N_4736);
nand U7705 (N_7705,N_5473,N_4832);
nor U7706 (N_7706,N_5485,N_5651);
or U7707 (N_7707,N_4317,N_5292);
or U7708 (N_7708,N_5447,N_5674);
nand U7709 (N_7709,N_4661,N_5638);
nand U7710 (N_7710,N_4731,N_4116);
xor U7711 (N_7711,N_4556,N_4736);
nor U7712 (N_7712,N_5379,N_4609);
nor U7713 (N_7713,N_4960,N_5740);
nor U7714 (N_7714,N_5287,N_4199);
or U7715 (N_7715,N_4469,N_4331);
or U7716 (N_7716,N_5805,N_5893);
or U7717 (N_7717,N_4789,N_4356);
nand U7718 (N_7718,N_4914,N_4923);
or U7719 (N_7719,N_4605,N_5214);
and U7720 (N_7720,N_5146,N_5995);
and U7721 (N_7721,N_4929,N_5917);
and U7722 (N_7722,N_5162,N_5355);
and U7723 (N_7723,N_4456,N_5824);
and U7724 (N_7724,N_4443,N_5733);
or U7725 (N_7725,N_4824,N_5226);
or U7726 (N_7726,N_4124,N_5450);
nand U7727 (N_7727,N_5353,N_5871);
or U7728 (N_7728,N_5693,N_5912);
and U7729 (N_7729,N_4263,N_5745);
and U7730 (N_7730,N_4488,N_5330);
nor U7731 (N_7731,N_5061,N_4467);
nor U7732 (N_7732,N_4590,N_4831);
nor U7733 (N_7733,N_5860,N_5587);
nor U7734 (N_7734,N_5303,N_5710);
nand U7735 (N_7735,N_5649,N_4123);
and U7736 (N_7736,N_5979,N_4475);
and U7737 (N_7737,N_4404,N_4722);
nor U7738 (N_7738,N_5250,N_4894);
and U7739 (N_7739,N_5871,N_4424);
or U7740 (N_7740,N_5312,N_4776);
nor U7741 (N_7741,N_5646,N_5968);
nand U7742 (N_7742,N_5453,N_5671);
nor U7743 (N_7743,N_4371,N_4451);
xnor U7744 (N_7744,N_5838,N_4016);
or U7745 (N_7745,N_4835,N_5830);
xor U7746 (N_7746,N_4015,N_5107);
nand U7747 (N_7747,N_5579,N_4876);
nor U7748 (N_7748,N_5541,N_4306);
or U7749 (N_7749,N_5129,N_4837);
nand U7750 (N_7750,N_4680,N_5677);
and U7751 (N_7751,N_5592,N_4121);
nand U7752 (N_7752,N_5144,N_4709);
and U7753 (N_7753,N_5271,N_5397);
nand U7754 (N_7754,N_5544,N_5321);
nor U7755 (N_7755,N_5188,N_4261);
nor U7756 (N_7756,N_5505,N_4342);
nand U7757 (N_7757,N_4186,N_5314);
or U7758 (N_7758,N_5088,N_4640);
nand U7759 (N_7759,N_4604,N_4711);
or U7760 (N_7760,N_4113,N_4803);
or U7761 (N_7761,N_5613,N_5060);
nor U7762 (N_7762,N_4006,N_4247);
nor U7763 (N_7763,N_4923,N_5415);
or U7764 (N_7764,N_5675,N_5776);
nand U7765 (N_7765,N_4510,N_4853);
xor U7766 (N_7766,N_5870,N_4026);
and U7767 (N_7767,N_4347,N_5841);
and U7768 (N_7768,N_5479,N_5344);
nand U7769 (N_7769,N_4319,N_5828);
nand U7770 (N_7770,N_4325,N_4108);
xor U7771 (N_7771,N_4233,N_4159);
nor U7772 (N_7772,N_4837,N_5367);
and U7773 (N_7773,N_4871,N_4543);
nand U7774 (N_7774,N_4698,N_4045);
and U7775 (N_7775,N_4516,N_4122);
or U7776 (N_7776,N_4354,N_5242);
and U7777 (N_7777,N_4217,N_4114);
or U7778 (N_7778,N_4958,N_5144);
xnor U7779 (N_7779,N_4844,N_5239);
and U7780 (N_7780,N_5375,N_4986);
and U7781 (N_7781,N_4466,N_4113);
nand U7782 (N_7782,N_4154,N_4668);
nor U7783 (N_7783,N_5622,N_4131);
and U7784 (N_7784,N_5228,N_4137);
and U7785 (N_7785,N_5795,N_5375);
or U7786 (N_7786,N_4176,N_4941);
nor U7787 (N_7787,N_5458,N_4574);
nor U7788 (N_7788,N_4863,N_4121);
or U7789 (N_7789,N_4459,N_4466);
xnor U7790 (N_7790,N_5189,N_5914);
or U7791 (N_7791,N_5009,N_4119);
xnor U7792 (N_7792,N_4007,N_5504);
or U7793 (N_7793,N_5688,N_4644);
and U7794 (N_7794,N_4878,N_5290);
nand U7795 (N_7795,N_5003,N_4952);
and U7796 (N_7796,N_4171,N_4326);
xnor U7797 (N_7797,N_5985,N_5491);
and U7798 (N_7798,N_4615,N_5055);
nor U7799 (N_7799,N_4323,N_5580);
or U7800 (N_7800,N_4071,N_4175);
and U7801 (N_7801,N_4124,N_4116);
nand U7802 (N_7802,N_5649,N_4508);
nor U7803 (N_7803,N_4422,N_5122);
and U7804 (N_7804,N_5668,N_4055);
nand U7805 (N_7805,N_4131,N_4795);
and U7806 (N_7806,N_5311,N_5491);
nor U7807 (N_7807,N_4201,N_5562);
nand U7808 (N_7808,N_5572,N_5350);
nor U7809 (N_7809,N_4525,N_5136);
and U7810 (N_7810,N_4406,N_4831);
nor U7811 (N_7811,N_5240,N_4813);
and U7812 (N_7812,N_4219,N_4162);
and U7813 (N_7813,N_5996,N_4550);
or U7814 (N_7814,N_5434,N_5492);
xor U7815 (N_7815,N_4150,N_5439);
xor U7816 (N_7816,N_5949,N_4704);
nor U7817 (N_7817,N_4855,N_5695);
or U7818 (N_7818,N_4595,N_4505);
and U7819 (N_7819,N_4660,N_5187);
or U7820 (N_7820,N_5468,N_5168);
and U7821 (N_7821,N_4298,N_4077);
and U7822 (N_7822,N_4989,N_5805);
nor U7823 (N_7823,N_4580,N_5210);
nor U7824 (N_7824,N_4644,N_5757);
and U7825 (N_7825,N_4963,N_4799);
nand U7826 (N_7826,N_5854,N_4400);
xor U7827 (N_7827,N_5507,N_5153);
nor U7828 (N_7828,N_5231,N_4849);
or U7829 (N_7829,N_4307,N_5612);
nor U7830 (N_7830,N_4108,N_4267);
and U7831 (N_7831,N_5172,N_4973);
nand U7832 (N_7832,N_4249,N_4281);
xnor U7833 (N_7833,N_5280,N_4757);
nand U7834 (N_7834,N_5284,N_4623);
nor U7835 (N_7835,N_4344,N_5242);
and U7836 (N_7836,N_5160,N_5128);
xor U7837 (N_7837,N_5315,N_4950);
nor U7838 (N_7838,N_4850,N_5316);
nor U7839 (N_7839,N_4596,N_5053);
and U7840 (N_7840,N_4922,N_5558);
or U7841 (N_7841,N_4813,N_5931);
nor U7842 (N_7842,N_5795,N_4371);
or U7843 (N_7843,N_4603,N_5124);
and U7844 (N_7844,N_5163,N_5443);
and U7845 (N_7845,N_4203,N_5703);
or U7846 (N_7846,N_5864,N_4367);
nand U7847 (N_7847,N_4530,N_4874);
and U7848 (N_7848,N_5626,N_5446);
or U7849 (N_7849,N_5122,N_4743);
and U7850 (N_7850,N_5403,N_5420);
nor U7851 (N_7851,N_4164,N_5475);
or U7852 (N_7852,N_5630,N_5335);
nand U7853 (N_7853,N_5702,N_5839);
nand U7854 (N_7854,N_5141,N_5398);
nand U7855 (N_7855,N_5542,N_4145);
nand U7856 (N_7856,N_5565,N_5078);
nor U7857 (N_7857,N_4530,N_5877);
and U7858 (N_7858,N_4126,N_5458);
nand U7859 (N_7859,N_5681,N_5806);
and U7860 (N_7860,N_5373,N_4002);
or U7861 (N_7861,N_5306,N_5081);
nand U7862 (N_7862,N_4400,N_5256);
or U7863 (N_7863,N_4261,N_4915);
and U7864 (N_7864,N_5286,N_4359);
and U7865 (N_7865,N_5453,N_4365);
or U7866 (N_7866,N_5907,N_4216);
or U7867 (N_7867,N_5653,N_5950);
or U7868 (N_7868,N_4042,N_5182);
or U7869 (N_7869,N_5186,N_5446);
and U7870 (N_7870,N_4741,N_4416);
nand U7871 (N_7871,N_5966,N_4878);
nor U7872 (N_7872,N_5135,N_4351);
or U7873 (N_7873,N_4547,N_5974);
nand U7874 (N_7874,N_4815,N_5794);
nor U7875 (N_7875,N_5905,N_5851);
xnor U7876 (N_7876,N_4209,N_5159);
nand U7877 (N_7877,N_4750,N_5205);
or U7878 (N_7878,N_5278,N_4587);
nand U7879 (N_7879,N_4844,N_4370);
and U7880 (N_7880,N_5942,N_5020);
nand U7881 (N_7881,N_4849,N_4705);
xnor U7882 (N_7882,N_4646,N_5848);
nand U7883 (N_7883,N_4429,N_5624);
or U7884 (N_7884,N_5348,N_4302);
nand U7885 (N_7885,N_4358,N_4602);
or U7886 (N_7886,N_4180,N_5611);
or U7887 (N_7887,N_4953,N_4691);
nand U7888 (N_7888,N_4680,N_4811);
nand U7889 (N_7889,N_5095,N_4876);
xnor U7890 (N_7890,N_5103,N_4554);
or U7891 (N_7891,N_5711,N_4303);
nor U7892 (N_7892,N_5841,N_4725);
or U7893 (N_7893,N_5956,N_4658);
nor U7894 (N_7894,N_4924,N_4344);
and U7895 (N_7895,N_5202,N_5086);
or U7896 (N_7896,N_5280,N_5527);
nand U7897 (N_7897,N_4141,N_4098);
or U7898 (N_7898,N_4106,N_5269);
and U7899 (N_7899,N_5685,N_5548);
xnor U7900 (N_7900,N_5572,N_5445);
and U7901 (N_7901,N_4727,N_4094);
nor U7902 (N_7902,N_4944,N_4308);
nand U7903 (N_7903,N_5362,N_4422);
nor U7904 (N_7904,N_5839,N_5802);
and U7905 (N_7905,N_4759,N_4529);
nand U7906 (N_7906,N_4307,N_4594);
nand U7907 (N_7907,N_5277,N_4338);
xnor U7908 (N_7908,N_4761,N_5711);
and U7909 (N_7909,N_4495,N_5851);
nand U7910 (N_7910,N_4250,N_5329);
or U7911 (N_7911,N_4941,N_5890);
and U7912 (N_7912,N_4809,N_4661);
nor U7913 (N_7913,N_5924,N_4888);
and U7914 (N_7914,N_5126,N_5362);
nor U7915 (N_7915,N_5086,N_5404);
or U7916 (N_7916,N_5233,N_4813);
and U7917 (N_7917,N_4972,N_4094);
nor U7918 (N_7918,N_5281,N_4647);
nor U7919 (N_7919,N_4383,N_5911);
and U7920 (N_7920,N_5392,N_5647);
xor U7921 (N_7921,N_4792,N_4357);
nor U7922 (N_7922,N_5628,N_4560);
and U7923 (N_7923,N_4969,N_5405);
or U7924 (N_7924,N_4955,N_4524);
or U7925 (N_7925,N_4655,N_4608);
and U7926 (N_7926,N_5000,N_5823);
nor U7927 (N_7927,N_5356,N_4549);
and U7928 (N_7928,N_4999,N_4660);
or U7929 (N_7929,N_4398,N_4372);
or U7930 (N_7930,N_5425,N_4645);
nand U7931 (N_7931,N_5995,N_4175);
and U7932 (N_7932,N_5993,N_4713);
nor U7933 (N_7933,N_5774,N_5324);
nor U7934 (N_7934,N_5639,N_4039);
or U7935 (N_7935,N_5513,N_5751);
and U7936 (N_7936,N_4277,N_5848);
and U7937 (N_7937,N_5042,N_4309);
nand U7938 (N_7938,N_4610,N_5044);
nor U7939 (N_7939,N_4586,N_4181);
xor U7940 (N_7940,N_4485,N_4122);
and U7941 (N_7941,N_4838,N_4677);
or U7942 (N_7942,N_5095,N_4560);
or U7943 (N_7943,N_4799,N_4275);
or U7944 (N_7944,N_5796,N_5149);
xor U7945 (N_7945,N_5532,N_4495);
nor U7946 (N_7946,N_4247,N_5337);
or U7947 (N_7947,N_4916,N_5007);
or U7948 (N_7948,N_4344,N_4151);
or U7949 (N_7949,N_5371,N_4610);
nand U7950 (N_7950,N_4103,N_4446);
or U7951 (N_7951,N_4872,N_5773);
or U7952 (N_7952,N_4926,N_4597);
xor U7953 (N_7953,N_4012,N_4271);
xnor U7954 (N_7954,N_4218,N_4775);
xnor U7955 (N_7955,N_4597,N_4258);
nor U7956 (N_7956,N_4868,N_5226);
or U7957 (N_7957,N_5549,N_5199);
xnor U7958 (N_7958,N_5939,N_5181);
nor U7959 (N_7959,N_4900,N_5728);
and U7960 (N_7960,N_5061,N_5778);
nand U7961 (N_7961,N_4186,N_5511);
nor U7962 (N_7962,N_5450,N_4145);
nand U7963 (N_7963,N_5025,N_5730);
nand U7964 (N_7964,N_4325,N_4427);
and U7965 (N_7965,N_4975,N_5287);
or U7966 (N_7966,N_5445,N_4670);
nand U7967 (N_7967,N_4360,N_4730);
or U7968 (N_7968,N_4896,N_5199);
nor U7969 (N_7969,N_5230,N_5231);
and U7970 (N_7970,N_4586,N_4951);
or U7971 (N_7971,N_5185,N_5681);
and U7972 (N_7972,N_4373,N_4853);
xor U7973 (N_7973,N_4755,N_5036);
and U7974 (N_7974,N_4511,N_4043);
nand U7975 (N_7975,N_4743,N_5133);
and U7976 (N_7976,N_5050,N_5268);
and U7977 (N_7977,N_5572,N_5621);
or U7978 (N_7978,N_5798,N_4577);
or U7979 (N_7979,N_5201,N_5053);
and U7980 (N_7980,N_4225,N_4558);
and U7981 (N_7981,N_5779,N_5034);
or U7982 (N_7982,N_5340,N_4719);
nor U7983 (N_7983,N_5686,N_5061);
xnor U7984 (N_7984,N_4174,N_5775);
nor U7985 (N_7985,N_4041,N_5029);
nand U7986 (N_7986,N_5863,N_5756);
nor U7987 (N_7987,N_5377,N_5362);
nor U7988 (N_7988,N_5552,N_5324);
nor U7989 (N_7989,N_5644,N_4163);
or U7990 (N_7990,N_4429,N_4672);
nand U7991 (N_7991,N_4678,N_4446);
or U7992 (N_7992,N_4273,N_4207);
nor U7993 (N_7993,N_5578,N_5177);
xor U7994 (N_7994,N_5716,N_4491);
or U7995 (N_7995,N_4567,N_4925);
xor U7996 (N_7996,N_4665,N_4724);
nor U7997 (N_7997,N_4204,N_4423);
or U7998 (N_7998,N_5124,N_5182);
or U7999 (N_7999,N_4884,N_5123);
and U8000 (N_8000,N_6022,N_6037);
and U8001 (N_8001,N_7019,N_6134);
and U8002 (N_8002,N_7041,N_6939);
nand U8003 (N_8003,N_6155,N_6408);
and U8004 (N_8004,N_6108,N_7875);
or U8005 (N_8005,N_7249,N_6757);
nor U8006 (N_8006,N_6700,N_7299);
xnor U8007 (N_8007,N_6528,N_6922);
nor U8008 (N_8008,N_7114,N_6925);
nand U8009 (N_8009,N_6815,N_7047);
or U8010 (N_8010,N_7971,N_6237);
nand U8011 (N_8011,N_6977,N_6906);
or U8012 (N_8012,N_7457,N_7731);
nand U8013 (N_8013,N_6090,N_6550);
and U8014 (N_8014,N_6872,N_6603);
and U8015 (N_8015,N_7310,N_6156);
nor U8016 (N_8016,N_6869,N_6904);
nor U8017 (N_8017,N_6209,N_6665);
nor U8018 (N_8018,N_6918,N_7754);
nand U8019 (N_8019,N_7077,N_7654);
nor U8020 (N_8020,N_6396,N_6173);
or U8021 (N_8021,N_6082,N_6505);
or U8022 (N_8022,N_6152,N_6766);
nand U8023 (N_8023,N_6667,N_6792);
or U8024 (N_8024,N_7984,N_7336);
nor U8025 (N_8025,N_6614,N_6126);
and U8026 (N_8026,N_6558,N_6067);
and U8027 (N_8027,N_6107,N_6187);
or U8028 (N_8028,N_7980,N_6099);
xnor U8029 (N_8029,N_6048,N_7843);
and U8030 (N_8030,N_6071,N_6739);
xor U8031 (N_8031,N_6199,N_7431);
nand U8032 (N_8032,N_7623,N_7451);
nor U8033 (N_8033,N_7831,N_6938);
xnor U8034 (N_8034,N_7344,N_6282);
nor U8035 (N_8035,N_7347,N_6125);
xor U8036 (N_8036,N_7696,N_6324);
or U8037 (N_8037,N_6449,N_7528);
xor U8038 (N_8038,N_6537,N_6901);
or U8039 (N_8039,N_6804,N_7750);
nor U8040 (N_8040,N_7246,N_7964);
nand U8041 (N_8041,N_7710,N_7278);
nand U8042 (N_8042,N_6623,N_7543);
nand U8043 (N_8043,N_6238,N_6086);
and U8044 (N_8044,N_7479,N_6276);
nand U8045 (N_8045,N_7008,N_6470);
or U8046 (N_8046,N_7178,N_6327);
nand U8047 (N_8047,N_7550,N_7760);
nand U8048 (N_8048,N_7301,N_6670);
nand U8049 (N_8049,N_7380,N_7179);
nand U8050 (N_8050,N_7627,N_6560);
and U8051 (N_8051,N_6926,N_7641);
nand U8052 (N_8052,N_6244,N_7507);
nand U8053 (N_8053,N_7578,N_7912);
and U8054 (N_8054,N_6229,N_7022);
nor U8055 (N_8055,N_7613,N_7144);
nand U8056 (N_8056,N_6095,N_6512);
or U8057 (N_8057,N_7902,N_6171);
or U8058 (N_8058,N_6932,N_7602);
nand U8059 (N_8059,N_7165,N_7872);
nor U8060 (N_8060,N_7481,N_6672);
and U8061 (N_8061,N_6378,N_6823);
nor U8062 (N_8062,N_6898,N_6930);
nand U8063 (N_8063,N_7597,N_6601);
and U8064 (N_8064,N_7515,N_6666);
nand U8065 (N_8065,N_7671,N_7115);
and U8066 (N_8066,N_7617,N_7261);
nor U8067 (N_8067,N_6397,N_6338);
xor U8068 (N_8068,N_6690,N_6681);
nor U8069 (N_8069,N_6159,N_6969);
nand U8070 (N_8070,N_7333,N_7498);
nand U8071 (N_8071,N_6629,N_6749);
or U8072 (N_8072,N_6120,N_7653);
nand U8073 (N_8073,N_7871,N_6006);
or U8074 (N_8074,N_6085,N_6825);
and U8075 (N_8075,N_7348,N_6363);
or U8076 (N_8076,N_7183,N_6870);
nand U8077 (N_8077,N_7109,N_6250);
nand U8078 (N_8078,N_7921,N_6440);
nor U8079 (N_8079,N_6599,N_7052);
and U8080 (N_8080,N_6060,N_7820);
and U8081 (N_8081,N_6716,N_7640);
and U8082 (N_8082,N_6389,N_6230);
and U8083 (N_8083,N_7462,N_6754);
and U8084 (N_8084,N_6794,N_6203);
and U8085 (N_8085,N_6343,N_7112);
or U8086 (N_8086,N_7447,N_6551);
or U8087 (N_8087,N_6542,N_7016);
or U8088 (N_8088,N_6581,N_7232);
xnor U8089 (N_8089,N_7535,N_6952);
and U8090 (N_8090,N_6758,N_7928);
and U8091 (N_8091,N_7706,N_6163);
and U8092 (N_8092,N_6136,N_7590);
and U8093 (N_8093,N_6088,N_7419);
and U8094 (N_8094,N_7588,N_7312);
and U8095 (N_8095,N_7197,N_7726);
nor U8096 (N_8096,N_7327,N_7734);
or U8097 (N_8097,N_6744,N_7905);
and U8098 (N_8098,N_7104,N_7832);
xnor U8099 (N_8099,N_7932,N_6101);
nand U8100 (N_8100,N_6721,N_7885);
nand U8101 (N_8101,N_7811,N_7961);
or U8102 (N_8102,N_7054,N_6308);
nand U8103 (N_8103,N_7725,N_7676);
and U8104 (N_8104,N_7199,N_7877);
nand U8105 (N_8105,N_6349,N_7445);
or U8106 (N_8106,N_7544,N_6764);
nand U8107 (N_8107,N_6046,N_7367);
nand U8108 (N_8108,N_6401,N_6944);
or U8109 (N_8109,N_6009,N_6236);
or U8110 (N_8110,N_7323,N_6279);
nand U8111 (N_8111,N_6717,N_7924);
nand U8112 (N_8112,N_6761,N_6169);
nor U8113 (N_8113,N_7596,N_6117);
and U8114 (N_8114,N_6743,N_7275);
and U8115 (N_8115,N_6891,N_6604);
or U8116 (N_8116,N_6856,N_6026);
nor U8117 (N_8117,N_7615,N_7945);
nor U8118 (N_8118,N_7709,N_6042);
or U8119 (N_8119,N_7252,N_6424);
or U8120 (N_8120,N_7891,N_7707);
nand U8121 (N_8121,N_6875,N_6049);
or U8122 (N_8122,N_6772,N_6266);
and U8123 (N_8123,N_6678,N_7430);
and U8124 (N_8124,N_7878,N_7659);
or U8125 (N_8125,N_7079,N_6927);
or U8126 (N_8126,N_6735,N_6121);
nor U8127 (N_8127,N_7700,N_7340);
nor U8128 (N_8128,N_7170,N_7120);
nor U8129 (N_8129,N_7857,N_6987);
or U8130 (N_8130,N_7387,N_6642);
and U8131 (N_8131,N_7014,N_6723);
and U8132 (N_8132,N_6016,N_6162);
or U8133 (N_8133,N_7386,N_6303);
and U8134 (N_8134,N_7744,N_6495);
or U8135 (N_8135,N_7551,N_6563);
or U8136 (N_8136,N_7554,N_7149);
and U8137 (N_8137,N_6083,N_7352);
and U8138 (N_8138,N_7258,N_6445);
or U8139 (N_8139,N_7168,N_6784);
or U8140 (N_8140,N_7009,N_7247);
or U8141 (N_8141,N_6168,N_7593);
nand U8142 (N_8142,N_6588,N_6684);
or U8143 (N_8143,N_6624,N_6316);
xor U8144 (N_8144,N_6641,N_7722);
and U8145 (N_8145,N_6334,N_6701);
nand U8146 (N_8146,N_7316,N_7791);
nor U8147 (N_8147,N_7856,N_7598);
nor U8148 (N_8148,N_6274,N_6552);
nor U8149 (N_8149,N_7089,N_6079);
and U8150 (N_8150,N_7043,N_7088);
or U8151 (N_8151,N_7600,N_6549);
nor U8152 (N_8152,N_6381,N_6267);
and U8153 (N_8153,N_7748,N_6142);
and U8154 (N_8154,N_7156,N_6995);
nand U8155 (N_8155,N_7205,N_7783);
or U8156 (N_8156,N_6834,N_7509);
or U8157 (N_8157,N_7682,N_7500);
nand U8158 (N_8158,N_6714,N_7514);
nor U8159 (N_8159,N_7879,N_7814);
nor U8160 (N_8160,N_7787,N_7901);
xor U8161 (N_8161,N_7440,N_7918);
nor U8162 (N_8162,N_7745,N_6565);
and U8163 (N_8163,N_6779,N_6135);
and U8164 (N_8164,N_6473,N_7495);
nand U8165 (N_8165,N_7582,N_6427);
nand U8166 (N_8166,N_6353,N_6269);
or U8167 (N_8167,N_7798,N_7675);
or U8168 (N_8168,N_6289,N_7473);
nor U8169 (N_8169,N_7045,N_6262);
nand U8170 (N_8170,N_6814,N_7900);
and U8171 (N_8171,N_6568,N_6184);
and U8172 (N_8172,N_6387,N_7240);
nor U8173 (N_8173,N_6265,N_7715);
or U8174 (N_8174,N_7066,N_6509);
or U8175 (N_8175,N_6727,N_6172);
and U8176 (N_8176,N_7632,N_6731);
or U8177 (N_8177,N_6031,N_6971);
and U8178 (N_8178,N_6688,N_6695);
or U8179 (N_8179,N_7753,N_6972);
and U8180 (N_8180,N_7191,N_6093);
nor U8181 (N_8181,N_7137,N_6076);
or U8182 (N_8182,N_6801,N_7893);
and U8183 (N_8183,N_6878,N_7307);
or U8184 (N_8184,N_7983,N_7095);
nor U8185 (N_8185,N_7004,N_7609);
and U8186 (N_8186,N_7525,N_7353);
and U8187 (N_8187,N_6294,N_6439);
or U8188 (N_8188,N_6531,N_6837);
and U8189 (N_8189,N_6907,N_7176);
nor U8190 (N_8190,N_7082,N_6235);
xnor U8191 (N_8191,N_7883,N_6617);
nand U8192 (N_8192,N_6242,N_7237);
nand U8193 (N_8193,N_7174,N_7434);
or U8194 (N_8194,N_6256,N_6566);
xor U8195 (N_8195,N_7011,N_7822);
or U8196 (N_8196,N_7366,N_6057);
or U8197 (N_8197,N_6021,N_6367);
and U8198 (N_8198,N_7889,N_7776);
or U8199 (N_8199,N_6336,N_7084);
nand U8200 (N_8200,N_7230,N_6973);
nor U8201 (N_8201,N_6065,N_6992);
and U8202 (N_8202,N_6354,N_6719);
nor U8203 (N_8203,N_6619,N_7086);
and U8204 (N_8204,N_7331,N_6506);
or U8205 (N_8205,N_7560,N_6207);
and U8206 (N_8206,N_6958,N_7000);
nor U8207 (N_8207,N_7920,N_6243);
and U8208 (N_8208,N_7134,N_6680);
or U8209 (N_8209,N_7127,N_7573);
nor U8210 (N_8210,N_7385,N_6945);
and U8211 (N_8211,N_6943,N_7839);
nand U8212 (N_8212,N_6472,N_7255);
or U8213 (N_8213,N_7061,N_7703);
nor U8214 (N_8214,N_7770,N_7780);
or U8215 (N_8215,N_7553,N_7250);
xor U8216 (N_8216,N_7065,N_6249);
and U8217 (N_8217,N_6188,N_7181);
or U8218 (N_8218,N_6544,N_6061);
xor U8219 (N_8219,N_6824,N_7136);
nand U8220 (N_8220,N_6038,N_6307);
or U8221 (N_8221,N_6051,N_7256);
and U8222 (N_8222,N_7827,N_6302);
and U8223 (N_8223,N_6423,N_7142);
or U8224 (N_8224,N_6632,N_7674);
and U8225 (N_8225,N_7332,N_6489);
or U8226 (N_8226,N_7433,N_6074);
nor U8227 (N_8227,N_6385,N_6287);
nand U8228 (N_8228,N_6379,N_7489);
nand U8229 (N_8229,N_7378,N_7542);
and U8230 (N_8230,N_7465,N_6131);
nand U8231 (N_8231,N_6689,N_7630);
nor U8232 (N_8232,N_7482,N_6477);
nand U8233 (N_8233,N_7953,N_6010);
nor U8234 (N_8234,N_6840,N_7098);
and U8235 (N_8235,N_7586,N_7665);
or U8236 (N_8236,N_6790,N_6193);
nor U8237 (N_8237,N_7618,N_7383);
or U8238 (N_8238,N_7412,N_7496);
nand U8239 (N_8239,N_7775,N_7846);
nand U8240 (N_8240,N_7037,N_7569);
and U8241 (N_8241,N_6948,N_6319);
nand U8242 (N_8242,N_7797,N_6015);
or U8243 (N_8243,N_6504,N_6873);
and U8244 (N_8244,N_7794,N_7155);
or U8245 (N_8245,N_6503,N_6756);
xnor U8246 (N_8246,N_6725,N_6127);
nor U8247 (N_8247,N_7426,N_7592);
xnor U8248 (N_8248,N_7202,N_6115);
nor U8249 (N_8249,N_7314,N_7030);
nor U8250 (N_8250,N_6584,N_6807);
nand U8251 (N_8251,N_6024,N_6874);
nand U8252 (N_8252,N_7666,N_7309);
and U8253 (N_8253,N_7313,N_6080);
or U8254 (N_8254,N_6299,N_6747);
xnor U8255 (N_8255,N_7979,N_7923);
and U8256 (N_8256,N_7236,N_7903);
and U8257 (N_8257,N_6218,N_6532);
and U8258 (N_8258,N_7097,N_6668);
nor U8259 (N_8259,N_6017,N_6377);
nor U8260 (N_8260,N_6315,N_7636);
nor U8261 (N_8261,N_6631,N_6774);
nor U8262 (N_8262,N_6194,N_7152);
nor U8263 (N_8263,N_7799,N_6803);
or U8264 (N_8264,N_6529,N_7954);
nor U8265 (N_8265,N_6593,N_6350);
and U8266 (N_8266,N_6097,N_6261);
or U8267 (N_8267,N_6252,N_7204);
and U8268 (N_8268,N_6114,N_7933);
nor U8269 (N_8269,N_6750,N_7420);
xor U8270 (N_8270,N_7015,N_6333);
nand U8271 (N_8271,N_7239,N_7169);
and U8272 (N_8272,N_6111,N_6513);
or U8273 (N_8273,N_7955,N_7616);
or U8274 (N_8274,N_7881,N_7716);
nand U8275 (N_8275,N_7579,N_7017);
and U8276 (N_8276,N_6166,N_7940);
nor U8277 (N_8277,N_6594,N_6443);
nand U8278 (N_8278,N_6459,N_6637);
and U8279 (N_8279,N_6070,N_7806);
xnor U8280 (N_8280,N_7994,N_6956);
nand U8281 (N_8281,N_7564,N_6069);
nor U8282 (N_8282,N_7439,N_6888);
nor U8283 (N_8283,N_7406,N_7192);
and U8284 (N_8284,N_6149,N_6013);
and U8285 (N_8285,N_6775,N_6094);
or U8286 (N_8286,N_6369,N_6933);
nand U8287 (N_8287,N_6413,N_7003);
or U8288 (N_8288,N_7294,N_7093);
or U8289 (N_8289,N_6182,N_6399);
or U8290 (N_8290,N_6283,N_7053);
and U8291 (N_8291,N_7742,N_6519);
xor U8292 (N_8292,N_6521,N_7492);
nor U8293 (N_8293,N_7375,N_6534);
or U8294 (N_8294,N_7849,N_7736);
nor U8295 (N_8295,N_7576,N_7391);
nor U8296 (N_8296,N_6292,N_7801);
and U8297 (N_8297,N_7935,N_6019);
nand U8298 (N_8298,N_6064,N_7215);
and U8299 (N_8299,N_6241,N_6795);
and U8300 (N_8300,N_6044,N_6966);
and U8301 (N_8301,N_6066,N_7368);
or U8302 (N_8302,N_7601,N_6452);
or U8303 (N_8303,N_6416,N_6373);
or U8304 (N_8304,N_6983,N_7823);
xnor U8305 (N_8305,N_7854,N_7096);
and U8306 (N_8306,N_7410,N_6596);
nand U8307 (N_8307,N_7010,N_7488);
nand U8308 (N_8308,N_7062,N_7511);
or U8309 (N_8309,N_7425,N_7999);
or U8310 (N_8310,N_7407,N_6818);
xnor U8311 (N_8311,N_7182,N_7944);
or U8312 (N_8312,N_6682,N_7946);
or U8313 (N_8313,N_7398,N_7397);
or U8314 (N_8314,N_6612,N_6417);
nor U8315 (N_8315,N_7159,N_7752);
nand U8316 (N_8316,N_7282,N_7677);
nand U8317 (N_8317,N_6540,N_6358);
or U8318 (N_8318,N_7860,N_7080);
and U8319 (N_8319,N_7619,N_7223);
nor U8320 (N_8320,N_7504,N_7289);
or U8321 (N_8321,N_7320,N_6579);
and U8322 (N_8322,N_7334,N_7816);
nand U8323 (N_8323,N_6164,N_7284);
nand U8324 (N_8324,N_6949,N_6909);
xor U8325 (N_8325,N_7468,N_6838);
nor U8326 (N_8326,N_7184,N_7886);
and U8327 (N_8327,N_7116,N_7241);
or U8328 (N_8328,N_6848,N_7264);
nor U8329 (N_8329,N_6635,N_6810);
nand U8330 (N_8330,N_7370,N_6778);
nand U8331 (N_8331,N_6900,N_6738);
xnor U8332 (N_8332,N_7563,N_6222);
xnor U8333 (N_8333,N_6616,N_6650);
nand U8334 (N_8334,N_7486,N_7304);
and U8335 (N_8335,N_7568,N_6864);
and U8336 (N_8336,N_7648,N_6997);
or U8337 (N_8337,N_7916,N_6685);
nor U8338 (N_8338,N_7911,N_7833);
nand U8339 (N_8339,N_7899,N_7807);
xor U8340 (N_8340,N_6102,N_7416);
or U8341 (N_8341,N_7638,N_6479);
nand U8342 (N_8342,N_6311,N_7730);
nor U8343 (N_8343,N_6760,N_6686);
and U8344 (N_8344,N_6862,N_7821);
and U8345 (N_8345,N_7975,N_7987);
nor U8346 (N_8346,N_6830,N_7728);
nand U8347 (N_8347,N_7358,N_6419);
or U8348 (N_8348,N_6465,N_6858);
nor U8349 (N_8349,N_6677,N_7941);
or U8350 (N_8350,N_7035,N_7478);
or U8351 (N_8351,N_6729,N_7669);
nand U8352 (N_8352,N_7122,N_7458);
and U8353 (N_8353,N_6713,N_7218);
nor U8354 (N_8354,N_6365,N_7529);
or U8355 (N_8355,N_6989,N_6897);
nor U8356 (N_8356,N_6857,N_6675);
nand U8357 (N_8357,N_6751,N_6454);
xnor U8358 (N_8358,N_6260,N_7540);
and U8359 (N_8359,N_7143,N_7815);
nor U8360 (N_8360,N_6105,N_6212);
nor U8361 (N_8361,N_7200,N_7896);
xnor U8362 (N_8362,N_6232,N_6765);
nor U8363 (N_8363,N_6482,N_7534);
and U8364 (N_8364,N_6518,N_7712);
nor U8365 (N_8365,N_7253,N_7063);
xor U8366 (N_8366,N_6297,N_7581);
and U8367 (N_8367,N_7664,N_7283);
and U8368 (N_8368,N_7865,N_6029);
nor U8369 (N_8369,N_7992,N_7271);
xnor U8370 (N_8370,N_6430,N_7888);
nand U8371 (N_8371,N_7698,N_6257);
nor U8372 (N_8372,N_7490,N_7840);
nor U8373 (N_8373,N_7138,N_7389);
nor U8374 (N_8374,N_7390,N_7296);
and U8375 (N_8375,N_7343,N_6598);
nand U8376 (N_8376,N_6447,N_6106);
or U8377 (N_8377,N_7652,N_6595);
nand U8378 (N_8378,N_7873,N_7032);
or U8379 (N_8379,N_7424,N_7107);
and U8380 (N_8380,N_7810,N_6174);
or U8381 (N_8381,N_6317,N_6640);
or U8382 (N_8382,N_6050,N_6915);
nor U8383 (N_8383,N_6457,N_7128);
and U8384 (N_8384,N_7910,N_7673);
xnor U8385 (N_8385,N_6411,N_7056);
or U8386 (N_8386,N_6832,N_6905);
and U8387 (N_8387,N_7245,N_6782);
nor U8388 (N_8388,N_7639,N_6696);
nor U8389 (N_8389,N_6376,N_6464);
or U8390 (N_8390,N_7476,N_6841);
and U8391 (N_8391,N_7020,N_7996);
xor U8392 (N_8392,N_6582,N_7771);
nor U8393 (N_8393,N_7235,N_7704);
xor U8394 (N_8394,N_7028,N_6546);
or U8395 (N_8395,N_6366,N_6177);
and U8396 (N_8396,N_6609,N_6318);
nor U8397 (N_8397,N_7790,N_7254);
nand U8398 (N_8398,N_6003,N_6910);
and U8399 (N_8399,N_7870,N_6104);
nor U8400 (N_8400,N_7546,N_7263);
and U8401 (N_8401,N_6855,N_6310);
nor U8402 (N_8402,N_7212,N_7038);
xor U8403 (N_8403,N_6895,N_7007);
nand U8404 (N_8404,N_6362,N_6852);
or U8405 (N_8405,N_7029,N_6762);
or U8406 (N_8406,N_7517,N_6705);
or U8407 (N_8407,N_7890,N_7354);
or U8408 (N_8408,N_6649,N_7147);
or U8409 (N_8409,N_6484,N_6781);
xnor U8410 (N_8410,N_6525,N_6660);
and U8411 (N_8411,N_6615,N_7637);
and U8412 (N_8412,N_7291,N_7758);
or U8413 (N_8413,N_7221,N_7683);
and U8414 (N_8414,N_7858,N_6920);
and U8415 (N_8415,N_7537,N_7303);
nor U8416 (N_8416,N_6979,N_6800);
and U8417 (N_8417,N_7025,N_7046);
and U8418 (N_8418,N_7161,N_6453);
nor U8419 (N_8419,N_6463,N_7982);
xnor U8420 (N_8420,N_6290,N_7772);
or U8421 (N_8421,N_7574,N_7269);
and U8422 (N_8422,N_7766,N_6089);
nor U8423 (N_8423,N_6331,N_7692);
and U8424 (N_8424,N_6217,N_7934);
xnor U8425 (N_8425,N_6109,N_6405);
and U8426 (N_8426,N_7119,N_6653);
nand U8427 (N_8427,N_6393,N_6293);
or U8428 (N_8428,N_7557,N_7219);
nand U8429 (N_8429,N_6154,N_6347);
and U8430 (N_8430,N_7552,N_7018);
nand U8431 (N_8431,N_6929,N_6985);
xor U8432 (N_8432,N_7057,N_7580);
or U8433 (N_8433,N_6081,N_6704);
or U8434 (N_8434,N_6842,N_6286);
or U8435 (N_8435,N_7085,N_7963);
and U8436 (N_8436,N_7251,N_6843);
nor U8437 (N_8437,N_7417,N_6715);
nor U8438 (N_8438,N_6388,N_7373);
and U8439 (N_8439,N_6570,N_6040);
nand U8440 (N_8440,N_7819,N_6968);
and U8441 (N_8441,N_6183,N_7157);
nor U8442 (N_8442,N_7413,N_6562);
nand U8443 (N_8443,N_7530,N_6889);
nand U8444 (N_8444,N_7297,N_7306);
and U8445 (N_8445,N_6718,N_7802);
nor U8446 (N_8446,N_6277,N_6702);
nor U8447 (N_8447,N_6755,N_6103);
nor U8448 (N_8448,N_7023,N_6697);
or U8449 (N_8449,N_7048,N_6198);
and U8450 (N_8450,N_6569,N_6763);
or U8451 (N_8451,N_6515,N_7699);
nand U8452 (N_8452,N_6543,N_7469);
nand U8453 (N_8453,N_6434,N_7837);
or U8454 (N_8454,N_7884,N_7670);
nor U8455 (N_8455,N_7864,N_7861);
nor U8456 (N_8456,N_7071,N_7985);
and U8457 (N_8457,N_6732,N_6863);
or U8458 (N_8458,N_6337,N_6881);
or U8459 (N_8459,N_7229,N_6191);
and U8460 (N_8460,N_6618,N_7555);
or U8461 (N_8461,N_6773,N_7188);
nand U8462 (N_8462,N_7915,N_7214);
nor U8463 (N_8463,N_7571,N_6545);
nand U8464 (N_8464,N_6662,N_7645);
nand U8465 (N_8465,N_6547,N_7091);
and U8466 (N_8466,N_7541,N_6630);
nand U8467 (N_8467,N_6567,N_6326);
or U8468 (N_8468,N_6935,N_6158);
or U8469 (N_8469,N_6428,N_7591);
xor U8470 (N_8470,N_6854,N_7759);
nand U8471 (N_8471,N_7943,N_6946);
or U8472 (N_8472,N_7527,N_7970);
and U8473 (N_8473,N_6124,N_7049);
and U8474 (N_8474,N_7210,N_7973);
nor U8475 (N_8475,N_6077,N_6435);
or U8476 (N_8476,N_6455,N_7863);
nor U8477 (N_8477,N_6817,N_7572);
nor U8478 (N_8478,N_6226,N_6627);
nand U8479 (N_8479,N_7190,N_6300);
nand U8480 (N_8480,N_6954,N_6959);
nor U8481 (N_8481,N_6986,N_7452);
and U8482 (N_8482,N_6110,N_6883);
or U8483 (N_8483,N_7624,N_7432);
nand U8484 (N_8484,N_6436,N_7012);
nand U8485 (N_8485,N_7950,N_7405);
xnor U8486 (N_8486,N_6309,N_6788);
nor U8487 (N_8487,N_6041,N_6960);
and U8488 (N_8488,N_7729,N_6524);
nor U8489 (N_8489,N_7384,N_7450);
nor U8490 (N_8490,N_7499,N_6175);
and U8491 (N_8491,N_7039,N_6228);
and U8492 (N_8492,N_7643,N_7548);
nand U8493 (N_8493,N_7164,N_6894);
nand U8494 (N_8494,N_6020,N_6391);
and U8495 (N_8495,N_7466,N_7101);
nand U8496 (N_8496,N_6144,N_6372);
nand U8497 (N_8497,N_6468,N_7850);
nand U8498 (N_8498,N_7907,N_7845);
nor U8499 (N_8499,N_7800,N_6500);
or U8500 (N_8500,N_7786,N_7939);
and U8501 (N_8501,N_7298,N_7809);
or U8502 (N_8502,N_7976,N_7453);
or U8503 (N_8503,N_7480,N_6777);
nand U8504 (N_8504,N_7732,N_7812);
or U8505 (N_8505,N_6053,N_7887);
or U8506 (N_8506,N_7828,N_6585);
nor U8507 (N_8507,N_6418,N_7997);
and U8508 (N_8508,N_6368,N_6119);
and U8509 (N_8509,N_6526,N_7634);
nand U8510 (N_8510,N_6113,N_7075);
nand U8511 (N_8511,N_6384,N_6305);
nor U8512 (N_8512,N_7936,N_7767);
nor U8513 (N_8513,N_7697,N_6831);
xnor U8514 (N_8514,N_7892,N_6734);
xnor U8515 (N_8515,N_6138,N_6708);
xor U8516 (N_8516,N_6027,N_7757);
nand U8517 (N_8517,N_7187,N_6112);
or U8518 (N_8518,N_7604,N_6556);
xnor U8519 (N_8519,N_7145,N_7050);
xor U8520 (N_8520,N_7092,N_6251);
nand U8521 (N_8521,N_7108,N_7033);
or U8522 (N_8522,N_7867,N_6055);
nand U8523 (N_8523,N_7171,N_7415);
or U8524 (N_8524,N_6380,N_7441);
nand U8525 (N_8525,N_6481,N_6431);
and U8526 (N_8526,N_6030,N_6056);
or U8527 (N_8527,N_6011,N_6098);
nor U8528 (N_8528,N_6263,N_7533);
nand U8529 (N_8529,N_6039,N_6255);
and U8530 (N_8530,N_6769,N_7599);
and U8531 (N_8531,N_6404,N_6247);
xnor U8532 (N_8532,N_7693,N_7605);
xor U8533 (N_8533,N_6023,N_7130);
nand U8534 (N_8534,N_7894,N_6383);
nand U8535 (N_8535,N_6984,N_7483);
or U8536 (N_8536,N_6942,N_7679);
nand U8537 (N_8537,N_7512,N_7224);
or U8538 (N_8538,N_6657,N_7100);
nor U8539 (N_8539,N_7656,N_7718);
or U8540 (N_8540,N_6047,N_7929);
and U8541 (N_8541,N_7140,N_7068);
or U8542 (N_8542,N_7160,N_6536);
nand U8543 (N_8543,N_7678,N_6698);
nor U8544 (N_8544,N_6160,N_6890);
and U8545 (N_8545,N_6796,N_6861);
xor U8546 (N_8546,N_7761,N_7993);
nand U8547 (N_8547,N_7244,N_6483);
and U8548 (N_8548,N_7668,N_6220);
nand U8549 (N_8549,N_7926,N_6970);
or U8550 (N_8550,N_6928,N_6737);
nand U8551 (N_8551,N_7455,N_6676);
and U8552 (N_8552,N_7520,N_7125);
nand U8553 (N_8553,N_7895,N_6032);
and U8554 (N_8554,N_7444,N_6474);
nand U8555 (N_8555,N_7379,N_6953);
nand U8556 (N_8556,N_6078,N_6306);
nor U8557 (N_8557,N_7981,N_6403);
and U8558 (N_8558,N_6882,N_6866);
or U8559 (N_8559,N_6190,N_7286);
nor U8560 (N_8560,N_7113,N_6916);
and U8561 (N_8561,N_7782,N_6167);
nand U8562 (N_8562,N_7974,N_6892);
or U8563 (N_8563,N_7565,N_7521);
or U8564 (N_8564,N_6441,N_7293);
nand U8565 (N_8565,N_7319,N_7471);
or U8566 (N_8566,N_7785,N_7154);
nand U8567 (N_8567,N_6264,N_7315);
nor U8568 (N_8568,N_6602,N_6605);
or U8569 (N_8569,N_7913,N_6555);
or U8570 (N_8570,N_6516,N_6461);
xor U8571 (N_8571,N_7106,N_6118);
or U8572 (N_8572,N_7629,N_7608);
nor U8573 (N_8573,N_6371,N_7908);
and U8574 (N_8574,N_6687,N_6370);
xor U8575 (N_8575,N_6146,N_7538);
nand U8576 (N_8576,N_7281,N_7382);
or U8577 (N_8577,N_7610,N_6153);
or U8578 (N_8578,N_7647,N_6432);
and U8579 (N_8579,N_6123,N_6829);
nor U8580 (N_8580,N_7268,N_6661);
nand U8581 (N_8581,N_7394,N_6975);
nand U8582 (N_8582,N_7614,N_6988);
and U8583 (N_8583,N_6991,N_7651);
or U8584 (N_8584,N_7222,N_7001);
nor U8585 (N_8585,N_7642,N_6375);
nor U8586 (N_8586,N_7305,N_6634);
xnor U8587 (N_8587,N_6091,N_6332);
xnor U8588 (N_8588,N_6215,N_7418);
nor U8589 (N_8589,N_7852,N_6390);
xnor U8590 (N_8590,N_7118,N_6225);
nor U8591 (N_8591,N_6143,N_6580);
and U8592 (N_8592,N_6493,N_7746);
and U8593 (N_8593,N_7723,N_6706);
nor U8594 (N_8594,N_6871,N_7295);
or U8595 (N_8595,N_6887,N_7603);
xnor U8596 (N_8596,N_7635,N_7260);
or U8597 (N_8597,N_6421,N_6996);
nand U8598 (N_8598,N_6643,N_7325);
nor U8599 (N_8599,N_6284,N_7720);
nand U8600 (N_8600,N_7139,N_6797);
nor U8601 (N_8601,N_7277,N_7403);
nand U8602 (N_8602,N_6776,N_6622);
nand U8603 (N_8603,N_6096,N_7328);
xnor U8604 (N_8604,N_7270,N_6137);
and U8605 (N_8605,N_6964,N_7408);
and U8606 (N_8606,N_6285,N_7285);
nand U8607 (N_8607,N_6410,N_6805);
or U8608 (N_8608,N_7141,N_6270);
or U8609 (N_8609,N_7667,N_7485);
or U8610 (N_8610,N_7702,N_6002);
or U8611 (N_8611,N_7942,N_7330);
and U8612 (N_8612,N_7060,N_6836);
nor U8613 (N_8613,N_7626,N_7769);
nand U8614 (N_8614,N_6941,N_7117);
or U8615 (N_8615,N_6176,N_7339);
or U8616 (N_8616,N_7189,N_7180);
xor U8617 (N_8617,N_6820,N_6406);
nor U8618 (N_8618,N_7813,N_7094);
nor U8619 (N_8619,N_6885,N_7562);
or U8620 (N_8620,N_6414,N_7393);
nand U8621 (N_8621,N_7349,N_6348);
xor U8622 (N_8622,N_6357,N_7743);
nor U8623 (N_8623,N_6899,N_7103);
nor U8624 (N_8624,N_7209,N_6912);
xnor U8625 (N_8625,N_7685,N_7317);
nand U8626 (N_8626,N_6412,N_7381);
nand U8627 (N_8627,N_6321,N_6819);
or U8628 (N_8628,N_6312,N_7531);
nor U8629 (N_8629,N_6007,N_6655);
nand U8630 (N_8630,N_6963,N_7904);
nor U8631 (N_8631,N_7721,N_7606);
xor U8632 (N_8632,N_6288,N_7949);
and U8633 (N_8633,N_6488,N_6448);
nor U8634 (N_8634,N_7672,N_7027);
nor U8635 (N_8635,N_7074,N_7036);
or U8636 (N_8636,N_7633,N_6679);
or U8637 (N_8637,N_6950,N_7927);
nand U8638 (N_8638,N_6768,N_6947);
and U8639 (N_8639,N_6221,N_7359);
xor U8640 (N_8640,N_7988,N_7459);
nand U8641 (N_8641,N_6273,N_6711);
and U8642 (N_8642,N_7404,N_7290);
nand U8643 (N_8643,N_6980,N_7751);
nor U8644 (N_8644,N_7829,N_7069);
or U8645 (N_8645,N_7991,N_7227);
nor U8646 (N_8646,N_7423,N_7694);
or U8647 (N_8647,N_7392,N_7414);
or U8648 (N_8648,N_6553,N_7962);
nand U8649 (N_8649,N_7194,N_6712);
nor U8650 (N_8650,N_6786,N_6012);
and U8651 (N_8651,N_7834,N_6564);
xor U8652 (N_8652,N_7688,N_7428);
nand U8653 (N_8653,N_6561,N_6005);
nor U8654 (N_8654,N_6740,N_7650);
xor U8655 (N_8655,N_6586,N_7859);
and U8656 (N_8656,N_7374,N_7919);
nor U8657 (N_8657,N_6342,N_7882);
and U8658 (N_8658,N_6771,N_6345);
or U8659 (N_8659,N_6798,N_7503);
or U8660 (N_8660,N_6133,N_7484);
and U8661 (N_8661,N_6498,N_7661);
or U8662 (N_8662,N_6523,N_6502);
nor U8663 (N_8663,N_7364,N_6202);
xor U8664 (N_8664,N_6458,N_6851);
nor U8665 (N_8665,N_6652,N_6785);
and U8666 (N_8666,N_6178,N_6062);
and U8667 (N_8667,N_7838,N_6940);
nand U8668 (N_8668,N_7522,N_7594);
nor U8669 (N_8669,N_6140,N_6054);
or U8670 (N_8670,N_6398,N_7166);
xor U8671 (N_8671,N_7595,N_7922);
or U8672 (N_8672,N_6908,N_6476);
nor U8673 (N_8673,N_6911,N_7880);
or U8674 (N_8674,N_6571,N_6692);
nand U8675 (N_8675,N_6196,N_7360);
or U8676 (N_8676,N_6382,N_6799);
or U8677 (N_8677,N_7708,N_6709);
and U8678 (N_8678,N_6210,N_6227);
and U8679 (N_8679,N_6141,N_7646);
or U8680 (N_8680,N_7549,N_6052);
nand U8681 (N_8681,N_7747,N_6967);
nand U8682 (N_8682,N_7040,N_7228);
nand U8683 (N_8683,N_7429,N_6787);
or U8684 (N_8684,N_7073,N_6246);
nand U8685 (N_8685,N_7539,N_7396);
nor U8686 (N_8686,N_7111,N_7585);
xor U8687 (N_8687,N_6998,N_7570);
nand U8688 (N_8688,N_7051,N_6607);
or U8689 (N_8689,N_6633,N_7989);
xor U8690 (N_8690,N_6278,N_6606);
nor U8691 (N_8691,N_6466,N_7369);
xnor U8692 (N_8692,N_7724,N_6186);
nand U8693 (N_8693,N_7427,N_6224);
nor U8694 (N_8694,N_6045,N_6344);
nor U8695 (N_8695,N_7288,N_6063);
nand U8696 (N_8696,N_7436,N_6780);
or U8697 (N_8697,N_6313,N_6620);
nor U8698 (N_8698,N_6296,N_6886);
nor U8699 (N_8699,N_6433,N_7207);
nor U8700 (N_8700,N_7841,N_6982);
nor U8701 (N_8701,N_6291,N_6320);
and U8702 (N_8702,N_6295,N_6339);
nor U8703 (N_8703,N_7220,N_7842);
nor U8704 (N_8704,N_7280,N_6018);
nand U8705 (N_8705,N_7739,N_7438);
nor U8706 (N_8706,N_7575,N_6497);
nor U8707 (N_8707,N_7361,N_6073);
xor U8708 (N_8708,N_6485,N_6025);
nor U8709 (N_8709,N_6189,N_6647);
and U8710 (N_8710,N_7474,N_6280);
xor U8711 (N_8711,N_7233,N_7276);
nand U8712 (N_8712,N_7267,N_6621);
and U8713 (N_8713,N_7611,N_7587);
or U8714 (N_8714,N_7493,N_6730);
nor U8715 (N_8715,N_6205,N_6033);
and U8716 (N_8716,N_7163,N_7449);
or U8717 (N_8717,N_6245,N_7217);
nand U8718 (N_8718,N_6919,N_6392);
xor U8719 (N_8719,N_7835,N_7078);
and U8720 (N_8720,N_6128,N_7705);
nand U8721 (N_8721,N_7972,N_7931);
nand U8722 (N_8722,N_7133,N_7897);
nand U8723 (N_8723,N_7847,N_6951);
or U8724 (N_8724,N_6407,N_6214);
and U8725 (N_8725,N_6589,N_6859);
or U8726 (N_8726,N_7701,N_6487);
and U8727 (N_8727,N_7526,N_7719);
or U8728 (N_8728,N_6646,N_7874);
nor U8729 (N_8729,N_7131,N_7826);
or U8730 (N_8730,N_6577,N_7978);
nor U8731 (N_8731,N_7818,N_6645);
xnor U8732 (N_8732,N_6034,N_6648);
or U8733 (N_8733,N_7242,N_6664);
nor U8734 (N_8734,N_6130,N_6301);
or U8735 (N_8735,N_7308,N_7435);
nand U8736 (N_8736,N_7365,N_7803);
nor U8737 (N_8737,N_6813,N_7185);
nand U8738 (N_8738,N_7081,N_7937);
or U8739 (N_8739,N_7649,N_6917);
or U8740 (N_8740,N_6444,N_7876);
xnor U8741 (N_8741,N_6736,N_6510);
and U8742 (N_8742,N_6877,N_6934);
nor U8743 (N_8743,N_6809,N_6703);
nor U8744 (N_8744,N_7266,N_7559);
xnor U8745 (N_8745,N_6644,N_7356);
nor U8746 (N_8746,N_6480,N_6575);
or U8747 (N_8747,N_7508,N_6360);
and U8748 (N_8748,N_7105,N_7442);
and U8749 (N_8749,N_6223,N_7848);
and U8750 (N_8750,N_7265,N_6921);
nor U8751 (N_8751,N_7561,N_7148);
nor U8752 (N_8752,N_7817,N_6583);
nor U8753 (N_8753,N_7764,N_7475);
or U8754 (N_8754,N_7513,N_7443);
or U8755 (N_8755,N_6351,N_6559);
and U8756 (N_8756,N_6201,N_7083);
nand U8757 (N_8757,N_6955,N_6508);
or U8758 (N_8758,N_6868,N_7566);
nor U8759 (N_8759,N_7660,N_6923);
xor U8760 (N_8760,N_7274,N_6669);
and U8761 (N_8761,N_6636,N_6231);
or U8762 (N_8762,N_6903,N_7342);
nand U8763 (N_8763,N_6213,N_7968);
or U8764 (N_8764,N_7167,N_7711);
nand U8765 (N_8765,N_7491,N_6879);
or U8766 (N_8766,N_6538,N_7567);
and U8767 (N_8767,N_7917,N_6976);
or U8768 (N_8768,N_6208,N_7625);
or U8769 (N_8769,N_6683,N_7681);
and U8770 (N_8770,N_6180,N_6161);
xor U8771 (N_8771,N_6352,N_6517);
xor U8772 (N_8772,N_7830,N_7733);
and U8773 (N_8773,N_7335,N_7345);
nand U8774 (N_8774,N_7395,N_7225);
nor U8775 (N_8775,N_6456,N_6965);
xor U8776 (N_8776,N_6961,N_7518);
or U8777 (N_8777,N_7658,N_7146);
nor U8778 (N_8778,N_7969,N_6720);
or U8779 (N_8779,N_7825,N_7690);
or U8780 (N_8780,N_7657,N_7741);
xnor U8781 (N_8781,N_7655,N_6554);
and U8782 (N_8782,N_6361,N_7351);
and U8783 (N_8783,N_6486,N_6304);
nor U8784 (N_8784,N_7713,N_6741);
nand U8785 (N_8785,N_7695,N_6268);
xnor U8786 (N_8786,N_7680,N_6844);
nor U8787 (N_8787,N_6185,N_6415);
or U8788 (N_8788,N_6752,N_7584);
and U8789 (N_8789,N_6671,N_7738);
xor U8790 (N_8790,N_7446,N_6359);
and U8791 (N_8791,N_6638,N_7059);
nor U8792 (N_8792,N_7763,N_7173);
nand U8793 (N_8793,N_7135,N_6822);
nand U8794 (N_8794,N_6139,N_6507);
nand U8795 (N_8795,N_6654,N_6658);
nor U8796 (N_8796,N_6722,N_6994);
xor U8797 (N_8797,N_6298,N_6329);
nand U8798 (N_8798,N_6145,N_6816);
nor U8799 (N_8799,N_7795,N_7960);
or U8800 (N_8800,N_6219,N_6590);
or U8801 (N_8801,N_6462,N_6587);
xnor U8802 (N_8802,N_7321,N_6846);
xor U8803 (N_8803,N_6557,N_6000);
nand U8804 (N_8804,N_6075,N_6707);
and U8805 (N_8805,N_7064,N_7755);
xnor U8806 (N_8806,N_6494,N_6748);
nand U8807 (N_8807,N_7067,N_6058);
and U8808 (N_8808,N_6460,N_7124);
and U8809 (N_8809,N_6402,N_7477);
nand U8810 (N_8810,N_7836,N_6422);
nand U8811 (N_8811,N_6710,N_7377);
and U8812 (N_8812,N_7956,N_7329);
nand U8813 (N_8813,N_7789,N_7322);
nor U8814 (N_8814,N_7958,N_6663);
nand U8815 (N_8815,N_6673,N_6420);
nor U8816 (N_8816,N_7620,N_6491);
nand U8817 (N_8817,N_6541,N_7914);
or U8818 (N_8818,N_6753,N_6084);
nand U8819 (N_8819,N_6693,N_6240);
nand U8820 (N_8820,N_7350,N_7151);
xnor U8821 (N_8821,N_7126,N_6129);
or U8822 (N_8822,N_6865,N_7622);
and U8823 (N_8823,N_7717,N_6323);
nor U8824 (N_8824,N_6913,N_6639);
nor U8825 (N_8825,N_6742,N_6004);
nor U8826 (N_8826,N_6608,N_6783);
nor U8827 (N_8827,N_7318,N_6087);
and U8828 (N_8828,N_7510,N_7226);
nor U8829 (N_8829,N_6597,N_7337);
xnor U8830 (N_8830,N_6200,N_7497);
and U8831 (N_8831,N_6386,N_6572);
and U8832 (N_8832,N_6514,N_6206);
or U8833 (N_8833,N_6179,N_7201);
nor U8834 (N_8834,N_6812,N_7198);
and U8835 (N_8835,N_7026,N_7487);
and U8836 (N_8836,N_6993,N_7607);
and U8837 (N_8837,N_6839,N_7338);
nand U8838 (N_8838,N_7257,N_6651);
or U8839 (N_8839,N_6699,N_7422);
or U8840 (N_8840,N_6409,N_6759);
and U8841 (N_8841,N_7957,N_6578);
nor U8842 (N_8842,N_7248,N_7102);
or U8843 (N_8843,N_6999,N_7042);
nor U8844 (N_8844,N_7362,N_7121);
xnor U8845 (N_8845,N_6849,N_6356);
or U8846 (N_8846,N_7302,N_7421);
nand U8847 (N_8847,N_6100,N_6530);
or U8848 (N_8848,N_6490,N_6471);
nand U8849 (N_8849,N_6394,N_7951);
nor U8850 (N_8850,N_6802,N_6467);
or U8851 (N_8851,N_6674,N_6036);
and U8852 (N_8852,N_7689,N_7357);
or U8853 (N_8853,N_7087,N_6122);
or U8854 (N_8854,N_7324,N_6008);
and U8855 (N_8855,N_6271,N_7238);
or U8856 (N_8856,N_7805,N_7628);
or U8857 (N_8857,N_7756,N_7388);
nand U8858 (N_8858,N_7013,N_6151);
and U8859 (N_8859,N_7005,N_6341);
and U8860 (N_8860,N_6437,N_6591);
nor U8861 (N_8861,N_6340,N_7909);
or U8862 (N_8862,N_7686,N_6535);
and U8863 (N_8863,N_6914,N_6527);
xor U8864 (N_8864,N_7400,N_6157);
nor U8865 (N_8865,N_6548,N_7532);
or U8866 (N_8866,N_6827,N_7583);
nor U8867 (N_8867,N_6847,N_7844);
nand U8868 (N_8868,N_7460,N_6746);
nand U8869 (N_8869,N_7262,N_6860);
nor U8870 (N_8870,N_6937,N_6811);
nand U8871 (N_8871,N_7524,N_6043);
nand U8872 (N_8872,N_7211,N_7851);
or U8873 (N_8873,N_6511,N_7862);
or U8874 (N_8874,N_6355,N_7464);
and U8875 (N_8875,N_6450,N_6478);
and U8876 (N_8876,N_7714,N_7687);
or U8877 (N_8877,N_7196,N_6197);
or U8878 (N_8878,N_7070,N_7990);
nor U8879 (N_8879,N_6659,N_7494);
or U8880 (N_8880,N_6148,N_6330);
and U8881 (N_8881,N_7123,N_7150);
and U8882 (N_8882,N_6850,N_7273);
xor U8883 (N_8883,N_6962,N_6981);
or U8884 (N_8884,N_7804,N_6902);
or U8885 (N_8885,N_6974,N_7612);
nand U8886 (N_8886,N_6691,N_6893);
or U8887 (N_8887,N_7099,N_7808);
nand U8888 (N_8888,N_6346,N_6656);
nand U8889 (N_8889,N_7995,N_7158);
nand U8890 (N_8890,N_6745,N_6726);
and U8891 (N_8891,N_7031,N_7792);
nor U8892 (N_8892,N_6165,N_7977);
or U8893 (N_8893,N_7855,N_6724);
and U8894 (N_8894,N_7577,N_7076);
and U8895 (N_8895,N_7663,N_7372);
and U8896 (N_8896,N_6014,N_6880);
nand U8897 (N_8897,N_6884,N_7778);
and U8898 (N_8898,N_6001,N_7172);
and U8899 (N_8899,N_7402,N_7773);
nand U8900 (N_8900,N_6446,N_7986);
or U8901 (N_8901,N_7234,N_7175);
nand U8902 (N_8902,N_7472,N_7193);
and U8903 (N_8903,N_7401,N_6248);
or U8904 (N_8904,N_7691,N_7055);
nand U8905 (N_8905,N_6828,N_6611);
nand U8906 (N_8906,N_6867,N_6116);
nor U8907 (N_8907,N_6791,N_7208);
and U8908 (N_8908,N_7998,N_6328);
nand U8909 (N_8909,N_7777,N_7621);
nand U8910 (N_8910,N_7545,N_6833);
nor U8911 (N_8911,N_7311,N_6767);
or U8912 (N_8912,N_7341,N_6924);
and U8913 (N_8913,N_6068,N_7506);
nand U8914 (N_8914,N_6451,N_6806);
nand U8915 (N_8915,N_7399,N_7967);
nor U8916 (N_8916,N_6613,N_7376);
and U8917 (N_8917,N_7409,N_6233);
or U8918 (N_8918,N_6374,N_7925);
nand U8919 (N_8919,N_7110,N_6694);
and U8920 (N_8920,N_6314,N_6576);
and U8921 (N_8921,N_7765,N_6400);
nor U8922 (N_8922,N_6808,N_7737);
nor U8923 (N_8923,N_7519,N_7461);
and U8924 (N_8924,N_7662,N_7132);
and U8925 (N_8925,N_6181,N_6931);
xor U8926 (N_8926,N_6426,N_6395);
nand U8927 (N_8927,N_7006,N_6957);
and U8928 (N_8928,N_7547,N_6573);
xor U8929 (N_8929,N_6600,N_7684);
nor U8930 (N_8930,N_6789,N_6896);
nor U8931 (N_8931,N_7948,N_7243);
or U8932 (N_8932,N_7727,N_7363);
and U8933 (N_8933,N_7774,N_7259);
nand U8934 (N_8934,N_7024,N_7788);
xor U8935 (N_8935,N_6501,N_6592);
nor U8936 (N_8936,N_6626,N_6092);
or U8937 (N_8937,N_6610,N_7002);
and U8938 (N_8938,N_6835,N_7186);
nor U8939 (N_8939,N_6574,N_7287);
nor U8940 (N_8940,N_6826,N_6793);
nor U8941 (N_8941,N_6496,N_7952);
nand U8942 (N_8942,N_7456,N_7272);
nor U8943 (N_8943,N_7231,N_7558);
and U8944 (N_8944,N_7501,N_7448);
or U8945 (N_8945,N_6072,N_6234);
and U8946 (N_8946,N_6325,N_7898);
nor U8947 (N_8947,N_7034,N_7796);
or U8948 (N_8948,N_7853,N_7784);
nor U8949 (N_8949,N_6628,N_7516);
xnor U8950 (N_8950,N_7213,N_6059);
nor U8951 (N_8951,N_6132,N_6853);
nor U8952 (N_8952,N_7463,N_6195);
xnor U8953 (N_8953,N_7930,N_6522);
xor U8954 (N_8954,N_7824,N_7502);
and U8955 (N_8955,N_6170,N_7470);
nand U8956 (N_8956,N_7644,N_6281);
nand U8957 (N_8957,N_7536,N_6275);
and U8958 (N_8958,N_6259,N_7326);
nor U8959 (N_8959,N_7906,N_7279);
or U8960 (N_8960,N_7735,N_7371);
xnor U8961 (N_8961,N_6364,N_7206);
or U8962 (N_8962,N_6429,N_7966);
nand U8963 (N_8963,N_6150,N_6335);
and U8964 (N_8964,N_6192,N_6438);
or U8965 (N_8965,N_7749,N_6216);
xnor U8966 (N_8966,N_7411,N_7216);
and U8967 (N_8967,N_6533,N_7869);
or U8968 (N_8968,N_7090,N_6499);
nand U8969 (N_8969,N_7947,N_7153);
nand U8970 (N_8970,N_6211,N_7300);
nor U8971 (N_8971,N_7454,N_6821);
or U8972 (N_8972,N_6442,N_6625);
xnor U8973 (N_8973,N_7177,N_6936);
or U8974 (N_8974,N_6254,N_6733);
nor U8975 (N_8975,N_7965,N_7781);
and U8976 (N_8976,N_6028,N_7195);
nand U8977 (N_8977,N_6990,N_7021);
nor U8978 (N_8978,N_6520,N_6770);
or U8979 (N_8979,N_6728,N_6035);
nor U8980 (N_8980,N_7740,N_6469);
nor U8981 (N_8981,N_6845,N_7959);
and U8982 (N_8982,N_7793,N_7938);
or U8983 (N_8983,N_7631,N_6239);
nand U8984 (N_8984,N_7203,N_7058);
nand U8985 (N_8985,N_7866,N_7505);
or U8986 (N_8986,N_7044,N_6322);
nor U8987 (N_8987,N_7868,N_6258);
and U8988 (N_8988,N_7523,N_6539);
and U8989 (N_8989,N_6492,N_7355);
nor U8990 (N_8990,N_7556,N_7129);
or U8991 (N_8991,N_7437,N_6978);
or U8992 (N_8992,N_6475,N_6204);
and U8993 (N_8993,N_7346,N_7072);
or U8994 (N_8994,N_6272,N_7589);
nand U8995 (N_8995,N_7467,N_7762);
or U8996 (N_8996,N_7162,N_7768);
nand U8997 (N_8997,N_6876,N_6147);
xnor U8998 (N_8998,N_6253,N_7292);
nor U8999 (N_8999,N_6425,N_7779);
nand U9000 (N_9000,N_7765,N_7841);
nand U9001 (N_9001,N_6963,N_7209);
and U9002 (N_9002,N_6096,N_6206);
xnor U9003 (N_9003,N_7660,N_7570);
nand U9004 (N_9004,N_6082,N_6660);
xor U9005 (N_9005,N_6250,N_6800);
nand U9006 (N_9006,N_7116,N_6345);
nor U9007 (N_9007,N_7570,N_6989);
nand U9008 (N_9008,N_6193,N_6379);
nand U9009 (N_9009,N_6573,N_6804);
xnor U9010 (N_9010,N_7647,N_7602);
nor U9011 (N_9011,N_6255,N_7610);
and U9012 (N_9012,N_7476,N_7893);
xor U9013 (N_9013,N_7585,N_6790);
or U9014 (N_9014,N_7118,N_7197);
nor U9015 (N_9015,N_6780,N_7354);
or U9016 (N_9016,N_7853,N_7794);
or U9017 (N_9017,N_7372,N_7340);
nand U9018 (N_9018,N_7097,N_6517);
xnor U9019 (N_9019,N_6957,N_7283);
nor U9020 (N_9020,N_7723,N_7851);
nand U9021 (N_9021,N_6831,N_6151);
nor U9022 (N_9022,N_6212,N_7539);
or U9023 (N_9023,N_6955,N_6768);
xnor U9024 (N_9024,N_6606,N_7126);
and U9025 (N_9025,N_7029,N_6190);
and U9026 (N_9026,N_6041,N_6889);
nor U9027 (N_9027,N_6215,N_7250);
or U9028 (N_9028,N_6375,N_7054);
xnor U9029 (N_9029,N_7462,N_6738);
and U9030 (N_9030,N_6717,N_7287);
or U9031 (N_9031,N_7975,N_6187);
nor U9032 (N_9032,N_6365,N_7264);
and U9033 (N_9033,N_7634,N_6904);
and U9034 (N_9034,N_6515,N_7916);
and U9035 (N_9035,N_6317,N_7181);
nor U9036 (N_9036,N_7595,N_6877);
nand U9037 (N_9037,N_7331,N_6378);
nand U9038 (N_9038,N_6332,N_7269);
nand U9039 (N_9039,N_6583,N_6975);
nand U9040 (N_9040,N_7598,N_6087);
and U9041 (N_9041,N_7809,N_7581);
and U9042 (N_9042,N_6952,N_7667);
and U9043 (N_9043,N_7131,N_7103);
nand U9044 (N_9044,N_7301,N_7453);
or U9045 (N_9045,N_6354,N_6375);
nand U9046 (N_9046,N_6812,N_6314);
or U9047 (N_9047,N_6677,N_7825);
or U9048 (N_9048,N_6525,N_7765);
and U9049 (N_9049,N_6234,N_6297);
or U9050 (N_9050,N_7099,N_6792);
nand U9051 (N_9051,N_6415,N_7952);
and U9052 (N_9052,N_6707,N_6514);
xnor U9053 (N_9053,N_7784,N_7513);
nor U9054 (N_9054,N_6211,N_7340);
or U9055 (N_9055,N_7725,N_7700);
and U9056 (N_9056,N_6747,N_7387);
or U9057 (N_9057,N_7829,N_6319);
and U9058 (N_9058,N_6474,N_7144);
nor U9059 (N_9059,N_7089,N_6020);
or U9060 (N_9060,N_7943,N_6327);
or U9061 (N_9061,N_6269,N_7587);
or U9062 (N_9062,N_6055,N_6538);
and U9063 (N_9063,N_6196,N_7856);
nor U9064 (N_9064,N_7830,N_6704);
or U9065 (N_9065,N_6990,N_7659);
and U9066 (N_9066,N_7741,N_7494);
nor U9067 (N_9067,N_7594,N_6889);
nor U9068 (N_9068,N_7388,N_6237);
and U9069 (N_9069,N_6002,N_6868);
nand U9070 (N_9070,N_6815,N_6044);
nand U9071 (N_9071,N_7105,N_6553);
nor U9072 (N_9072,N_6059,N_6643);
or U9073 (N_9073,N_6773,N_7860);
nor U9074 (N_9074,N_6117,N_7987);
nand U9075 (N_9075,N_6881,N_7245);
nand U9076 (N_9076,N_6375,N_7301);
and U9077 (N_9077,N_7456,N_6432);
and U9078 (N_9078,N_6848,N_6415);
nor U9079 (N_9079,N_6252,N_6304);
nor U9080 (N_9080,N_6208,N_6258);
nor U9081 (N_9081,N_7019,N_6480);
nand U9082 (N_9082,N_6433,N_6136);
nor U9083 (N_9083,N_6082,N_6031);
or U9084 (N_9084,N_6819,N_7933);
or U9085 (N_9085,N_6732,N_7490);
nand U9086 (N_9086,N_6340,N_6100);
nand U9087 (N_9087,N_6942,N_6507);
and U9088 (N_9088,N_6773,N_7896);
nand U9089 (N_9089,N_7349,N_6206);
nand U9090 (N_9090,N_7171,N_6169);
or U9091 (N_9091,N_6507,N_6251);
xnor U9092 (N_9092,N_7122,N_7562);
nand U9093 (N_9093,N_6000,N_7038);
and U9094 (N_9094,N_7516,N_7043);
and U9095 (N_9095,N_6506,N_7336);
nor U9096 (N_9096,N_7241,N_6398);
or U9097 (N_9097,N_6737,N_7114);
nor U9098 (N_9098,N_7568,N_7610);
or U9099 (N_9099,N_7523,N_6024);
nand U9100 (N_9100,N_6151,N_6113);
or U9101 (N_9101,N_6657,N_6468);
or U9102 (N_9102,N_7871,N_7578);
nor U9103 (N_9103,N_6860,N_6889);
nor U9104 (N_9104,N_7208,N_7073);
xnor U9105 (N_9105,N_7990,N_7736);
and U9106 (N_9106,N_6429,N_6913);
or U9107 (N_9107,N_6974,N_7231);
nor U9108 (N_9108,N_6912,N_6553);
nor U9109 (N_9109,N_7256,N_6217);
and U9110 (N_9110,N_7788,N_7553);
nor U9111 (N_9111,N_7727,N_6912);
nand U9112 (N_9112,N_7649,N_6446);
or U9113 (N_9113,N_7560,N_6684);
nor U9114 (N_9114,N_7118,N_7313);
nand U9115 (N_9115,N_6445,N_6390);
or U9116 (N_9116,N_6951,N_7886);
nor U9117 (N_9117,N_6966,N_6596);
and U9118 (N_9118,N_6733,N_7303);
nor U9119 (N_9119,N_7687,N_6518);
and U9120 (N_9120,N_6694,N_6517);
nor U9121 (N_9121,N_6913,N_7485);
and U9122 (N_9122,N_6121,N_7780);
nor U9123 (N_9123,N_6682,N_7702);
and U9124 (N_9124,N_7124,N_7817);
and U9125 (N_9125,N_6396,N_6854);
or U9126 (N_9126,N_7527,N_6819);
and U9127 (N_9127,N_6275,N_7584);
nand U9128 (N_9128,N_7914,N_7415);
nor U9129 (N_9129,N_6528,N_7742);
xor U9130 (N_9130,N_7350,N_6833);
nand U9131 (N_9131,N_6080,N_6999);
and U9132 (N_9132,N_6297,N_6609);
nand U9133 (N_9133,N_6327,N_6286);
or U9134 (N_9134,N_6158,N_7065);
nor U9135 (N_9135,N_7921,N_7578);
and U9136 (N_9136,N_6890,N_6342);
xnor U9137 (N_9137,N_6714,N_6055);
nand U9138 (N_9138,N_7388,N_6447);
xor U9139 (N_9139,N_7629,N_7286);
and U9140 (N_9140,N_6613,N_7131);
nor U9141 (N_9141,N_7254,N_6978);
and U9142 (N_9142,N_7329,N_7463);
or U9143 (N_9143,N_7990,N_6798);
xor U9144 (N_9144,N_6007,N_7160);
and U9145 (N_9145,N_7199,N_7126);
or U9146 (N_9146,N_7019,N_7327);
nor U9147 (N_9147,N_6200,N_6761);
and U9148 (N_9148,N_7784,N_7277);
and U9149 (N_9149,N_6363,N_6596);
nor U9150 (N_9150,N_7085,N_6043);
or U9151 (N_9151,N_6699,N_7661);
or U9152 (N_9152,N_6570,N_7721);
nand U9153 (N_9153,N_6182,N_6657);
or U9154 (N_9154,N_6243,N_7760);
xnor U9155 (N_9155,N_6226,N_6756);
xor U9156 (N_9156,N_6803,N_7819);
nand U9157 (N_9157,N_7089,N_6524);
or U9158 (N_9158,N_6256,N_6749);
nor U9159 (N_9159,N_7051,N_6534);
or U9160 (N_9160,N_7831,N_6058);
and U9161 (N_9161,N_6196,N_7167);
or U9162 (N_9162,N_7239,N_6237);
xnor U9163 (N_9163,N_6374,N_6603);
or U9164 (N_9164,N_6417,N_6091);
or U9165 (N_9165,N_7873,N_7950);
nand U9166 (N_9166,N_6410,N_7387);
nand U9167 (N_9167,N_6329,N_7828);
nor U9168 (N_9168,N_6292,N_7962);
nand U9169 (N_9169,N_7381,N_6799);
and U9170 (N_9170,N_7560,N_7216);
nand U9171 (N_9171,N_7783,N_7556);
and U9172 (N_9172,N_7563,N_6643);
nand U9173 (N_9173,N_7688,N_7355);
or U9174 (N_9174,N_6386,N_6901);
or U9175 (N_9175,N_7495,N_7078);
or U9176 (N_9176,N_7212,N_7885);
nor U9177 (N_9177,N_7870,N_7627);
nand U9178 (N_9178,N_6902,N_7589);
nand U9179 (N_9179,N_6419,N_7127);
and U9180 (N_9180,N_7422,N_7491);
nand U9181 (N_9181,N_6437,N_7694);
or U9182 (N_9182,N_7177,N_7306);
or U9183 (N_9183,N_6915,N_6679);
nor U9184 (N_9184,N_7881,N_6008);
and U9185 (N_9185,N_6762,N_7637);
and U9186 (N_9186,N_7653,N_7899);
and U9187 (N_9187,N_6649,N_6066);
or U9188 (N_9188,N_6524,N_7863);
nand U9189 (N_9189,N_7356,N_7620);
and U9190 (N_9190,N_7002,N_6492);
nand U9191 (N_9191,N_6013,N_7598);
or U9192 (N_9192,N_7767,N_7406);
or U9193 (N_9193,N_6677,N_7644);
or U9194 (N_9194,N_7754,N_6634);
nor U9195 (N_9195,N_7229,N_6026);
and U9196 (N_9196,N_6937,N_6993);
nand U9197 (N_9197,N_7639,N_7120);
or U9198 (N_9198,N_7185,N_7420);
nand U9199 (N_9199,N_6161,N_7867);
nand U9200 (N_9200,N_6665,N_7761);
xnor U9201 (N_9201,N_6052,N_6413);
nor U9202 (N_9202,N_6677,N_6627);
and U9203 (N_9203,N_6674,N_7013);
nor U9204 (N_9204,N_6034,N_6081);
nor U9205 (N_9205,N_6423,N_6484);
xnor U9206 (N_9206,N_7024,N_7882);
and U9207 (N_9207,N_7181,N_7350);
nand U9208 (N_9208,N_6691,N_7232);
and U9209 (N_9209,N_7563,N_6112);
nand U9210 (N_9210,N_6221,N_7940);
and U9211 (N_9211,N_7258,N_6604);
nor U9212 (N_9212,N_7697,N_6654);
nand U9213 (N_9213,N_6738,N_7051);
nand U9214 (N_9214,N_6836,N_6720);
nor U9215 (N_9215,N_7408,N_7775);
nor U9216 (N_9216,N_6130,N_6232);
and U9217 (N_9217,N_7634,N_7831);
nor U9218 (N_9218,N_7947,N_6094);
nor U9219 (N_9219,N_7504,N_7682);
nand U9220 (N_9220,N_7109,N_7488);
nand U9221 (N_9221,N_6223,N_7550);
nor U9222 (N_9222,N_7301,N_6594);
or U9223 (N_9223,N_6922,N_7286);
and U9224 (N_9224,N_7661,N_6437);
or U9225 (N_9225,N_7669,N_7457);
nor U9226 (N_9226,N_6988,N_7637);
or U9227 (N_9227,N_6588,N_7117);
or U9228 (N_9228,N_7998,N_7048);
nand U9229 (N_9229,N_7788,N_6584);
or U9230 (N_9230,N_7533,N_7210);
or U9231 (N_9231,N_7823,N_6388);
nand U9232 (N_9232,N_7333,N_7646);
nor U9233 (N_9233,N_7444,N_7238);
and U9234 (N_9234,N_6470,N_7800);
xor U9235 (N_9235,N_6752,N_7957);
and U9236 (N_9236,N_6105,N_7952);
nand U9237 (N_9237,N_7786,N_7343);
and U9238 (N_9238,N_6649,N_7855);
nand U9239 (N_9239,N_7109,N_7003);
or U9240 (N_9240,N_6157,N_7638);
or U9241 (N_9241,N_7040,N_6386);
or U9242 (N_9242,N_6087,N_6456);
or U9243 (N_9243,N_6991,N_6087);
nor U9244 (N_9244,N_7284,N_6160);
nor U9245 (N_9245,N_6702,N_6527);
or U9246 (N_9246,N_6643,N_6982);
nor U9247 (N_9247,N_6148,N_7082);
nand U9248 (N_9248,N_7684,N_7581);
or U9249 (N_9249,N_6850,N_6842);
nor U9250 (N_9250,N_6950,N_7449);
nor U9251 (N_9251,N_7870,N_6845);
or U9252 (N_9252,N_6474,N_7160);
or U9253 (N_9253,N_6705,N_6490);
nor U9254 (N_9254,N_7846,N_7226);
and U9255 (N_9255,N_7092,N_7325);
xnor U9256 (N_9256,N_6885,N_7195);
xor U9257 (N_9257,N_6143,N_6118);
nand U9258 (N_9258,N_6621,N_6355);
and U9259 (N_9259,N_7414,N_6945);
nand U9260 (N_9260,N_7367,N_7417);
nor U9261 (N_9261,N_6985,N_6873);
or U9262 (N_9262,N_7461,N_7840);
and U9263 (N_9263,N_7686,N_6960);
or U9264 (N_9264,N_7501,N_6516);
nand U9265 (N_9265,N_7456,N_6192);
nand U9266 (N_9266,N_7310,N_6318);
nor U9267 (N_9267,N_7096,N_6787);
and U9268 (N_9268,N_7137,N_6423);
nand U9269 (N_9269,N_6518,N_7640);
and U9270 (N_9270,N_7607,N_7946);
nor U9271 (N_9271,N_7924,N_6235);
nor U9272 (N_9272,N_6693,N_6947);
or U9273 (N_9273,N_6952,N_6018);
or U9274 (N_9274,N_7904,N_7193);
nand U9275 (N_9275,N_7853,N_7602);
nor U9276 (N_9276,N_7317,N_6654);
and U9277 (N_9277,N_7546,N_7452);
or U9278 (N_9278,N_7052,N_7138);
and U9279 (N_9279,N_6368,N_7125);
nand U9280 (N_9280,N_6031,N_6917);
xor U9281 (N_9281,N_6707,N_6053);
xnor U9282 (N_9282,N_6830,N_7420);
or U9283 (N_9283,N_7989,N_6601);
and U9284 (N_9284,N_7421,N_7060);
nor U9285 (N_9285,N_7223,N_7536);
nor U9286 (N_9286,N_6148,N_7732);
nand U9287 (N_9287,N_6388,N_6260);
nand U9288 (N_9288,N_7867,N_6002);
nand U9289 (N_9289,N_7323,N_6715);
xnor U9290 (N_9290,N_6910,N_6699);
nand U9291 (N_9291,N_7664,N_7253);
nand U9292 (N_9292,N_7542,N_7304);
or U9293 (N_9293,N_6546,N_7674);
and U9294 (N_9294,N_7104,N_7601);
nand U9295 (N_9295,N_7231,N_7975);
nand U9296 (N_9296,N_7794,N_7735);
nor U9297 (N_9297,N_6551,N_7966);
nand U9298 (N_9298,N_7799,N_7607);
nor U9299 (N_9299,N_7340,N_6076);
nor U9300 (N_9300,N_6739,N_7613);
nand U9301 (N_9301,N_6496,N_6914);
and U9302 (N_9302,N_6620,N_6454);
and U9303 (N_9303,N_6088,N_7973);
nand U9304 (N_9304,N_7796,N_6943);
nor U9305 (N_9305,N_7395,N_6102);
and U9306 (N_9306,N_6057,N_7517);
nand U9307 (N_9307,N_7928,N_6371);
or U9308 (N_9308,N_6856,N_6470);
or U9309 (N_9309,N_6258,N_6237);
xnor U9310 (N_9310,N_6526,N_7152);
or U9311 (N_9311,N_7177,N_7626);
or U9312 (N_9312,N_6445,N_7753);
nand U9313 (N_9313,N_6209,N_7560);
or U9314 (N_9314,N_7103,N_6328);
nor U9315 (N_9315,N_7882,N_7416);
and U9316 (N_9316,N_6221,N_6591);
and U9317 (N_9317,N_6517,N_7446);
and U9318 (N_9318,N_7403,N_6223);
nor U9319 (N_9319,N_7325,N_6936);
nor U9320 (N_9320,N_6752,N_6994);
nand U9321 (N_9321,N_7891,N_6630);
nand U9322 (N_9322,N_7508,N_6641);
and U9323 (N_9323,N_6892,N_7717);
or U9324 (N_9324,N_6872,N_7550);
or U9325 (N_9325,N_6687,N_6648);
nor U9326 (N_9326,N_7442,N_6965);
or U9327 (N_9327,N_7781,N_6722);
and U9328 (N_9328,N_7612,N_7904);
nand U9329 (N_9329,N_7911,N_6654);
or U9330 (N_9330,N_7397,N_6059);
nand U9331 (N_9331,N_7249,N_6583);
nand U9332 (N_9332,N_6000,N_7202);
or U9333 (N_9333,N_7654,N_7785);
and U9334 (N_9334,N_6335,N_6564);
and U9335 (N_9335,N_7808,N_7068);
nor U9336 (N_9336,N_7781,N_7010);
nand U9337 (N_9337,N_6720,N_6117);
nand U9338 (N_9338,N_7000,N_6473);
xor U9339 (N_9339,N_6102,N_6777);
or U9340 (N_9340,N_6594,N_6726);
nand U9341 (N_9341,N_6899,N_6497);
or U9342 (N_9342,N_6994,N_7236);
nor U9343 (N_9343,N_6916,N_6356);
and U9344 (N_9344,N_7760,N_6003);
nor U9345 (N_9345,N_7762,N_6875);
nand U9346 (N_9346,N_7198,N_7819);
nor U9347 (N_9347,N_6040,N_7304);
and U9348 (N_9348,N_7378,N_7065);
xor U9349 (N_9349,N_7390,N_6978);
nor U9350 (N_9350,N_7826,N_6180);
and U9351 (N_9351,N_7922,N_7593);
or U9352 (N_9352,N_6339,N_6209);
nand U9353 (N_9353,N_6715,N_6036);
or U9354 (N_9354,N_6829,N_6623);
and U9355 (N_9355,N_6040,N_6695);
nand U9356 (N_9356,N_7830,N_6920);
and U9357 (N_9357,N_7559,N_6406);
and U9358 (N_9358,N_6359,N_7954);
nand U9359 (N_9359,N_6616,N_6349);
and U9360 (N_9360,N_7981,N_7150);
or U9361 (N_9361,N_7074,N_6224);
nand U9362 (N_9362,N_6981,N_7723);
nand U9363 (N_9363,N_7789,N_7304);
and U9364 (N_9364,N_6911,N_6982);
or U9365 (N_9365,N_7303,N_6664);
and U9366 (N_9366,N_6861,N_7543);
xor U9367 (N_9367,N_6077,N_6053);
xnor U9368 (N_9368,N_6520,N_6234);
or U9369 (N_9369,N_7312,N_7311);
or U9370 (N_9370,N_7728,N_7397);
xnor U9371 (N_9371,N_6465,N_7564);
nand U9372 (N_9372,N_6042,N_6435);
nor U9373 (N_9373,N_7052,N_6562);
nand U9374 (N_9374,N_6451,N_7299);
xor U9375 (N_9375,N_6438,N_6207);
nor U9376 (N_9376,N_6156,N_6628);
nor U9377 (N_9377,N_6667,N_7753);
or U9378 (N_9378,N_6191,N_7558);
or U9379 (N_9379,N_6909,N_6708);
nor U9380 (N_9380,N_7139,N_6828);
or U9381 (N_9381,N_6163,N_6405);
nor U9382 (N_9382,N_6194,N_7941);
nor U9383 (N_9383,N_7574,N_6535);
and U9384 (N_9384,N_6630,N_6906);
nand U9385 (N_9385,N_6330,N_7043);
or U9386 (N_9386,N_6220,N_6935);
or U9387 (N_9387,N_7461,N_6803);
nor U9388 (N_9388,N_7618,N_6313);
and U9389 (N_9389,N_6062,N_6223);
nand U9390 (N_9390,N_6008,N_6242);
nor U9391 (N_9391,N_7085,N_6913);
and U9392 (N_9392,N_7919,N_6498);
nand U9393 (N_9393,N_7237,N_6648);
xnor U9394 (N_9394,N_7122,N_7111);
nor U9395 (N_9395,N_7277,N_6505);
xnor U9396 (N_9396,N_7922,N_6778);
nor U9397 (N_9397,N_6504,N_7666);
and U9398 (N_9398,N_6123,N_6733);
nor U9399 (N_9399,N_7672,N_7889);
nand U9400 (N_9400,N_7763,N_6859);
or U9401 (N_9401,N_7607,N_6090);
and U9402 (N_9402,N_6706,N_6783);
and U9403 (N_9403,N_6227,N_7056);
and U9404 (N_9404,N_6893,N_7015);
nand U9405 (N_9405,N_6235,N_7723);
or U9406 (N_9406,N_6129,N_7332);
nand U9407 (N_9407,N_7711,N_7095);
and U9408 (N_9408,N_6392,N_7667);
or U9409 (N_9409,N_7478,N_6636);
nor U9410 (N_9410,N_6988,N_7053);
nand U9411 (N_9411,N_7551,N_6862);
xnor U9412 (N_9412,N_6806,N_6135);
xnor U9413 (N_9413,N_7599,N_6379);
xnor U9414 (N_9414,N_7499,N_6904);
and U9415 (N_9415,N_7147,N_6580);
or U9416 (N_9416,N_7435,N_7098);
and U9417 (N_9417,N_7086,N_7577);
nor U9418 (N_9418,N_6031,N_7271);
nor U9419 (N_9419,N_6128,N_7517);
nand U9420 (N_9420,N_6273,N_6458);
and U9421 (N_9421,N_7773,N_6967);
nor U9422 (N_9422,N_7918,N_6887);
and U9423 (N_9423,N_7890,N_7391);
or U9424 (N_9424,N_7972,N_6757);
and U9425 (N_9425,N_7612,N_6278);
xor U9426 (N_9426,N_7983,N_6183);
or U9427 (N_9427,N_7215,N_7909);
nand U9428 (N_9428,N_6794,N_6219);
or U9429 (N_9429,N_7574,N_7526);
or U9430 (N_9430,N_7759,N_7915);
nor U9431 (N_9431,N_7588,N_6232);
nand U9432 (N_9432,N_6611,N_6926);
nand U9433 (N_9433,N_7370,N_7174);
nand U9434 (N_9434,N_7129,N_6931);
nor U9435 (N_9435,N_7862,N_7873);
nor U9436 (N_9436,N_7102,N_7329);
nor U9437 (N_9437,N_7495,N_6791);
or U9438 (N_9438,N_7521,N_7289);
and U9439 (N_9439,N_7670,N_7419);
nor U9440 (N_9440,N_6978,N_6770);
or U9441 (N_9441,N_6154,N_6689);
and U9442 (N_9442,N_7997,N_6426);
xor U9443 (N_9443,N_6723,N_7657);
or U9444 (N_9444,N_6258,N_7398);
or U9445 (N_9445,N_6108,N_6118);
nand U9446 (N_9446,N_6019,N_6373);
or U9447 (N_9447,N_6502,N_6646);
and U9448 (N_9448,N_6211,N_6997);
nor U9449 (N_9449,N_7075,N_7396);
or U9450 (N_9450,N_6619,N_6467);
nor U9451 (N_9451,N_7472,N_6938);
or U9452 (N_9452,N_6970,N_7090);
and U9453 (N_9453,N_7919,N_6122);
nand U9454 (N_9454,N_6015,N_7190);
and U9455 (N_9455,N_7561,N_6676);
nand U9456 (N_9456,N_6942,N_7948);
and U9457 (N_9457,N_6655,N_6331);
nor U9458 (N_9458,N_7978,N_7845);
nand U9459 (N_9459,N_6464,N_6239);
nor U9460 (N_9460,N_6634,N_7916);
nor U9461 (N_9461,N_6176,N_6480);
and U9462 (N_9462,N_6002,N_6951);
nor U9463 (N_9463,N_7337,N_7568);
or U9464 (N_9464,N_6356,N_7758);
and U9465 (N_9465,N_6132,N_6512);
nor U9466 (N_9466,N_7136,N_7319);
nor U9467 (N_9467,N_6801,N_6649);
or U9468 (N_9468,N_6090,N_7102);
nand U9469 (N_9469,N_7788,N_7055);
and U9470 (N_9470,N_7871,N_6020);
and U9471 (N_9471,N_6876,N_7096);
nand U9472 (N_9472,N_6008,N_7936);
or U9473 (N_9473,N_6483,N_7863);
nor U9474 (N_9474,N_7189,N_7322);
xnor U9475 (N_9475,N_7166,N_6938);
nand U9476 (N_9476,N_6863,N_6276);
nor U9477 (N_9477,N_6416,N_7556);
nor U9478 (N_9478,N_7997,N_6885);
and U9479 (N_9479,N_7151,N_6949);
and U9480 (N_9480,N_6853,N_7837);
xnor U9481 (N_9481,N_7105,N_7152);
nor U9482 (N_9482,N_6132,N_6993);
nor U9483 (N_9483,N_7879,N_7733);
nor U9484 (N_9484,N_7008,N_7073);
or U9485 (N_9485,N_6971,N_6137);
xor U9486 (N_9486,N_6920,N_7762);
nand U9487 (N_9487,N_7982,N_6225);
and U9488 (N_9488,N_7216,N_7378);
or U9489 (N_9489,N_6094,N_7400);
nor U9490 (N_9490,N_7444,N_6541);
nor U9491 (N_9491,N_6416,N_7251);
nand U9492 (N_9492,N_6804,N_6338);
nor U9493 (N_9493,N_6023,N_7960);
nor U9494 (N_9494,N_7287,N_7554);
or U9495 (N_9495,N_6231,N_6583);
xnor U9496 (N_9496,N_7114,N_7804);
xor U9497 (N_9497,N_6591,N_7491);
and U9498 (N_9498,N_7880,N_7530);
nor U9499 (N_9499,N_7643,N_7058);
and U9500 (N_9500,N_7187,N_6635);
nor U9501 (N_9501,N_6720,N_7459);
nor U9502 (N_9502,N_6388,N_7326);
xnor U9503 (N_9503,N_7430,N_7770);
xnor U9504 (N_9504,N_7370,N_7693);
or U9505 (N_9505,N_7678,N_7689);
or U9506 (N_9506,N_6247,N_6234);
nor U9507 (N_9507,N_6734,N_6180);
or U9508 (N_9508,N_6160,N_7186);
nor U9509 (N_9509,N_7702,N_6107);
or U9510 (N_9510,N_6250,N_6304);
and U9511 (N_9511,N_6116,N_7431);
nor U9512 (N_9512,N_7264,N_7706);
xnor U9513 (N_9513,N_6605,N_7731);
nor U9514 (N_9514,N_7048,N_6238);
nand U9515 (N_9515,N_6405,N_7368);
nor U9516 (N_9516,N_7326,N_6799);
or U9517 (N_9517,N_7765,N_7964);
nor U9518 (N_9518,N_6957,N_7879);
and U9519 (N_9519,N_6675,N_6649);
nor U9520 (N_9520,N_6919,N_7666);
nand U9521 (N_9521,N_6327,N_7873);
nand U9522 (N_9522,N_7178,N_6456);
or U9523 (N_9523,N_7236,N_6672);
or U9524 (N_9524,N_6598,N_6988);
nand U9525 (N_9525,N_6894,N_7049);
nand U9526 (N_9526,N_6134,N_7868);
or U9527 (N_9527,N_6581,N_7716);
nor U9528 (N_9528,N_7948,N_6522);
nor U9529 (N_9529,N_6045,N_7400);
nand U9530 (N_9530,N_6705,N_6571);
and U9531 (N_9531,N_7739,N_7874);
or U9532 (N_9532,N_7549,N_7800);
xnor U9533 (N_9533,N_6362,N_7195);
and U9534 (N_9534,N_7698,N_6306);
nor U9535 (N_9535,N_6800,N_7286);
nor U9536 (N_9536,N_7926,N_7243);
or U9537 (N_9537,N_7545,N_6503);
nor U9538 (N_9538,N_7030,N_7119);
and U9539 (N_9539,N_7127,N_7966);
xnor U9540 (N_9540,N_6686,N_7162);
and U9541 (N_9541,N_7270,N_6144);
and U9542 (N_9542,N_6982,N_6471);
or U9543 (N_9543,N_6980,N_7543);
nor U9544 (N_9544,N_7983,N_7206);
and U9545 (N_9545,N_7679,N_7401);
or U9546 (N_9546,N_7443,N_7710);
nand U9547 (N_9547,N_7509,N_7034);
nor U9548 (N_9548,N_7678,N_7581);
nor U9549 (N_9549,N_6797,N_7022);
or U9550 (N_9550,N_7934,N_7987);
and U9551 (N_9551,N_6361,N_6931);
or U9552 (N_9552,N_6209,N_6546);
or U9553 (N_9553,N_6768,N_7617);
xor U9554 (N_9554,N_6275,N_6125);
nand U9555 (N_9555,N_6055,N_6525);
nor U9556 (N_9556,N_6988,N_7409);
nor U9557 (N_9557,N_7339,N_6607);
nor U9558 (N_9558,N_7732,N_6757);
and U9559 (N_9559,N_7044,N_6835);
xnor U9560 (N_9560,N_6925,N_6567);
nor U9561 (N_9561,N_6822,N_6296);
nor U9562 (N_9562,N_6514,N_6786);
nor U9563 (N_9563,N_7364,N_7756);
or U9564 (N_9564,N_7812,N_7067);
nand U9565 (N_9565,N_7541,N_7517);
nor U9566 (N_9566,N_7255,N_6034);
xnor U9567 (N_9567,N_6890,N_6834);
or U9568 (N_9568,N_7294,N_7070);
and U9569 (N_9569,N_6158,N_6203);
and U9570 (N_9570,N_7168,N_6304);
and U9571 (N_9571,N_7576,N_6996);
xnor U9572 (N_9572,N_6435,N_7823);
nand U9573 (N_9573,N_6526,N_7890);
nor U9574 (N_9574,N_6428,N_7899);
nand U9575 (N_9575,N_7180,N_7267);
and U9576 (N_9576,N_7939,N_7682);
or U9577 (N_9577,N_7498,N_6541);
or U9578 (N_9578,N_7037,N_7014);
or U9579 (N_9579,N_6210,N_6149);
xnor U9580 (N_9580,N_6457,N_7058);
nand U9581 (N_9581,N_7969,N_6675);
or U9582 (N_9582,N_6684,N_7803);
and U9583 (N_9583,N_7495,N_6832);
and U9584 (N_9584,N_6451,N_7559);
and U9585 (N_9585,N_7665,N_6990);
or U9586 (N_9586,N_7964,N_6056);
or U9587 (N_9587,N_7701,N_6578);
nor U9588 (N_9588,N_6009,N_7505);
xnor U9589 (N_9589,N_6121,N_7733);
xnor U9590 (N_9590,N_7688,N_6781);
and U9591 (N_9591,N_6167,N_6419);
nor U9592 (N_9592,N_6327,N_7288);
xnor U9593 (N_9593,N_6872,N_7243);
nand U9594 (N_9594,N_7980,N_7099);
or U9595 (N_9595,N_6901,N_7038);
nor U9596 (N_9596,N_6032,N_7640);
or U9597 (N_9597,N_7317,N_7739);
nor U9598 (N_9598,N_7578,N_7033);
nor U9599 (N_9599,N_6668,N_6140);
xor U9600 (N_9600,N_6042,N_6393);
or U9601 (N_9601,N_7523,N_6097);
nand U9602 (N_9602,N_7711,N_7565);
or U9603 (N_9603,N_6060,N_7097);
nand U9604 (N_9604,N_7982,N_6544);
or U9605 (N_9605,N_7681,N_7918);
nor U9606 (N_9606,N_7161,N_7144);
and U9607 (N_9607,N_7245,N_7011);
or U9608 (N_9608,N_6903,N_6832);
and U9609 (N_9609,N_7020,N_7195);
and U9610 (N_9610,N_7133,N_6966);
and U9611 (N_9611,N_7072,N_7778);
nand U9612 (N_9612,N_7502,N_7262);
and U9613 (N_9613,N_6533,N_6708);
or U9614 (N_9614,N_6445,N_6652);
xnor U9615 (N_9615,N_6018,N_7482);
nor U9616 (N_9616,N_6818,N_7798);
xor U9617 (N_9617,N_6902,N_7592);
nor U9618 (N_9618,N_7005,N_6455);
or U9619 (N_9619,N_6997,N_7562);
and U9620 (N_9620,N_7135,N_7433);
nand U9621 (N_9621,N_6717,N_6489);
nor U9622 (N_9622,N_7097,N_7090);
and U9623 (N_9623,N_6384,N_6675);
nand U9624 (N_9624,N_6650,N_7549);
or U9625 (N_9625,N_7530,N_7857);
or U9626 (N_9626,N_7241,N_6812);
nand U9627 (N_9627,N_6340,N_7828);
and U9628 (N_9628,N_7371,N_6517);
and U9629 (N_9629,N_7399,N_6835);
xnor U9630 (N_9630,N_7939,N_7437);
and U9631 (N_9631,N_6593,N_7510);
nand U9632 (N_9632,N_7116,N_7593);
nand U9633 (N_9633,N_7638,N_7337);
nor U9634 (N_9634,N_6403,N_6472);
or U9635 (N_9635,N_6086,N_6057);
nand U9636 (N_9636,N_7076,N_6845);
or U9637 (N_9637,N_6905,N_7984);
and U9638 (N_9638,N_7837,N_6526);
and U9639 (N_9639,N_6236,N_7507);
nand U9640 (N_9640,N_6560,N_7609);
or U9641 (N_9641,N_6457,N_6771);
nor U9642 (N_9642,N_7177,N_7096);
nor U9643 (N_9643,N_6543,N_7648);
and U9644 (N_9644,N_7292,N_6369);
nand U9645 (N_9645,N_6881,N_7086);
nor U9646 (N_9646,N_7567,N_7786);
xnor U9647 (N_9647,N_7038,N_6746);
or U9648 (N_9648,N_6450,N_7022);
xnor U9649 (N_9649,N_7114,N_7749);
nand U9650 (N_9650,N_7388,N_6313);
nand U9651 (N_9651,N_6085,N_7733);
and U9652 (N_9652,N_6334,N_6820);
xnor U9653 (N_9653,N_6426,N_7341);
xnor U9654 (N_9654,N_7095,N_7606);
xor U9655 (N_9655,N_6651,N_6392);
nor U9656 (N_9656,N_7371,N_7298);
nand U9657 (N_9657,N_7149,N_7781);
nand U9658 (N_9658,N_6188,N_7748);
or U9659 (N_9659,N_7323,N_7045);
nor U9660 (N_9660,N_7532,N_7661);
xnor U9661 (N_9661,N_6023,N_6066);
nor U9662 (N_9662,N_6590,N_7860);
or U9663 (N_9663,N_7523,N_7832);
or U9664 (N_9664,N_7593,N_6555);
xnor U9665 (N_9665,N_7425,N_6206);
nand U9666 (N_9666,N_6332,N_7373);
and U9667 (N_9667,N_6710,N_6817);
nand U9668 (N_9668,N_6952,N_7191);
nand U9669 (N_9669,N_7929,N_7241);
nand U9670 (N_9670,N_6131,N_6282);
nor U9671 (N_9671,N_7202,N_7895);
and U9672 (N_9672,N_7063,N_6167);
xnor U9673 (N_9673,N_6937,N_7875);
xor U9674 (N_9674,N_6184,N_6368);
nand U9675 (N_9675,N_7828,N_7934);
nand U9676 (N_9676,N_7348,N_6293);
and U9677 (N_9677,N_6617,N_7586);
or U9678 (N_9678,N_6926,N_6768);
nand U9679 (N_9679,N_7787,N_6773);
nand U9680 (N_9680,N_7941,N_7169);
nor U9681 (N_9681,N_6682,N_7916);
nand U9682 (N_9682,N_7587,N_7683);
and U9683 (N_9683,N_7640,N_6006);
and U9684 (N_9684,N_6997,N_6900);
or U9685 (N_9685,N_7171,N_7249);
and U9686 (N_9686,N_7051,N_6942);
and U9687 (N_9687,N_7436,N_7550);
and U9688 (N_9688,N_6748,N_6305);
and U9689 (N_9689,N_7399,N_7935);
nor U9690 (N_9690,N_6448,N_6091);
and U9691 (N_9691,N_7274,N_6502);
nand U9692 (N_9692,N_7648,N_7187);
nor U9693 (N_9693,N_7034,N_6659);
nor U9694 (N_9694,N_6771,N_6214);
nand U9695 (N_9695,N_7449,N_7206);
or U9696 (N_9696,N_7231,N_7343);
and U9697 (N_9697,N_6358,N_7042);
nand U9698 (N_9698,N_6449,N_7540);
nand U9699 (N_9699,N_6628,N_6294);
or U9700 (N_9700,N_7144,N_7280);
or U9701 (N_9701,N_6835,N_6062);
or U9702 (N_9702,N_6343,N_6864);
and U9703 (N_9703,N_7112,N_7640);
nor U9704 (N_9704,N_7327,N_7457);
or U9705 (N_9705,N_6313,N_6861);
and U9706 (N_9706,N_7951,N_6917);
xor U9707 (N_9707,N_7843,N_7352);
xor U9708 (N_9708,N_7494,N_7696);
or U9709 (N_9709,N_6561,N_7149);
or U9710 (N_9710,N_7774,N_6477);
or U9711 (N_9711,N_7314,N_6842);
and U9712 (N_9712,N_6714,N_6846);
nand U9713 (N_9713,N_7213,N_6702);
and U9714 (N_9714,N_6831,N_7733);
nand U9715 (N_9715,N_6053,N_6209);
nand U9716 (N_9716,N_6289,N_6581);
xnor U9717 (N_9717,N_7585,N_6825);
or U9718 (N_9718,N_6056,N_6652);
xnor U9719 (N_9719,N_6297,N_7964);
or U9720 (N_9720,N_7809,N_7450);
nor U9721 (N_9721,N_6907,N_7016);
nand U9722 (N_9722,N_7656,N_6646);
nand U9723 (N_9723,N_7476,N_7985);
nor U9724 (N_9724,N_6623,N_6465);
or U9725 (N_9725,N_7981,N_7498);
nand U9726 (N_9726,N_6327,N_7675);
nor U9727 (N_9727,N_6270,N_7956);
nor U9728 (N_9728,N_6368,N_6556);
or U9729 (N_9729,N_6671,N_6002);
and U9730 (N_9730,N_7939,N_7302);
xnor U9731 (N_9731,N_6389,N_7833);
or U9732 (N_9732,N_7140,N_7109);
and U9733 (N_9733,N_7428,N_7793);
or U9734 (N_9734,N_7857,N_6269);
nor U9735 (N_9735,N_6512,N_6694);
or U9736 (N_9736,N_7696,N_6528);
or U9737 (N_9737,N_7765,N_7436);
or U9738 (N_9738,N_7679,N_6399);
nand U9739 (N_9739,N_7943,N_7768);
and U9740 (N_9740,N_6609,N_7595);
xnor U9741 (N_9741,N_7918,N_7132);
nor U9742 (N_9742,N_6999,N_6354);
and U9743 (N_9743,N_7116,N_7037);
and U9744 (N_9744,N_6435,N_7008);
nand U9745 (N_9745,N_7073,N_7461);
nor U9746 (N_9746,N_6281,N_7003);
and U9747 (N_9747,N_6564,N_6312);
nor U9748 (N_9748,N_6913,N_7690);
nand U9749 (N_9749,N_6861,N_7567);
nor U9750 (N_9750,N_6630,N_7729);
or U9751 (N_9751,N_6336,N_7187);
and U9752 (N_9752,N_7196,N_7719);
or U9753 (N_9753,N_6047,N_7572);
nor U9754 (N_9754,N_6192,N_6983);
nor U9755 (N_9755,N_6286,N_7358);
or U9756 (N_9756,N_6693,N_6310);
and U9757 (N_9757,N_7693,N_7552);
or U9758 (N_9758,N_7353,N_7840);
or U9759 (N_9759,N_6539,N_7196);
nand U9760 (N_9760,N_6436,N_7808);
nand U9761 (N_9761,N_7413,N_6529);
or U9762 (N_9762,N_6071,N_6554);
or U9763 (N_9763,N_7579,N_6432);
nor U9764 (N_9764,N_7582,N_6221);
and U9765 (N_9765,N_7400,N_6532);
and U9766 (N_9766,N_7307,N_7495);
or U9767 (N_9767,N_7588,N_6074);
nand U9768 (N_9768,N_6722,N_6753);
and U9769 (N_9769,N_6858,N_6265);
nor U9770 (N_9770,N_6049,N_7653);
nand U9771 (N_9771,N_6261,N_7907);
nor U9772 (N_9772,N_6332,N_6172);
or U9773 (N_9773,N_6826,N_7496);
and U9774 (N_9774,N_6999,N_6551);
or U9775 (N_9775,N_6711,N_6735);
and U9776 (N_9776,N_7486,N_6911);
nor U9777 (N_9777,N_6937,N_7144);
nor U9778 (N_9778,N_7751,N_6627);
or U9779 (N_9779,N_6661,N_7383);
or U9780 (N_9780,N_7745,N_6666);
nand U9781 (N_9781,N_7470,N_6534);
and U9782 (N_9782,N_6283,N_7715);
and U9783 (N_9783,N_6609,N_7363);
nand U9784 (N_9784,N_7992,N_6452);
or U9785 (N_9785,N_7756,N_7405);
or U9786 (N_9786,N_6130,N_6155);
nor U9787 (N_9787,N_6493,N_7876);
xnor U9788 (N_9788,N_6787,N_6631);
or U9789 (N_9789,N_7799,N_6886);
nand U9790 (N_9790,N_7952,N_7332);
nor U9791 (N_9791,N_6353,N_7121);
xnor U9792 (N_9792,N_6195,N_7494);
or U9793 (N_9793,N_7362,N_6325);
and U9794 (N_9794,N_6959,N_6161);
and U9795 (N_9795,N_6153,N_6203);
nand U9796 (N_9796,N_6058,N_6818);
nor U9797 (N_9797,N_7730,N_7075);
nor U9798 (N_9798,N_7546,N_6146);
nor U9799 (N_9799,N_7867,N_7437);
nand U9800 (N_9800,N_6832,N_7373);
nor U9801 (N_9801,N_6010,N_7587);
nor U9802 (N_9802,N_6142,N_6500);
nand U9803 (N_9803,N_7369,N_7411);
nor U9804 (N_9804,N_7423,N_6423);
and U9805 (N_9805,N_6528,N_7229);
nand U9806 (N_9806,N_7437,N_6945);
or U9807 (N_9807,N_6609,N_6714);
nand U9808 (N_9808,N_6663,N_7559);
or U9809 (N_9809,N_7776,N_6895);
xor U9810 (N_9810,N_7487,N_6404);
or U9811 (N_9811,N_7204,N_7628);
and U9812 (N_9812,N_6027,N_6257);
and U9813 (N_9813,N_7457,N_6660);
nor U9814 (N_9814,N_7045,N_7897);
xor U9815 (N_9815,N_6363,N_6358);
nand U9816 (N_9816,N_6168,N_6546);
xnor U9817 (N_9817,N_6675,N_7441);
nand U9818 (N_9818,N_6518,N_7870);
and U9819 (N_9819,N_6841,N_6561);
nor U9820 (N_9820,N_7257,N_7585);
nand U9821 (N_9821,N_7072,N_7841);
and U9822 (N_9822,N_6461,N_6561);
and U9823 (N_9823,N_7509,N_7335);
nor U9824 (N_9824,N_6407,N_7715);
or U9825 (N_9825,N_6271,N_6534);
or U9826 (N_9826,N_7266,N_7831);
or U9827 (N_9827,N_6397,N_6284);
nand U9828 (N_9828,N_6813,N_7186);
and U9829 (N_9829,N_6705,N_7925);
nand U9830 (N_9830,N_7601,N_6883);
and U9831 (N_9831,N_6879,N_6190);
nor U9832 (N_9832,N_7554,N_6038);
nor U9833 (N_9833,N_6640,N_7427);
or U9834 (N_9834,N_6964,N_7174);
and U9835 (N_9835,N_7100,N_6839);
nand U9836 (N_9836,N_7646,N_7852);
xnor U9837 (N_9837,N_7486,N_6774);
or U9838 (N_9838,N_7979,N_6054);
nand U9839 (N_9839,N_6997,N_6799);
nor U9840 (N_9840,N_6471,N_7544);
nor U9841 (N_9841,N_7590,N_7823);
nor U9842 (N_9842,N_7797,N_6336);
or U9843 (N_9843,N_7530,N_6154);
or U9844 (N_9844,N_7482,N_7518);
or U9845 (N_9845,N_6848,N_7334);
and U9846 (N_9846,N_7104,N_6996);
or U9847 (N_9847,N_6509,N_6909);
nor U9848 (N_9848,N_6635,N_7306);
or U9849 (N_9849,N_6748,N_7163);
and U9850 (N_9850,N_7708,N_7214);
or U9851 (N_9851,N_6820,N_7725);
and U9852 (N_9852,N_7597,N_7680);
xnor U9853 (N_9853,N_7842,N_7455);
nand U9854 (N_9854,N_6237,N_7919);
nand U9855 (N_9855,N_7240,N_6699);
and U9856 (N_9856,N_7266,N_6695);
and U9857 (N_9857,N_7173,N_6696);
nor U9858 (N_9858,N_7895,N_7488);
nor U9859 (N_9859,N_7436,N_6507);
and U9860 (N_9860,N_7767,N_6702);
or U9861 (N_9861,N_6410,N_6274);
nor U9862 (N_9862,N_7251,N_6904);
or U9863 (N_9863,N_6696,N_7702);
xor U9864 (N_9864,N_6061,N_6102);
xnor U9865 (N_9865,N_7500,N_7692);
and U9866 (N_9866,N_7064,N_7730);
and U9867 (N_9867,N_6250,N_7718);
xor U9868 (N_9868,N_6795,N_6361);
nor U9869 (N_9869,N_6653,N_6896);
nor U9870 (N_9870,N_7440,N_7372);
nand U9871 (N_9871,N_7624,N_7214);
or U9872 (N_9872,N_7424,N_7363);
nand U9873 (N_9873,N_7669,N_6386);
and U9874 (N_9874,N_7818,N_7807);
or U9875 (N_9875,N_7242,N_6088);
xor U9876 (N_9876,N_6061,N_6910);
or U9877 (N_9877,N_7608,N_6460);
nor U9878 (N_9878,N_6495,N_6793);
nand U9879 (N_9879,N_6544,N_6948);
nor U9880 (N_9880,N_7361,N_7015);
or U9881 (N_9881,N_7947,N_7113);
nand U9882 (N_9882,N_6885,N_7846);
or U9883 (N_9883,N_6233,N_7877);
or U9884 (N_9884,N_7250,N_7550);
nor U9885 (N_9885,N_7912,N_7951);
and U9886 (N_9886,N_6122,N_6463);
xor U9887 (N_9887,N_6611,N_6185);
nand U9888 (N_9888,N_6106,N_7421);
or U9889 (N_9889,N_7549,N_6149);
or U9890 (N_9890,N_7628,N_6341);
nand U9891 (N_9891,N_7988,N_7299);
or U9892 (N_9892,N_6873,N_6949);
nor U9893 (N_9893,N_6170,N_7027);
nand U9894 (N_9894,N_7661,N_7630);
nand U9895 (N_9895,N_6058,N_7372);
nand U9896 (N_9896,N_7567,N_7799);
nor U9897 (N_9897,N_7940,N_6671);
nor U9898 (N_9898,N_7554,N_7168);
or U9899 (N_9899,N_6674,N_6060);
nor U9900 (N_9900,N_6669,N_7052);
xnor U9901 (N_9901,N_6084,N_7990);
and U9902 (N_9902,N_6483,N_7966);
or U9903 (N_9903,N_7475,N_7335);
xor U9904 (N_9904,N_7017,N_6440);
nand U9905 (N_9905,N_7924,N_7143);
and U9906 (N_9906,N_7035,N_6146);
xnor U9907 (N_9907,N_6834,N_7313);
nor U9908 (N_9908,N_7123,N_6849);
or U9909 (N_9909,N_6082,N_7642);
nand U9910 (N_9910,N_6919,N_7695);
and U9911 (N_9911,N_6067,N_7732);
xor U9912 (N_9912,N_7540,N_6353);
or U9913 (N_9913,N_6714,N_7202);
nand U9914 (N_9914,N_6320,N_6775);
or U9915 (N_9915,N_7200,N_6219);
nor U9916 (N_9916,N_6968,N_7586);
or U9917 (N_9917,N_7393,N_6778);
and U9918 (N_9918,N_7183,N_7180);
nor U9919 (N_9919,N_7228,N_7646);
and U9920 (N_9920,N_6678,N_7628);
and U9921 (N_9921,N_6416,N_7829);
nor U9922 (N_9922,N_7593,N_6662);
nor U9923 (N_9923,N_7274,N_7225);
and U9924 (N_9924,N_7168,N_6035);
nor U9925 (N_9925,N_6349,N_7269);
and U9926 (N_9926,N_7201,N_6305);
and U9927 (N_9927,N_7739,N_6080);
and U9928 (N_9928,N_6984,N_7594);
nand U9929 (N_9929,N_6395,N_7656);
and U9930 (N_9930,N_7920,N_7662);
or U9931 (N_9931,N_6268,N_6219);
nor U9932 (N_9932,N_7424,N_6306);
or U9933 (N_9933,N_6039,N_7748);
nor U9934 (N_9934,N_6944,N_7655);
nor U9935 (N_9935,N_6342,N_7757);
nand U9936 (N_9936,N_7775,N_6895);
or U9937 (N_9937,N_7864,N_6489);
and U9938 (N_9938,N_6780,N_6540);
and U9939 (N_9939,N_6962,N_6171);
and U9940 (N_9940,N_6608,N_6135);
xnor U9941 (N_9941,N_7690,N_7269);
nand U9942 (N_9942,N_6122,N_7243);
and U9943 (N_9943,N_6809,N_7295);
nand U9944 (N_9944,N_7051,N_6963);
and U9945 (N_9945,N_7535,N_6308);
or U9946 (N_9946,N_6871,N_7445);
nor U9947 (N_9947,N_7734,N_7114);
nor U9948 (N_9948,N_7522,N_7281);
nand U9949 (N_9949,N_6377,N_7612);
nor U9950 (N_9950,N_7876,N_6531);
nor U9951 (N_9951,N_7518,N_6362);
and U9952 (N_9952,N_7590,N_7009);
or U9953 (N_9953,N_6032,N_7139);
xor U9954 (N_9954,N_7176,N_7132);
or U9955 (N_9955,N_6387,N_7604);
and U9956 (N_9956,N_7705,N_6686);
xor U9957 (N_9957,N_6273,N_7478);
or U9958 (N_9958,N_7491,N_7011);
and U9959 (N_9959,N_7012,N_6122);
and U9960 (N_9960,N_7086,N_6265);
nor U9961 (N_9961,N_6937,N_7076);
nand U9962 (N_9962,N_6777,N_7352);
nand U9963 (N_9963,N_7096,N_6381);
nand U9964 (N_9964,N_7943,N_7139);
and U9965 (N_9965,N_6842,N_6930);
xor U9966 (N_9966,N_6762,N_7274);
and U9967 (N_9967,N_6796,N_6081);
nor U9968 (N_9968,N_6235,N_7647);
nand U9969 (N_9969,N_7027,N_6990);
nor U9970 (N_9970,N_6652,N_7269);
nor U9971 (N_9971,N_6508,N_6220);
or U9972 (N_9972,N_6638,N_7252);
nor U9973 (N_9973,N_6032,N_7524);
nor U9974 (N_9974,N_6299,N_7732);
nand U9975 (N_9975,N_6990,N_6399);
nor U9976 (N_9976,N_6351,N_7816);
nor U9977 (N_9977,N_7745,N_7685);
or U9978 (N_9978,N_7409,N_6489);
and U9979 (N_9979,N_6389,N_6004);
and U9980 (N_9980,N_6097,N_6140);
and U9981 (N_9981,N_7871,N_6953);
nand U9982 (N_9982,N_6758,N_6669);
nor U9983 (N_9983,N_7241,N_7035);
nor U9984 (N_9984,N_6342,N_6739);
xnor U9985 (N_9985,N_7037,N_6742);
nor U9986 (N_9986,N_7983,N_6455);
nor U9987 (N_9987,N_6498,N_7297);
nand U9988 (N_9988,N_6713,N_6250);
nand U9989 (N_9989,N_7826,N_6014);
and U9990 (N_9990,N_7339,N_6669);
and U9991 (N_9991,N_6102,N_6216);
or U9992 (N_9992,N_7464,N_7661);
nand U9993 (N_9993,N_7489,N_7388);
nor U9994 (N_9994,N_7634,N_7350);
nand U9995 (N_9995,N_6168,N_6149);
or U9996 (N_9996,N_6822,N_6006);
nand U9997 (N_9997,N_6979,N_7744);
and U9998 (N_9998,N_7311,N_6258);
and U9999 (N_9999,N_7683,N_7146);
nand U10000 (N_10000,N_8169,N_8266);
or U10001 (N_10001,N_9319,N_9865);
and U10002 (N_10002,N_9476,N_9818);
xnor U10003 (N_10003,N_8999,N_9913);
and U10004 (N_10004,N_9722,N_8708);
nor U10005 (N_10005,N_9196,N_8632);
or U10006 (N_10006,N_8384,N_9915);
nor U10007 (N_10007,N_9153,N_9210);
and U10008 (N_10008,N_9683,N_9755);
nand U10009 (N_10009,N_9531,N_9439);
or U10010 (N_10010,N_8642,N_9647);
nand U10011 (N_10011,N_8952,N_8785);
and U10012 (N_10012,N_8457,N_9745);
or U10013 (N_10013,N_8887,N_8964);
nand U10014 (N_10014,N_8331,N_9332);
or U10015 (N_10015,N_8661,N_9864);
nand U10016 (N_10016,N_8564,N_9374);
and U10017 (N_10017,N_8637,N_8685);
and U10018 (N_10018,N_9324,N_8795);
nor U10019 (N_10019,N_8680,N_8627);
or U10020 (N_10020,N_9856,N_9232);
and U10021 (N_10021,N_9654,N_9260);
and U10022 (N_10022,N_8601,N_8466);
or U10023 (N_10023,N_9455,N_8065);
and U10024 (N_10024,N_8376,N_9958);
or U10025 (N_10025,N_9699,N_8584);
nor U10026 (N_10026,N_9032,N_9488);
nor U10027 (N_10027,N_9806,N_9621);
or U10028 (N_10028,N_8748,N_8617);
nand U10029 (N_10029,N_9545,N_9307);
nand U10030 (N_10030,N_8890,N_9892);
and U10031 (N_10031,N_9614,N_8934);
or U10032 (N_10032,N_8931,N_8888);
nor U10033 (N_10033,N_8421,N_8413);
nand U10034 (N_10034,N_9199,N_8358);
or U10035 (N_10035,N_9570,N_9867);
xnor U10036 (N_10036,N_8396,N_8096);
nand U10037 (N_10037,N_9236,N_9036);
nor U10038 (N_10038,N_8310,N_8140);
nand U10039 (N_10039,N_8416,N_9623);
xor U10040 (N_10040,N_8640,N_8092);
nand U10041 (N_10041,N_8225,N_8148);
nand U10042 (N_10042,N_8390,N_8268);
xnor U10043 (N_10043,N_9854,N_9300);
xnor U10044 (N_10044,N_9747,N_9180);
nand U10045 (N_10045,N_9428,N_8496);
nand U10046 (N_10046,N_8633,N_8389);
or U10047 (N_10047,N_8347,N_8136);
and U10048 (N_10048,N_8075,N_8764);
and U10049 (N_10049,N_8700,N_9471);
nand U10050 (N_10050,N_8976,N_9863);
nor U10051 (N_10051,N_8682,N_9167);
or U10052 (N_10052,N_9100,N_8377);
and U10053 (N_10053,N_9157,N_8525);
nor U10054 (N_10054,N_9228,N_8497);
nor U10055 (N_10055,N_8248,N_8908);
and U10056 (N_10056,N_9619,N_8520);
or U10057 (N_10057,N_8866,N_9787);
nor U10058 (N_10058,N_9861,N_8307);
xor U10059 (N_10059,N_9390,N_8769);
nand U10060 (N_10060,N_9530,N_9600);
and U10061 (N_10061,N_8287,N_9959);
nand U10062 (N_10062,N_9176,N_8158);
nor U10063 (N_10063,N_9447,N_8576);
and U10064 (N_10064,N_8464,N_9487);
or U10065 (N_10065,N_8736,N_8926);
nor U10066 (N_10066,N_8198,N_9509);
nor U10067 (N_10067,N_8154,N_9386);
nand U10068 (N_10068,N_9443,N_9735);
nand U10069 (N_10069,N_8130,N_8654);
nand U10070 (N_10070,N_9110,N_8300);
or U10071 (N_10071,N_9879,N_8545);
xnor U10072 (N_10072,N_9342,N_8765);
nand U10073 (N_10073,N_9172,N_8181);
nand U10074 (N_10074,N_8998,N_8082);
nand U10075 (N_10075,N_9967,N_9022);
and U10076 (N_10076,N_8492,N_8155);
nor U10077 (N_10077,N_8216,N_9721);
nand U10078 (N_10078,N_9508,N_8361);
nand U10079 (N_10079,N_9523,N_8005);
or U10080 (N_10080,N_8556,N_8345);
xor U10081 (N_10081,N_9785,N_8949);
nand U10082 (N_10082,N_8339,N_8600);
nor U10083 (N_10083,N_8873,N_8652);
and U10084 (N_10084,N_8730,N_9966);
or U10085 (N_10085,N_9952,N_9568);
or U10086 (N_10086,N_9125,N_8176);
or U10087 (N_10087,N_8230,N_8021);
nand U10088 (N_10088,N_8774,N_8575);
or U10089 (N_10089,N_9177,N_9204);
nand U10090 (N_10090,N_8656,N_8288);
and U10091 (N_10091,N_9645,N_8137);
and U10092 (N_10092,N_8244,N_9298);
nor U10093 (N_10093,N_9174,N_8441);
and U10094 (N_10094,N_8966,N_8537);
and U10095 (N_10095,N_9908,N_9610);
nor U10096 (N_10096,N_9451,N_9123);
nand U10097 (N_10097,N_9077,N_8067);
and U10098 (N_10098,N_8916,N_9766);
nor U10099 (N_10099,N_9019,N_8740);
nor U10100 (N_10100,N_9944,N_8606);
nand U10101 (N_10101,N_8157,N_8337);
or U10102 (N_10102,N_9823,N_8049);
nor U10103 (N_10103,N_8684,N_9928);
nand U10104 (N_10104,N_8552,N_8052);
nand U10105 (N_10105,N_8024,N_8603);
or U10106 (N_10106,N_9895,N_9395);
nand U10107 (N_10107,N_9789,N_9387);
or U10108 (N_10108,N_8591,N_8479);
and U10109 (N_10109,N_8110,N_9831);
nor U10110 (N_10110,N_8104,N_8593);
xnor U10111 (N_10111,N_9763,N_9992);
nand U10112 (N_10112,N_9408,N_8720);
nor U10113 (N_10113,N_9760,N_9905);
or U10114 (N_10114,N_8679,N_9957);
and U10115 (N_10115,N_9611,N_9556);
xor U10116 (N_10116,N_8876,N_8835);
or U10117 (N_10117,N_9676,N_8753);
or U10118 (N_10118,N_9783,N_8779);
nand U10119 (N_10119,N_8983,N_8105);
and U10120 (N_10120,N_9977,N_9575);
xor U10121 (N_10121,N_9999,N_8256);
nor U10122 (N_10122,N_9802,N_8463);
nor U10123 (N_10123,N_8234,N_8459);
or U10124 (N_10124,N_8078,N_9657);
nand U10125 (N_10125,N_9423,N_9014);
and U10126 (N_10126,N_9564,N_8484);
or U10127 (N_10127,N_9986,N_9881);
nand U10128 (N_10128,N_9279,N_9033);
nand U10129 (N_10129,N_9811,N_9758);
nand U10130 (N_10130,N_8804,N_9127);
and U10131 (N_10131,N_9672,N_8532);
or U10132 (N_10132,N_8750,N_9883);
and U10133 (N_10133,N_8846,N_9026);
xor U10134 (N_10134,N_8311,N_8222);
nor U10135 (N_10135,N_9283,N_8508);
nand U10136 (N_10136,N_8605,N_8102);
and U10137 (N_10137,N_8710,N_8566);
nand U10138 (N_10138,N_8906,N_9420);
nor U10139 (N_10139,N_8536,N_9063);
or U10140 (N_10140,N_9261,N_8385);
and U10141 (N_10141,N_8841,N_9808);
nor U10142 (N_10142,N_8927,N_9713);
nor U10143 (N_10143,N_9477,N_8073);
nor U10144 (N_10144,N_8480,N_9891);
nor U10145 (N_10145,N_9354,N_8123);
or U10146 (N_10146,N_9138,N_8852);
and U10147 (N_10147,N_8335,N_9490);
xor U10148 (N_10148,N_9248,N_9130);
nand U10149 (N_10149,N_8206,N_9414);
xor U10150 (N_10150,N_9532,N_8410);
nor U10151 (N_10151,N_9468,N_8868);
nor U10152 (N_10152,N_8238,N_9500);
and U10153 (N_10153,N_9886,N_8151);
nand U10154 (N_10154,N_8387,N_8871);
and U10155 (N_10155,N_8917,N_8639);
and U10156 (N_10156,N_8121,N_9356);
or U10157 (N_10157,N_9616,N_9059);
nor U10158 (N_10158,N_8970,N_8109);
xor U10159 (N_10159,N_9540,N_9947);
nand U10160 (N_10160,N_8086,N_8296);
and U10161 (N_10161,N_9842,N_9862);
xor U10162 (N_10162,N_9137,N_9853);
nor U10163 (N_10163,N_9179,N_8395);
or U10164 (N_10164,N_9027,N_8364);
nand U10165 (N_10165,N_9045,N_8099);
and U10166 (N_10166,N_9517,N_8574);
nor U10167 (N_10167,N_8760,N_9569);
and U10168 (N_10168,N_9285,N_9371);
and U10169 (N_10169,N_9296,N_9695);
nor U10170 (N_10170,N_9475,N_8360);
and U10171 (N_10171,N_8408,N_9376);
nand U10172 (N_10172,N_9572,N_8167);
nand U10173 (N_10173,N_8735,N_9074);
nand U10174 (N_10174,N_8382,N_8514);
nor U10175 (N_10175,N_9466,N_8269);
nand U10176 (N_10176,N_8636,N_8319);
or U10177 (N_10177,N_8861,N_9360);
and U10178 (N_10178,N_8418,N_9843);
nand U10179 (N_10179,N_8539,N_9410);
or U10180 (N_10180,N_9230,N_9046);
nand U10181 (N_10181,N_8722,N_8996);
nand U10182 (N_10182,N_9561,N_9761);
nor U10183 (N_10183,N_9639,N_8895);
nand U10184 (N_10184,N_9281,N_8659);
xnor U10185 (N_10185,N_9929,N_9768);
nor U10186 (N_10186,N_9698,N_8793);
and U10187 (N_10187,N_9121,N_8678);
nand U10188 (N_10188,N_8451,N_9229);
nand U10189 (N_10189,N_9933,N_8759);
nor U10190 (N_10190,N_8783,N_8404);
and U10191 (N_10191,N_8276,N_8456);
and U10192 (N_10192,N_8405,N_8341);
nand U10193 (N_10193,N_8942,N_9028);
or U10194 (N_10194,N_8303,N_9023);
nand U10195 (N_10195,N_9797,N_9786);
or U10196 (N_10196,N_8941,N_8281);
or U10197 (N_10197,N_8056,N_9227);
or U10198 (N_10198,N_9331,N_9144);
and U10199 (N_10199,N_8796,N_8038);
and U10200 (N_10200,N_8721,N_9953);
nor U10201 (N_10201,N_9193,N_9717);
nand U10202 (N_10202,N_8257,N_8126);
and U10203 (N_10203,N_9921,N_8233);
xnor U10204 (N_10204,N_9772,N_9636);
or U10205 (N_10205,N_8899,N_9963);
nor U10206 (N_10206,N_9813,N_9163);
or U10207 (N_10207,N_8443,N_9497);
nand U10208 (N_10208,N_9827,N_9764);
and U10209 (N_10209,N_9962,N_8320);
nor U10210 (N_10210,N_8840,N_9334);
and U10211 (N_10211,N_9994,N_8587);
nor U10212 (N_10212,N_8589,N_9494);
nor U10213 (N_10213,N_9529,N_9311);
and U10214 (N_10214,N_9080,N_9914);
nand U10215 (N_10215,N_9025,N_8313);
nor U10216 (N_10216,N_9094,N_9543);
nand U10217 (N_10217,N_9112,N_8438);
nand U10218 (N_10218,N_9613,N_8623);
or U10219 (N_10219,N_9218,N_9235);
nand U10220 (N_10220,N_9800,N_9712);
nand U10221 (N_10221,N_9799,N_9264);
and U10222 (N_10222,N_9678,N_9377);
nor U10223 (N_10223,N_8006,N_8100);
nand U10224 (N_10224,N_9277,N_8582);
or U10225 (N_10225,N_9478,N_9780);
or U10226 (N_10226,N_9980,N_8351);
nor U10227 (N_10227,N_8815,N_8950);
xor U10228 (N_10228,N_9159,N_8935);
nor U10229 (N_10229,N_8184,N_9852);
or U10230 (N_10230,N_9051,N_9784);
xor U10231 (N_10231,N_8848,N_9057);
or U10232 (N_10232,N_9140,N_8820);
nand U10233 (N_10233,N_8943,N_9979);
nor U10234 (N_10234,N_8164,N_8144);
xor U10235 (N_10235,N_8663,N_8170);
nor U10236 (N_10236,N_9492,N_9456);
nand U10237 (N_10237,N_8139,N_9859);
nand U10238 (N_10238,N_9788,N_9981);
and U10239 (N_10239,N_9837,N_9079);
nand U10240 (N_10240,N_8106,N_9774);
or U10241 (N_10241,N_8650,N_9520);
nand U10242 (N_10242,N_9486,N_9397);
nand U10243 (N_10243,N_8305,N_8077);
and U10244 (N_10244,N_9591,N_8084);
nor U10245 (N_10245,N_9348,N_8229);
nand U10246 (N_10246,N_8235,N_8207);
and U10247 (N_10247,N_8485,N_9058);
nor U10248 (N_10248,N_8547,N_9208);
or U10249 (N_10249,N_8429,N_9048);
xor U10250 (N_10250,N_8910,N_9113);
and U10251 (N_10251,N_9716,N_8677);
nor U10252 (N_10252,N_8784,N_9688);
and U10253 (N_10253,N_8366,N_9133);
and U10254 (N_10254,N_8565,N_8285);
and U10255 (N_10255,N_8754,N_9782);
or U10256 (N_10256,N_8322,N_8488);
xnor U10257 (N_10257,N_8669,N_8428);
or U10258 (N_10258,N_9732,N_9481);
and U10259 (N_10259,N_9271,N_9171);
xnor U10260 (N_10260,N_8977,N_8008);
and U10261 (N_10261,N_8019,N_9313);
xor U10262 (N_10262,N_9887,N_8128);
and U10263 (N_10263,N_8426,N_9373);
or U10264 (N_10264,N_8780,N_8010);
nand U10265 (N_10265,N_9554,N_9544);
nor U10266 (N_10266,N_8521,N_9906);
nand U10267 (N_10267,N_8041,N_8433);
or U10268 (N_10268,N_9701,N_8023);
nor U10269 (N_10269,N_9352,N_8187);
or U10270 (N_10270,N_8286,N_8746);
xnor U10271 (N_10271,N_9649,N_8930);
nor U10272 (N_10272,N_9555,N_9485);
and U10273 (N_10273,N_8517,N_8057);
or U10274 (N_10274,N_8007,N_9803);
nand U10275 (N_10275,N_8321,N_9590);
and U10276 (N_10276,N_8353,N_9987);
nand U10277 (N_10277,N_8686,N_9625);
xnor U10278 (N_10278,N_9347,N_8262);
and U10279 (N_10279,N_8417,N_9539);
or U10280 (N_10280,N_8424,N_8775);
nand U10281 (N_10281,N_9918,N_9253);
and U10282 (N_10282,N_9320,N_9946);
or U10283 (N_10283,N_8701,N_9156);
nand U10284 (N_10284,N_9875,N_9630);
nand U10285 (N_10285,N_8694,N_9652);
or U10286 (N_10286,N_8132,N_9696);
and U10287 (N_10287,N_9426,N_8847);
nand U10288 (N_10288,N_9441,N_8491);
nor U10289 (N_10289,N_8355,N_8756);
or U10290 (N_10290,N_9017,N_8274);
nor U10291 (N_10291,N_8218,N_9744);
and U10292 (N_10292,N_8020,N_8602);
or U10293 (N_10293,N_8315,N_9375);
nor U10294 (N_10294,N_9927,N_8743);
nand U10295 (N_10295,N_8114,N_9437);
nand U10296 (N_10296,N_9359,N_8690);
xor U10297 (N_10297,N_8612,N_8088);
nor U10298 (N_10298,N_8246,N_8211);
nand U10299 (N_10299,N_9850,N_8912);
nor U10300 (N_10300,N_8833,N_8245);
nor U10301 (N_10301,N_9909,N_8432);
xnor U10302 (N_10302,N_9793,N_8280);
nor U10303 (N_10303,N_8069,N_8597);
and U10304 (N_10304,N_9824,N_8634);
and U10305 (N_10305,N_8250,N_8548);
or U10306 (N_10306,N_9038,N_8383);
or U10307 (N_10307,N_8853,N_9935);
xor U10308 (N_10308,N_8261,N_9646);
nand U10309 (N_10309,N_9065,N_8791);
or U10310 (N_10310,N_8001,N_8881);
nand U10311 (N_10311,N_9241,N_8995);
nand U10312 (N_10312,N_8658,N_9270);
or U10313 (N_10313,N_8452,N_8357);
and U10314 (N_10314,N_8987,N_8431);
or U10315 (N_10315,N_8131,N_8503);
or U10316 (N_10316,N_9162,N_9995);
and U10317 (N_10317,N_8440,N_8919);
or U10318 (N_10318,N_8975,N_8558);
and U10319 (N_10319,N_9286,N_9629);
nand U10320 (N_10320,N_8732,N_8772);
nand U10321 (N_10321,N_9366,N_8299);
nand U10322 (N_10322,N_8519,N_9617);
nand U10323 (N_10323,N_8688,N_8516);
nor U10324 (N_10324,N_8778,N_9226);
nand U10325 (N_10325,N_9974,N_8204);
or U10326 (N_10326,N_9409,N_8394);
and U10327 (N_10327,N_8925,N_8034);
and U10328 (N_10328,N_8118,N_8079);
nor U10329 (N_10329,N_9593,N_8146);
nand U10330 (N_10330,N_9249,N_8878);
nand U10331 (N_10331,N_9432,N_8338);
or U10332 (N_10332,N_9693,N_9391);
or U10333 (N_10333,N_9463,N_8427);
and U10334 (N_10334,N_8651,N_9009);
nor U10335 (N_10335,N_8270,N_9641);
and U10336 (N_10336,N_8186,N_8924);
nor U10337 (N_10337,N_9724,N_9413);
nand U10338 (N_10338,N_9637,N_8553);
xor U10339 (N_10339,N_8107,N_9430);
xor U10340 (N_10340,N_8398,N_9679);
nor U10341 (N_10341,N_8009,N_9147);
and U10342 (N_10342,N_9299,N_9495);
or U10343 (N_10343,N_8854,N_9644);
nor U10344 (N_10344,N_9658,N_8900);
or U10345 (N_10345,N_8255,N_8407);
xnor U10346 (N_10346,N_8371,N_9247);
nor U10347 (N_10347,N_9779,N_8501);
or U10348 (N_10348,N_8568,N_9493);
xnor U10349 (N_10349,N_8716,N_8450);
or U10350 (N_10350,N_9663,N_8807);
nor U10351 (N_10351,N_8051,N_9706);
nand U10352 (N_10352,N_8115,N_9815);
nand U10353 (N_10353,N_9107,N_8972);
nand U10354 (N_10354,N_8253,N_8369);
nor U10355 (N_10355,N_9343,N_8318);
and U10356 (N_10356,N_9627,N_8555);
nor U10357 (N_10357,N_8523,N_9002);
and U10358 (N_10358,N_9075,N_9052);
or U10359 (N_10359,N_8857,N_8757);
nand U10360 (N_10360,N_8787,N_8546);
or U10361 (N_10361,N_9985,N_8411);
or U10362 (N_10362,N_9405,N_8557);
or U10363 (N_10363,N_8609,N_8201);
nor U10364 (N_10364,N_9422,N_8055);
or U10365 (N_10365,N_9207,N_8786);
nand U10366 (N_10366,N_9438,N_9118);
or U10367 (N_10367,N_8290,N_9982);
and U10368 (N_10368,N_9234,N_8448);
nor U10369 (N_10369,N_9584,N_8435);
nor U10370 (N_10370,N_8048,N_8015);
and U10371 (N_10371,N_9445,N_8097);
or U10372 (N_10372,N_8346,N_8692);
and U10373 (N_10373,N_9665,N_9257);
nand U10374 (N_10374,N_8535,N_8192);
or U10375 (N_10375,N_8168,N_8018);
and U10376 (N_10376,N_9361,N_9911);
nor U10377 (N_10377,N_8724,N_9469);
or U10378 (N_10378,N_8141,N_8837);
nor U10379 (N_10379,N_8241,N_8742);
nand U10380 (N_10380,N_8209,N_8162);
or U10381 (N_10381,N_9381,N_8821);
nor U10382 (N_10382,N_9704,N_9379);
xor U10383 (N_10383,N_9898,N_8607);
nand U10384 (N_10384,N_8089,N_9727);
or U10385 (N_10385,N_8227,N_8909);
or U10386 (N_10386,N_8664,N_8037);
and U10387 (N_10387,N_9700,N_9511);
nor U10388 (N_10388,N_9551,N_9903);
nor U10389 (N_10389,N_8326,N_8892);
nor U10390 (N_10390,N_8402,N_9276);
or U10391 (N_10391,N_9835,N_9514);
nor U10392 (N_10392,N_9925,N_8190);
nand U10393 (N_10393,N_9690,N_8709);
or U10394 (N_10394,N_8240,N_9588);
nand U10395 (N_10395,N_8884,N_8430);
and U10396 (N_10396,N_8135,N_8819);
xor U10397 (N_10397,N_9503,N_8094);
or U10398 (N_10398,N_9563,N_8348);
nor U10399 (N_10399,N_8344,N_8777);
and U10400 (N_10400,N_9444,N_9740);
nor U10401 (N_10401,N_9145,N_9450);
and U10402 (N_10402,N_9301,N_8153);
nor U10403 (N_10403,N_9015,N_9128);
nand U10404 (N_10404,N_8687,N_9845);
and U10405 (N_10405,N_9804,N_8482);
nor U10406 (N_10406,N_8367,N_8862);
or U10407 (N_10407,N_9734,N_9369);
and U10408 (N_10408,N_9836,N_8472);
nor U10409 (N_10409,N_8028,N_9245);
or U10410 (N_10410,N_8763,N_9817);
or U10411 (N_10411,N_9192,N_8812);
or U10412 (N_10412,N_8505,N_9238);
nand U10413 (N_10413,N_9501,N_9305);
nand U10414 (N_10414,N_9686,N_8328);
and U10415 (N_10415,N_9007,N_8000);
and U10416 (N_10416,N_8495,N_8570);
or U10417 (N_10417,N_8622,N_9039);
nor U10418 (N_10418,N_8208,N_8766);
or U10419 (N_10419,N_8239,N_8932);
and U10420 (N_10420,N_9188,N_9765);
and U10421 (N_10421,N_8386,N_9607);
and U10422 (N_10422,N_9560,N_8544);
nand U10423 (N_10423,N_9233,N_9323);
and U10424 (N_10424,N_9976,N_8843);
xor U10425 (N_10425,N_8254,N_9525);
nand U10426 (N_10426,N_8631,N_9090);
nand U10427 (N_10427,N_9383,N_8493);
xnor U10428 (N_10428,N_9435,N_9295);
nand U10429 (N_10429,N_9718,N_9129);
nor U10430 (N_10430,N_8327,N_9938);
or U10431 (N_10431,N_8827,N_8272);
nand U10432 (N_10432,N_9589,N_9904);
nand U10433 (N_10433,N_8611,N_8231);
and U10434 (N_10434,N_8524,N_8188);
or U10435 (N_10435,N_9060,N_8683);
or U10436 (N_10436,N_8989,N_9858);
and U10437 (N_10437,N_8583,N_8666);
or U10438 (N_10438,N_9655,N_8236);
nor U10439 (N_10439,N_8436,N_8896);
xnor U10440 (N_10440,N_9189,N_9930);
and U10441 (N_10441,N_8380,N_8956);
nor U10442 (N_10442,N_8053,N_8112);
and U10443 (N_10443,N_9205,N_9198);
xor U10444 (N_10444,N_9834,N_8907);
nand U10445 (N_10445,N_9306,N_9526);
nand U10446 (N_10446,N_8798,N_9223);
or U10447 (N_10447,N_9459,N_9703);
or U10448 (N_10448,N_8180,N_9567);
or U10449 (N_10449,N_9132,N_8074);
nand U10450 (N_10450,N_9175,N_8044);
nor U10451 (N_10451,N_8711,N_8414);
or U10452 (N_10452,N_8646,N_8210);
nor U10453 (N_10453,N_8071,N_9728);
nor U10454 (N_10454,N_8704,N_8745);
xor U10455 (N_10455,N_9689,N_8226);
xor U10456 (N_10456,N_8586,N_8595);
nor U10457 (N_10457,N_9183,N_9993);
xor U10458 (N_10458,N_9884,N_9510);
nand U10459 (N_10459,N_9282,N_9416);
xor U10460 (N_10460,N_9626,N_9341);
nor U10461 (N_10461,N_9328,N_9220);
and U10462 (N_10462,N_9622,N_8585);
or U10463 (N_10463,N_9338,N_8033);
nor U10464 (N_10464,N_9515,N_9832);
nand U10465 (N_10465,N_8461,N_9290);
and U10466 (N_10466,N_8422,N_8567);
nand U10467 (N_10467,N_8620,N_9874);
nor U10468 (N_10468,N_9384,N_8946);
or U10469 (N_10469,N_8026,N_9603);
or U10470 (N_10470,N_9085,N_9329);
nor U10471 (N_10471,N_8969,N_8391);
nor U10472 (N_10472,N_8036,N_8984);
nor U10473 (N_10473,N_8737,N_9458);
nand U10474 (N_10474,N_9934,N_9767);
nor U10475 (N_10475,N_8196,N_8771);
nor U10476 (N_10476,N_9651,N_9237);
nand U10477 (N_10477,N_9425,N_9304);
nor U10478 (N_10478,N_9961,N_9134);
nand U10479 (N_10479,N_9418,N_9008);
or U10480 (N_10480,N_8551,N_9098);
nand U10481 (N_10481,N_8668,N_8808);
nor U10482 (N_10482,N_8992,N_8867);
or U10483 (N_10483,N_8403,N_9166);
nor U10484 (N_10484,N_8799,N_8083);
or U10485 (N_10485,N_9615,N_9096);
nand U10486 (N_10486,N_8506,N_9239);
nor U10487 (N_10487,N_9535,N_8062);
nor U10488 (N_10488,N_8166,N_9926);
nor U10489 (N_10489,N_8279,N_8309);
nand U10490 (N_10490,N_9321,N_9365);
xnor U10491 (N_10491,N_8193,N_9103);
or U10492 (N_10492,N_9792,N_8502);
nand U10493 (N_10493,N_9392,N_9573);
or U10494 (N_10494,N_8581,N_8260);
nand U10495 (N_10495,N_8076,N_8149);
nor U10496 (N_10496,N_8093,N_8629);
xor U10497 (N_10497,N_9541,N_9604);
nor U10498 (N_10498,N_8965,N_9880);
or U10499 (N_10499,N_9889,N_9412);
nor U10500 (N_10500,N_8671,N_8836);
nor U10501 (N_10501,N_8295,N_8674);
and U10502 (N_10502,N_8951,N_9200);
nand U10503 (N_10503,N_9116,N_8706);
nand U10504 (N_10504,N_9656,N_9566);
nor U10505 (N_10505,N_8973,N_8696);
or U10506 (N_10506,N_8043,N_9505);
nand U10507 (N_10507,N_9442,N_9585);
nor U10508 (N_10508,N_9970,N_8013);
or U10509 (N_10509,N_9243,N_9099);
and U10510 (N_10510,N_8165,N_9355);
nor U10511 (N_10511,N_8904,N_9291);
nand U10512 (N_10512,N_9246,N_8259);
nand U10513 (N_10513,N_8194,N_9664);
or U10514 (N_10514,N_8554,N_8571);
or U10515 (N_10515,N_9833,N_9221);
and U10516 (N_10516,N_9095,N_8813);
nand U10517 (N_10517,N_8676,N_8381);
nand U10518 (N_10518,N_8200,N_9968);
or U10519 (N_10519,N_9794,N_9809);
nor U10520 (N_10520,N_9093,N_8662);
xor U10521 (N_10521,N_9807,N_9733);
or U10522 (N_10522,N_9258,N_8462);
xnor U10523 (N_10523,N_8985,N_8726);
or U10524 (N_10524,N_9109,N_9901);
and U10525 (N_10525,N_9460,N_8247);
or U10526 (N_10526,N_8275,N_8393);
xor U10527 (N_10527,N_9310,N_9349);
or U10528 (N_10528,N_8362,N_8865);
xor U10529 (N_10529,N_9710,N_8824);
and U10530 (N_10530,N_9870,N_9344);
xor U10531 (N_10531,N_8834,N_9565);
or U10532 (N_10532,N_8070,N_8042);
nor U10533 (N_10533,N_9989,N_8522);
or U10534 (N_10534,N_9484,N_9729);
or U10535 (N_10535,N_8027,N_9840);
nor U10536 (N_10536,N_9991,N_9576);
nand U10537 (N_10537,N_8370,N_9671);
nor U10538 (N_10538,N_9920,N_8598);
or U10539 (N_10539,N_9762,N_9771);
and U10540 (N_10540,N_8755,N_8509);
nand U10541 (N_10541,N_9070,N_9294);
nand U10542 (N_10542,N_9149,N_8660);
nor U10543 (N_10543,N_9066,N_8481);
nor U10544 (N_10544,N_8147,N_9940);
nor U10545 (N_10545,N_9602,N_9043);
xor U10546 (N_10546,N_9393,N_9292);
nand U10547 (N_10547,N_8838,N_9297);
xor U10548 (N_10548,N_8399,N_8822);
and U10549 (N_10549,N_8359,N_8872);
nand U10550 (N_10550,N_9050,N_8205);
or U10551 (N_10551,N_9433,N_8714);
and U10552 (N_10552,N_9574,N_8047);
nand U10553 (N_10553,N_8897,N_8752);
nand U10554 (N_10554,N_8308,N_8974);
or U10555 (N_10555,N_9709,N_8016);
nor U10556 (N_10556,N_9582,N_8050);
and U10557 (N_10557,N_8372,N_8185);
nor U10558 (N_10558,N_9150,N_9333);
or U10559 (N_10559,N_9857,N_9819);
or U10560 (N_10560,N_8171,N_9708);
nand U10561 (N_10561,N_9446,N_9491);
xnor U10562 (N_10562,N_9773,N_8526);
or U10563 (N_10563,N_9669,N_8845);
or U10564 (N_10564,N_8022,N_8947);
or U10565 (N_10565,N_8529,N_8641);
nor U10566 (N_10566,N_8080,N_8343);
or U10567 (N_10567,N_9846,N_8446);
and U10568 (N_10568,N_9326,N_8738);
nand U10569 (N_10569,N_8449,N_9368);
and U10570 (N_10570,N_8915,N_8921);
or U10571 (N_10571,N_8090,N_8979);
and U10572 (N_10572,N_8352,N_8850);
and U10573 (N_10573,N_8844,N_8292);
and U10574 (N_10574,N_8487,N_9869);
nand U10575 (N_10575,N_8439,N_8729);
xnor U10576 (N_10576,N_9984,N_9579);
nor U10577 (N_10577,N_8619,N_9830);
or U10578 (N_10578,N_9062,N_9251);
nor U10579 (N_10579,N_9597,N_9715);
nor U10580 (N_10580,N_8616,N_9364);
nor U10581 (N_10581,N_8849,N_9756);
or U10582 (N_10582,N_9752,N_9860);
and U10583 (N_10583,N_9231,N_9978);
or U10584 (N_10584,N_8954,N_8776);
and U10585 (N_10585,N_9083,N_9751);
nor U10586 (N_10586,N_9262,N_8792);
nand U10587 (N_10587,N_9169,N_8938);
and U10588 (N_10588,N_8767,N_9996);
and U10589 (N_10589,N_8068,N_8826);
nand U10590 (N_10590,N_9164,N_8797);
nand U10591 (N_10591,N_8478,N_8761);
or U10592 (N_10592,N_8810,N_8948);
nor U10593 (N_10593,N_9769,N_9796);
and U10594 (N_10594,N_9201,N_8643);
nor U10595 (N_10595,N_9217,N_9191);
xnor U10596 (N_10596,N_8271,N_8788);
nand U10597 (N_10597,N_9424,N_9273);
nor U10598 (N_10598,N_9668,N_9866);
nand U10599 (N_10599,N_9778,N_9049);
nor U10600 (N_10600,N_9449,N_8356);
and U10601 (N_10601,N_8374,N_8874);
nand U10602 (N_10602,N_8278,N_9838);
and U10603 (N_10603,N_8731,N_9142);
or U10604 (N_10604,N_9548,N_9315);
nor U10605 (N_10605,N_9631,N_8415);
nand U10606 (N_10606,N_8699,N_8569);
nor U10607 (N_10607,N_8045,N_9370);
nor U10608 (N_10608,N_9650,N_9346);
nor U10609 (N_10609,N_9960,N_9101);
nand U10610 (N_10610,N_9464,N_8202);
and U10611 (N_10611,N_9667,N_8990);
nand U10612 (N_10612,N_8717,N_9448);
nand U10613 (N_10613,N_9399,N_9224);
nand U10614 (N_10614,N_8423,N_8842);
nor U10615 (N_10615,N_9136,N_8301);
and U10616 (N_10616,N_9115,N_9126);
or U10617 (N_10617,N_9440,N_8773);
or U10618 (N_10618,N_8626,N_8425);
xor U10619 (N_10619,N_8101,N_9473);
nor U10620 (N_10620,N_9470,N_9798);
and U10621 (N_10621,N_8875,N_9878);
or U10622 (N_10622,N_9907,N_8098);
nand U10623 (N_10623,N_9882,N_8997);
and U10624 (N_10624,N_9632,N_9010);
or U10625 (N_10625,N_8091,N_9902);
and U10626 (N_10626,N_9087,N_9351);
or U10627 (N_10627,N_8528,N_8111);
nor U10628 (N_10628,N_8739,N_9244);
nor U10629 (N_10629,N_9064,N_8940);
nand U10630 (N_10630,N_8217,N_9211);
and U10631 (N_10631,N_8624,N_9599);
nor U10632 (N_10632,N_9499,N_8511);
or U10633 (N_10633,N_8510,N_8373);
and U10634 (N_10634,N_9182,N_8851);
xor U10635 (N_10635,N_8143,N_8025);
xor U10636 (N_10636,N_9474,N_9436);
and U10637 (N_10637,N_8725,N_8647);
or U10638 (N_10638,N_9972,N_9685);
nor U10639 (N_10639,N_9922,N_9011);
nor U10640 (N_10640,N_9362,N_8794);
nor U10641 (N_10641,N_9741,N_9997);
nor U10642 (N_10642,N_9628,N_8455);
or U10643 (N_10643,N_9367,N_8312);
nand U10644 (N_10644,N_8465,N_9759);
or U10645 (N_10645,N_9820,N_9462);
nand U10646 (N_10646,N_9702,N_8534);
and U10647 (N_10647,N_9350,N_9000);
or U10648 (N_10648,N_8142,N_8902);
nand U10649 (N_10649,N_9124,N_9791);
nor U10650 (N_10650,N_9106,N_9941);
nand U10651 (N_10651,N_8499,N_9849);
and U10652 (N_10652,N_8284,N_8961);
xnor U10653 (N_10653,N_8014,N_9102);
nand U10654 (N_10654,N_8060,N_8476);
nor U10655 (N_10655,N_8434,N_8809);
nand U10656 (N_10656,N_9053,N_9512);
nor U10657 (N_10657,N_8003,N_9047);
and U10658 (N_10658,N_9775,N_8474);
nor U10659 (N_10659,N_8648,N_8713);
and U10660 (N_10660,N_9202,N_9919);
or U10661 (N_10661,N_9661,N_9814);
and U10662 (N_10662,N_8273,N_8538);
nor U10663 (N_10663,N_8507,N_9104);
and U10664 (N_10664,N_8665,N_9691);
or U10665 (N_10665,N_8831,N_9951);
xnor U10666 (N_10666,N_8420,N_9146);
nand U10667 (N_10667,N_8032,N_8175);
nand U10668 (N_10668,N_8458,N_8213);
nor U10669 (N_10669,N_8653,N_8957);
nor U10670 (N_10670,N_9078,N_8573);
and U10671 (N_10671,N_8630,N_9398);
nand U10672 (N_10672,N_9680,N_9916);
or U10673 (N_10673,N_9923,N_9673);
and U10674 (N_10674,N_8830,N_9161);
or U10675 (N_10675,N_8963,N_8058);
and U10676 (N_10676,N_9097,N_9948);
nor U10677 (N_10677,N_8596,N_8453);
or U10678 (N_10678,N_9452,N_8727);
xor U10679 (N_10679,N_9403,N_9917);
nor U10680 (N_10680,N_8560,N_8885);
nand U10681 (N_10681,N_9461,N_9594);
nor U10682 (N_10682,N_8733,N_9844);
or U10683 (N_10683,N_9314,N_8470);
nor U10684 (N_10684,N_8504,N_9380);
nand U10685 (N_10685,N_9417,N_8294);
nand U10686 (N_10686,N_8442,N_9421);
or U10687 (N_10687,N_8182,N_8264);
and U10688 (N_10688,N_9533,N_8803);
nand U10689 (N_10689,N_9431,N_8823);
and U10690 (N_10690,N_8249,N_8649);
nand U10691 (N_10691,N_9472,N_8922);
and U10692 (N_10692,N_9583,N_8723);
or U10693 (N_10693,N_8599,N_8498);
nand U10694 (N_10694,N_9197,N_8030);
or U10695 (N_10695,N_8197,N_9893);
and U10696 (N_10696,N_8901,N_8937);
and U10697 (N_10697,N_9847,N_9003);
and U10698 (N_10698,N_8031,N_8012);
nand U10699 (N_10699,N_8805,N_9971);
and U10700 (N_10700,N_8981,N_8297);
xor U10701 (N_10701,N_8400,N_8002);
nand U10702 (N_10702,N_9897,N_8122);
and U10703 (N_10703,N_9031,N_8886);
nand U10704 (N_10704,N_8342,N_8475);
nand U10705 (N_10705,N_8697,N_9120);
or U10706 (N_10706,N_8323,N_9677);
or U10707 (N_10707,N_9284,N_8252);
nor U10708 (N_10708,N_9562,N_8316);
and U10709 (N_10709,N_8445,N_9318);
nand U10710 (N_10710,N_8768,N_9670);
nand U10711 (N_10711,N_8929,N_9581);
xor U10712 (N_10712,N_9801,N_9945);
and U10713 (N_10713,N_8689,N_8156);
nor U10714 (N_10714,N_8336,N_9939);
nor U10715 (N_10715,N_8419,N_8460);
and U10716 (N_10716,N_8959,N_9816);
nor U10717 (N_10717,N_9552,N_8734);
and U10718 (N_10718,N_9694,N_9666);
or U10719 (N_10719,N_8707,N_9363);
and U10720 (N_10720,N_8258,N_9580);
xor U10721 (N_10721,N_9293,N_8471);
or U10722 (N_10722,N_9692,N_9073);
nand U10723 (N_10723,N_9072,N_8512);
or U10724 (N_10724,N_9212,N_8944);
and U10725 (N_10725,N_9730,N_9404);
nor U10726 (N_10726,N_9634,N_9682);
and U10727 (N_10727,N_9067,N_8718);
nand U10728 (N_10728,N_9267,N_9018);
nand U10729 (N_10729,N_8855,N_8818);
nor U10730 (N_10730,N_8863,N_8693);
or U10731 (N_10731,N_8265,N_9558);
or U10732 (N_10732,N_8263,N_8066);
or U10733 (N_10733,N_8409,N_9983);
nor U10734 (N_10734,N_8800,N_9578);
nand U10735 (N_10735,N_9143,N_9746);
nand U10736 (N_10736,N_8040,N_9170);
and U10737 (N_10737,N_8749,N_8172);
or U10738 (N_10738,N_9044,N_8945);
or U10739 (N_10739,N_9148,N_9871);
xnor U10740 (N_10740,N_9937,N_8349);
xnor U10741 (N_10741,N_9309,N_8215);
or U10742 (N_10742,N_9549,N_9119);
nor U10743 (N_10743,N_9571,N_8980);
and U10744 (N_10744,N_8869,N_9822);
nand U10745 (N_10745,N_8673,N_8968);
nor U10746 (N_10746,N_9624,N_9899);
and U10747 (N_10747,N_8982,N_9810);
and U10748 (N_10748,N_9184,N_9012);
and U10749 (N_10749,N_8173,N_9034);
nor U10750 (N_10750,N_9742,N_9757);
and U10751 (N_10751,N_9020,N_8454);
nand U10752 (N_10752,N_9402,N_9605);
or U10753 (N_10753,N_8046,N_8406);
nor U10754 (N_10754,N_9252,N_9949);
xnor U10755 (N_10755,N_9389,N_9542);
or U10756 (N_10756,N_9165,N_8183);
nand U10757 (N_10757,N_8635,N_9086);
or U10758 (N_10758,N_9269,N_8392);
and U10759 (N_10759,N_8563,N_9419);
or U10760 (N_10760,N_9587,N_8177);
and U10761 (N_10761,N_8133,N_9705);
nor U10762 (N_10762,N_9973,N_9805);
and U10763 (N_10763,N_8802,N_9821);
xor U10764 (N_10764,N_9738,N_8579);
nor U10765 (N_10765,N_9158,N_9187);
nand U10766 (N_10766,N_8816,N_9675);
nor U10767 (N_10767,N_8081,N_8712);
nor U10768 (N_10768,N_8978,N_8447);
nor U10769 (N_10769,N_9454,N_8870);
nand U10770 (N_10770,N_9518,N_9139);
xnor U10771 (N_10771,N_9330,N_8604);
or U10772 (N_10772,N_8304,N_9055);
or U10773 (N_10773,N_9900,N_8561);
and U10774 (N_10774,N_9723,N_9648);
nand U10775 (N_10775,N_8859,N_9910);
and U10776 (N_10776,N_8741,N_8103);
or U10777 (N_10777,N_9737,N_9482);
or U10778 (N_10778,N_9592,N_9339);
and U10779 (N_10779,N_8543,N_9242);
and U10780 (N_10780,N_8914,N_8129);
nor U10781 (N_10781,N_9776,N_8789);
and U10782 (N_10782,N_9839,N_8251);
or U10783 (N_10783,N_9965,N_9178);
and U10784 (N_10784,N_9557,N_8333);
or U10785 (N_10785,N_8655,N_9105);
nand U10786 (N_10786,N_9890,N_9483);
and U10787 (N_10787,N_8814,N_8388);
or U10788 (N_10788,N_9640,N_8150);
nor U10789 (N_10789,N_9071,N_9633);
and U10790 (N_10790,N_8054,N_8469);
nand U10791 (N_10791,N_8317,N_8298);
nor U10792 (N_10792,N_8702,N_8087);
nor U10793 (N_10793,N_8883,N_8594);
xor U10794 (N_10794,N_8334,N_8762);
nand U10795 (N_10795,N_9005,N_9618);
xor U10796 (N_10796,N_8437,N_9595);
nor U10797 (N_10797,N_9606,N_9894);
nor U10798 (N_10798,N_9553,N_9479);
and U10799 (N_10799,N_9209,N_9795);
and U10800 (N_10800,N_8243,N_8124);
nand U10801 (N_10801,N_9586,N_8293);
nand U10802 (N_10802,N_9457,N_9707);
and U10803 (N_10803,N_8986,N_9240);
nand U10804 (N_10804,N_8125,N_9988);
or U10805 (N_10805,N_9082,N_9004);
nand U10806 (N_10806,N_9037,N_9340);
and U10807 (N_10807,N_8728,N_9598);
or U10808 (N_10808,N_8061,N_8747);
nor U10809 (N_10809,N_9131,N_9826);
nor U10810 (N_10810,N_8879,N_9825);
or U10811 (N_10811,N_9215,N_8119);
or U10812 (N_10812,N_9194,N_9855);
and U10813 (N_10813,N_9851,N_8282);
nand U10814 (N_10814,N_8939,N_8490);
nand U10815 (N_10815,N_9620,N_8203);
or U10816 (N_10816,N_9868,N_9195);
or U10817 (N_10817,N_8578,N_9275);
nand U10818 (N_10818,N_8513,N_8220);
or U10819 (N_10819,N_8127,N_8541);
and U10820 (N_10820,N_9942,N_8039);
nand U10821 (N_10821,N_9400,N_9069);
nand U10822 (N_10822,N_9537,N_9272);
or U10823 (N_10823,N_8117,N_8199);
nor U10824 (N_10824,N_8267,N_8681);
or U10825 (N_10825,N_9117,N_9108);
and U10826 (N_10826,N_9638,N_9006);
or U10827 (N_10827,N_9396,N_8913);
and U10828 (N_10828,N_9635,N_8988);
xnor U10829 (N_10829,N_8324,N_9681);
or U10830 (N_10830,N_8645,N_8179);
or U10831 (N_10831,N_9660,N_9029);
nor U10832 (N_10832,N_9042,N_9714);
nand U10833 (N_10833,N_8379,N_9527);
nand U10834 (N_10834,N_9280,N_9092);
or U10835 (N_10835,N_9335,N_9091);
xor U10836 (N_10836,N_8223,N_8332);
and U10837 (N_10837,N_8811,N_8638);
or U10838 (N_10838,N_8219,N_8891);
or U10839 (N_10839,N_9061,N_9496);
nor U10840 (N_10840,N_9185,N_9739);
or U10841 (N_10841,N_8580,N_8960);
nand U10842 (N_10842,N_9111,N_8903);
nor U10843 (N_10843,N_8483,N_9931);
or U10844 (N_10844,N_9506,N_9711);
and U10845 (N_10845,N_8214,N_9250);
nand U10846 (N_10846,N_9203,N_9325);
or U10847 (N_10847,N_9829,N_8991);
or U10848 (N_10848,N_9308,N_9480);
and U10849 (N_10849,N_8839,N_8667);
nor U10850 (N_10850,N_8242,N_9256);
or U10851 (N_10851,N_9943,N_8494);
or U10852 (N_10852,N_9266,N_9538);
xor U10853 (N_10853,N_8614,N_9336);
and U10854 (N_10854,N_9577,N_8542);
or U10855 (N_10855,N_8590,N_9749);
nor U10856 (N_10856,N_8159,N_8953);
xnor U10857 (N_10857,N_9743,N_8134);
nor U10858 (N_10858,N_8923,N_9302);
xnor U10859 (N_10859,N_9068,N_8152);
xnor U10860 (N_10860,N_8306,N_9219);
nand U10861 (N_10861,N_9385,N_8350);
nor U10862 (N_10862,N_8911,N_8889);
and U10863 (N_10863,N_8468,N_8703);
xor U10864 (N_10864,N_9378,N_8163);
nor U10865 (N_10865,N_8825,N_8189);
or U10866 (N_10866,N_9114,N_8368);
nand U10867 (N_10867,N_8232,N_8577);
nand U10868 (N_10868,N_9662,N_9522);
xnor U10869 (N_10869,N_8675,N_9056);
nand U10870 (N_10870,N_9547,N_9001);
and U10871 (N_10871,N_9674,N_9225);
nand U10872 (N_10872,N_9596,N_8486);
nor U10873 (N_10873,N_8397,N_9429);
nand U10874 (N_10874,N_9750,N_8017);
and U10875 (N_10875,N_8195,N_8955);
nor U10876 (N_10876,N_9337,N_9601);
nor U10877 (N_10877,N_9777,N_9502);
and U10878 (N_10878,N_8363,N_8325);
nand U10879 (N_10879,N_9841,N_9975);
and U10880 (N_10880,N_8628,N_8059);
or U10881 (N_10881,N_9173,N_9382);
nor U10882 (N_10882,N_9719,N_9322);
or U10883 (N_10883,N_8212,N_9912);
and U10884 (N_10884,N_8518,N_9088);
nor U10885 (N_10885,N_8828,N_8064);
xor U10886 (N_10886,N_9190,N_9726);
nand U10887 (N_10887,N_8790,N_8615);
nor U10888 (N_10888,N_8004,N_9394);
nand U10889 (N_10889,N_9612,N_9041);
xnor U10890 (N_10890,N_8531,N_8365);
or U10891 (N_10891,N_8354,N_9528);
nand U10892 (N_10892,N_9154,N_8289);
nand U10893 (N_10893,N_9265,N_9358);
or U10894 (N_10894,N_8549,N_9885);
xnor U10895 (N_10895,N_9507,N_9642);
and U10896 (N_10896,N_8113,N_9213);
nor U10897 (N_10897,N_9754,N_8877);
or U10898 (N_10898,N_8967,N_9609);
and U10899 (N_10899,N_9550,N_9254);
nand U10900 (N_10900,N_8618,N_8625);
nor U10901 (N_10901,N_9312,N_8228);
nor U10902 (N_10902,N_9030,N_9181);
and U10903 (N_10903,N_9214,N_9932);
xnor U10904 (N_10904,N_8657,N_9054);
or U10905 (N_10905,N_8829,N_8145);
nor U10906 (N_10906,N_9415,N_8515);
nor U10907 (N_10907,N_9697,N_9206);
or U10908 (N_10908,N_8936,N_8744);
nand U10909 (N_10909,N_8613,N_8527);
or U10910 (N_10910,N_9084,N_8806);
nor U10911 (N_10911,N_9089,N_9504);
nand U10912 (N_10912,N_8029,N_9289);
and U10913 (N_10913,N_8644,N_9155);
or U10914 (N_10914,N_8610,N_8237);
and U10915 (N_10915,N_9021,N_9687);
xor U10916 (N_10916,N_9465,N_8933);
nor U10917 (N_10917,N_9372,N_9954);
or U10918 (N_10918,N_8072,N_8378);
and U10919 (N_10919,N_9781,N_8928);
nor U10920 (N_10920,N_9828,N_9720);
and U10921 (N_10921,N_8864,N_8758);
and U10922 (N_10922,N_9877,N_8856);
nand U10923 (N_10923,N_8715,N_8291);
or U10924 (N_10924,N_9872,N_8801);
nor U10925 (N_10925,N_9731,N_8882);
xnor U10926 (N_10926,N_8905,N_8500);
nand U10927 (N_10927,N_8550,N_9186);
and U10928 (N_10928,N_8592,N_9263);
and U10929 (N_10929,N_9160,N_8473);
and U10930 (N_10930,N_9151,N_8174);
or U10931 (N_10931,N_8178,N_9406);
nand U10932 (N_10932,N_8489,N_9748);
and U10933 (N_10933,N_9998,N_9259);
xor U10934 (N_10934,N_9453,N_9888);
or U10935 (N_10935,N_8719,N_8994);
and U10936 (N_10936,N_8314,N_9725);
xnor U10937 (N_10937,N_8302,N_8958);
nor U10938 (N_10938,N_8095,N_9345);
nor U10939 (N_10939,N_8562,N_9955);
and U10940 (N_10940,N_8329,N_8221);
or U10941 (N_10941,N_8695,N_9790);
xnor U10942 (N_10942,N_9040,N_8920);
nand U10943 (N_10943,N_8085,N_9255);
and U10944 (N_10944,N_9035,N_8138);
xnor U10945 (N_10945,N_9513,N_9317);
nor U10946 (N_10946,N_9141,N_9467);
nor U10947 (N_10947,N_9608,N_9643);
nor U10948 (N_10948,N_9316,N_8108);
nor U10949 (N_10949,N_8672,N_9659);
xor U10950 (N_10950,N_8751,N_8698);
nand U10951 (N_10951,N_9407,N_8277);
or U10952 (N_10952,N_8971,N_9924);
or U10953 (N_10953,N_8540,N_9969);
or U10954 (N_10954,N_9873,N_8621);
nand U10955 (N_10955,N_9135,N_9519);
nand U10956 (N_10956,N_8340,N_8412);
nor U10957 (N_10957,N_9956,N_9770);
nor U10958 (N_10958,N_8191,N_9327);
or U10959 (N_10959,N_8375,N_9812);
or U10960 (N_10960,N_8401,N_9848);
xor U10961 (N_10961,N_8782,N_9303);
or U10962 (N_10962,N_9288,N_9950);
and U10963 (N_10963,N_8283,N_8467);
and U10964 (N_10964,N_9990,N_8608);
and U10965 (N_10965,N_9546,N_8116);
xnor U10966 (N_10966,N_9896,N_9287);
nor U10967 (N_10967,N_9081,N_9736);
or U10968 (N_10968,N_8993,N_8893);
or U10969 (N_10969,N_9411,N_8035);
nand U10970 (N_10970,N_9076,N_9278);
nand U10971 (N_10971,N_9427,N_9401);
or U10972 (N_10972,N_9489,N_9964);
or U10973 (N_10973,N_9684,N_8860);
or U10974 (N_10974,N_8120,N_8161);
nor U10975 (N_10975,N_9536,N_9388);
nand U10976 (N_10976,N_9753,N_8533);
nor U10977 (N_10977,N_8588,N_9516);
and U10978 (N_10978,N_8770,N_8224);
nor U10979 (N_10979,N_9936,N_9434);
xor U10980 (N_10980,N_9122,N_8330);
and U10981 (N_10981,N_8530,N_8670);
and U10982 (N_10982,N_8880,N_9268);
nor U10983 (N_10983,N_9222,N_8559);
or U10984 (N_10984,N_9876,N_8962);
nand U10985 (N_10985,N_8918,N_8817);
or U10986 (N_10986,N_9013,N_9353);
nand U10987 (N_10987,N_8781,N_8572);
nand U10988 (N_10988,N_9024,N_9534);
and U10989 (N_10989,N_8894,N_9152);
nor U10990 (N_10990,N_8858,N_8063);
nor U10991 (N_10991,N_8705,N_9274);
nand U10992 (N_10992,N_8444,N_8898);
and U10993 (N_10993,N_9357,N_8011);
or U10994 (N_10994,N_8691,N_9559);
xnor U10995 (N_10995,N_9653,N_9521);
or U10996 (N_10996,N_8477,N_9498);
and U10997 (N_10997,N_9524,N_8160);
and U10998 (N_10998,N_8832,N_9016);
nor U10999 (N_10999,N_9168,N_9216);
nor U11000 (N_11000,N_8629,N_9543);
nor U11001 (N_11001,N_9231,N_9372);
xnor U11002 (N_11002,N_8692,N_8295);
and U11003 (N_11003,N_8083,N_8076);
and U11004 (N_11004,N_8698,N_8411);
nand U11005 (N_11005,N_8662,N_9348);
or U11006 (N_11006,N_8555,N_9616);
and U11007 (N_11007,N_8763,N_8998);
nand U11008 (N_11008,N_8418,N_8130);
and U11009 (N_11009,N_8401,N_9358);
or U11010 (N_11010,N_8950,N_8958);
or U11011 (N_11011,N_9124,N_8979);
and U11012 (N_11012,N_9547,N_8901);
and U11013 (N_11013,N_9590,N_8138);
nand U11014 (N_11014,N_8432,N_8343);
and U11015 (N_11015,N_9960,N_8801);
nor U11016 (N_11016,N_8896,N_8301);
or U11017 (N_11017,N_9090,N_9176);
nand U11018 (N_11018,N_9238,N_8413);
nand U11019 (N_11019,N_8901,N_9437);
or U11020 (N_11020,N_8021,N_9210);
nor U11021 (N_11021,N_9265,N_8722);
or U11022 (N_11022,N_9115,N_8274);
and U11023 (N_11023,N_9454,N_9833);
nor U11024 (N_11024,N_8109,N_8633);
nand U11025 (N_11025,N_8115,N_8640);
and U11026 (N_11026,N_8260,N_8962);
nor U11027 (N_11027,N_8487,N_9800);
xnor U11028 (N_11028,N_8617,N_9611);
nand U11029 (N_11029,N_8049,N_8725);
and U11030 (N_11030,N_9061,N_8539);
and U11031 (N_11031,N_8240,N_8718);
nand U11032 (N_11032,N_8117,N_9251);
or U11033 (N_11033,N_8678,N_9722);
or U11034 (N_11034,N_8087,N_8536);
or U11035 (N_11035,N_8567,N_9103);
and U11036 (N_11036,N_8963,N_9283);
nor U11037 (N_11037,N_9188,N_9374);
nor U11038 (N_11038,N_8769,N_8653);
nand U11039 (N_11039,N_8741,N_8104);
or U11040 (N_11040,N_9637,N_9841);
xor U11041 (N_11041,N_8967,N_9364);
and U11042 (N_11042,N_8639,N_8816);
or U11043 (N_11043,N_8197,N_8068);
and U11044 (N_11044,N_9718,N_9251);
nand U11045 (N_11045,N_9903,N_9963);
or U11046 (N_11046,N_9868,N_8093);
nand U11047 (N_11047,N_8301,N_9735);
nand U11048 (N_11048,N_8764,N_8279);
and U11049 (N_11049,N_8093,N_9632);
and U11050 (N_11050,N_8237,N_9425);
and U11051 (N_11051,N_8121,N_8515);
nand U11052 (N_11052,N_8539,N_9993);
and U11053 (N_11053,N_8920,N_9144);
nand U11054 (N_11054,N_8669,N_8564);
nor U11055 (N_11055,N_8578,N_8554);
and U11056 (N_11056,N_9659,N_9934);
or U11057 (N_11057,N_8721,N_8937);
nor U11058 (N_11058,N_8386,N_8821);
nand U11059 (N_11059,N_8088,N_8053);
and U11060 (N_11060,N_9725,N_9647);
and U11061 (N_11061,N_9860,N_8758);
or U11062 (N_11062,N_8405,N_8505);
nand U11063 (N_11063,N_9932,N_9938);
xnor U11064 (N_11064,N_9391,N_9234);
nor U11065 (N_11065,N_8381,N_9324);
and U11066 (N_11066,N_8768,N_9342);
nor U11067 (N_11067,N_9705,N_8922);
or U11068 (N_11068,N_9420,N_8584);
or U11069 (N_11069,N_8112,N_9197);
and U11070 (N_11070,N_9223,N_9359);
nor U11071 (N_11071,N_9203,N_8434);
xnor U11072 (N_11072,N_8624,N_9073);
and U11073 (N_11073,N_9002,N_8732);
xnor U11074 (N_11074,N_9274,N_9174);
xnor U11075 (N_11075,N_8617,N_8849);
nand U11076 (N_11076,N_9610,N_8786);
nand U11077 (N_11077,N_9469,N_9288);
or U11078 (N_11078,N_8503,N_8541);
nor U11079 (N_11079,N_9822,N_8300);
nor U11080 (N_11080,N_8694,N_9899);
nor U11081 (N_11081,N_8841,N_9480);
nand U11082 (N_11082,N_8789,N_8659);
nand U11083 (N_11083,N_9879,N_9272);
nand U11084 (N_11084,N_8466,N_9846);
and U11085 (N_11085,N_9981,N_8137);
or U11086 (N_11086,N_8897,N_8219);
xor U11087 (N_11087,N_9510,N_9516);
nand U11088 (N_11088,N_8955,N_9903);
nor U11089 (N_11089,N_8676,N_8553);
and U11090 (N_11090,N_8273,N_8036);
nor U11091 (N_11091,N_8948,N_9993);
and U11092 (N_11092,N_8158,N_8885);
nor U11093 (N_11093,N_8643,N_8223);
nand U11094 (N_11094,N_8300,N_8626);
xnor U11095 (N_11095,N_9918,N_9567);
nor U11096 (N_11096,N_8386,N_8697);
nor U11097 (N_11097,N_8083,N_9033);
nor U11098 (N_11098,N_8324,N_8182);
nand U11099 (N_11099,N_9453,N_9909);
nand U11100 (N_11100,N_8985,N_8859);
nand U11101 (N_11101,N_8754,N_8551);
nand U11102 (N_11102,N_8572,N_9580);
or U11103 (N_11103,N_8202,N_8360);
or U11104 (N_11104,N_9097,N_8147);
nor U11105 (N_11105,N_9351,N_8725);
nor U11106 (N_11106,N_9654,N_9661);
xor U11107 (N_11107,N_8044,N_8941);
and U11108 (N_11108,N_9375,N_9264);
nand U11109 (N_11109,N_9867,N_9927);
nand U11110 (N_11110,N_8115,N_9624);
nand U11111 (N_11111,N_8353,N_8709);
or U11112 (N_11112,N_8380,N_9080);
and U11113 (N_11113,N_9236,N_8037);
nor U11114 (N_11114,N_8015,N_8701);
and U11115 (N_11115,N_9440,N_8844);
nor U11116 (N_11116,N_9342,N_9169);
or U11117 (N_11117,N_9209,N_8842);
nor U11118 (N_11118,N_9764,N_8582);
or U11119 (N_11119,N_9626,N_9652);
and U11120 (N_11120,N_8812,N_8545);
nor U11121 (N_11121,N_9326,N_9669);
nor U11122 (N_11122,N_9760,N_8190);
and U11123 (N_11123,N_9309,N_9629);
nand U11124 (N_11124,N_8395,N_8516);
nand U11125 (N_11125,N_9729,N_9415);
nor U11126 (N_11126,N_8866,N_9223);
or U11127 (N_11127,N_8392,N_8346);
nand U11128 (N_11128,N_8720,N_9369);
or U11129 (N_11129,N_9482,N_8191);
or U11130 (N_11130,N_8039,N_9274);
or U11131 (N_11131,N_8734,N_9009);
nor U11132 (N_11132,N_9874,N_9095);
or U11133 (N_11133,N_9788,N_8189);
nor U11134 (N_11134,N_8941,N_9605);
nor U11135 (N_11135,N_9569,N_8389);
nor U11136 (N_11136,N_9592,N_8407);
nor U11137 (N_11137,N_8414,N_9436);
nand U11138 (N_11138,N_8145,N_8934);
xor U11139 (N_11139,N_8889,N_9657);
or U11140 (N_11140,N_8567,N_8007);
or U11141 (N_11141,N_9810,N_9522);
nor U11142 (N_11142,N_8012,N_8784);
nand U11143 (N_11143,N_8176,N_9674);
nor U11144 (N_11144,N_8482,N_8937);
nor U11145 (N_11145,N_8114,N_9076);
nand U11146 (N_11146,N_8641,N_9026);
xor U11147 (N_11147,N_8656,N_8401);
or U11148 (N_11148,N_8083,N_8760);
nor U11149 (N_11149,N_9794,N_8909);
or U11150 (N_11150,N_9597,N_9157);
nor U11151 (N_11151,N_9011,N_8751);
or U11152 (N_11152,N_8875,N_9683);
or U11153 (N_11153,N_8911,N_8473);
nand U11154 (N_11154,N_8599,N_8092);
xor U11155 (N_11155,N_8959,N_9187);
and U11156 (N_11156,N_9070,N_9511);
or U11157 (N_11157,N_9191,N_8796);
and U11158 (N_11158,N_9025,N_8399);
and U11159 (N_11159,N_9049,N_9930);
nor U11160 (N_11160,N_8029,N_9437);
nor U11161 (N_11161,N_8806,N_8240);
xnor U11162 (N_11162,N_8226,N_8566);
nor U11163 (N_11163,N_9432,N_9968);
nand U11164 (N_11164,N_8908,N_9658);
xor U11165 (N_11165,N_9311,N_8016);
nand U11166 (N_11166,N_8309,N_9378);
and U11167 (N_11167,N_9472,N_9608);
nor U11168 (N_11168,N_8383,N_9700);
nor U11169 (N_11169,N_8826,N_8859);
nand U11170 (N_11170,N_9803,N_9344);
or U11171 (N_11171,N_8112,N_9139);
or U11172 (N_11172,N_9048,N_8987);
nor U11173 (N_11173,N_9164,N_9868);
xnor U11174 (N_11174,N_9649,N_8365);
or U11175 (N_11175,N_8798,N_8208);
or U11176 (N_11176,N_9928,N_8204);
or U11177 (N_11177,N_8479,N_9559);
and U11178 (N_11178,N_8505,N_8611);
nor U11179 (N_11179,N_9046,N_9852);
and U11180 (N_11180,N_9890,N_9185);
nand U11181 (N_11181,N_9512,N_9546);
nand U11182 (N_11182,N_9324,N_9666);
and U11183 (N_11183,N_9944,N_9391);
and U11184 (N_11184,N_9047,N_9363);
nor U11185 (N_11185,N_9095,N_8146);
nor U11186 (N_11186,N_8792,N_9497);
or U11187 (N_11187,N_9195,N_9669);
nand U11188 (N_11188,N_9236,N_9507);
and U11189 (N_11189,N_8037,N_8508);
or U11190 (N_11190,N_9376,N_8124);
and U11191 (N_11191,N_8002,N_9146);
nand U11192 (N_11192,N_9764,N_8674);
nor U11193 (N_11193,N_8426,N_9957);
nand U11194 (N_11194,N_9248,N_8574);
nor U11195 (N_11195,N_8973,N_8597);
nor U11196 (N_11196,N_9237,N_9667);
or U11197 (N_11197,N_8633,N_8711);
nor U11198 (N_11198,N_8780,N_8936);
or U11199 (N_11199,N_8739,N_9264);
nand U11200 (N_11200,N_9540,N_9417);
and U11201 (N_11201,N_9418,N_8787);
or U11202 (N_11202,N_9525,N_8141);
nor U11203 (N_11203,N_8316,N_8487);
xnor U11204 (N_11204,N_8529,N_9184);
or U11205 (N_11205,N_8357,N_9950);
and U11206 (N_11206,N_8148,N_8872);
nand U11207 (N_11207,N_8849,N_9599);
and U11208 (N_11208,N_9987,N_8378);
or U11209 (N_11209,N_8019,N_9230);
nand U11210 (N_11210,N_9292,N_8046);
xnor U11211 (N_11211,N_9492,N_8352);
or U11212 (N_11212,N_8474,N_8149);
nand U11213 (N_11213,N_8879,N_9051);
nor U11214 (N_11214,N_8377,N_9582);
nor U11215 (N_11215,N_8484,N_9013);
nand U11216 (N_11216,N_8916,N_9328);
nand U11217 (N_11217,N_9003,N_8183);
and U11218 (N_11218,N_9761,N_9406);
nor U11219 (N_11219,N_9417,N_8585);
nor U11220 (N_11220,N_8608,N_8230);
nand U11221 (N_11221,N_8562,N_9195);
or U11222 (N_11222,N_9064,N_8285);
and U11223 (N_11223,N_8264,N_9442);
nand U11224 (N_11224,N_8834,N_8535);
nor U11225 (N_11225,N_8353,N_8017);
and U11226 (N_11226,N_9377,N_8101);
nor U11227 (N_11227,N_8756,N_9517);
xor U11228 (N_11228,N_8795,N_9842);
nor U11229 (N_11229,N_9722,N_9553);
nand U11230 (N_11230,N_9371,N_9122);
or U11231 (N_11231,N_9856,N_8961);
nor U11232 (N_11232,N_8458,N_8820);
nor U11233 (N_11233,N_8770,N_9662);
nor U11234 (N_11234,N_8751,N_8797);
xnor U11235 (N_11235,N_8317,N_9730);
nand U11236 (N_11236,N_8902,N_8944);
nor U11237 (N_11237,N_9661,N_9177);
nor U11238 (N_11238,N_8350,N_8447);
and U11239 (N_11239,N_8696,N_8437);
nor U11240 (N_11240,N_8673,N_9821);
and U11241 (N_11241,N_8344,N_8798);
or U11242 (N_11242,N_9857,N_9863);
or U11243 (N_11243,N_9981,N_9349);
xnor U11244 (N_11244,N_9007,N_8808);
or U11245 (N_11245,N_9884,N_8176);
nor U11246 (N_11246,N_9288,N_8281);
nor U11247 (N_11247,N_8482,N_8432);
and U11248 (N_11248,N_9261,N_9785);
nor U11249 (N_11249,N_9425,N_9051);
nor U11250 (N_11250,N_9151,N_8272);
nand U11251 (N_11251,N_8897,N_9037);
nor U11252 (N_11252,N_9836,N_9457);
or U11253 (N_11253,N_9387,N_8570);
and U11254 (N_11254,N_8050,N_9557);
and U11255 (N_11255,N_8297,N_8083);
nand U11256 (N_11256,N_9527,N_8444);
nor U11257 (N_11257,N_9944,N_9889);
or U11258 (N_11258,N_9650,N_9724);
nand U11259 (N_11259,N_9757,N_9043);
or U11260 (N_11260,N_8132,N_9981);
and U11261 (N_11261,N_8242,N_8701);
nor U11262 (N_11262,N_8949,N_9123);
nor U11263 (N_11263,N_9556,N_9822);
nand U11264 (N_11264,N_9501,N_8513);
nand U11265 (N_11265,N_9860,N_8151);
nand U11266 (N_11266,N_9898,N_9644);
and U11267 (N_11267,N_8959,N_9331);
and U11268 (N_11268,N_8160,N_8099);
nand U11269 (N_11269,N_9455,N_9524);
nor U11270 (N_11270,N_8151,N_9613);
xor U11271 (N_11271,N_8587,N_9447);
and U11272 (N_11272,N_8232,N_8354);
or U11273 (N_11273,N_9278,N_9203);
or U11274 (N_11274,N_9360,N_9034);
or U11275 (N_11275,N_9779,N_8461);
nand U11276 (N_11276,N_9820,N_9861);
xnor U11277 (N_11277,N_9360,N_8739);
and U11278 (N_11278,N_9206,N_9228);
and U11279 (N_11279,N_8323,N_9394);
and U11280 (N_11280,N_9745,N_9780);
nand U11281 (N_11281,N_8544,N_8695);
nor U11282 (N_11282,N_8638,N_8784);
and U11283 (N_11283,N_8997,N_9893);
or U11284 (N_11284,N_8831,N_9570);
nand U11285 (N_11285,N_8208,N_9769);
or U11286 (N_11286,N_9008,N_8563);
or U11287 (N_11287,N_8251,N_9067);
nand U11288 (N_11288,N_8614,N_9758);
and U11289 (N_11289,N_9278,N_8223);
and U11290 (N_11290,N_9206,N_8909);
xor U11291 (N_11291,N_9635,N_9699);
and U11292 (N_11292,N_9867,N_9035);
and U11293 (N_11293,N_8953,N_8864);
and U11294 (N_11294,N_8024,N_9516);
nor U11295 (N_11295,N_9005,N_9284);
or U11296 (N_11296,N_9916,N_9722);
or U11297 (N_11297,N_8581,N_9801);
or U11298 (N_11298,N_8742,N_9148);
and U11299 (N_11299,N_8356,N_9511);
and U11300 (N_11300,N_8725,N_9390);
nor U11301 (N_11301,N_9752,N_9344);
and U11302 (N_11302,N_8820,N_8569);
nand U11303 (N_11303,N_8070,N_8282);
nand U11304 (N_11304,N_8339,N_9425);
nor U11305 (N_11305,N_9531,N_8155);
nand U11306 (N_11306,N_8725,N_8230);
nand U11307 (N_11307,N_9592,N_8495);
nand U11308 (N_11308,N_9686,N_8102);
nand U11309 (N_11309,N_8012,N_8712);
nand U11310 (N_11310,N_9215,N_9548);
nand U11311 (N_11311,N_9422,N_9455);
or U11312 (N_11312,N_9372,N_9676);
and U11313 (N_11313,N_9911,N_9227);
xnor U11314 (N_11314,N_9433,N_8153);
and U11315 (N_11315,N_9072,N_8945);
or U11316 (N_11316,N_9824,N_8998);
and U11317 (N_11317,N_9408,N_9980);
nor U11318 (N_11318,N_8277,N_8934);
xor U11319 (N_11319,N_9931,N_8017);
nand U11320 (N_11320,N_9844,N_8289);
or U11321 (N_11321,N_8123,N_9776);
or U11322 (N_11322,N_8599,N_8368);
nand U11323 (N_11323,N_8251,N_9215);
and U11324 (N_11324,N_9343,N_8731);
xnor U11325 (N_11325,N_8171,N_9284);
and U11326 (N_11326,N_9215,N_9701);
or U11327 (N_11327,N_9998,N_8547);
nor U11328 (N_11328,N_8267,N_9512);
nand U11329 (N_11329,N_9895,N_8096);
nand U11330 (N_11330,N_8546,N_9582);
or U11331 (N_11331,N_8757,N_8479);
nand U11332 (N_11332,N_9804,N_9979);
nand U11333 (N_11333,N_9198,N_9286);
or U11334 (N_11334,N_9746,N_9201);
nand U11335 (N_11335,N_9058,N_8008);
nand U11336 (N_11336,N_9694,N_8477);
and U11337 (N_11337,N_8712,N_9546);
nor U11338 (N_11338,N_9378,N_8579);
nand U11339 (N_11339,N_8414,N_8007);
and U11340 (N_11340,N_9015,N_9040);
nand U11341 (N_11341,N_9403,N_9339);
and U11342 (N_11342,N_8784,N_9044);
nand U11343 (N_11343,N_8237,N_8337);
and U11344 (N_11344,N_8771,N_9349);
or U11345 (N_11345,N_9459,N_8908);
nor U11346 (N_11346,N_9218,N_8349);
or U11347 (N_11347,N_8322,N_9270);
nand U11348 (N_11348,N_9943,N_8259);
nand U11349 (N_11349,N_8423,N_9148);
and U11350 (N_11350,N_8140,N_8689);
nand U11351 (N_11351,N_9708,N_9306);
and U11352 (N_11352,N_9111,N_9373);
nor U11353 (N_11353,N_8842,N_9919);
and U11354 (N_11354,N_8883,N_8645);
or U11355 (N_11355,N_8324,N_8342);
xor U11356 (N_11356,N_8375,N_9370);
nand U11357 (N_11357,N_8111,N_8224);
xnor U11358 (N_11358,N_8072,N_9953);
nor U11359 (N_11359,N_9573,N_9398);
xnor U11360 (N_11360,N_8949,N_8733);
nor U11361 (N_11361,N_8916,N_8607);
or U11362 (N_11362,N_9174,N_8521);
xnor U11363 (N_11363,N_9892,N_8794);
or U11364 (N_11364,N_9502,N_9519);
nor U11365 (N_11365,N_9162,N_8322);
nand U11366 (N_11366,N_8996,N_8590);
and U11367 (N_11367,N_8815,N_8093);
nor U11368 (N_11368,N_9300,N_8428);
or U11369 (N_11369,N_8041,N_9957);
nand U11370 (N_11370,N_8783,N_9653);
nand U11371 (N_11371,N_8459,N_9513);
or U11372 (N_11372,N_9806,N_9118);
or U11373 (N_11373,N_9573,N_8739);
or U11374 (N_11374,N_9390,N_8976);
and U11375 (N_11375,N_9632,N_8902);
or U11376 (N_11376,N_8117,N_8019);
and U11377 (N_11377,N_8704,N_9894);
or U11378 (N_11378,N_9175,N_8854);
xor U11379 (N_11379,N_9325,N_9347);
and U11380 (N_11380,N_8510,N_9969);
or U11381 (N_11381,N_9237,N_8802);
or U11382 (N_11382,N_9131,N_9140);
or U11383 (N_11383,N_9306,N_9540);
nor U11384 (N_11384,N_8269,N_8130);
xnor U11385 (N_11385,N_9341,N_8442);
xnor U11386 (N_11386,N_9493,N_9035);
or U11387 (N_11387,N_8596,N_9200);
and U11388 (N_11388,N_8806,N_8846);
and U11389 (N_11389,N_9295,N_9907);
and U11390 (N_11390,N_8143,N_9113);
nand U11391 (N_11391,N_9068,N_9582);
or U11392 (N_11392,N_8540,N_9508);
nand U11393 (N_11393,N_8309,N_9942);
and U11394 (N_11394,N_9588,N_8893);
nor U11395 (N_11395,N_9396,N_8704);
nand U11396 (N_11396,N_8485,N_9575);
nor U11397 (N_11397,N_9441,N_8376);
or U11398 (N_11398,N_9945,N_8308);
or U11399 (N_11399,N_8570,N_9150);
and U11400 (N_11400,N_8942,N_9633);
and U11401 (N_11401,N_9541,N_9413);
xor U11402 (N_11402,N_9538,N_8093);
and U11403 (N_11403,N_9105,N_8510);
or U11404 (N_11404,N_9058,N_8616);
nor U11405 (N_11405,N_8793,N_9206);
xnor U11406 (N_11406,N_9571,N_9716);
nor U11407 (N_11407,N_8038,N_8831);
nor U11408 (N_11408,N_8879,N_8804);
and U11409 (N_11409,N_8316,N_9150);
or U11410 (N_11410,N_8013,N_8422);
and U11411 (N_11411,N_8368,N_8625);
nand U11412 (N_11412,N_8138,N_9374);
nor U11413 (N_11413,N_8140,N_8947);
and U11414 (N_11414,N_9703,N_9936);
and U11415 (N_11415,N_9470,N_8515);
nor U11416 (N_11416,N_8932,N_8223);
nand U11417 (N_11417,N_9283,N_9999);
nand U11418 (N_11418,N_8513,N_9731);
nor U11419 (N_11419,N_8827,N_8902);
or U11420 (N_11420,N_9630,N_9960);
or U11421 (N_11421,N_8729,N_8603);
nor U11422 (N_11422,N_8866,N_8709);
and U11423 (N_11423,N_9783,N_8260);
and U11424 (N_11424,N_8919,N_8948);
or U11425 (N_11425,N_9644,N_8022);
nor U11426 (N_11426,N_8819,N_8506);
xor U11427 (N_11427,N_9037,N_8185);
nand U11428 (N_11428,N_8836,N_8834);
and U11429 (N_11429,N_9422,N_9300);
nor U11430 (N_11430,N_8408,N_9786);
nand U11431 (N_11431,N_8265,N_8385);
or U11432 (N_11432,N_9080,N_9128);
xnor U11433 (N_11433,N_9492,N_9947);
or U11434 (N_11434,N_9668,N_9308);
nand U11435 (N_11435,N_9374,N_8036);
and U11436 (N_11436,N_9588,N_8867);
or U11437 (N_11437,N_9344,N_8605);
and U11438 (N_11438,N_8998,N_9740);
xnor U11439 (N_11439,N_9273,N_8774);
and U11440 (N_11440,N_8580,N_8481);
xor U11441 (N_11441,N_8911,N_9788);
nor U11442 (N_11442,N_9506,N_9264);
nor U11443 (N_11443,N_8350,N_9607);
or U11444 (N_11444,N_8691,N_9645);
nor U11445 (N_11445,N_9037,N_9573);
or U11446 (N_11446,N_9604,N_9840);
and U11447 (N_11447,N_9719,N_9029);
and U11448 (N_11448,N_8994,N_8300);
xor U11449 (N_11449,N_9886,N_8810);
nand U11450 (N_11450,N_9767,N_9045);
nand U11451 (N_11451,N_9106,N_8843);
or U11452 (N_11452,N_9823,N_9696);
nor U11453 (N_11453,N_9585,N_9200);
nand U11454 (N_11454,N_9551,N_8212);
nand U11455 (N_11455,N_9572,N_8542);
and U11456 (N_11456,N_9234,N_8663);
nor U11457 (N_11457,N_9597,N_8529);
nor U11458 (N_11458,N_9199,N_9224);
and U11459 (N_11459,N_8733,N_8476);
xnor U11460 (N_11460,N_9995,N_8784);
and U11461 (N_11461,N_8877,N_8864);
nand U11462 (N_11462,N_9541,N_9251);
xor U11463 (N_11463,N_8036,N_9419);
or U11464 (N_11464,N_9161,N_9463);
nand U11465 (N_11465,N_9950,N_9819);
xnor U11466 (N_11466,N_8228,N_8677);
and U11467 (N_11467,N_8077,N_9425);
nor U11468 (N_11468,N_8858,N_8321);
nand U11469 (N_11469,N_9501,N_8986);
and U11470 (N_11470,N_8164,N_8443);
or U11471 (N_11471,N_9747,N_8866);
nor U11472 (N_11472,N_8345,N_9066);
or U11473 (N_11473,N_9581,N_9392);
nor U11474 (N_11474,N_9094,N_8649);
or U11475 (N_11475,N_8721,N_9324);
and U11476 (N_11476,N_8164,N_9069);
xor U11477 (N_11477,N_8010,N_8235);
nor U11478 (N_11478,N_8001,N_8605);
and U11479 (N_11479,N_8459,N_9256);
nand U11480 (N_11480,N_9705,N_8346);
nor U11481 (N_11481,N_8008,N_8913);
or U11482 (N_11482,N_9059,N_8883);
or U11483 (N_11483,N_9978,N_9515);
xnor U11484 (N_11484,N_9286,N_9212);
xor U11485 (N_11485,N_9450,N_8735);
and U11486 (N_11486,N_8627,N_8297);
nor U11487 (N_11487,N_9463,N_8732);
nand U11488 (N_11488,N_9762,N_9813);
nor U11489 (N_11489,N_9437,N_8679);
nor U11490 (N_11490,N_9789,N_9118);
or U11491 (N_11491,N_8822,N_8537);
xnor U11492 (N_11492,N_8349,N_8447);
xor U11493 (N_11493,N_8460,N_9867);
nand U11494 (N_11494,N_9648,N_9844);
or U11495 (N_11495,N_8056,N_8780);
or U11496 (N_11496,N_9349,N_9372);
or U11497 (N_11497,N_8265,N_9872);
and U11498 (N_11498,N_8122,N_9675);
xnor U11499 (N_11499,N_8620,N_8380);
or U11500 (N_11500,N_9449,N_9560);
nand U11501 (N_11501,N_8017,N_8674);
nand U11502 (N_11502,N_8247,N_8492);
xor U11503 (N_11503,N_8645,N_8893);
or U11504 (N_11504,N_9436,N_8011);
or U11505 (N_11505,N_8792,N_8668);
nor U11506 (N_11506,N_8585,N_8985);
and U11507 (N_11507,N_9485,N_8512);
nor U11508 (N_11508,N_8181,N_8511);
and U11509 (N_11509,N_9135,N_9634);
xor U11510 (N_11510,N_8446,N_8069);
or U11511 (N_11511,N_9858,N_9596);
or U11512 (N_11512,N_9960,N_9798);
nor U11513 (N_11513,N_9432,N_8050);
nor U11514 (N_11514,N_8631,N_9283);
or U11515 (N_11515,N_8362,N_9695);
or U11516 (N_11516,N_8056,N_8407);
nor U11517 (N_11517,N_9327,N_8713);
nand U11518 (N_11518,N_9862,N_9188);
or U11519 (N_11519,N_8091,N_8270);
or U11520 (N_11520,N_9196,N_8561);
nand U11521 (N_11521,N_8574,N_9636);
nand U11522 (N_11522,N_8557,N_8602);
nor U11523 (N_11523,N_9682,N_9468);
nand U11524 (N_11524,N_8713,N_9094);
and U11525 (N_11525,N_9686,N_8454);
nor U11526 (N_11526,N_9113,N_8557);
nor U11527 (N_11527,N_8420,N_9075);
or U11528 (N_11528,N_9539,N_8797);
xnor U11529 (N_11529,N_9537,N_8270);
xnor U11530 (N_11530,N_9300,N_9892);
nor U11531 (N_11531,N_8678,N_8033);
or U11532 (N_11532,N_9719,N_8098);
nand U11533 (N_11533,N_9591,N_8857);
nand U11534 (N_11534,N_9759,N_8858);
nand U11535 (N_11535,N_9160,N_8081);
and U11536 (N_11536,N_9049,N_8738);
xor U11537 (N_11537,N_9340,N_8402);
and U11538 (N_11538,N_8022,N_8846);
and U11539 (N_11539,N_8803,N_9653);
and U11540 (N_11540,N_9434,N_9508);
xnor U11541 (N_11541,N_9389,N_9297);
nor U11542 (N_11542,N_8619,N_8147);
and U11543 (N_11543,N_9962,N_9645);
or U11544 (N_11544,N_9271,N_8519);
and U11545 (N_11545,N_9747,N_9665);
nand U11546 (N_11546,N_8698,N_9758);
or U11547 (N_11547,N_9125,N_8026);
nor U11548 (N_11548,N_8091,N_8166);
nand U11549 (N_11549,N_9462,N_8274);
nor U11550 (N_11550,N_8377,N_8189);
and U11551 (N_11551,N_8470,N_9810);
or U11552 (N_11552,N_9260,N_8440);
xnor U11553 (N_11553,N_8848,N_8318);
nor U11554 (N_11554,N_9657,N_9749);
and U11555 (N_11555,N_9481,N_8287);
nor U11556 (N_11556,N_8800,N_9249);
nand U11557 (N_11557,N_9949,N_8172);
nor U11558 (N_11558,N_9532,N_9281);
nand U11559 (N_11559,N_8092,N_9896);
and U11560 (N_11560,N_8524,N_9502);
nand U11561 (N_11561,N_9837,N_8203);
nand U11562 (N_11562,N_9207,N_8964);
or U11563 (N_11563,N_9112,N_8311);
nand U11564 (N_11564,N_9881,N_8297);
nand U11565 (N_11565,N_9447,N_9894);
and U11566 (N_11566,N_9860,N_9434);
or U11567 (N_11567,N_9479,N_8992);
and U11568 (N_11568,N_9794,N_9344);
xnor U11569 (N_11569,N_9540,N_9826);
nor U11570 (N_11570,N_9058,N_9133);
or U11571 (N_11571,N_8545,N_8817);
nand U11572 (N_11572,N_8981,N_8478);
and U11573 (N_11573,N_8258,N_8824);
and U11574 (N_11574,N_9086,N_8357);
nand U11575 (N_11575,N_8454,N_9842);
or U11576 (N_11576,N_9369,N_8167);
nor U11577 (N_11577,N_8231,N_8044);
or U11578 (N_11578,N_8758,N_9514);
nor U11579 (N_11579,N_9040,N_8943);
nor U11580 (N_11580,N_9937,N_8289);
or U11581 (N_11581,N_9015,N_8268);
nand U11582 (N_11582,N_8494,N_8698);
nand U11583 (N_11583,N_8863,N_8298);
nor U11584 (N_11584,N_9255,N_8871);
or U11585 (N_11585,N_9350,N_8900);
nor U11586 (N_11586,N_8830,N_8276);
and U11587 (N_11587,N_8752,N_8557);
and U11588 (N_11588,N_8371,N_8917);
or U11589 (N_11589,N_8633,N_8272);
nand U11590 (N_11590,N_9855,N_8429);
nand U11591 (N_11591,N_9306,N_8010);
and U11592 (N_11592,N_9507,N_8590);
nand U11593 (N_11593,N_9575,N_9108);
nand U11594 (N_11594,N_8889,N_8535);
or U11595 (N_11595,N_8656,N_9227);
nor U11596 (N_11596,N_9577,N_9040);
or U11597 (N_11597,N_9801,N_8142);
nor U11598 (N_11598,N_8205,N_9764);
nor U11599 (N_11599,N_9762,N_8783);
and U11600 (N_11600,N_9746,N_8758);
and U11601 (N_11601,N_9835,N_8813);
and U11602 (N_11602,N_8397,N_8664);
and U11603 (N_11603,N_9240,N_9236);
or U11604 (N_11604,N_8948,N_8180);
or U11605 (N_11605,N_8412,N_8202);
and U11606 (N_11606,N_9678,N_8591);
nor U11607 (N_11607,N_8117,N_9812);
nand U11608 (N_11608,N_9070,N_8053);
nand U11609 (N_11609,N_9469,N_9247);
xor U11610 (N_11610,N_9081,N_9237);
and U11611 (N_11611,N_9650,N_9471);
and U11612 (N_11612,N_8571,N_8671);
nor U11613 (N_11613,N_8850,N_9681);
nor U11614 (N_11614,N_8183,N_9873);
xnor U11615 (N_11615,N_9239,N_8491);
nor U11616 (N_11616,N_8529,N_9003);
or U11617 (N_11617,N_8767,N_9253);
xor U11618 (N_11618,N_8601,N_9863);
nor U11619 (N_11619,N_8893,N_9826);
xnor U11620 (N_11620,N_8469,N_9639);
nand U11621 (N_11621,N_8271,N_8282);
or U11622 (N_11622,N_8573,N_8152);
nand U11623 (N_11623,N_8011,N_9254);
nand U11624 (N_11624,N_9286,N_9033);
nand U11625 (N_11625,N_8199,N_8182);
nor U11626 (N_11626,N_8071,N_8079);
and U11627 (N_11627,N_8965,N_9267);
and U11628 (N_11628,N_8438,N_9741);
nor U11629 (N_11629,N_9106,N_8027);
nor U11630 (N_11630,N_8823,N_8567);
nand U11631 (N_11631,N_8928,N_8572);
or U11632 (N_11632,N_9068,N_9041);
nand U11633 (N_11633,N_9335,N_9195);
and U11634 (N_11634,N_9017,N_8373);
nand U11635 (N_11635,N_9433,N_9125);
nor U11636 (N_11636,N_8342,N_8167);
or U11637 (N_11637,N_8207,N_8657);
xnor U11638 (N_11638,N_9809,N_9332);
and U11639 (N_11639,N_8907,N_9963);
and U11640 (N_11640,N_9923,N_8668);
nor U11641 (N_11641,N_9635,N_9027);
xor U11642 (N_11642,N_9847,N_9161);
and U11643 (N_11643,N_9477,N_9118);
nand U11644 (N_11644,N_9182,N_8492);
and U11645 (N_11645,N_9168,N_8115);
or U11646 (N_11646,N_9713,N_9569);
nor U11647 (N_11647,N_9892,N_8964);
or U11648 (N_11648,N_8880,N_8741);
and U11649 (N_11649,N_9907,N_8933);
nand U11650 (N_11650,N_9618,N_8666);
and U11651 (N_11651,N_8425,N_9900);
or U11652 (N_11652,N_9230,N_9895);
nor U11653 (N_11653,N_8311,N_8185);
and U11654 (N_11654,N_9942,N_8414);
and U11655 (N_11655,N_9606,N_8151);
or U11656 (N_11656,N_9493,N_8365);
and U11657 (N_11657,N_9117,N_9092);
xor U11658 (N_11658,N_8423,N_9018);
nand U11659 (N_11659,N_8135,N_8764);
nand U11660 (N_11660,N_8738,N_9622);
xnor U11661 (N_11661,N_9198,N_9967);
xnor U11662 (N_11662,N_8000,N_8953);
nand U11663 (N_11663,N_8382,N_9488);
xor U11664 (N_11664,N_9471,N_9402);
nor U11665 (N_11665,N_8276,N_9900);
nand U11666 (N_11666,N_8654,N_9432);
or U11667 (N_11667,N_9742,N_8990);
and U11668 (N_11668,N_8756,N_9565);
nor U11669 (N_11669,N_9516,N_9584);
or U11670 (N_11670,N_9398,N_9199);
nand U11671 (N_11671,N_9032,N_8819);
or U11672 (N_11672,N_8462,N_8447);
nor U11673 (N_11673,N_8716,N_8763);
or U11674 (N_11674,N_8393,N_9324);
nand U11675 (N_11675,N_9730,N_8279);
xor U11676 (N_11676,N_8987,N_9738);
nand U11677 (N_11677,N_9198,N_8945);
and U11678 (N_11678,N_9257,N_8446);
nand U11679 (N_11679,N_8033,N_9708);
nand U11680 (N_11680,N_8663,N_9028);
nand U11681 (N_11681,N_8176,N_9878);
and U11682 (N_11682,N_9533,N_9703);
xor U11683 (N_11683,N_9038,N_8701);
or U11684 (N_11684,N_9264,N_9183);
or U11685 (N_11685,N_8938,N_8940);
nor U11686 (N_11686,N_9583,N_9154);
and U11687 (N_11687,N_8784,N_8004);
or U11688 (N_11688,N_8140,N_8454);
nand U11689 (N_11689,N_8353,N_8247);
or U11690 (N_11690,N_9341,N_9676);
nor U11691 (N_11691,N_9637,N_8396);
nand U11692 (N_11692,N_9624,N_9155);
nand U11693 (N_11693,N_8796,N_8600);
nor U11694 (N_11694,N_8534,N_8261);
nand U11695 (N_11695,N_8097,N_8651);
or U11696 (N_11696,N_9814,N_9989);
nand U11697 (N_11697,N_9772,N_9349);
xnor U11698 (N_11698,N_9767,N_9312);
and U11699 (N_11699,N_9143,N_8348);
or U11700 (N_11700,N_8195,N_8023);
and U11701 (N_11701,N_9496,N_8165);
nor U11702 (N_11702,N_8697,N_8753);
nand U11703 (N_11703,N_9076,N_9462);
nand U11704 (N_11704,N_9402,N_9748);
xnor U11705 (N_11705,N_8573,N_8402);
nor U11706 (N_11706,N_9641,N_9377);
nand U11707 (N_11707,N_9443,N_8881);
and U11708 (N_11708,N_9619,N_8377);
nand U11709 (N_11709,N_9723,N_9465);
xor U11710 (N_11710,N_9184,N_9835);
or U11711 (N_11711,N_8845,N_8732);
nand U11712 (N_11712,N_9288,N_9750);
nand U11713 (N_11713,N_9534,N_8753);
nor U11714 (N_11714,N_9442,N_8158);
and U11715 (N_11715,N_8216,N_8051);
nand U11716 (N_11716,N_8133,N_9167);
nand U11717 (N_11717,N_8916,N_8207);
nand U11718 (N_11718,N_8071,N_8823);
and U11719 (N_11719,N_9870,N_9523);
or U11720 (N_11720,N_9447,N_9634);
nand U11721 (N_11721,N_8562,N_8568);
or U11722 (N_11722,N_9457,N_8120);
nand U11723 (N_11723,N_9834,N_8284);
and U11724 (N_11724,N_8717,N_8027);
xnor U11725 (N_11725,N_8276,N_8773);
nand U11726 (N_11726,N_8290,N_9264);
nand U11727 (N_11727,N_8083,N_8123);
nor U11728 (N_11728,N_8611,N_8731);
and U11729 (N_11729,N_9054,N_8173);
nand U11730 (N_11730,N_8029,N_9114);
xnor U11731 (N_11731,N_9528,N_8870);
nor U11732 (N_11732,N_9186,N_9262);
nor U11733 (N_11733,N_9225,N_9756);
and U11734 (N_11734,N_8640,N_9216);
or U11735 (N_11735,N_8824,N_9056);
or U11736 (N_11736,N_9153,N_9368);
and U11737 (N_11737,N_9653,N_9766);
and U11738 (N_11738,N_8044,N_8996);
and U11739 (N_11739,N_8671,N_8953);
or U11740 (N_11740,N_8607,N_8446);
xor U11741 (N_11741,N_9041,N_8097);
nor U11742 (N_11742,N_9200,N_8945);
and U11743 (N_11743,N_8593,N_9456);
xnor U11744 (N_11744,N_9389,N_9609);
nor U11745 (N_11745,N_9406,N_9161);
nor U11746 (N_11746,N_8187,N_9358);
nor U11747 (N_11747,N_9856,N_9421);
or U11748 (N_11748,N_9790,N_9396);
nand U11749 (N_11749,N_8271,N_8456);
or U11750 (N_11750,N_8805,N_8539);
or U11751 (N_11751,N_9048,N_8581);
and U11752 (N_11752,N_9879,N_9855);
xor U11753 (N_11753,N_9693,N_9161);
nand U11754 (N_11754,N_8010,N_9537);
or U11755 (N_11755,N_9217,N_9018);
or U11756 (N_11756,N_8186,N_9508);
nand U11757 (N_11757,N_9089,N_8116);
nand U11758 (N_11758,N_9156,N_9034);
nand U11759 (N_11759,N_9026,N_9657);
or U11760 (N_11760,N_8920,N_9183);
nor U11761 (N_11761,N_9108,N_9740);
and U11762 (N_11762,N_8730,N_8577);
nand U11763 (N_11763,N_9033,N_9065);
and U11764 (N_11764,N_9619,N_8608);
nor U11765 (N_11765,N_9355,N_8363);
or U11766 (N_11766,N_8641,N_9747);
and U11767 (N_11767,N_9765,N_9406);
and U11768 (N_11768,N_9148,N_9422);
nand U11769 (N_11769,N_8590,N_9161);
nand U11770 (N_11770,N_9782,N_9254);
xnor U11771 (N_11771,N_8370,N_9556);
nand U11772 (N_11772,N_9063,N_9343);
or U11773 (N_11773,N_9542,N_8452);
or U11774 (N_11774,N_9679,N_9964);
xnor U11775 (N_11775,N_8245,N_9031);
xnor U11776 (N_11776,N_8668,N_9399);
nand U11777 (N_11777,N_8496,N_8998);
and U11778 (N_11778,N_8811,N_9913);
and U11779 (N_11779,N_8299,N_8197);
nand U11780 (N_11780,N_8688,N_9543);
nand U11781 (N_11781,N_9137,N_8604);
and U11782 (N_11782,N_8445,N_9829);
xor U11783 (N_11783,N_8930,N_9685);
or U11784 (N_11784,N_8648,N_9141);
nor U11785 (N_11785,N_9677,N_8809);
and U11786 (N_11786,N_9744,N_8400);
nand U11787 (N_11787,N_9255,N_8324);
nand U11788 (N_11788,N_8810,N_9295);
nor U11789 (N_11789,N_9279,N_8260);
nand U11790 (N_11790,N_9872,N_9785);
xnor U11791 (N_11791,N_8167,N_9202);
or U11792 (N_11792,N_9530,N_9583);
nor U11793 (N_11793,N_9238,N_8008);
nand U11794 (N_11794,N_8601,N_9285);
nand U11795 (N_11795,N_9966,N_8872);
and U11796 (N_11796,N_8958,N_8594);
nor U11797 (N_11797,N_8846,N_9016);
and U11798 (N_11798,N_9144,N_8772);
and U11799 (N_11799,N_9183,N_8721);
nor U11800 (N_11800,N_8786,N_8787);
nand U11801 (N_11801,N_9265,N_8757);
nand U11802 (N_11802,N_8702,N_8347);
and U11803 (N_11803,N_8321,N_9941);
or U11804 (N_11804,N_9637,N_9985);
or U11805 (N_11805,N_9714,N_8346);
nand U11806 (N_11806,N_9865,N_8880);
nor U11807 (N_11807,N_8501,N_8463);
or U11808 (N_11808,N_9463,N_9937);
or U11809 (N_11809,N_9795,N_9762);
and U11810 (N_11810,N_8383,N_9608);
nor U11811 (N_11811,N_9867,N_8154);
nand U11812 (N_11812,N_8222,N_8626);
or U11813 (N_11813,N_9689,N_8908);
and U11814 (N_11814,N_9479,N_8201);
and U11815 (N_11815,N_8406,N_9163);
or U11816 (N_11816,N_8814,N_8130);
nand U11817 (N_11817,N_9651,N_9849);
and U11818 (N_11818,N_8036,N_9517);
nand U11819 (N_11819,N_9352,N_9025);
and U11820 (N_11820,N_9365,N_9161);
nor U11821 (N_11821,N_8049,N_9542);
xor U11822 (N_11822,N_8984,N_9157);
xor U11823 (N_11823,N_9517,N_8597);
and U11824 (N_11824,N_8986,N_9171);
and U11825 (N_11825,N_8949,N_9031);
and U11826 (N_11826,N_9857,N_8237);
nand U11827 (N_11827,N_8302,N_9905);
nand U11828 (N_11828,N_9604,N_9016);
and U11829 (N_11829,N_8301,N_8160);
nor U11830 (N_11830,N_8748,N_8960);
nand U11831 (N_11831,N_9145,N_8864);
nor U11832 (N_11832,N_9373,N_9034);
xor U11833 (N_11833,N_9028,N_9776);
and U11834 (N_11834,N_8735,N_9226);
nand U11835 (N_11835,N_8334,N_9658);
or U11836 (N_11836,N_8265,N_9601);
xnor U11837 (N_11837,N_9534,N_8453);
xnor U11838 (N_11838,N_8821,N_9205);
nand U11839 (N_11839,N_8766,N_9186);
nand U11840 (N_11840,N_9803,N_8042);
nor U11841 (N_11841,N_8131,N_8261);
and U11842 (N_11842,N_9200,N_8738);
and U11843 (N_11843,N_9443,N_9316);
and U11844 (N_11844,N_9281,N_9175);
nand U11845 (N_11845,N_9140,N_8762);
or U11846 (N_11846,N_8418,N_9115);
nor U11847 (N_11847,N_8151,N_9260);
xnor U11848 (N_11848,N_8088,N_9072);
nand U11849 (N_11849,N_8931,N_8448);
and U11850 (N_11850,N_8969,N_8857);
or U11851 (N_11851,N_8091,N_8549);
and U11852 (N_11852,N_8605,N_8000);
and U11853 (N_11853,N_8866,N_9896);
nor U11854 (N_11854,N_9198,N_9369);
or U11855 (N_11855,N_9205,N_8000);
or U11856 (N_11856,N_9700,N_8931);
nor U11857 (N_11857,N_9575,N_8338);
nor U11858 (N_11858,N_9648,N_9443);
and U11859 (N_11859,N_8676,N_9389);
nand U11860 (N_11860,N_9530,N_8118);
or U11861 (N_11861,N_8100,N_9573);
and U11862 (N_11862,N_9311,N_9827);
and U11863 (N_11863,N_9043,N_8976);
xor U11864 (N_11864,N_9792,N_8156);
or U11865 (N_11865,N_8539,N_8402);
and U11866 (N_11866,N_8015,N_9643);
and U11867 (N_11867,N_9413,N_8875);
nor U11868 (N_11868,N_8736,N_9639);
and U11869 (N_11869,N_9480,N_8047);
and U11870 (N_11870,N_9381,N_8021);
xnor U11871 (N_11871,N_8780,N_8440);
nor U11872 (N_11872,N_8749,N_9241);
and U11873 (N_11873,N_8101,N_9754);
nand U11874 (N_11874,N_8882,N_8697);
nor U11875 (N_11875,N_8874,N_9816);
or U11876 (N_11876,N_8369,N_8384);
or U11877 (N_11877,N_8403,N_9261);
or U11878 (N_11878,N_9054,N_9186);
nand U11879 (N_11879,N_8632,N_8642);
nand U11880 (N_11880,N_9263,N_9597);
nor U11881 (N_11881,N_9459,N_8508);
and U11882 (N_11882,N_8658,N_9047);
and U11883 (N_11883,N_8521,N_8534);
nor U11884 (N_11884,N_8122,N_8415);
nor U11885 (N_11885,N_8415,N_8632);
nand U11886 (N_11886,N_9294,N_9702);
or U11887 (N_11887,N_8144,N_8411);
and U11888 (N_11888,N_8269,N_8592);
xor U11889 (N_11889,N_8241,N_9654);
or U11890 (N_11890,N_9428,N_9498);
or U11891 (N_11891,N_9493,N_8932);
xor U11892 (N_11892,N_9020,N_8469);
nor U11893 (N_11893,N_9812,N_8624);
or U11894 (N_11894,N_8307,N_9182);
or U11895 (N_11895,N_9947,N_9164);
nand U11896 (N_11896,N_9786,N_8733);
nor U11897 (N_11897,N_9175,N_9841);
or U11898 (N_11898,N_9219,N_8897);
nor U11899 (N_11899,N_8667,N_8271);
nand U11900 (N_11900,N_8312,N_9149);
and U11901 (N_11901,N_8936,N_9064);
or U11902 (N_11902,N_8861,N_9994);
xnor U11903 (N_11903,N_8885,N_9104);
nor U11904 (N_11904,N_9565,N_9785);
nand U11905 (N_11905,N_8929,N_8540);
nor U11906 (N_11906,N_9752,N_9465);
and U11907 (N_11907,N_8864,N_8691);
or U11908 (N_11908,N_9673,N_9310);
nand U11909 (N_11909,N_9925,N_9976);
nor U11910 (N_11910,N_8468,N_8327);
and U11911 (N_11911,N_9564,N_8304);
or U11912 (N_11912,N_8799,N_8098);
nand U11913 (N_11913,N_9528,N_8331);
or U11914 (N_11914,N_8988,N_8280);
nor U11915 (N_11915,N_8178,N_9952);
xor U11916 (N_11916,N_9112,N_9407);
nor U11917 (N_11917,N_9483,N_8589);
nor U11918 (N_11918,N_8495,N_8791);
nor U11919 (N_11919,N_8185,N_9551);
nand U11920 (N_11920,N_9653,N_9299);
or U11921 (N_11921,N_9936,N_8691);
nor U11922 (N_11922,N_8805,N_8812);
nand U11923 (N_11923,N_8761,N_9673);
nand U11924 (N_11924,N_8393,N_9631);
nor U11925 (N_11925,N_9489,N_9077);
or U11926 (N_11926,N_9873,N_9845);
or U11927 (N_11927,N_8790,N_9133);
and U11928 (N_11928,N_9912,N_9169);
and U11929 (N_11929,N_9975,N_9658);
nor U11930 (N_11930,N_9372,N_8588);
nor U11931 (N_11931,N_8167,N_9282);
nand U11932 (N_11932,N_8137,N_8000);
and U11933 (N_11933,N_8141,N_9020);
nand U11934 (N_11934,N_9367,N_9908);
or U11935 (N_11935,N_9768,N_8603);
nor U11936 (N_11936,N_8423,N_8168);
nor U11937 (N_11937,N_8096,N_9348);
nor U11938 (N_11938,N_8153,N_8754);
nor U11939 (N_11939,N_9696,N_8616);
and U11940 (N_11940,N_9476,N_9551);
nand U11941 (N_11941,N_9932,N_9153);
xor U11942 (N_11942,N_9479,N_9164);
nand U11943 (N_11943,N_9057,N_8722);
nand U11944 (N_11944,N_8484,N_9082);
nor U11945 (N_11945,N_8523,N_8520);
and U11946 (N_11946,N_8647,N_8847);
or U11947 (N_11947,N_8891,N_9320);
and U11948 (N_11948,N_8061,N_9109);
nand U11949 (N_11949,N_9568,N_9455);
and U11950 (N_11950,N_8809,N_9292);
nor U11951 (N_11951,N_9905,N_8341);
and U11952 (N_11952,N_9514,N_9233);
nand U11953 (N_11953,N_8893,N_9327);
and U11954 (N_11954,N_9544,N_9182);
nor U11955 (N_11955,N_9189,N_9075);
xnor U11956 (N_11956,N_9570,N_8253);
and U11957 (N_11957,N_8598,N_9680);
nor U11958 (N_11958,N_9211,N_9115);
nand U11959 (N_11959,N_8001,N_8642);
or U11960 (N_11960,N_9948,N_8863);
and U11961 (N_11961,N_8238,N_9586);
or U11962 (N_11962,N_9576,N_8684);
and U11963 (N_11963,N_8195,N_8289);
xnor U11964 (N_11964,N_9208,N_9533);
nor U11965 (N_11965,N_9218,N_8442);
nand U11966 (N_11966,N_8925,N_9846);
xnor U11967 (N_11967,N_9883,N_9203);
nor U11968 (N_11968,N_8163,N_9468);
and U11969 (N_11969,N_9219,N_9847);
nand U11970 (N_11970,N_8359,N_8960);
or U11971 (N_11971,N_8552,N_8714);
nand U11972 (N_11972,N_9613,N_9008);
or U11973 (N_11973,N_9516,N_9336);
nor U11974 (N_11974,N_8328,N_8808);
and U11975 (N_11975,N_8895,N_9347);
nor U11976 (N_11976,N_9215,N_9299);
or U11977 (N_11977,N_8565,N_9537);
nand U11978 (N_11978,N_8126,N_9655);
xor U11979 (N_11979,N_9500,N_9543);
nor U11980 (N_11980,N_8668,N_8016);
nor U11981 (N_11981,N_9593,N_8112);
or U11982 (N_11982,N_8432,N_9375);
and U11983 (N_11983,N_9693,N_8333);
nand U11984 (N_11984,N_8176,N_8156);
or U11985 (N_11985,N_9478,N_9178);
and U11986 (N_11986,N_8121,N_9470);
nand U11987 (N_11987,N_8316,N_9465);
or U11988 (N_11988,N_8250,N_8658);
xnor U11989 (N_11989,N_9969,N_9884);
nand U11990 (N_11990,N_9593,N_8841);
nand U11991 (N_11991,N_8613,N_9081);
nor U11992 (N_11992,N_8428,N_9044);
and U11993 (N_11993,N_8472,N_8401);
and U11994 (N_11994,N_9191,N_9248);
nand U11995 (N_11995,N_9733,N_8155);
or U11996 (N_11996,N_9509,N_9679);
xor U11997 (N_11997,N_9169,N_8994);
nand U11998 (N_11998,N_9782,N_9435);
and U11999 (N_11999,N_9976,N_8113);
nor U12000 (N_12000,N_10969,N_11431);
or U12001 (N_12001,N_10463,N_11892);
nand U12002 (N_12002,N_11032,N_10519);
nor U12003 (N_12003,N_10116,N_11517);
nor U12004 (N_12004,N_10595,N_10728);
or U12005 (N_12005,N_11300,N_11659);
or U12006 (N_12006,N_10311,N_11419);
or U12007 (N_12007,N_10660,N_11863);
or U12008 (N_12008,N_11026,N_11034);
nand U12009 (N_12009,N_11769,N_11317);
nor U12010 (N_12010,N_11741,N_11004);
xor U12011 (N_12011,N_11212,N_11726);
nand U12012 (N_12012,N_10177,N_10924);
xnor U12013 (N_12013,N_10146,N_10062);
nand U12014 (N_12014,N_10475,N_11414);
nor U12015 (N_12015,N_11422,N_10798);
and U12016 (N_12016,N_10037,N_11530);
nand U12017 (N_12017,N_11228,N_10920);
and U12018 (N_12018,N_10200,N_11861);
and U12019 (N_12019,N_11194,N_11233);
nor U12020 (N_12020,N_11258,N_11661);
or U12021 (N_12021,N_11810,N_10716);
or U12022 (N_12022,N_10398,N_10726);
or U12023 (N_12023,N_11943,N_10386);
or U12024 (N_12024,N_11471,N_11203);
and U12025 (N_12025,N_10316,N_11293);
nor U12026 (N_12026,N_10459,N_11591);
and U12027 (N_12027,N_10497,N_10906);
xnor U12028 (N_12028,N_11296,N_10259);
nor U12029 (N_12029,N_11149,N_11724);
nand U12030 (N_12030,N_10941,N_10529);
nand U12031 (N_12031,N_10206,N_11276);
and U12032 (N_12032,N_10397,N_11041);
or U12033 (N_12033,N_10372,N_11039);
nor U12034 (N_12034,N_10283,N_11397);
xnor U12035 (N_12035,N_11833,N_10006);
nor U12036 (N_12036,N_10354,N_10488);
or U12037 (N_12037,N_10710,N_10773);
and U12038 (N_12038,N_11009,N_11989);
or U12039 (N_12039,N_11054,N_11786);
nor U12040 (N_12040,N_11177,N_10778);
nor U12041 (N_12041,N_11027,N_11285);
nand U12042 (N_12042,N_10676,N_11230);
nand U12043 (N_12043,N_10277,N_10167);
and U12044 (N_12044,N_11541,N_10797);
nor U12045 (N_12045,N_11209,N_11898);
nand U12046 (N_12046,N_10000,N_11876);
and U12047 (N_12047,N_10958,N_11208);
xnor U12048 (N_12048,N_10059,N_10912);
nand U12049 (N_12049,N_11796,N_10182);
or U12050 (N_12050,N_11988,N_11868);
nand U12051 (N_12051,N_11959,N_10988);
nand U12052 (N_12052,N_11494,N_10426);
or U12053 (N_12053,N_11660,N_10455);
or U12054 (N_12054,N_11896,N_10885);
nor U12055 (N_12055,N_10799,N_10703);
nor U12056 (N_12056,N_11901,N_11284);
nor U12057 (N_12057,N_11062,N_10980);
nand U12058 (N_12058,N_11337,N_10026);
or U12059 (N_12059,N_11515,N_10262);
and U12060 (N_12060,N_10528,N_11506);
nor U12061 (N_12061,N_11475,N_11050);
nand U12062 (N_12062,N_10496,N_10091);
nand U12063 (N_12063,N_11218,N_10139);
nor U12064 (N_12064,N_11392,N_10827);
nand U12065 (N_12065,N_11335,N_11148);
and U12066 (N_12066,N_11634,N_10966);
nand U12067 (N_12067,N_10217,N_10098);
or U12068 (N_12068,N_10466,N_10141);
and U12069 (N_12069,N_10093,N_10585);
nand U12070 (N_12070,N_11927,N_10701);
nor U12071 (N_12071,N_11622,N_10044);
xnor U12072 (N_12072,N_10298,N_11791);
nor U12073 (N_12073,N_11491,N_11639);
nand U12074 (N_12074,N_10396,N_11060);
nand U12075 (N_12075,N_10263,N_11339);
nand U12076 (N_12076,N_10084,N_10584);
nand U12077 (N_12077,N_11836,N_11525);
nand U12078 (N_12078,N_11554,N_11484);
nor U12079 (N_12079,N_10057,N_11320);
or U12080 (N_12080,N_11520,N_11731);
and U12081 (N_12081,N_10621,N_11464);
nand U12082 (N_12082,N_11559,N_10190);
and U12083 (N_12083,N_11937,N_10881);
nand U12084 (N_12084,N_11082,N_11888);
nor U12085 (N_12085,N_11438,N_10117);
and U12086 (N_12086,N_11749,N_10154);
and U12087 (N_12087,N_11151,N_11167);
xor U12088 (N_12088,N_11692,N_10166);
nor U12089 (N_12089,N_11220,N_11911);
nor U12090 (N_12090,N_11044,N_11845);
and U12091 (N_12091,N_10563,N_10597);
or U12092 (N_12092,N_10013,N_10187);
and U12093 (N_12093,N_11254,N_11941);
and U12094 (N_12094,N_10744,N_11906);
nor U12095 (N_12095,N_10504,N_10122);
nor U12096 (N_12096,N_10367,N_11578);
or U12097 (N_12097,N_10658,N_10695);
or U12098 (N_12098,N_10168,N_10108);
or U12099 (N_12099,N_10685,N_11547);
nand U12100 (N_12100,N_10754,N_10417);
nor U12101 (N_12101,N_10602,N_10382);
nand U12102 (N_12102,N_11432,N_11206);
xor U12103 (N_12103,N_11684,N_10423);
or U12104 (N_12104,N_11568,N_10617);
xor U12105 (N_12105,N_11925,N_11608);
nor U12106 (N_12106,N_11991,N_11361);
and U12107 (N_12107,N_10665,N_11222);
nand U12108 (N_12108,N_11664,N_10952);
and U12109 (N_12109,N_10739,N_10300);
nor U12110 (N_12110,N_11002,N_11346);
or U12111 (N_12111,N_10564,N_11827);
nor U12112 (N_12112,N_11150,N_11662);
nor U12113 (N_12113,N_11116,N_10219);
or U12114 (N_12114,N_10930,N_11821);
or U12115 (N_12115,N_10434,N_11739);
nor U12116 (N_12116,N_10207,N_10979);
and U12117 (N_12117,N_10982,N_10048);
nand U12118 (N_12118,N_10087,N_10285);
and U12119 (N_12119,N_11262,N_10853);
xnor U12120 (N_12120,N_11118,N_11366);
nor U12121 (N_12121,N_10025,N_10557);
and U12122 (N_12122,N_10272,N_10032);
or U12123 (N_12123,N_10607,N_10295);
and U12124 (N_12124,N_11294,N_11129);
nor U12125 (N_12125,N_11143,N_10641);
or U12126 (N_12126,N_11020,N_11918);
or U12127 (N_12127,N_11882,N_10990);
and U12128 (N_12128,N_10713,N_11881);
nand U12129 (N_12129,N_11866,N_11385);
nand U12130 (N_12130,N_11446,N_10513);
and U12131 (N_12131,N_10593,N_11486);
or U12132 (N_12132,N_10137,N_10222);
or U12133 (N_12133,N_10944,N_10619);
nor U12134 (N_12134,N_11737,N_11519);
or U12135 (N_12135,N_10800,N_11551);
or U12136 (N_12136,N_10796,N_10771);
nand U12137 (N_12137,N_10101,N_10369);
nand U12138 (N_12138,N_11632,N_10391);
nor U12139 (N_12139,N_10140,N_11711);
nor U12140 (N_12140,N_11008,N_10229);
or U12141 (N_12141,N_11204,N_11500);
and U12142 (N_12142,N_10942,N_11405);
nor U12143 (N_12143,N_11755,N_11123);
and U12144 (N_12144,N_11685,N_11072);
and U12145 (N_12145,N_11862,N_10258);
nor U12146 (N_12146,N_10544,N_11606);
or U12147 (N_12147,N_11449,N_11127);
nand U12148 (N_12148,N_11428,N_10293);
xnor U12149 (N_12149,N_11156,N_10839);
or U12150 (N_12150,N_10679,N_10786);
nand U12151 (N_12151,N_10787,N_11847);
nand U12152 (N_12152,N_10095,N_10393);
and U12153 (N_12153,N_11185,N_10824);
and U12154 (N_12154,N_10075,N_11552);
nor U12155 (N_12155,N_11899,N_11994);
or U12156 (N_12156,N_11101,N_10317);
nor U12157 (N_12157,N_11553,N_10169);
and U12158 (N_12158,N_10702,N_10536);
nand U12159 (N_12159,N_10805,N_11736);
and U12160 (N_12160,N_10629,N_10869);
xnor U12161 (N_12161,N_10202,N_10662);
xnor U12162 (N_12162,N_11990,N_11012);
or U12163 (N_12163,N_10905,N_10724);
and U12164 (N_12164,N_10943,N_10668);
nor U12165 (N_12165,N_10416,N_10440);
nor U12166 (N_12166,N_11409,N_10254);
and U12167 (N_12167,N_11851,N_11281);
and U12168 (N_12168,N_10681,N_10328);
and U12169 (N_12169,N_10748,N_10014);
nand U12170 (N_12170,N_11213,N_11670);
nor U12171 (N_12171,N_11891,N_11113);
and U12172 (N_12172,N_10368,N_11939);
xnor U12173 (N_12173,N_10663,N_11013);
nand U12174 (N_12174,N_11135,N_10851);
nand U12175 (N_12175,N_10307,N_10763);
xnor U12176 (N_12176,N_11858,N_11406);
or U12177 (N_12177,N_11426,N_11586);
nor U12178 (N_12178,N_10768,N_10226);
nor U12179 (N_12179,N_10633,N_10170);
nand U12180 (N_12180,N_11442,N_10600);
and U12181 (N_12181,N_10001,N_11681);
nor U12182 (N_12182,N_10596,N_10238);
and U12183 (N_12183,N_11631,N_11915);
nand U12184 (N_12184,N_10220,N_10056);
nand U12185 (N_12185,N_10845,N_11114);
nand U12186 (N_12186,N_10953,N_11318);
nand U12187 (N_12187,N_10365,N_11964);
or U12188 (N_12188,N_10627,N_11125);
or U12189 (N_12189,N_10592,N_10591);
nor U12190 (N_12190,N_11751,N_11745);
xor U12191 (N_12191,N_11652,N_11313);
and U12192 (N_12192,N_10162,N_11037);
xor U12193 (N_12193,N_11248,N_10541);
nor U12194 (N_12194,N_11945,N_10446);
and U12195 (N_12195,N_11526,N_11534);
nand U12196 (N_12196,N_10189,N_10073);
or U12197 (N_12197,N_11727,N_10118);
or U12198 (N_12198,N_10828,N_11017);
nor U12199 (N_12199,N_11562,N_11638);
or U12200 (N_12200,N_10718,N_10212);
nor U12201 (N_12201,N_10394,N_11869);
nor U12202 (N_12202,N_11056,N_10068);
nor U12203 (N_12203,N_11473,N_10089);
xnor U12204 (N_12204,N_10256,N_11987);
or U12205 (N_12205,N_10740,N_10558);
or U12206 (N_12206,N_10246,N_11815);
or U12207 (N_12207,N_11415,N_10358);
nand U12208 (N_12208,N_11225,N_10264);
nand U12209 (N_12209,N_11818,N_10896);
nor U12210 (N_12210,N_11495,N_10045);
and U12211 (N_12211,N_11504,N_10331);
and U12212 (N_12212,N_10100,N_10576);
nand U12213 (N_12213,N_10871,N_11158);
nor U12214 (N_12214,N_11391,N_11761);
nand U12215 (N_12215,N_10181,N_11132);
xnor U12216 (N_12216,N_10691,N_11919);
xor U12217 (N_12217,N_10659,N_10554);
and U12218 (N_12218,N_11133,N_10986);
and U12219 (N_12219,N_11970,N_10537);
nor U12220 (N_12220,N_10147,N_11059);
nor U12221 (N_12221,N_10961,N_11055);
xnor U12222 (N_12222,N_11908,N_10337);
and U12223 (N_12223,N_10491,N_11688);
nor U12224 (N_12224,N_11333,N_11721);
nand U12225 (N_12225,N_10506,N_11253);
nor U12226 (N_12226,N_10092,N_10543);
nand U12227 (N_12227,N_11347,N_11732);
and U12228 (N_12228,N_11903,N_11718);
xor U12229 (N_12229,N_10292,N_11386);
nand U12230 (N_12230,N_11913,N_10461);
xor U12231 (N_12231,N_10735,N_11878);
xnor U12232 (N_12232,N_10155,N_11252);
nand U12233 (N_12233,N_10872,N_11673);
and U12234 (N_12234,N_10775,N_10329);
and U12235 (N_12235,N_10962,N_11413);
or U12236 (N_12236,N_11676,N_11752);
nand U12237 (N_12237,N_10965,N_10379);
or U12238 (N_12238,N_10344,N_11802);
nand U12239 (N_12239,N_10042,N_11563);
nor U12240 (N_12240,N_10188,N_11649);
nand U12241 (N_12241,N_11348,N_11326);
nand U12242 (N_12242,N_11665,N_11794);
nor U12243 (N_12243,N_11329,N_11617);
and U12244 (N_12244,N_11592,N_10430);
and U12245 (N_12245,N_10086,N_11493);
xor U12246 (N_12246,N_11641,N_10039);
nor U12247 (N_12247,N_11668,N_10255);
and U12248 (N_12248,N_11453,N_10268);
xor U12249 (N_12249,N_10575,N_11340);
and U12250 (N_12250,N_11308,N_10931);
nand U12251 (N_12251,N_10034,N_11687);
nor U12252 (N_12252,N_11816,N_11250);
nand U12253 (N_12253,N_11689,N_11324);
xor U12254 (N_12254,N_10485,N_11202);
nor U12255 (N_12255,N_11544,N_10489);
or U12256 (N_12256,N_10811,N_11207);
or U12257 (N_12257,N_11289,N_11619);
nor U12258 (N_12258,N_11146,N_10677);
nor U12259 (N_12259,N_11587,N_10227);
xor U12260 (N_12260,N_11672,N_10992);
or U12261 (N_12261,N_10359,N_10035);
xor U12262 (N_12262,N_11540,N_11773);
nor U12263 (N_12263,N_11932,N_11140);
and U12264 (N_12264,N_10243,N_10149);
and U12265 (N_12265,N_11644,N_11266);
xor U12266 (N_12266,N_11275,N_11051);
and U12267 (N_12267,N_10825,N_10630);
nor U12268 (N_12268,N_11443,N_10556);
nand U12269 (N_12269,N_10566,N_10049);
xnor U12270 (N_12270,N_10671,N_11934);
nand U12271 (N_12271,N_11098,N_10644);
and U12272 (N_12272,N_10405,N_10927);
nor U12273 (N_12273,N_11338,N_10050);
and U12274 (N_12274,N_10736,N_11165);
nand U12275 (N_12275,N_10051,N_10016);
or U12276 (N_12276,N_11772,N_10891);
xor U12277 (N_12277,N_10484,N_10102);
and U12278 (N_12278,N_10814,N_10517);
or U12279 (N_12279,N_10836,N_10892);
xor U12280 (N_12280,N_11246,N_10785);
and U12281 (N_12281,N_10682,N_11283);
xor U12282 (N_12282,N_10864,N_11826);
or U12283 (N_12283,N_10545,N_10464);
nor U12284 (N_12284,N_11837,N_11537);
nor U12285 (N_12285,N_11097,N_11066);
and U12286 (N_12286,N_11679,N_11249);
nor U12287 (N_12287,N_10751,N_10109);
and U12288 (N_12288,N_10589,N_11311);
xor U12289 (N_12289,N_11374,N_11977);
nor U12290 (N_12290,N_11314,N_10737);
and U12291 (N_12291,N_10360,N_10078);
nand U12292 (N_12292,N_11956,N_11709);
or U12293 (N_12293,N_10571,N_10572);
or U12294 (N_12294,N_10288,N_10395);
nand U12295 (N_12295,N_10901,N_10581);
nor U12296 (N_12296,N_11890,N_10631);
and U12297 (N_12297,N_11877,N_10830);
and U12298 (N_12298,N_11395,N_10082);
and U12299 (N_12299,N_11425,N_10474);
xnor U12300 (N_12300,N_11677,N_10435);
or U12301 (N_12301,N_11912,N_11190);
nor U12302 (N_12302,N_11403,N_11920);
nand U12303 (N_12303,N_10303,N_10144);
nor U12304 (N_12304,N_11897,N_11434);
nand U12305 (N_12305,N_10722,N_10721);
nand U12306 (N_12306,N_11611,N_10165);
nand U12307 (N_12307,N_11089,N_11393);
and U12308 (N_12308,N_10664,N_11109);
or U12309 (N_12309,N_10085,N_11560);
nand U12310 (N_12310,N_10192,N_10613);
xor U12311 (N_12311,N_11226,N_11260);
nor U12312 (N_12312,N_11463,N_10302);
nor U12313 (N_12313,N_11105,N_11949);
xor U12314 (N_12314,N_10250,N_11297);
and U12315 (N_12315,N_11503,N_11229);
nor U12316 (N_12316,N_11838,N_11141);
nor U12317 (N_12317,N_11119,N_10547);
nor U12318 (N_12318,N_11079,N_11624);
or U12319 (N_12319,N_10636,N_10401);
xnor U12320 (N_12320,N_10291,N_10080);
or U12321 (N_12321,N_10729,N_10819);
nand U12322 (N_12322,N_11223,N_11380);
and U12323 (N_12323,N_10112,N_10539);
xor U12324 (N_12324,N_10984,N_10625);
nand U12325 (N_12325,N_10333,N_10088);
nor U12326 (N_12326,N_10985,N_11136);
nor U12327 (N_12327,N_10148,N_11690);
nor U12328 (N_12328,N_10950,N_10741);
nor U12329 (N_12329,N_11103,N_11299);
nand U12330 (N_12330,N_11214,N_10289);
nand U12331 (N_12331,N_11086,N_10041);
nor U12332 (N_12332,N_11459,N_10060);
nand U12333 (N_12333,N_10209,N_10647);
and U12334 (N_12334,N_11754,N_11000);
xnor U12335 (N_12335,N_10308,N_10770);
nand U12336 (N_12336,N_11981,N_11510);
nor U12337 (N_12337,N_11930,N_11699);
or U12338 (N_12338,N_10947,N_10176);
or U12339 (N_12339,N_10287,N_10387);
nand U12340 (N_12340,N_10015,N_10483);
and U12341 (N_12341,N_10420,N_10530);
nor U12342 (N_12342,N_11458,N_10903);
and U12343 (N_12343,N_10119,N_10234);
nand U12344 (N_12344,N_10479,N_11478);
or U12345 (N_12345,N_10348,N_10204);
or U12346 (N_12346,N_10731,N_10138);
and U12347 (N_12347,N_10829,N_11880);
nand U12348 (N_12348,N_11159,N_10477);
or U12349 (N_12349,N_10454,N_11518);
and U12350 (N_12350,N_10708,N_10332);
nor U12351 (N_12351,N_10764,N_10507);
or U12352 (N_12352,N_11369,N_11963);
or U12353 (N_12353,N_11049,N_11697);
nand U12354 (N_12354,N_11470,N_11744);
nor U12355 (N_12355,N_10590,N_11024);
nor U12356 (N_12356,N_10527,N_11774);
and U12357 (N_12357,N_10555,N_11251);
nand U12358 (N_12358,N_10862,N_10327);
nand U12359 (N_12359,N_10347,N_10094);
nand U12360 (N_12360,N_11144,N_10253);
or U12361 (N_12361,N_10526,N_11775);
nand U12362 (N_12362,N_11543,N_11196);
and U12363 (N_12363,N_11788,N_10606);
nor U12364 (N_12364,N_11843,N_11356);
and U12365 (N_12365,N_11479,N_10179);
nor U12366 (N_12366,N_11444,N_10550);
nor U12367 (N_12367,N_11753,N_10481);
xnor U12368 (N_12368,N_11485,N_10486);
xor U12369 (N_12369,N_10216,N_10514);
or U12370 (N_12370,N_11698,N_11407);
nor U12371 (N_12371,N_10723,N_11035);
nor U12372 (N_12372,N_10193,N_10462);
xnor U12373 (N_12373,N_10419,N_10058);
nor U12374 (N_12374,N_11033,N_10542);
nor U12375 (N_12375,N_11860,N_11975);
xnor U12376 (N_12376,N_10587,N_11567);
or U12377 (N_12377,N_11354,N_10615);
or U12378 (N_12378,N_11789,N_10399);
nand U12379 (N_12379,N_11045,N_11723);
and U12380 (N_12380,N_10650,N_10503);
nor U12381 (N_12381,N_11278,N_10275);
nand U12382 (N_12382,N_11872,N_11870);
nor U12383 (N_12383,N_11342,N_10833);
or U12384 (N_12384,N_10714,N_11581);
and U12385 (N_12385,N_11855,N_11798);
or U12386 (N_12386,N_11694,N_11390);
xnor U12387 (N_12387,N_10579,N_10410);
nor U12388 (N_12388,N_11474,N_10011);
xor U12389 (N_12389,N_11865,N_10110);
and U12390 (N_12390,N_11131,N_10172);
nand U12391 (N_12391,N_11383,N_10588);
and U12392 (N_12392,N_11487,N_10652);
nor U12393 (N_12393,N_11336,N_10335);
nand U12394 (N_12394,N_11957,N_11653);
nand U12395 (N_12395,N_11005,N_10628);
and U12396 (N_12396,N_10404,N_11256);
or U12397 (N_12397,N_10334,N_11725);
nand U12398 (N_12398,N_10473,N_10578);
nor U12399 (N_12399,N_10767,N_11671);
nor U12400 (N_12400,N_11169,N_11613);
nand U12401 (N_12401,N_10433,N_11738);
nand U12402 (N_12402,N_10377,N_11070);
or U12403 (N_12403,N_10928,N_10698);
nor U12404 (N_12404,N_11467,N_10351);
nor U12405 (N_12405,N_10447,N_10028);
nor U12406 (N_12406,N_10126,N_11747);
and U12407 (N_12407,N_11588,N_10183);
or U12408 (N_12408,N_11388,N_10760);
nor U12409 (N_12409,N_11936,N_10910);
nand U12410 (N_12410,N_11481,N_10349);
nand U12411 (N_12411,N_10330,N_11823);
nor U12412 (N_12412,N_11511,N_10495);
nor U12413 (N_12413,N_10601,N_11931);
or U12414 (N_12414,N_10390,N_10709);
nor U12415 (N_12415,N_10705,N_10946);
nand U12416 (N_12416,N_10002,N_10801);
and U12417 (N_12417,N_11603,N_10129);
xnor U12418 (N_12418,N_10626,N_11763);
or U12419 (N_12419,N_11978,N_10371);
and U12420 (N_12420,N_10790,N_10104);
nand U12421 (N_12421,N_11923,N_10231);
nand U12422 (N_12422,N_11379,N_11628);
nor U12423 (N_12423,N_11776,N_11658);
and U12424 (N_12424,N_11087,N_10225);
and U12425 (N_12425,N_11714,N_11768);
nor U12426 (N_12426,N_11015,N_11824);
nor U12427 (N_12427,N_10346,N_10239);
nor U12428 (N_12428,N_10673,N_11359);
and U12429 (N_12429,N_10776,N_11242);
nand U12430 (N_12430,N_11437,N_10022);
nand U12431 (N_12431,N_10657,N_11236);
nand U12432 (N_12432,N_11411,N_10551);
and U12433 (N_12433,N_11468,N_10996);
and U12434 (N_12434,N_11536,N_10321);
or U12435 (N_12435,N_10971,N_11344);
nor U12436 (N_12436,N_10772,N_11656);
nand U12437 (N_12437,N_11655,N_10968);
or U12438 (N_12438,N_11166,N_11601);
xor U12439 (N_12439,N_11535,N_10294);
xor U12440 (N_12440,N_11408,N_10727);
nor U12441 (N_12441,N_11371,N_11269);
and U12442 (N_12442,N_11549,N_10815);
xor U12443 (N_12443,N_11599,N_11512);
or U12444 (N_12444,N_10224,N_10849);
or U12445 (N_12445,N_10339,N_11382);
or U12446 (N_12446,N_11439,N_11580);
nor U12447 (N_12447,N_10128,N_10918);
nand U12448 (N_12448,N_11040,N_10977);
and U12449 (N_12449,N_11343,N_10686);
and U12450 (N_12450,N_11322,N_10598);
and U12451 (N_12451,N_10687,N_11436);
or U12452 (N_12452,N_11889,N_11175);
xnor U12453 (N_12453,N_10970,N_10732);
and U12454 (N_12454,N_10866,N_10645);
and U12455 (N_12455,N_10840,N_11234);
nand U12456 (N_12456,N_10052,N_10750);
nor U12457 (N_12457,N_11704,N_10717);
nand U12458 (N_12458,N_11982,N_10418);
nor U12459 (N_12459,N_11701,N_11178);
nor U12460 (N_12460,N_10194,N_11492);
and U12461 (N_12461,N_11304,N_10765);
xnor U12462 (N_12462,N_11594,N_11106);
or U12463 (N_12463,N_11951,N_10949);
nor U12464 (N_12464,N_10789,N_11351);
nand U12465 (N_12465,N_11451,N_10392);
nor U12466 (N_12466,N_11996,N_11910);
nand U12467 (N_12467,N_10638,N_10762);
nor U12468 (N_12468,N_10055,N_10421);
or U12469 (N_12469,N_11528,N_11952);
or U12470 (N_12470,N_11799,N_10184);
or U12471 (N_12471,N_11983,N_10568);
or U12472 (N_12472,N_10411,N_11716);
or U12473 (N_12473,N_10983,N_11929);
nand U12474 (N_12474,N_11122,N_11968);
nor U12475 (N_12475,N_11227,N_11669);
xor U12476 (N_12476,N_11092,N_10995);
nand U12477 (N_12477,N_11813,N_11364);
nand U12478 (N_12478,N_11315,N_10646);
and U12479 (N_12479,N_10338,N_11466);
xor U12480 (N_12480,N_10323,N_11573);
xor U12481 (N_12481,N_11812,N_10385);
nand U12482 (N_12482,N_10005,N_11967);
or U12483 (N_12483,N_11245,N_10780);
or U12484 (N_12484,N_11272,N_10859);
and U12485 (N_12485,N_11874,N_11782);
nand U12486 (N_12486,N_10614,N_11235);
nor U12487 (N_12487,N_11871,N_10221);
or U12488 (N_12488,N_10604,N_10260);
nor U12489 (N_12489,N_10546,N_10911);
or U12490 (N_12490,N_11678,N_11427);
nor U12491 (N_12491,N_11680,N_10063);
and U12492 (N_12492,N_11186,N_11130);
nand U12493 (N_12493,N_10487,N_10637);
and U12494 (N_12494,N_10704,N_10175);
or U12495 (N_12495,N_11508,N_11593);
nand U12496 (N_12496,N_10569,N_11216);
xnor U12497 (N_12497,N_10700,N_11244);
or U12498 (N_12498,N_10935,N_10934);
nor U12499 (N_12499,N_10929,N_10838);
nand U12500 (N_12500,N_11757,N_10185);
or U12501 (N_12501,N_11400,N_11433);
or U12502 (N_12502,N_11507,N_11334);
nor U12503 (N_12503,N_10832,N_10009);
or U12504 (N_12504,N_11971,N_10047);
and U12505 (N_12505,N_11846,N_11305);
or U12506 (N_12506,N_11734,N_11188);
and U12507 (N_12507,N_10355,N_10973);
nand U12508 (N_12508,N_11145,N_10672);
and U12509 (N_12509,N_10043,N_11396);
xor U12510 (N_12510,N_11084,N_11465);
or U12511 (N_12511,N_10922,N_11328);
xor U12512 (N_12512,N_11582,N_10867);
nand U12513 (N_12513,N_11985,N_10689);
nand U12514 (N_12514,N_10898,N_10053);
or U12515 (N_12515,N_10612,N_11088);
nand U12516 (N_12516,N_10567,N_10019);
nand U12517 (N_12517,N_11490,N_11924);
and U12518 (N_12518,N_11946,N_10813);
or U12519 (N_12519,N_11955,N_10795);
nand U12520 (N_12520,N_11268,N_11839);
and U12521 (N_12521,N_10916,N_11729);
or U12522 (N_12522,N_10257,N_10653);
nand U12523 (N_12523,N_11288,N_11712);
and U12524 (N_12524,N_10214,N_10573);
nor U12525 (N_12525,N_10743,N_11155);
or U12526 (N_12526,N_11488,N_10939);
or U12527 (N_12527,N_11640,N_10450);
and U12528 (N_12528,N_10356,N_11025);
xnor U12529 (N_12529,N_11999,N_11091);
or U12530 (N_12530,N_10694,N_11501);
nand U12531 (N_12531,N_10492,N_10081);
xor U12532 (N_12532,N_11533,N_10870);
or U12533 (N_12533,N_11513,N_10161);
nor U12534 (N_12534,N_11856,N_11247);
and U12535 (N_12535,N_10402,N_11938);
or U12536 (N_12536,N_10880,N_10997);
and U12537 (N_12537,N_11111,N_11550);
and U12538 (N_12538,N_11976,N_11349);
or U12539 (N_12539,N_10875,N_10326);
or U12540 (N_12540,N_10794,N_11509);
and U12541 (N_12541,N_10560,N_11979);
xor U12542 (N_12542,N_11829,N_11625);
xnor U12543 (N_12543,N_11094,N_11270);
or U12544 (N_12544,N_10549,N_11505);
nor U12545 (N_12545,N_11642,N_10413);
and U12546 (N_12546,N_11590,N_10376);
or U12547 (N_12547,N_10914,N_10877);
xor U12548 (N_12548,N_10297,N_10817);
nor U12549 (N_12549,N_10810,N_11210);
and U12550 (N_12550,N_11394,N_10915);
or U12551 (N_12551,N_11596,N_11237);
nand U12552 (N_12552,N_10639,N_11189);
nand U12553 (N_12553,N_11046,N_11372);
nand U12554 (N_12554,N_10444,N_11489);
xnor U12555 (N_12555,N_10675,N_10299);
or U12556 (N_12556,N_10908,N_10400);
and U12557 (N_12557,N_11884,N_11997);
or U12558 (N_12558,N_10610,N_10133);
or U12559 (N_12559,N_10561,N_10834);
nand U12560 (N_12560,N_10023,N_11817);
nand U12561 (N_12561,N_10759,N_11139);
and U12562 (N_12562,N_11651,N_10074);
and U12563 (N_12563,N_10756,N_10707);
and U12564 (N_12564,N_10265,N_11445);
and U12565 (N_12565,N_10024,N_10114);
xor U12566 (N_12566,N_10123,N_11793);
nand U12567 (N_12567,N_10437,N_11454);
nor U12568 (N_12568,N_10111,N_10690);
nor U12569 (N_12569,N_11398,N_11373);
nand U12570 (N_12570,N_11038,N_10067);
and U12571 (N_12571,N_10804,N_11523);
xnor U12572 (N_12572,N_11461,N_11389);
or U12573 (N_12573,N_11820,N_11630);
nor U12574 (N_12574,N_11900,N_10213);
and U12575 (N_12575,N_10203,N_11287);
and U12576 (N_12576,N_11496,N_11646);
nor U12577 (N_12577,N_10820,N_11683);
xor U12578 (N_12578,N_10315,N_10314);
nor U12579 (N_12579,N_11864,N_10522);
or U12580 (N_12580,N_11853,N_10963);
nand U12581 (N_12581,N_10163,N_10065);
and U12582 (N_12582,N_11241,N_10252);
nor U12583 (N_12583,N_10917,N_11643);
nand U12584 (N_12584,N_10310,N_10808);
xor U12585 (N_12585,N_10622,N_11401);
xnor U12586 (N_12586,N_10964,N_10186);
nand U12587 (N_12587,N_10684,N_11472);
xnor U12588 (N_12588,N_11341,N_11693);
and U12589 (N_12589,N_10223,N_10431);
nand U12590 (N_12590,N_11597,N_11110);
or U12591 (N_12591,N_10749,N_10432);
or U12592 (N_12592,N_11455,N_10670);
nand U12593 (N_12593,N_11261,N_10976);
nand U12594 (N_12594,N_11561,N_10124);
or U12595 (N_12595,N_10150,N_11053);
nor U12596 (N_12596,N_11147,N_10651);
or U12597 (N_12597,N_11748,N_11654);
xnor U12598 (N_12598,N_11264,N_11663);
nand U12599 (N_12599,N_11695,N_10648);
nand U12600 (N_12600,N_11857,N_10407);
and U12601 (N_12601,N_11809,N_10784);
and U12602 (N_12602,N_10467,N_10649);
and U12603 (N_12603,N_10296,N_11514);
or U12604 (N_12604,N_10279,N_11265);
nand U12605 (N_12605,N_10027,N_11362);
nor U12606 (N_12606,N_11984,N_10937);
and U12607 (N_12607,N_10957,N_10244);
or U12608 (N_12608,N_11023,N_10769);
and U12609 (N_12609,N_10125,N_10199);
nor U12610 (N_12610,N_11521,N_11102);
xor U12611 (N_12611,N_11303,N_10548);
and U12612 (N_12612,N_10070,N_10594);
nor U12613 (N_12613,N_10196,N_11043);
nand U12614 (N_12614,N_10616,N_11569);
nand U12615 (N_12615,N_11875,N_11352);
nor U12616 (N_12616,N_10201,N_11279);
xnor U12617 (N_12617,N_11200,N_11947);
or U12618 (N_12618,N_10251,N_10734);
or U12619 (N_12619,N_11424,N_10017);
nor U12620 (N_12620,N_10064,N_11355);
nor U12621 (N_12621,N_10151,N_10974);
or U12622 (N_12622,N_10079,N_10809);
nand U12623 (N_12623,N_11031,N_11370);
nand U12624 (N_12624,N_10021,N_11168);
and U12625 (N_12625,N_11933,N_11061);
nand U12626 (N_12626,N_11367,N_10136);
and U12627 (N_12627,N_11844,N_11179);
nand U12628 (N_12628,N_10697,N_11879);
and U12629 (N_12629,N_10991,N_11153);
and U12630 (N_12630,N_10174,N_11052);
xor U12631 (N_12631,N_10847,N_10159);
nand U12632 (N_12632,N_10624,N_11267);
nand U12633 (N_12633,N_10443,N_11014);
and U12634 (N_12634,N_10375,N_11499);
nor U12635 (N_12635,N_11350,N_10211);
or U12636 (N_12636,N_11327,N_10902);
nand U12637 (N_12637,N_10007,N_10515);
nand U12638 (N_12638,N_11616,N_11421);
nor U12639 (N_12639,N_10499,N_10846);
or U12640 (N_12640,N_10951,N_10843);
and U12641 (N_12641,N_10425,N_11047);
nor U12642 (N_12642,N_11441,N_10868);
or U12643 (N_12643,N_11986,N_10907);
and U12644 (N_12644,N_11781,N_10720);
xnor U12645 (N_12645,N_11211,N_10856);
nor U12646 (N_12646,N_11399,N_11719);
and U12647 (N_12647,N_11006,N_11579);
nand U12648 (N_12648,N_10178,N_11330);
or U12649 (N_12649,N_11312,N_11702);
nor U12650 (N_12650,N_10456,N_10198);
or U12651 (N_12651,N_11476,N_10887);
or U12652 (N_12652,N_11310,N_11615);
nand U12653 (N_12653,N_11529,N_11360);
xnor U12654 (N_12654,N_10097,N_11965);
or U12655 (N_12655,N_11614,N_11787);
and U12656 (N_12656,N_11539,N_11585);
and U12657 (N_12657,N_10706,N_10448);
and U12658 (N_12658,N_11764,N_10683);
or U12659 (N_12659,N_11565,N_11435);
nor U12660 (N_12660,N_10975,N_10955);
or U12661 (N_12661,N_10956,N_11790);
or U12662 (N_12662,N_11605,N_11859);
or U12663 (N_12663,N_11609,N_11792);
or U12664 (N_12664,N_10069,N_11353);
nor U12665 (N_12665,N_10132,N_10618);
xnor U12666 (N_12666,N_11080,N_10270);
nand U12667 (N_12667,N_10010,N_11286);
nor U12668 (N_12668,N_10533,N_10978);
or U12669 (N_12669,N_10583,N_10472);
nor U12670 (N_12670,N_10197,N_10353);
or U12671 (N_12671,N_11576,N_11161);
nand U12672 (N_12672,N_11626,N_11064);
and U12673 (N_12673,N_11618,N_11610);
or U12674 (N_12674,N_10103,N_10895);
nor U12675 (N_12675,N_10501,N_11595);
or U12676 (N_12676,N_10428,N_10030);
nand U12677 (N_12677,N_11807,N_11003);
and U12678 (N_12678,N_10696,N_11691);
or U12679 (N_12679,N_11176,N_11076);
and U12680 (N_12680,N_11274,N_11375);
nand U12681 (N_12681,N_10274,N_11730);
nor U12682 (N_12682,N_11715,N_11733);
xor U12683 (N_12683,N_10524,N_10266);
nor U12684 (N_12684,N_11325,N_11602);
xnor U12685 (N_12685,N_10863,N_10445);
or U12686 (N_12686,N_11700,N_10115);
and U12687 (N_12687,N_11778,N_11058);
nand U12688 (N_12688,N_10823,N_11307);
or U12689 (N_12689,N_10841,N_11566);
nor U12690 (N_12690,N_11173,N_11182);
nor U12691 (N_12691,N_11516,N_11163);
nand U12692 (N_12692,N_10054,N_10033);
or U12693 (N_12693,N_11538,N_11822);
nand U12694 (N_12694,N_11108,N_11377);
nand U12695 (N_12695,N_10510,N_11068);
or U12696 (N_12696,N_10999,N_11477);
or U12697 (N_12697,N_11848,N_11420);
nand U12698 (N_12698,N_10712,N_11765);
and U12699 (N_12699,N_10458,N_10281);
and U12700 (N_12700,N_10883,N_11332);
and U12701 (N_12701,N_11808,N_10020);
nand U12702 (N_12702,N_11825,N_11124);
xnor U12703 (N_12703,N_10654,N_10678);
and U12704 (N_12704,N_10500,N_11128);
or U12705 (N_12705,N_10127,N_10669);
xor U12706 (N_12706,N_10158,N_10782);
nor U12707 (N_12707,N_11797,N_10855);
nand U12708 (N_12708,N_10306,N_11240);
nor U12709 (N_12709,N_11546,N_10807);
nand U12710 (N_12710,N_10923,N_11029);
or U12711 (N_12711,N_11572,N_11958);
and U12712 (N_12712,N_10318,N_11482);
and U12713 (N_12713,N_10874,N_10725);
nor U12714 (N_12714,N_10336,N_11886);
or U12715 (N_12715,N_10886,N_10465);
nor U12716 (N_12716,N_10309,N_11647);
xnor U12717 (N_12717,N_10342,N_10076);
and U12718 (N_12718,N_11604,N_10498);
nand U12719 (N_12719,N_10688,N_10438);
nor U12720 (N_12720,N_11071,N_11319);
nor U12721 (N_12721,N_10171,N_10180);
xor U12722 (N_12722,N_11942,N_11450);
or U12723 (N_12723,N_11722,N_10083);
or U12724 (N_12724,N_10656,N_10460);
nor U12725 (N_12725,N_10381,N_11090);
or U12726 (N_12726,N_10821,N_11779);
nand U12727 (N_12727,N_10313,N_11584);
and U12728 (N_12728,N_11814,N_10884);
nor U12729 (N_12729,N_11423,N_11365);
or U12730 (N_12730,N_10959,N_11854);
or U12731 (N_12731,N_11703,N_11995);
or U12732 (N_12732,N_10004,N_10666);
and U12733 (N_12733,N_11960,N_11357);
xor U12734 (N_12734,N_10861,N_11558);
nor U12735 (N_12735,N_11429,N_11972);
nor U12736 (N_12736,N_10107,N_10468);
or U12737 (N_12737,N_10692,N_11831);
or U12738 (N_12738,N_10562,N_10046);
nand U12739 (N_12739,N_11650,N_11612);
nor U12740 (N_12740,N_10304,N_10844);
or U12741 (N_12741,N_11717,N_11800);
nand U12742 (N_12742,N_10777,N_11635);
nand U12743 (N_12743,N_10142,N_11187);
nor U12744 (N_12744,N_10812,N_11830);
and U12745 (N_12745,N_11331,N_11221);
nand U12746 (N_12746,N_10531,N_11527);
nand U12747 (N_12747,N_10781,N_11121);
and U12748 (N_12748,N_11667,N_10897);
nand U12749 (N_12749,N_10130,N_11785);
or U12750 (N_12750,N_11416,N_11440);
nor U12751 (N_12751,N_11713,N_10860);
nand U12752 (N_12752,N_11457,N_10439);
or U12753 (N_12753,N_10452,N_11921);
or U12754 (N_12754,N_10090,N_11570);
nor U12755 (N_12755,N_10793,N_10758);
nor U12756 (N_12756,N_11452,N_11806);
nor U12757 (N_12757,N_11627,N_10040);
and U12758 (N_12758,N_10890,N_10989);
and U12759 (N_12759,N_10135,N_10143);
nand U12760 (N_12760,N_10987,N_10469);
nor U12761 (N_12761,N_11805,N_10512);
or U12762 (N_12762,N_11633,N_11104);
xor U12763 (N_12763,N_10494,N_11771);
nand U12764 (N_12764,N_11885,N_11232);
nand U12765 (N_12765,N_11928,N_11197);
and U12766 (N_12766,N_10818,N_11706);
or U12767 (N_12767,N_11172,N_11301);
and U12768 (N_12768,N_10609,N_11637);
or U12769 (N_12769,N_10424,N_10711);
and U12770 (N_12770,N_10699,N_10882);
and U12771 (N_12771,N_11935,N_11735);
xnor U12772 (N_12772,N_10230,N_10852);
or U12773 (N_12773,N_11171,N_11542);
or U12774 (N_12774,N_11740,N_10921);
and U12775 (N_12775,N_10284,N_10301);
or U12776 (N_12776,N_11181,N_11917);
nand U12777 (N_12777,N_10889,N_10945);
or U12778 (N_12778,N_11598,N_11948);
nand U12779 (N_12779,N_10981,N_10378);
nand U12780 (N_12780,N_10061,N_11083);
or U12781 (N_12781,N_11001,N_10783);
or U12782 (N_12782,N_10490,N_10909);
nand U12783 (N_12783,N_11069,N_10746);
nor U12784 (N_12784,N_10345,N_11803);
xnor U12785 (N_12785,N_10012,N_10632);
xor U12786 (N_12786,N_10343,N_11907);
and U12787 (N_12787,N_10406,N_11674);
nand U12788 (N_12788,N_11524,N_10516);
nor U12789 (N_12789,N_10570,N_11462);
and U12790 (N_12790,N_11358,N_10357);
nand U12791 (N_12791,N_11832,N_11483);
nand U12792 (N_12792,N_10029,N_11522);
nand U12793 (N_12793,N_11387,N_10322);
and U12794 (N_12794,N_11497,N_10954);
or U12795 (N_12795,N_10948,N_11840);
nor U12796 (N_12796,N_10441,N_10470);
nor U12797 (N_12797,N_11993,N_10228);
xor U12798 (N_12798,N_11404,N_10620);
or U12799 (N_12799,N_10374,N_11620);
nand U12800 (N_12800,N_11022,N_10240);
xnor U12801 (N_12801,N_10312,N_10873);
or U12802 (N_12802,N_10099,N_10156);
or U12803 (N_12803,N_10894,N_11909);
nor U12804 (N_12804,N_10538,N_10635);
and U12805 (N_12805,N_11239,N_10403);
and U12806 (N_12806,N_10865,N_11746);
or U12807 (N_12807,N_10153,N_10320);
or U12808 (N_12808,N_10215,N_10940);
nor U12809 (N_12809,N_10457,N_10998);
xor U12810 (N_12810,N_11564,N_11780);
nor U12811 (N_12811,N_11969,N_10553);
and U12812 (N_12812,N_11766,N_10565);
and U12813 (N_12813,N_10608,N_10453);
or U12814 (N_12814,N_10031,N_10802);
and U12815 (N_12815,N_10241,N_10480);
nor U12816 (N_12816,N_10071,N_10850);
or U12817 (N_12817,N_11795,N_11448);
and U12818 (N_12818,N_11456,N_11783);
xor U12819 (N_12819,N_10774,N_11954);
nand U12820 (N_12820,N_10857,N_11096);
or U12821 (N_12821,N_10634,N_10640);
nand U12822 (N_12822,N_11224,N_10267);
xnor U12823 (N_12823,N_10878,N_11777);
nand U12824 (N_12824,N_11160,N_11545);
nand U12825 (N_12825,N_11074,N_11756);
nand U12826 (N_12826,N_11666,N_10325);
xor U12827 (N_12827,N_11750,N_10449);
and U12828 (N_12828,N_11974,N_10237);
or U12829 (N_12829,N_11368,N_11743);
nor U12830 (N_12830,N_11902,N_11728);
and U12831 (N_12831,N_11944,N_11447);
or U12832 (N_12832,N_11556,N_11112);
and U12833 (N_12833,N_10661,N_11021);
nor U12834 (N_12834,N_11174,N_11291);
or U12835 (N_12835,N_10559,N_10451);
and U12836 (N_12836,N_11238,N_10837);
or U12837 (N_12837,N_10157,N_11126);
nor U12838 (N_12838,N_10208,N_10747);
or U12839 (N_12839,N_10408,N_10791);
or U12840 (N_12840,N_11904,N_11767);
and U12841 (N_12841,N_10967,N_10236);
or U12842 (N_12842,N_10752,N_11036);
or U12843 (N_12843,N_11378,N_10429);
nor U12844 (N_12844,N_10858,N_11381);
and U12845 (N_12845,N_10120,N_10730);
or U12846 (N_12846,N_10072,N_10271);
nor U12847 (N_12847,N_11217,N_11193);
and U12848 (N_12848,N_10008,N_10733);
or U12849 (N_12849,N_10535,N_10933);
nor U12850 (N_12850,N_11645,N_11418);
or U12851 (N_12851,N_11195,N_11257);
and U12852 (N_12852,N_10248,N_10534);
nor U12853 (N_12853,N_11093,N_11600);
nand U12854 (N_12854,N_10580,N_10574);
nor U12855 (N_12855,N_11295,N_11804);
nor U12856 (N_12856,N_10210,N_10106);
nor U12857 (N_12857,N_10925,N_11922);
nand U12858 (N_12858,N_11762,N_11940);
or U12859 (N_12859,N_11302,N_10899);
xnor U12860 (N_12860,N_11784,N_11583);
and U12861 (N_12861,N_11410,N_10173);
nor U12862 (N_12862,N_10520,N_10131);
xor U12863 (N_12863,N_11243,N_11316);
nor U12864 (N_12864,N_11215,N_11219);
nand U12865 (N_12865,N_10121,N_10761);
nand U12866 (N_12866,N_10938,N_10427);
or U12867 (N_12867,N_10113,N_11095);
xor U12868 (N_12868,N_11117,N_11081);
or U12869 (N_12869,N_11648,N_10442);
nand U12870 (N_12870,N_10384,N_11961);
and U12871 (N_12871,N_11115,N_10822);
nor U12872 (N_12872,N_11914,N_11905);
nor U12873 (N_12873,N_11028,N_10972);
or U12874 (N_12874,N_11120,N_10164);
and U12875 (N_12875,N_11201,N_11417);
and U12876 (N_12876,N_10757,N_10235);
nand U12877 (N_12877,N_11621,N_10278);
nand U12878 (N_12878,N_10876,N_10904);
or U12879 (N_12879,N_10362,N_10742);
or U12880 (N_12880,N_11010,N_10412);
nand U12881 (N_12881,N_10509,N_11770);
nand U12882 (N_12882,N_11557,N_11555);
or U12883 (N_12883,N_10893,N_10680);
or U12884 (N_12884,N_11078,N_10247);
nor U12885 (N_12885,N_10195,N_11280);
nand U12886 (N_12886,N_11460,N_11199);
nor U12887 (N_12887,N_10245,N_11306);
or U12888 (N_12888,N_11134,N_11019);
nor U12889 (N_12889,N_11152,N_11142);
or U12890 (N_12890,N_10269,N_10273);
nand U12891 (N_12891,N_11231,N_10409);
nor U12892 (N_12892,N_10364,N_10994);
or U12893 (N_12893,N_11742,N_10586);
or U12894 (N_12894,N_10389,N_10693);
xor U12895 (N_12895,N_11271,N_11137);
nand U12896 (N_12896,N_11384,N_11498);
and U12897 (N_12897,N_11292,N_10831);
or U12898 (N_12898,N_10766,N_11363);
nor U12899 (N_12899,N_11255,N_10205);
nand U12900 (N_12900,N_11842,N_11067);
and U12901 (N_12901,N_10476,N_10505);
nor U12902 (N_12902,N_11623,N_10018);
or U12903 (N_12903,N_11048,N_11893);
nor U12904 (N_12904,N_10745,N_10835);
nand U12905 (N_12905,N_10482,N_10478);
or U12906 (N_12906,N_11402,N_11480);
or U12907 (N_12907,N_11164,N_10261);
or U12908 (N_12908,N_10415,N_11290);
nor U12909 (N_12909,N_11916,N_11998);
or U12910 (N_12910,N_11531,N_10152);
or U12911 (N_12911,N_11873,N_10919);
or U12912 (N_12912,N_11011,N_10848);
nand U12913 (N_12913,N_11309,N_11205);
and U12914 (N_12914,N_10232,N_10370);
xor U12915 (N_12915,N_10932,N_10003);
or U12916 (N_12916,N_11085,N_11259);
or U12917 (N_12917,N_11042,N_10674);
and U12918 (N_12918,N_11852,N_11323);
or U12919 (N_12919,N_10319,N_11077);
nor U12920 (N_12920,N_10066,N_10788);
xnor U12921 (N_12921,N_10038,N_10577);
nor U12922 (N_12922,N_11636,N_10363);
xor U12923 (N_12923,N_11834,N_10715);
or U12924 (N_12924,N_10373,N_10900);
nand U12925 (N_12925,N_10324,N_10511);
or U12926 (N_12926,N_10879,N_10249);
and U12927 (N_12927,N_11030,N_11170);
nand U12928 (N_12928,N_10826,N_10842);
and U12929 (N_12929,N_10096,N_11841);
nand U12930 (N_12930,N_10508,N_11469);
and U12931 (N_12931,N_10936,N_11007);
or U12932 (N_12932,N_10242,N_11696);
nand U12933 (N_12933,N_10350,N_10361);
nand U12934 (N_12934,N_10599,N_11867);
nand U12935 (N_12935,N_10290,N_11263);
xnor U12936 (N_12936,N_10719,N_11629);
nand U12937 (N_12937,N_11894,N_10816);
nand U12938 (N_12938,N_10105,N_10388);
or U12939 (N_12939,N_11707,N_10502);
and U12940 (N_12940,N_10792,N_11980);
xor U12941 (N_12941,N_10960,N_10623);
and U12942 (N_12942,N_10493,N_10605);
nand U12943 (N_12943,N_11162,N_11574);
nand U12944 (N_12944,N_11710,N_11950);
and U12945 (N_12945,N_11657,N_10383);
nand U12946 (N_12946,N_10134,N_11835);
nor U12947 (N_12947,N_10523,N_11502);
nor U12948 (N_12948,N_11198,N_11191);
and U12949 (N_12949,N_10160,N_10806);
nand U12950 (N_12950,N_11321,N_11277);
and U12951 (N_12951,N_10854,N_10305);
nand U12952 (N_12952,N_11298,N_10993);
nand U12953 (N_12953,N_11345,N_11887);
and U12954 (N_12954,N_10280,N_11926);
and U12955 (N_12955,N_10518,N_11850);
nand U12956 (N_12956,N_11607,N_10282);
nand U12957 (N_12957,N_11107,N_10755);
nand U12958 (N_12958,N_10436,N_11686);
xnor U12959 (N_12959,N_10341,N_11180);
nor U12960 (N_12960,N_10414,N_11801);
and U12961 (N_12961,N_11057,N_11953);
nor U12962 (N_12962,N_10233,N_10642);
and U12963 (N_12963,N_11675,N_10471);
nor U12964 (N_12964,N_11430,N_10380);
or U12965 (N_12965,N_10077,N_11883);
nor U12966 (N_12966,N_11720,N_10422);
nor U12967 (N_12967,N_11192,N_11895);
and U12968 (N_12968,N_11548,N_10738);
nor U12969 (N_12969,N_11966,N_10888);
or U12970 (N_12970,N_11577,N_10603);
nand U12971 (N_12971,N_10036,N_11376);
nand U12972 (N_12972,N_11065,N_10532);
nand U12973 (N_12973,N_11575,N_11811);
or U12974 (N_12974,N_11154,N_10276);
or U12975 (N_12975,N_11682,N_10611);
xor U12976 (N_12976,N_10352,N_11849);
xor U12977 (N_12977,N_11589,N_10753);
nor U12978 (N_12978,N_11073,N_11705);
and U12979 (N_12979,N_11183,N_11100);
nor U12980 (N_12980,N_11532,N_11973);
or U12981 (N_12981,N_11099,N_10779);
nor U12982 (N_12982,N_11758,N_10926);
xor U12983 (N_12983,N_11571,N_10667);
xnor U12984 (N_12984,N_11282,N_10286);
xor U12985 (N_12985,N_10913,N_10540);
and U12986 (N_12986,N_11075,N_10340);
or U12987 (N_12987,N_11760,N_10366);
nand U12988 (N_12988,N_10218,N_10582);
nand U12989 (N_12989,N_11759,N_11138);
and U12990 (N_12990,N_10552,N_10191);
nor U12991 (N_12991,N_11063,N_11184);
nand U12992 (N_12992,N_11992,N_11157);
nand U12993 (N_12993,N_11412,N_10525);
nor U12994 (N_12994,N_11819,N_10655);
or U12995 (N_12995,N_11018,N_11962);
or U12996 (N_12996,N_11828,N_10803);
and U12997 (N_12997,N_11273,N_11016);
nor U12998 (N_12998,N_11708,N_10643);
or U12999 (N_12999,N_10521,N_10145);
nor U13000 (N_13000,N_10104,N_10820);
or U13001 (N_13001,N_10158,N_10991);
and U13002 (N_13002,N_10785,N_10113);
and U13003 (N_13003,N_11687,N_10517);
and U13004 (N_13004,N_11998,N_10837);
or U13005 (N_13005,N_10937,N_10290);
or U13006 (N_13006,N_11651,N_11250);
nor U13007 (N_13007,N_10062,N_11377);
xor U13008 (N_13008,N_10369,N_11261);
nor U13009 (N_13009,N_11182,N_11964);
nor U13010 (N_13010,N_11996,N_11745);
or U13011 (N_13011,N_11676,N_10409);
or U13012 (N_13012,N_10472,N_11822);
nand U13013 (N_13013,N_11922,N_11688);
nand U13014 (N_13014,N_10979,N_11363);
or U13015 (N_13015,N_11436,N_11625);
or U13016 (N_13016,N_10317,N_11366);
or U13017 (N_13017,N_11548,N_11051);
and U13018 (N_13018,N_11500,N_11123);
and U13019 (N_13019,N_10995,N_11895);
nor U13020 (N_13020,N_10089,N_10169);
nor U13021 (N_13021,N_11867,N_11101);
and U13022 (N_13022,N_11995,N_11994);
xnor U13023 (N_13023,N_11168,N_10115);
xor U13024 (N_13024,N_11880,N_11460);
nand U13025 (N_13025,N_11633,N_10549);
and U13026 (N_13026,N_11495,N_10337);
nor U13027 (N_13027,N_11008,N_10877);
nand U13028 (N_13028,N_11491,N_10975);
and U13029 (N_13029,N_10539,N_11269);
nand U13030 (N_13030,N_10266,N_11537);
nand U13031 (N_13031,N_11791,N_11582);
nor U13032 (N_13032,N_10481,N_10407);
nor U13033 (N_13033,N_10506,N_10848);
xnor U13034 (N_13034,N_10895,N_10424);
or U13035 (N_13035,N_10970,N_11700);
or U13036 (N_13036,N_11516,N_11100);
xor U13037 (N_13037,N_11078,N_10221);
and U13038 (N_13038,N_10812,N_10049);
and U13039 (N_13039,N_11105,N_10795);
nor U13040 (N_13040,N_10386,N_11270);
or U13041 (N_13041,N_10800,N_10375);
or U13042 (N_13042,N_11845,N_11590);
or U13043 (N_13043,N_10990,N_10096);
nor U13044 (N_13044,N_11314,N_11845);
or U13045 (N_13045,N_11516,N_10657);
nor U13046 (N_13046,N_10197,N_11932);
nand U13047 (N_13047,N_10039,N_11661);
xnor U13048 (N_13048,N_10712,N_10434);
nand U13049 (N_13049,N_10595,N_10630);
and U13050 (N_13050,N_11727,N_11729);
nand U13051 (N_13051,N_11951,N_10570);
nor U13052 (N_13052,N_11051,N_11728);
nor U13053 (N_13053,N_11874,N_11224);
or U13054 (N_13054,N_10585,N_10428);
and U13055 (N_13055,N_10328,N_11714);
or U13056 (N_13056,N_10774,N_11108);
or U13057 (N_13057,N_10680,N_11120);
and U13058 (N_13058,N_11214,N_10884);
xnor U13059 (N_13059,N_11834,N_11378);
nor U13060 (N_13060,N_11960,N_10606);
nand U13061 (N_13061,N_10255,N_10820);
xnor U13062 (N_13062,N_11289,N_11583);
or U13063 (N_13063,N_10300,N_10715);
xor U13064 (N_13064,N_10760,N_11213);
or U13065 (N_13065,N_10915,N_10602);
nand U13066 (N_13066,N_11852,N_10467);
or U13067 (N_13067,N_11912,N_10104);
and U13068 (N_13068,N_11303,N_10283);
nor U13069 (N_13069,N_11655,N_10731);
nor U13070 (N_13070,N_10478,N_10346);
and U13071 (N_13071,N_10373,N_11565);
nor U13072 (N_13072,N_11195,N_10590);
or U13073 (N_13073,N_10568,N_11499);
and U13074 (N_13074,N_11663,N_11649);
or U13075 (N_13075,N_11667,N_10562);
or U13076 (N_13076,N_11113,N_11150);
and U13077 (N_13077,N_11778,N_11373);
xnor U13078 (N_13078,N_11263,N_10548);
nor U13079 (N_13079,N_11765,N_11647);
nand U13080 (N_13080,N_11335,N_11847);
or U13081 (N_13081,N_10096,N_11713);
or U13082 (N_13082,N_10486,N_11625);
or U13083 (N_13083,N_11152,N_10598);
nor U13084 (N_13084,N_11979,N_11021);
and U13085 (N_13085,N_10412,N_11358);
and U13086 (N_13086,N_11826,N_11788);
nor U13087 (N_13087,N_10352,N_11516);
nor U13088 (N_13088,N_10721,N_10312);
xnor U13089 (N_13089,N_10418,N_10747);
nand U13090 (N_13090,N_11150,N_11810);
nand U13091 (N_13091,N_10751,N_10778);
nand U13092 (N_13092,N_10541,N_11100);
or U13093 (N_13093,N_11905,N_10550);
nand U13094 (N_13094,N_11352,N_10628);
nor U13095 (N_13095,N_10656,N_10564);
and U13096 (N_13096,N_11354,N_11838);
or U13097 (N_13097,N_11845,N_10445);
or U13098 (N_13098,N_10296,N_11981);
nor U13099 (N_13099,N_10017,N_10051);
xor U13100 (N_13100,N_11879,N_11956);
or U13101 (N_13101,N_10627,N_10649);
or U13102 (N_13102,N_10235,N_10490);
nor U13103 (N_13103,N_11817,N_10734);
or U13104 (N_13104,N_10949,N_11071);
or U13105 (N_13105,N_10082,N_11094);
nor U13106 (N_13106,N_11598,N_11663);
nand U13107 (N_13107,N_11819,N_10933);
and U13108 (N_13108,N_10091,N_10834);
and U13109 (N_13109,N_10054,N_11774);
nand U13110 (N_13110,N_11061,N_11911);
and U13111 (N_13111,N_10747,N_10209);
nand U13112 (N_13112,N_10127,N_11088);
and U13113 (N_13113,N_10630,N_10535);
nor U13114 (N_13114,N_11671,N_11876);
xor U13115 (N_13115,N_11751,N_10744);
nor U13116 (N_13116,N_11001,N_10219);
or U13117 (N_13117,N_10397,N_10026);
nand U13118 (N_13118,N_10213,N_11841);
or U13119 (N_13119,N_10910,N_11194);
xnor U13120 (N_13120,N_11179,N_11331);
nor U13121 (N_13121,N_11614,N_10021);
or U13122 (N_13122,N_11148,N_10276);
and U13123 (N_13123,N_11808,N_11784);
and U13124 (N_13124,N_11789,N_11480);
xor U13125 (N_13125,N_11669,N_11381);
nand U13126 (N_13126,N_10661,N_11241);
and U13127 (N_13127,N_10252,N_11912);
nor U13128 (N_13128,N_10421,N_10907);
or U13129 (N_13129,N_11797,N_10028);
and U13130 (N_13130,N_11713,N_10287);
nor U13131 (N_13131,N_11402,N_10687);
or U13132 (N_13132,N_10548,N_11867);
xnor U13133 (N_13133,N_10007,N_11927);
nor U13134 (N_13134,N_10785,N_11540);
nand U13135 (N_13135,N_11869,N_10371);
and U13136 (N_13136,N_10203,N_10217);
nand U13137 (N_13137,N_11028,N_11898);
or U13138 (N_13138,N_10465,N_11252);
nor U13139 (N_13139,N_11011,N_10886);
nand U13140 (N_13140,N_10722,N_10756);
xnor U13141 (N_13141,N_11717,N_11301);
and U13142 (N_13142,N_10994,N_11687);
nor U13143 (N_13143,N_11431,N_11926);
xor U13144 (N_13144,N_11667,N_10182);
or U13145 (N_13145,N_11737,N_10188);
nand U13146 (N_13146,N_10349,N_11545);
xor U13147 (N_13147,N_10988,N_11728);
nor U13148 (N_13148,N_10742,N_11759);
nor U13149 (N_13149,N_10743,N_10600);
or U13150 (N_13150,N_11426,N_11787);
nand U13151 (N_13151,N_10199,N_11118);
and U13152 (N_13152,N_10646,N_10972);
or U13153 (N_13153,N_10320,N_11682);
nand U13154 (N_13154,N_11522,N_11340);
nand U13155 (N_13155,N_11537,N_10741);
or U13156 (N_13156,N_10117,N_11061);
and U13157 (N_13157,N_10283,N_11285);
and U13158 (N_13158,N_10639,N_10185);
and U13159 (N_13159,N_11439,N_11423);
or U13160 (N_13160,N_11400,N_10825);
or U13161 (N_13161,N_11822,N_11355);
and U13162 (N_13162,N_10224,N_10834);
or U13163 (N_13163,N_10695,N_10022);
nand U13164 (N_13164,N_11701,N_10275);
or U13165 (N_13165,N_10630,N_10208);
nand U13166 (N_13166,N_11788,N_11714);
or U13167 (N_13167,N_11608,N_10419);
nor U13168 (N_13168,N_11813,N_10748);
nand U13169 (N_13169,N_10085,N_11035);
and U13170 (N_13170,N_11781,N_10099);
nand U13171 (N_13171,N_11514,N_11014);
nor U13172 (N_13172,N_11945,N_10346);
nand U13173 (N_13173,N_10578,N_10316);
or U13174 (N_13174,N_11787,N_11513);
nand U13175 (N_13175,N_10977,N_10571);
or U13176 (N_13176,N_10536,N_10317);
nand U13177 (N_13177,N_11924,N_10196);
nand U13178 (N_13178,N_10587,N_11453);
or U13179 (N_13179,N_11312,N_11115);
and U13180 (N_13180,N_10900,N_11046);
nand U13181 (N_13181,N_10433,N_10393);
nor U13182 (N_13182,N_10696,N_11359);
xor U13183 (N_13183,N_11071,N_11910);
nor U13184 (N_13184,N_11804,N_11914);
or U13185 (N_13185,N_10186,N_11742);
nand U13186 (N_13186,N_10406,N_10307);
nor U13187 (N_13187,N_10250,N_10552);
or U13188 (N_13188,N_11530,N_11779);
or U13189 (N_13189,N_10131,N_10491);
or U13190 (N_13190,N_10388,N_11888);
xnor U13191 (N_13191,N_11258,N_10403);
nand U13192 (N_13192,N_10071,N_10385);
or U13193 (N_13193,N_10350,N_10719);
nor U13194 (N_13194,N_10232,N_10999);
or U13195 (N_13195,N_10572,N_11239);
nor U13196 (N_13196,N_11254,N_10353);
and U13197 (N_13197,N_11419,N_10668);
or U13198 (N_13198,N_11973,N_11074);
or U13199 (N_13199,N_10576,N_11318);
and U13200 (N_13200,N_10689,N_10953);
xor U13201 (N_13201,N_11865,N_10618);
xnor U13202 (N_13202,N_11285,N_10285);
and U13203 (N_13203,N_11569,N_11338);
nor U13204 (N_13204,N_10858,N_10650);
nand U13205 (N_13205,N_11818,N_10530);
nand U13206 (N_13206,N_10703,N_10782);
and U13207 (N_13207,N_11544,N_10453);
or U13208 (N_13208,N_11796,N_11399);
or U13209 (N_13209,N_10015,N_10434);
nand U13210 (N_13210,N_10163,N_11286);
and U13211 (N_13211,N_10154,N_10192);
xnor U13212 (N_13212,N_10301,N_10434);
nand U13213 (N_13213,N_11460,N_11070);
nand U13214 (N_13214,N_10752,N_10602);
or U13215 (N_13215,N_11249,N_11134);
or U13216 (N_13216,N_10527,N_10036);
or U13217 (N_13217,N_10512,N_10612);
or U13218 (N_13218,N_11680,N_11087);
nor U13219 (N_13219,N_11312,N_10712);
or U13220 (N_13220,N_10417,N_11176);
nand U13221 (N_13221,N_11916,N_11471);
nor U13222 (N_13222,N_11684,N_10926);
or U13223 (N_13223,N_10348,N_11200);
and U13224 (N_13224,N_10686,N_10454);
and U13225 (N_13225,N_10076,N_11879);
nand U13226 (N_13226,N_10300,N_11177);
and U13227 (N_13227,N_11621,N_10548);
or U13228 (N_13228,N_10078,N_11667);
nand U13229 (N_13229,N_10271,N_11489);
nor U13230 (N_13230,N_10997,N_10076);
and U13231 (N_13231,N_11421,N_11781);
and U13232 (N_13232,N_11188,N_10174);
xor U13233 (N_13233,N_11743,N_10046);
or U13234 (N_13234,N_10508,N_10434);
nand U13235 (N_13235,N_10892,N_10225);
or U13236 (N_13236,N_11350,N_10589);
nand U13237 (N_13237,N_10205,N_11651);
or U13238 (N_13238,N_11354,N_10909);
and U13239 (N_13239,N_11322,N_11472);
nand U13240 (N_13240,N_10967,N_11204);
or U13241 (N_13241,N_10335,N_10000);
nand U13242 (N_13242,N_10512,N_11069);
or U13243 (N_13243,N_10023,N_10661);
or U13244 (N_13244,N_11938,N_10375);
and U13245 (N_13245,N_11198,N_11630);
or U13246 (N_13246,N_11287,N_10191);
and U13247 (N_13247,N_10271,N_11293);
nand U13248 (N_13248,N_10758,N_11261);
nand U13249 (N_13249,N_11843,N_10691);
or U13250 (N_13250,N_10859,N_11644);
or U13251 (N_13251,N_10957,N_10452);
nand U13252 (N_13252,N_11607,N_10187);
or U13253 (N_13253,N_11004,N_10906);
and U13254 (N_13254,N_10778,N_10990);
or U13255 (N_13255,N_11929,N_11467);
and U13256 (N_13256,N_10340,N_11330);
or U13257 (N_13257,N_11720,N_11314);
nor U13258 (N_13258,N_10399,N_10856);
xnor U13259 (N_13259,N_11682,N_11581);
or U13260 (N_13260,N_10466,N_10058);
and U13261 (N_13261,N_11764,N_11083);
nand U13262 (N_13262,N_11535,N_10429);
nand U13263 (N_13263,N_10425,N_11162);
nor U13264 (N_13264,N_10841,N_10445);
xnor U13265 (N_13265,N_11058,N_11860);
xor U13266 (N_13266,N_11178,N_11442);
or U13267 (N_13267,N_11335,N_10778);
nor U13268 (N_13268,N_10000,N_10566);
nor U13269 (N_13269,N_10645,N_10876);
or U13270 (N_13270,N_11698,N_10467);
nor U13271 (N_13271,N_11580,N_10997);
or U13272 (N_13272,N_11051,N_11828);
and U13273 (N_13273,N_10152,N_10082);
nand U13274 (N_13274,N_10617,N_10957);
nor U13275 (N_13275,N_11319,N_10339);
and U13276 (N_13276,N_10468,N_11781);
and U13277 (N_13277,N_11366,N_11015);
xor U13278 (N_13278,N_10123,N_11482);
and U13279 (N_13279,N_10261,N_11353);
and U13280 (N_13280,N_11436,N_10049);
or U13281 (N_13281,N_11679,N_10258);
or U13282 (N_13282,N_10894,N_10544);
or U13283 (N_13283,N_10913,N_10584);
nand U13284 (N_13284,N_11692,N_10538);
nor U13285 (N_13285,N_11309,N_10521);
and U13286 (N_13286,N_10517,N_11534);
nand U13287 (N_13287,N_11878,N_11918);
nand U13288 (N_13288,N_10290,N_11283);
and U13289 (N_13289,N_11486,N_10273);
nand U13290 (N_13290,N_11934,N_10445);
and U13291 (N_13291,N_10389,N_10526);
or U13292 (N_13292,N_10876,N_10019);
nor U13293 (N_13293,N_11825,N_11862);
nor U13294 (N_13294,N_10460,N_11039);
nor U13295 (N_13295,N_10278,N_10308);
nand U13296 (N_13296,N_10848,N_11553);
or U13297 (N_13297,N_11539,N_10696);
nand U13298 (N_13298,N_11166,N_10881);
nor U13299 (N_13299,N_11048,N_11028);
nand U13300 (N_13300,N_10135,N_10005);
and U13301 (N_13301,N_10635,N_11528);
nor U13302 (N_13302,N_10242,N_10890);
and U13303 (N_13303,N_10313,N_11371);
and U13304 (N_13304,N_10073,N_11056);
or U13305 (N_13305,N_10240,N_11202);
and U13306 (N_13306,N_10951,N_11300);
nand U13307 (N_13307,N_10069,N_10059);
nand U13308 (N_13308,N_10589,N_10865);
and U13309 (N_13309,N_11449,N_10142);
and U13310 (N_13310,N_11518,N_11460);
xnor U13311 (N_13311,N_11454,N_10530);
nor U13312 (N_13312,N_11502,N_10146);
nand U13313 (N_13313,N_10063,N_11786);
or U13314 (N_13314,N_11879,N_10483);
and U13315 (N_13315,N_11514,N_11353);
nor U13316 (N_13316,N_11294,N_10853);
nand U13317 (N_13317,N_10694,N_11154);
and U13318 (N_13318,N_10014,N_11009);
and U13319 (N_13319,N_10846,N_10271);
or U13320 (N_13320,N_11612,N_10901);
nand U13321 (N_13321,N_11171,N_11807);
and U13322 (N_13322,N_10749,N_10641);
nand U13323 (N_13323,N_11107,N_10514);
nand U13324 (N_13324,N_11438,N_10260);
or U13325 (N_13325,N_10676,N_10120);
or U13326 (N_13326,N_10370,N_10322);
and U13327 (N_13327,N_10573,N_10361);
and U13328 (N_13328,N_11698,N_11685);
and U13329 (N_13329,N_10582,N_11890);
and U13330 (N_13330,N_10544,N_10373);
xnor U13331 (N_13331,N_10923,N_10168);
and U13332 (N_13332,N_11005,N_11809);
or U13333 (N_13333,N_11030,N_11940);
nand U13334 (N_13334,N_11896,N_11146);
nand U13335 (N_13335,N_10574,N_11297);
nor U13336 (N_13336,N_10641,N_10172);
or U13337 (N_13337,N_10663,N_11343);
xor U13338 (N_13338,N_10346,N_11360);
and U13339 (N_13339,N_11190,N_11164);
and U13340 (N_13340,N_11721,N_10152);
and U13341 (N_13341,N_11136,N_11342);
nand U13342 (N_13342,N_11271,N_10630);
or U13343 (N_13343,N_11268,N_11949);
and U13344 (N_13344,N_10964,N_10794);
nor U13345 (N_13345,N_10289,N_11991);
nand U13346 (N_13346,N_11603,N_10981);
nand U13347 (N_13347,N_10927,N_10178);
or U13348 (N_13348,N_10758,N_11140);
or U13349 (N_13349,N_11733,N_11351);
nand U13350 (N_13350,N_11305,N_11148);
xnor U13351 (N_13351,N_10637,N_11511);
nand U13352 (N_13352,N_11503,N_11623);
and U13353 (N_13353,N_10346,N_10240);
or U13354 (N_13354,N_11588,N_11223);
or U13355 (N_13355,N_11754,N_10748);
and U13356 (N_13356,N_10214,N_11852);
nand U13357 (N_13357,N_10838,N_11209);
nand U13358 (N_13358,N_11058,N_10050);
or U13359 (N_13359,N_10468,N_10664);
nand U13360 (N_13360,N_11289,N_11336);
nor U13361 (N_13361,N_11606,N_10836);
xnor U13362 (N_13362,N_11213,N_10733);
or U13363 (N_13363,N_11285,N_11774);
nand U13364 (N_13364,N_11253,N_10932);
nor U13365 (N_13365,N_11436,N_10659);
and U13366 (N_13366,N_11245,N_10274);
xor U13367 (N_13367,N_10833,N_10823);
and U13368 (N_13368,N_11417,N_11381);
nand U13369 (N_13369,N_10881,N_11157);
xor U13370 (N_13370,N_11162,N_10505);
nor U13371 (N_13371,N_10589,N_11571);
nor U13372 (N_13372,N_11330,N_10223);
xnor U13373 (N_13373,N_11412,N_11180);
and U13374 (N_13374,N_11453,N_11500);
nor U13375 (N_13375,N_11359,N_10305);
nor U13376 (N_13376,N_10711,N_10212);
or U13377 (N_13377,N_10842,N_10609);
nor U13378 (N_13378,N_10614,N_11234);
xnor U13379 (N_13379,N_10529,N_11355);
or U13380 (N_13380,N_11271,N_11050);
or U13381 (N_13381,N_11201,N_10052);
xor U13382 (N_13382,N_10093,N_11787);
and U13383 (N_13383,N_10580,N_10250);
and U13384 (N_13384,N_10577,N_11455);
or U13385 (N_13385,N_11660,N_10761);
nand U13386 (N_13386,N_11143,N_11132);
nand U13387 (N_13387,N_10783,N_11552);
nor U13388 (N_13388,N_10633,N_11955);
nor U13389 (N_13389,N_10459,N_11126);
or U13390 (N_13390,N_11264,N_10026);
xor U13391 (N_13391,N_11565,N_11287);
and U13392 (N_13392,N_11039,N_10569);
or U13393 (N_13393,N_10341,N_10452);
or U13394 (N_13394,N_11587,N_10666);
nand U13395 (N_13395,N_11850,N_10574);
or U13396 (N_13396,N_11150,N_11779);
or U13397 (N_13397,N_11294,N_10142);
and U13398 (N_13398,N_10919,N_10726);
xnor U13399 (N_13399,N_10215,N_10423);
nand U13400 (N_13400,N_10603,N_11852);
or U13401 (N_13401,N_10745,N_10843);
and U13402 (N_13402,N_11648,N_11490);
nor U13403 (N_13403,N_11752,N_11182);
and U13404 (N_13404,N_10787,N_11063);
and U13405 (N_13405,N_11548,N_10593);
nor U13406 (N_13406,N_11339,N_11349);
and U13407 (N_13407,N_11674,N_10781);
and U13408 (N_13408,N_11718,N_11817);
nand U13409 (N_13409,N_11862,N_10595);
nor U13410 (N_13410,N_10532,N_11944);
and U13411 (N_13411,N_10309,N_11373);
nor U13412 (N_13412,N_10110,N_10496);
nor U13413 (N_13413,N_11038,N_11329);
nor U13414 (N_13414,N_10578,N_10025);
or U13415 (N_13415,N_10619,N_11964);
nor U13416 (N_13416,N_10867,N_10488);
nand U13417 (N_13417,N_10793,N_10233);
and U13418 (N_13418,N_10165,N_10512);
nand U13419 (N_13419,N_10600,N_10248);
nor U13420 (N_13420,N_11108,N_10049);
nor U13421 (N_13421,N_10072,N_10137);
or U13422 (N_13422,N_11530,N_11341);
nor U13423 (N_13423,N_10770,N_11328);
nor U13424 (N_13424,N_10834,N_10712);
or U13425 (N_13425,N_11113,N_11249);
nand U13426 (N_13426,N_11418,N_11689);
or U13427 (N_13427,N_10403,N_10480);
nand U13428 (N_13428,N_11377,N_10907);
nor U13429 (N_13429,N_10746,N_10856);
and U13430 (N_13430,N_11456,N_10910);
or U13431 (N_13431,N_10220,N_11694);
or U13432 (N_13432,N_11840,N_10067);
nand U13433 (N_13433,N_10263,N_10394);
and U13434 (N_13434,N_11396,N_10932);
and U13435 (N_13435,N_11644,N_11220);
nand U13436 (N_13436,N_10783,N_11321);
nand U13437 (N_13437,N_11809,N_11524);
and U13438 (N_13438,N_10404,N_11924);
and U13439 (N_13439,N_11437,N_10148);
xor U13440 (N_13440,N_10902,N_10599);
or U13441 (N_13441,N_11540,N_10492);
nor U13442 (N_13442,N_10730,N_11772);
or U13443 (N_13443,N_11202,N_11195);
nand U13444 (N_13444,N_11804,N_11311);
and U13445 (N_13445,N_10295,N_10498);
xnor U13446 (N_13446,N_11968,N_11159);
or U13447 (N_13447,N_10032,N_11319);
and U13448 (N_13448,N_10440,N_11187);
nor U13449 (N_13449,N_10046,N_11166);
nand U13450 (N_13450,N_11909,N_10447);
nand U13451 (N_13451,N_11038,N_10704);
or U13452 (N_13452,N_10218,N_10143);
nand U13453 (N_13453,N_11164,N_10439);
and U13454 (N_13454,N_11586,N_10473);
and U13455 (N_13455,N_10037,N_10832);
nor U13456 (N_13456,N_10825,N_10735);
nor U13457 (N_13457,N_11281,N_10389);
nand U13458 (N_13458,N_10352,N_11476);
nor U13459 (N_13459,N_10319,N_11139);
nand U13460 (N_13460,N_11779,N_10995);
nand U13461 (N_13461,N_10516,N_10906);
nor U13462 (N_13462,N_10549,N_11566);
nand U13463 (N_13463,N_10755,N_11260);
nor U13464 (N_13464,N_10373,N_10365);
nand U13465 (N_13465,N_10899,N_10273);
nor U13466 (N_13466,N_10343,N_11840);
and U13467 (N_13467,N_11065,N_11437);
or U13468 (N_13468,N_10048,N_11755);
and U13469 (N_13469,N_10320,N_10135);
or U13470 (N_13470,N_11929,N_11709);
or U13471 (N_13471,N_10249,N_11921);
and U13472 (N_13472,N_10635,N_10071);
xnor U13473 (N_13473,N_11583,N_11810);
or U13474 (N_13474,N_10839,N_11356);
nand U13475 (N_13475,N_10551,N_10794);
or U13476 (N_13476,N_10377,N_10895);
nor U13477 (N_13477,N_10950,N_10581);
nor U13478 (N_13478,N_10584,N_11218);
nor U13479 (N_13479,N_11955,N_11768);
xor U13480 (N_13480,N_10734,N_10197);
nand U13481 (N_13481,N_10271,N_11232);
nor U13482 (N_13482,N_11874,N_11097);
nand U13483 (N_13483,N_11361,N_10165);
or U13484 (N_13484,N_11082,N_11354);
or U13485 (N_13485,N_10758,N_11620);
nand U13486 (N_13486,N_10455,N_10921);
nand U13487 (N_13487,N_10021,N_10653);
and U13488 (N_13488,N_10290,N_11735);
xor U13489 (N_13489,N_11109,N_11407);
or U13490 (N_13490,N_10613,N_10740);
nand U13491 (N_13491,N_10245,N_11369);
nor U13492 (N_13492,N_10384,N_10752);
or U13493 (N_13493,N_10592,N_10306);
and U13494 (N_13494,N_11030,N_11247);
or U13495 (N_13495,N_11206,N_10553);
nand U13496 (N_13496,N_10407,N_10792);
nand U13497 (N_13497,N_11590,N_11890);
nor U13498 (N_13498,N_11652,N_10135);
nor U13499 (N_13499,N_10958,N_10770);
and U13500 (N_13500,N_10209,N_11695);
nand U13501 (N_13501,N_11662,N_10100);
or U13502 (N_13502,N_10839,N_10364);
or U13503 (N_13503,N_11407,N_10022);
nor U13504 (N_13504,N_10428,N_11444);
or U13505 (N_13505,N_11212,N_11917);
and U13506 (N_13506,N_11436,N_10600);
nor U13507 (N_13507,N_10898,N_10261);
and U13508 (N_13508,N_11084,N_10085);
xor U13509 (N_13509,N_10063,N_10226);
nand U13510 (N_13510,N_11861,N_10073);
nor U13511 (N_13511,N_11222,N_11046);
or U13512 (N_13512,N_11514,N_10310);
nand U13513 (N_13513,N_11880,N_10572);
xor U13514 (N_13514,N_10668,N_11543);
nor U13515 (N_13515,N_10814,N_10503);
nor U13516 (N_13516,N_11914,N_10801);
and U13517 (N_13517,N_10656,N_11974);
and U13518 (N_13518,N_10063,N_11354);
nor U13519 (N_13519,N_10766,N_10715);
nand U13520 (N_13520,N_10276,N_11985);
or U13521 (N_13521,N_10887,N_11284);
or U13522 (N_13522,N_10466,N_10012);
xnor U13523 (N_13523,N_11403,N_10353);
xnor U13524 (N_13524,N_10028,N_10199);
or U13525 (N_13525,N_10618,N_10556);
nor U13526 (N_13526,N_11527,N_11768);
nor U13527 (N_13527,N_10567,N_11034);
nand U13528 (N_13528,N_10534,N_11629);
nand U13529 (N_13529,N_11627,N_11875);
or U13530 (N_13530,N_10817,N_11231);
and U13531 (N_13531,N_10026,N_10831);
nor U13532 (N_13532,N_10326,N_11050);
nor U13533 (N_13533,N_11425,N_10851);
nand U13534 (N_13534,N_11157,N_11715);
nand U13535 (N_13535,N_10470,N_10778);
or U13536 (N_13536,N_11922,N_11369);
xnor U13537 (N_13537,N_10274,N_11719);
and U13538 (N_13538,N_10478,N_10621);
nor U13539 (N_13539,N_11716,N_10421);
or U13540 (N_13540,N_11161,N_10158);
nor U13541 (N_13541,N_10525,N_10781);
or U13542 (N_13542,N_11312,N_10888);
nand U13543 (N_13543,N_10006,N_10713);
nand U13544 (N_13544,N_10129,N_11783);
xor U13545 (N_13545,N_10528,N_11248);
xor U13546 (N_13546,N_10584,N_11425);
and U13547 (N_13547,N_11561,N_11604);
and U13548 (N_13548,N_10199,N_10336);
nor U13549 (N_13549,N_11442,N_10772);
nand U13550 (N_13550,N_10258,N_11621);
and U13551 (N_13551,N_11275,N_10092);
and U13552 (N_13552,N_10018,N_10690);
xnor U13553 (N_13553,N_10400,N_11428);
and U13554 (N_13554,N_11444,N_11225);
nand U13555 (N_13555,N_10592,N_10403);
and U13556 (N_13556,N_10681,N_10178);
or U13557 (N_13557,N_10337,N_11640);
nand U13558 (N_13558,N_11656,N_11141);
nand U13559 (N_13559,N_11818,N_11336);
nand U13560 (N_13560,N_10642,N_10836);
nand U13561 (N_13561,N_11633,N_11154);
nor U13562 (N_13562,N_10306,N_10787);
or U13563 (N_13563,N_11626,N_11924);
and U13564 (N_13564,N_10423,N_10536);
or U13565 (N_13565,N_10190,N_10474);
and U13566 (N_13566,N_10731,N_11065);
nor U13567 (N_13567,N_11265,N_10980);
or U13568 (N_13568,N_10455,N_10492);
or U13569 (N_13569,N_10757,N_11661);
nor U13570 (N_13570,N_10906,N_10663);
nand U13571 (N_13571,N_10498,N_10602);
nor U13572 (N_13572,N_11136,N_11544);
or U13573 (N_13573,N_11444,N_10109);
nor U13574 (N_13574,N_11145,N_10547);
and U13575 (N_13575,N_10488,N_10161);
nor U13576 (N_13576,N_10747,N_10276);
nand U13577 (N_13577,N_11523,N_10782);
nand U13578 (N_13578,N_10970,N_10173);
nor U13579 (N_13579,N_11158,N_11133);
nand U13580 (N_13580,N_11265,N_10814);
and U13581 (N_13581,N_10908,N_10770);
nand U13582 (N_13582,N_11295,N_10414);
or U13583 (N_13583,N_11460,N_10624);
nand U13584 (N_13584,N_11369,N_11718);
nor U13585 (N_13585,N_11459,N_11941);
or U13586 (N_13586,N_11250,N_10579);
nor U13587 (N_13587,N_10030,N_10724);
nor U13588 (N_13588,N_10690,N_11597);
and U13589 (N_13589,N_11641,N_11601);
nand U13590 (N_13590,N_10790,N_10377);
nand U13591 (N_13591,N_10366,N_11789);
or U13592 (N_13592,N_10128,N_11954);
or U13593 (N_13593,N_10393,N_10613);
or U13594 (N_13594,N_10605,N_11659);
nand U13595 (N_13595,N_10373,N_10378);
nor U13596 (N_13596,N_10769,N_10723);
nand U13597 (N_13597,N_11528,N_11512);
nand U13598 (N_13598,N_10302,N_10905);
or U13599 (N_13599,N_11732,N_10605);
xnor U13600 (N_13600,N_11611,N_10074);
and U13601 (N_13601,N_10956,N_11722);
nand U13602 (N_13602,N_10615,N_11258);
or U13603 (N_13603,N_10804,N_11830);
and U13604 (N_13604,N_10044,N_10765);
and U13605 (N_13605,N_10017,N_11633);
and U13606 (N_13606,N_10173,N_10395);
xnor U13607 (N_13607,N_11033,N_10567);
and U13608 (N_13608,N_11464,N_11807);
xnor U13609 (N_13609,N_11406,N_10756);
nor U13610 (N_13610,N_11942,N_10448);
nand U13611 (N_13611,N_11603,N_11730);
nor U13612 (N_13612,N_10488,N_11400);
or U13613 (N_13613,N_11087,N_11060);
and U13614 (N_13614,N_10539,N_10014);
xnor U13615 (N_13615,N_10748,N_11070);
and U13616 (N_13616,N_10695,N_11470);
or U13617 (N_13617,N_11768,N_10260);
nand U13618 (N_13618,N_10225,N_11581);
xnor U13619 (N_13619,N_10956,N_11281);
or U13620 (N_13620,N_11199,N_11491);
nor U13621 (N_13621,N_11072,N_10512);
or U13622 (N_13622,N_10452,N_11814);
nor U13623 (N_13623,N_11685,N_11890);
and U13624 (N_13624,N_10143,N_11764);
xnor U13625 (N_13625,N_11289,N_11047);
nand U13626 (N_13626,N_10060,N_10810);
nor U13627 (N_13627,N_11987,N_10321);
nor U13628 (N_13628,N_11610,N_10851);
and U13629 (N_13629,N_10394,N_10571);
nand U13630 (N_13630,N_10526,N_10625);
nor U13631 (N_13631,N_11657,N_10726);
nor U13632 (N_13632,N_11415,N_10585);
and U13633 (N_13633,N_11920,N_11118);
and U13634 (N_13634,N_11138,N_11067);
xnor U13635 (N_13635,N_10831,N_11077);
nor U13636 (N_13636,N_11393,N_11463);
and U13637 (N_13637,N_10057,N_10920);
xnor U13638 (N_13638,N_11726,N_10357);
and U13639 (N_13639,N_11329,N_11198);
nor U13640 (N_13640,N_10427,N_11300);
or U13641 (N_13641,N_11540,N_11344);
or U13642 (N_13642,N_11427,N_10484);
or U13643 (N_13643,N_11682,N_10885);
nor U13644 (N_13644,N_11049,N_10355);
nor U13645 (N_13645,N_11076,N_11892);
or U13646 (N_13646,N_11108,N_10354);
or U13647 (N_13647,N_10881,N_10906);
and U13648 (N_13648,N_11960,N_10385);
nor U13649 (N_13649,N_10503,N_10185);
or U13650 (N_13650,N_11433,N_10125);
and U13651 (N_13651,N_10991,N_10106);
and U13652 (N_13652,N_11774,N_11003);
xnor U13653 (N_13653,N_11441,N_11050);
or U13654 (N_13654,N_10948,N_11897);
or U13655 (N_13655,N_11380,N_10557);
nand U13656 (N_13656,N_10780,N_11993);
nand U13657 (N_13657,N_10655,N_11191);
nor U13658 (N_13658,N_10561,N_11979);
or U13659 (N_13659,N_10545,N_10727);
nor U13660 (N_13660,N_10188,N_10484);
or U13661 (N_13661,N_10986,N_10127);
xnor U13662 (N_13662,N_11593,N_10208);
nand U13663 (N_13663,N_11100,N_10864);
and U13664 (N_13664,N_10494,N_11026);
or U13665 (N_13665,N_11068,N_11963);
nor U13666 (N_13666,N_10157,N_11698);
nor U13667 (N_13667,N_10354,N_11633);
and U13668 (N_13668,N_10229,N_10966);
nor U13669 (N_13669,N_11994,N_11061);
and U13670 (N_13670,N_11311,N_11416);
nor U13671 (N_13671,N_11374,N_10912);
xnor U13672 (N_13672,N_10849,N_10229);
nand U13673 (N_13673,N_10496,N_10156);
xnor U13674 (N_13674,N_11575,N_11684);
or U13675 (N_13675,N_11837,N_11279);
or U13676 (N_13676,N_11969,N_10262);
or U13677 (N_13677,N_10801,N_11819);
and U13678 (N_13678,N_10270,N_11959);
xnor U13679 (N_13679,N_11299,N_10043);
and U13680 (N_13680,N_11889,N_11136);
nor U13681 (N_13681,N_10088,N_10080);
nor U13682 (N_13682,N_10085,N_10202);
nor U13683 (N_13683,N_10097,N_10353);
or U13684 (N_13684,N_11614,N_10550);
or U13685 (N_13685,N_10426,N_10098);
nand U13686 (N_13686,N_10764,N_10343);
or U13687 (N_13687,N_10295,N_11993);
xnor U13688 (N_13688,N_11099,N_10010);
and U13689 (N_13689,N_11265,N_10808);
and U13690 (N_13690,N_11432,N_11177);
or U13691 (N_13691,N_10570,N_10528);
or U13692 (N_13692,N_10984,N_11294);
xnor U13693 (N_13693,N_11393,N_10823);
nand U13694 (N_13694,N_11065,N_11547);
nand U13695 (N_13695,N_11646,N_10217);
nand U13696 (N_13696,N_10930,N_10912);
nand U13697 (N_13697,N_11484,N_10406);
nor U13698 (N_13698,N_10859,N_11898);
nand U13699 (N_13699,N_10340,N_10520);
nor U13700 (N_13700,N_10249,N_10014);
nor U13701 (N_13701,N_10628,N_11902);
nor U13702 (N_13702,N_11797,N_11860);
or U13703 (N_13703,N_10974,N_10022);
or U13704 (N_13704,N_11517,N_10997);
or U13705 (N_13705,N_10028,N_10229);
and U13706 (N_13706,N_10354,N_11833);
or U13707 (N_13707,N_11197,N_11471);
and U13708 (N_13708,N_11486,N_10732);
and U13709 (N_13709,N_10100,N_11316);
nand U13710 (N_13710,N_11042,N_11272);
nor U13711 (N_13711,N_11638,N_11312);
xnor U13712 (N_13712,N_10388,N_10939);
and U13713 (N_13713,N_11241,N_10275);
nor U13714 (N_13714,N_11504,N_11140);
or U13715 (N_13715,N_11582,N_11712);
nand U13716 (N_13716,N_11512,N_10371);
nand U13717 (N_13717,N_10514,N_11608);
nor U13718 (N_13718,N_11302,N_11759);
nor U13719 (N_13719,N_11122,N_10878);
xor U13720 (N_13720,N_10786,N_11747);
or U13721 (N_13721,N_11214,N_10539);
xnor U13722 (N_13722,N_11448,N_10771);
xnor U13723 (N_13723,N_10703,N_11003);
nand U13724 (N_13724,N_10311,N_10695);
nand U13725 (N_13725,N_10727,N_10131);
xor U13726 (N_13726,N_11504,N_11830);
nand U13727 (N_13727,N_10011,N_11321);
or U13728 (N_13728,N_10407,N_11275);
or U13729 (N_13729,N_10955,N_11753);
and U13730 (N_13730,N_10150,N_10033);
nand U13731 (N_13731,N_10190,N_10146);
nand U13732 (N_13732,N_10547,N_10061);
and U13733 (N_13733,N_11358,N_10820);
nand U13734 (N_13734,N_11865,N_10125);
xor U13735 (N_13735,N_11486,N_10248);
nor U13736 (N_13736,N_10171,N_11476);
and U13737 (N_13737,N_11636,N_11579);
nand U13738 (N_13738,N_10284,N_10091);
or U13739 (N_13739,N_10385,N_10909);
and U13740 (N_13740,N_10441,N_10457);
nand U13741 (N_13741,N_10985,N_10287);
nor U13742 (N_13742,N_10818,N_11188);
xor U13743 (N_13743,N_11460,N_11047);
nand U13744 (N_13744,N_11305,N_11042);
nand U13745 (N_13745,N_11485,N_11586);
nor U13746 (N_13746,N_11732,N_11617);
or U13747 (N_13747,N_11135,N_11308);
and U13748 (N_13748,N_10090,N_11758);
nand U13749 (N_13749,N_10218,N_11358);
and U13750 (N_13750,N_11329,N_11056);
nand U13751 (N_13751,N_11144,N_10270);
nor U13752 (N_13752,N_10095,N_10586);
nor U13753 (N_13753,N_11972,N_11941);
and U13754 (N_13754,N_10943,N_11767);
nand U13755 (N_13755,N_10931,N_10199);
nor U13756 (N_13756,N_10162,N_11152);
nand U13757 (N_13757,N_10481,N_11918);
or U13758 (N_13758,N_10841,N_10640);
nor U13759 (N_13759,N_11302,N_11972);
and U13760 (N_13760,N_11311,N_11716);
nand U13761 (N_13761,N_10065,N_11159);
and U13762 (N_13762,N_10081,N_11020);
nand U13763 (N_13763,N_11081,N_11816);
nand U13764 (N_13764,N_11145,N_11933);
nand U13765 (N_13765,N_10097,N_10066);
nand U13766 (N_13766,N_11373,N_10616);
nand U13767 (N_13767,N_11681,N_10225);
nand U13768 (N_13768,N_10465,N_10100);
and U13769 (N_13769,N_11781,N_10843);
nor U13770 (N_13770,N_11463,N_11557);
or U13771 (N_13771,N_10064,N_10949);
and U13772 (N_13772,N_11899,N_11865);
xor U13773 (N_13773,N_11345,N_10652);
or U13774 (N_13774,N_11166,N_10056);
nand U13775 (N_13775,N_11543,N_10622);
or U13776 (N_13776,N_11535,N_10616);
and U13777 (N_13777,N_11379,N_10305);
xor U13778 (N_13778,N_10446,N_11315);
or U13779 (N_13779,N_10956,N_11100);
and U13780 (N_13780,N_10342,N_10554);
xor U13781 (N_13781,N_11335,N_10814);
and U13782 (N_13782,N_11294,N_11411);
nand U13783 (N_13783,N_11878,N_10802);
nor U13784 (N_13784,N_10173,N_11300);
or U13785 (N_13785,N_11873,N_10853);
or U13786 (N_13786,N_11554,N_11614);
and U13787 (N_13787,N_10595,N_10222);
and U13788 (N_13788,N_10462,N_11561);
nand U13789 (N_13789,N_10168,N_10714);
and U13790 (N_13790,N_11698,N_10478);
or U13791 (N_13791,N_10739,N_11001);
nor U13792 (N_13792,N_10558,N_10956);
xor U13793 (N_13793,N_11890,N_11995);
xnor U13794 (N_13794,N_10506,N_10298);
and U13795 (N_13795,N_10186,N_11964);
and U13796 (N_13796,N_11281,N_10200);
or U13797 (N_13797,N_11161,N_10428);
or U13798 (N_13798,N_11017,N_11281);
or U13799 (N_13799,N_11337,N_11000);
and U13800 (N_13800,N_10831,N_10748);
and U13801 (N_13801,N_10090,N_11680);
and U13802 (N_13802,N_10054,N_10878);
or U13803 (N_13803,N_10689,N_10118);
or U13804 (N_13804,N_10742,N_10461);
and U13805 (N_13805,N_10280,N_10510);
or U13806 (N_13806,N_11586,N_11237);
or U13807 (N_13807,N_11799,N_11379);
nor U13808 (N_13808,N_10180,N_11027);
nor U13809 (N_13809,N_11072,N_11160);
nand U13810 (N_13810,N_10987,N_11393);
nor U13811 (N_13811,N_11991,N_11697);
nand U13812 (N_13812,N_10412,N_11616);
nor U13813 (N_13813,N_10653,N_10950);
or U13814 (N_13814,N_11833,N_10755);
or U13815 (N_13815,N_11536,N_10589);
or U13816 (N_13816,N_11825,N_11487);
or U13817 (N_13817,N_10886,N_11246);
xor U13818 (N_13818,N_11518,N_11378);
nand U13819 (N_13819,N_11638,N_11789);
nor U13820 (N_13820,N_10494,N_11192);
or U13821 (N_13821,N_11941,N_10543);
nor U13822 (N_13822,N_11905,N_10750);
nor U13823 (N_13823,N_11115,N_10857);
nand U13824 (N_13824,N_11712,N_10944);
nor U13825 (N_13825,N_11073,N_11974);
xnor U13826 (N_13826,N_11714,N_10625);
nand U13827 (N_13827,N_10067,N_10518);
or U13828 (N_13828,N_11286,N_11502);
nor U13829 (N_13829,N_11779,N_10302);
nor U13830 (N_13830,N_11451,N_10742);
and U13831 (N_13831,N_10575,N_10833);
or U13832 (N_13832,N_10820,N_10811);
and U13833 (N_13833,N_10835,N_11447);
and U13834 (N_13834,N_11022,N_11724);
nand U13835 (N_13835,N_10897,N_11492);
nand U13836 (N_13836,N_10512,N_11008);
nand U13837 (N_13837,N_10690,N_10785);
xor U13838 (N_13838,N_11907,N_10088);
nor U13839 (N_13839,N_11188,N_10475);
or U13840 (N_13840,N_10691,N_11923);
and U13841 (N_13841,N_11062,N_11515);
nand U13842 (N_13842,N_11534,N_10356);
nor U13843 (N_13843,N_11017,N_11918);
and U13844 (N_13844,N_11048,N_11334);
nor U13845 (N_13845,N_10851,N_10080);
nand U13846 (N_13846,N_10354,N_11012);
nand U13847 (N_13847,N_10344,N_10259);
nor U13848 (N_13848,N_11470,N_10840);
or U13849 (N_13849,N_11086,N_11279);
nor U13850 (N_13850,N_11684,N_11421);
or U13851 (N_13851,N_10875,N_11671);
nor U13852 (N_13852,N_10974,N_10498);
and U13853 (N_13853,N_10840,N_11361);
and U13854 (N_13854,N_10633,N_10366);
nand U13855 (N_13855,N_10952,N_10966);
xnor U13856 (N_13856,N_10128,N_10776);
or U13857 (N_13857,N_11617,N_11574);
and U13858 (N_13858,N_10438,N_10584);
and U13859 (N_13859,N_11679,N_10746);
or U13860 (N_13860,N_11810,N_10088);
nor U13861 (N_13861,N_10040,N_10303);
and U13862 (N_13862,N_11435,N_10763);
or U13863 (N_13863,N_10004,N_10864);
nor U13864 (N_13864,N_10958,N_11005);
and U13865 (N_13865,N_11280,N_11312);
nor U13866 (N_13866,N_10954,N_11533);
xor U13867 (N_13867,N_11405,N_11086);
and U13868 (N_13868,N_11091,N_11224);
xnor U13869 (N_13869,N_11564,N_11823);
nor U13870 (N_13870,N_11224,N_10410);
and U13871 (N_13871,N_10470,N_11052);
or U13872 (N_13872,N_10471,N_10729);
nor U13873 (N_13873,N_11236,N_10175);
or U13874 (N_13874,N_11848,N_11785);
xor U13875 (N_13875,N_11404,N_10198);
nand U13876 (N_13876,N_10101,N_11405);
xor U13877 (N_13877,N_10891,N_10439);
or U13878 (N_13878,N_11026,N_10084);
xor U13879 (N_13879,N_10888,N_11484);
nand U13880 (N_13880,N_10894,N_11127);
xor U13881 (N_13881,N_10844,N_10280);
or U13882 (N_13882,N_10264,N_11480);
and U13883 (N_13883,N_10231,N_10954);
or U13884 (N_13884,N_10740,N_10811);
nor U13885 (N_13885,N_11137,N_11580);
nand U13886 (N_13886,N_11994,N_10173);
nand U13887 (N_13887,N_11201,N_11377);
nor U13888 (N_13888,N_11156,N_11603);
and U13889 (N_13889,N_11345,N_11475);
and U13890 (N_13890,N_10962,N_10395);
nor U13891 (N_13891,N_11933,N_10928);
nor U13892 (N_13892,N_11128,N_11996);
or U13893 (N_13893,N_11699,N_11799);
nand U13894 (N_13894,N_10584,N_10086);
and U13895 (N_13895,N_10243,N_11622);
and U13896 (N_13896,N_11299,N_11689);
nor U13897 (N_13897,N_10657,N_10111);
nand U13898 (N_13898,N_10494,N_11191);
and U13899 (N_13899,N_10119,N_10320);
and U13900 (N_13900,N_10447,N_10913);
and U13901 (N_13901,N_11082,N_10500);
or U13902 (N_13902,N_10293,N_10010);
or U13903 (N_13903,N_11872,N_10542);
xnor U13904 (N_13904,N_11269,N_10237);
nor U13905 (N_13905,N_11061,N_10958);
nor U13906 (N_13906,N_11607,N_11684);
nand U13907 (N_13907,N_11241,N_11126);
or U13908 (N_13908,N_11710,N_11739);
and U13909 (N_13909,N_10573,N_11602);
and U13910 (N_13910,N_10270,N_11388);
nand U13911 (N_13911,N_10934,N_11258);
nand U13912 (N_13912,N_11547,N_10501);
and U13913 (N_13913,N_11203,N_11365);
or U13914 (N_13914,N_11946,N_10637);
or U13915 (N_13915,N_11800,N_10370);
and U13916 (N_13916,N_11983,N_11024);
nor U13917 (N_13917,N_11067,N_11224);
and U13918 (N_13918,N_11109,N_10526);
or U13919 (N_13919,N_10187,N_10345);
nand U13920 (N_13920,N_11462,N_10267);
or U13921 (N_13921,N_10277,N_11750);
nor U13922 (N_13922,N_11494,N_10174);
xnor U13923 (N_13923,N_10392,N_10457);
nand U13924 (N_13924,N_11168,N_11700);
nor U13925 (N_13925,N_10088,N_11888);
or U13926 (N_13926,N_11491,N_10939);
or U13927 (N_13927,N_11137,N_10871);
and U13928 (N_13928,N_10868,N_10891);
nor U13929 (N_13929,N_10186,N_11416);
nand U13930 (N_13930,N_11462,N_11922);
nor U13931 (N_13931,N_11435,N_11772);
or U13932 (N_13932,N_10286,N_10339);
and U13933 (N_13933,N_11237,N_11173);
nand U13934 (N_13934,N_11274,N_11903);
and U13935 (N_13935,N_10382,N_10105);
or U13936 (N_13936,N_11403,N_11625);
or U13937 (N_13937,N_11037,N_11769);
nand U13938 (N_13938,N_10328,N_11199);
nand U13939 (N_13939,N_10784,N_10394);
and U13940 (N_13940,N_11642,N_10563);
nor U13941 (N_13941,N_10611,N_11361);
nand U13942 (N_13942,N_11431,N_11928);
and U13943 (N_13943,N_10268,N_11220);
and U13944 (N_13944,N_10146,N_10807);
and U13945 (N_13945,N_10973,N_10310);
nor U13946 (N_13946,N_11951,N_10601);
nor U13947 (N_13947,N_10375,N_10193);
nor U13948 (N_13948,N_11651,N_11112);
nand U13949 (N_13949,N_11195,N_11054);
or U13950 (N_13950,N_11563,N_10071);
or U13951 (N_13951,N_11118,N_10770);
nor U13952 (N_13952,N_10087,N_10993);
or U13953 (N_13953,N_10130,N_10334);
and U13954 (N_13954,N_10530,N_11418);
nor U13955 (N_13955,N_10435,N_11153);
xor U13956 (N_13956,N_11218,N_10406);
nor U13957 (N_13957,N_10709,N_11995);
and U13958 (N_13958,N_10841,N_10013);
nand U13959 (N_13959,N_10396,N_10353);
nor U13960 (N_13960,N_10247,N_11142);
nand U13961 (N_13961,N_11622,N_11225);
xnor U13962 (N_13962,N_10634,N_10722);
and U13963 (N_13963,N_11935,N_10611);
or U13964 (N_13964,N_11287,N_11350);
nor U13965 (N_13965,N_11784,N_10696);
and U13966 (N_13966,N_11448,N_10582);
xor U13967 (N_13967,N_10934,N_11643);
and U13968 (N_13968,N_10195,N_11552);
or U13969 (N_13969,N_10316,N_10296);
and U13970 (N_13970,N_11774,N_11563);
nor U13971 (N_13971,N_10819,N_10710);
or U13972 (N_13972,N_10865,N_10164);
xnor U13973 (N_13973,N_11118,N_10010);
nand U13974 (N_13974,N_10199,N_11483);
or U13975 (N_13975,N_10850,N_10043);
or U13976 (N_13976,N_10269,N_11096);
and U13977 (N_13977,N_10556,N_11384);
nand U13978 (N_13978,N_11242,N_10442);
or U13979 (N_13979,N_10474,N_10533);
and U13980 (N_13980,N_11688,N_10700);
nand U13981 (N_13981,N_10989,N_11932);
nor U13982 (N_13982,N_10519,N_11276);
or U13983 (N_13983,N_11176,N_10501);
nand U13984 (N_13984,N_10182,N_11600);
and U13985 (N_13985,N_10657,N_11693);
or U13986 (N_13986,N_11049,N_10381);
nor U13987 (N_13987,N_11764,N_10925);
and U13988 (N_13988,N_10773,N_10409);
nor U13989 (N_13989,N_10559,N_11721);
nor U13990 (N_13990,N_10688,N_11811);
nor U13991 (N_13991,N_11816,N_10381);
and U13992 (N_13992,N_10983,N_11777);
and U13993 (N_13993,N_10597,N_11742);
nand U13994 (N_13994,N_11996,N_10903);
nand U13995 (N_13995,N_10899,N_10121);
nand U13996 (N_13996,N_10704,N_10248);
or U13997 (N_13997,N_11200,N_11882);
or U13998 (N_13998,N_10582,N_11930);
nor U13999 (N_13999,N_10626,N_11094);
and U14000 (N_14000,N_13818,N_12016);
nand U14001 (N_14001,N_12646,N_12076);
and U14002 (N_14002,N_12958,N_12576);
and U14003 (N_14003,N_13232,N_13666);
nor U14004 (N_14004,N_12173,N_13813);
nand U14005 (N_14005,N_13983,N_13571);
xor U14006 (N_14006,N_13941,N_13411);
or U14007 (N_14007,N_12867,N_13884);
and U14008 (N_14008,N_13976,N_13268);
and U14009 (N_14009,N_12056,N_13673);
xnor U14010 (N_14010,N_12081,N_13606);
and U14011 (N_14011,N_12654,N_13706);
nor U14012 (N_14012,N_13497,N_13070);
and U14013 (N_14013,N_12024,N_13780);
or U14014 (N_14014,N_12542,N_13504);
nor U14015 (N_14015,N_12157,N_13208);
and U14016 (N_14016,N_12652,N_13811);
xor U14017 (N_14017,N_13942,N_12405);
and U14018 (N_14018,N_13972,N_13175);
and U14019 (N_14019,N_12154,N_13836);
nand U14020 (N_14020,N_13763,N_13808);
nor U14021 (N_14021,N_13547,N_13069);
xnor U14022 (N_14022,N_13735,N_13262);
xnor U14023 (N_14023,N_12120,N_12351);
and U14024 (N_14024,N_13801,N_13546);
and U14025 (N_14025,N_12860,N_12788);
xor U14026 (N_14026,N_12094,N_13099);
nor U14027 (N_14027,N_12194,N_13889);
or U14028 (N_14028,N_13775,N_13021);
nand U14029 (N_14029,N_13985,N_12767);
nand U14030 (N_14030,N_13251,N_13198);
nor U14031 (N_14031,N_12544,N_13226);
nor U14032 (N_14032,N_12805,N_13404);
and U14033 (N_14033,N_12978,N_13211);
nor U14034 (N_14034,N_12192,N_13587);
and U14035 (N_14035,N_13594,N_12772);
nor U14036 (N_14036,N_13974,N_13943);
nand U14037 (N_14037,N_13352,N_13905);
or U14038 (N_14038,N_13957,N_13533);
and U14039 (N_14039,N_13375,N_12782);
nor U14040 (N_14040,N_13691,N_12730);
or U14041 (N_14041,N_13241,N_13168);
or U14042 (N_14042,N_12326,N_13598);
nand U14043 (N_14043,N_13576,N_12315);
nor U14044 (N_14044,N_13769,N_12493);
and U14045 (N_14045,N_12831,N_12815);
nor U14046 (N_14046,N_12577,N_12611);
nor U14047 (N_14047,N_12383,N_13559);
nand U14048 (N_14048,N_12262,N_13630);
or U14049 (N_14049,N_12986,N_12321);
or U14050 (N_14050,N_13124,N_13341);
nand U14051 (N_14051,N_13939,N_12913);
nand U14052 (N_14052,N_13442,N_13906);
nor U14053 (N_14053,N_13311,N_13878);
or U14054 (N_14054,N_13409,N_13724);
and U14055 (N_14055,N_13540,N_12446);
nand U14056 (N_14056,N_12539,N_12711);
nand U14057 (N_14057,N_12002,N_12172);
nor U14058 (N_14058,N_13414,N_12503);
and U14059 (N_14059,N_13891,N_13144);
nand U14060 (N_14060,N_12047,N_12840);
and U14061 (N_14061,N_12655,N_13862);
or U14062 (N_14062,N_12416,N_13339);
nor U14063 (N_14063,N_13350,N_12995);
nand U14064 (N_14064,N_12130,N_13291);
nor U14065 (N_14065,N_13066,N_12828);
nand U14066 (N_14066,N_13892,N_12530);
and U14067 (N_14067,N_13730,N_13383);
nand U14068 (N_14068,N_12472,N_12944);
nand U14069 (N_14069,N_12448,N_13233);
and U14070 (N_14070,N_12255,N_12293);
nand U14071 (N_14071,N_12987,N_12393);
nand U14072 (N_14072,N_12042,N_13385);
xnor U14073 (N_14073,N_13090,N_12115);
xor U14074 (N_14074,N_13574,N_13776);
and U14075 (N_14075,N_13652,N_13096);
and U14076 (N_14076,N_12318,N_13745);
xnor U14077 (N_14077,N_12842,N_13035);
nand U14078 (N_14078,N_12689,N_12701);
or U14079 (N_14079,N_13732,N_13543);
or U14080 (N_14080,N_13524,N_12093);
nand U14081 (N_14081,N_13025,N_12070);
nor U14082 (N_14082,N_13555,N_13402);
nor U14083 (N_14083,N_12594,N_13223);
nand U14084 (N_14084,N_13231,N_13687);
nor U14085 (N_14085,N_13662,N_12686);
and U14086 (N_14086,N_13683,N_12792);
or U14087 (N_14087,N_12350,N_12159);
or U14088 (N_14088,N_13931,N_13933);
or U14089 (N_14089,N_13966,N_12078);
nor U14090 (N_14090,N_13212,N_12495);
or U14091 (N_14091,N_12642,N_13969);
nor U14092 (N_14092,N_12160,N_12325);
nor U14093 (N_14093,N_13838,N_12011);
xnor U14094 (N_14094,N_13167,N_12625);
xnor U14095 (N_14095,N_12851,N_12905);
and U14096 (N_14096,N_12934,N_13716);
or U14097 (N_14097,N_13823,N_13756);
nor U14098 (N_14098,N_12531,N_12339);
nand U14099 (N_14099,N_13016,N_13253);
nand U14100 (N_14100,N_12897,N_13807);
nor U14101 (N_14101,N_12122,N_13050);
nand U14102 (N_14102,N_13705,N_12813);
and U14103 (N_14103,N_13292,N_12209);
nor U14104 (N_14104,N_12796,N_12486);
nor U14105 (N_14105,N_12358,N_12514);
xor U14106 (N_14106,N_12196,N_13249);
nand U14107 (N_14107,N_13114,N_12227);
or U14108 (N_14108,N_12640,N_13484);
and U14109 (N_14109,N_13234,N_13703);
and U14110 (N_14110,N_12754,N_13370);
or U14111 (N_14111,N_13216,N_13992);
nand U14112 (N_14112,N_12785,N_12459);
xnor U14113 (N_14113,N_13179,N_13213);
or U14114 (N_14114,N_13004,N_13270);
and U14115 (N_14115,N_12907,N_12957);
and U14116 (N_14116,N_12604,N_12764);
or U14117 (N_14117,N_13174,N_13772);
and U14118 (N_14118,N_13516,N_13834);
xor U14119 (N_14119,N_13796,N_13815);
xnor U14120 (N_14120,N_13954,N_12869);
nand U14121 (N_14121,N_13827,N_13786);
nand U14122 (N_14122,N_13554,N_12881);
nand U14123 (N_14123,N_13399,N_13420);
or U14124 (N_14124,N_13464,N_12932);
nand U14125 (N_14125,N_12487,N_13087);
and U14126 (N_14126,N_13798,N_13681);
or U14127 (N_14127,N_13723,N_12908);
and U14128 (N_14128,N_12770,N_13742);
and U14129 (N_14129,N_12397,N_12543);
nand U14130 (N_14130,N_12829,N_13449);
and U14131 (N_14131,N_12456,N_13721);
and U14132 (N_14132,N_13828,N_12494);
nand U14133 (N_14133,N_13577,N_12036);
and U14134 (N_14134,N_12273,N_12302);
xor U14135 (N_14135,N_13659,N_13619);
xor U14136 (N_14136,N_13201,N_12210);
or U14137 (N_14137,N_12352,N_12034);
or U14138 (N_14138,N_12187,N_12454);
nor U14139 (N_14139,N_12880,N_12850);
and U14140 (N_14140,N_12832,N_12801);
nand U14141 (N_14141,N_12497,N_12281);
or U14142 (N_14142,N_13169,N_12375);
and U14143 (N_14143,N_12362,N_12233);
nor U14144 (N_14144,N_13100,N_12463);
nand U14145 (N_14145,N_12031,N_13867);
xor U14146 (N_14146,N_12774,N_12526);
or U14147 (N_14147,N_13572,N_13145);
xnor U14148 (N_14148,N_12877,N_13837);
nand U14149 (N_14149,N_13416,N_13845);
and U14150 (N_14150,N_13355,N_12866);
and U14151 (N_14151,N_12716,N_13015);
nand U14152 (N_14152,N_13346,N_13890);
nor U14153 (N_14153,N_13782,N_13645);
nor U14154 (N_14154,N_12875,N_13315);
or U14155 (N_14155,N_12690,N_12521);
or U14156 (N_14156,N_13215,N_12311);
xnor U14157 (N_14157,N_12170,N_13075);
and U14158 (N_14158,N_13508,N_12569);
or U14159 (N_14159,N_13443,N_12385);
xnor U14160 (N_14160,N_12954,N_12677);
nor U14161 (N_14161,N_12142,N_13709);
nor U14162 (N_14162,N_12341,N_13266);
or U14163 (N_14163,N_13754,N_13479);
or U14164 (N_14164,N_12606,N_13258);
nand U14165 (N_14165,N_13427,N_12335);
or U14166 (N_14166,N_12516,N_13582);
and U14167 (N_14167,N_13435,N_13230);
nand U14168 (N_14168,N_12660,N_12040);
nor U14169 (N_14169,N_13365,N_13136);
or U14170 (N_14170,N_13738,N_13515);
nand U14171 (N_14171,N_13600,N_12798);
nor U14172 (N_14172,N_12663,N_12125);
nor U14173 (N_14173,N_12438,N_13461);
xnor U14174 (N_14174,N_13332,N_13601);
xnor U14175 (N_14175,N_12280,N_12347);
nor U14176 (N_14176,N_12753,N_12166);
nand U14177 (N_14177,N_13084,N_13789);
nand U14178 (N_14178,N_12901,N_13679);
nand U14179 (N_14179,N_13254,N_12799);
or U14180 (N_14180,N_13044,N_12938);
nand U14181 (N_14181,N_13558,N_12052);
or U14182 (N_14182,N_12023,N_13613);
nor U14183 (N_14183,N_13312,N_12119);
nor U14184 (N_14184,N_13200,N_12478);
nand U14185 (N_14185,N_12030,N_13887);
nor U14186 (N_14186,N_13809,N_13591);
and U14187 (N_14187,N_12557,N_13736);
and U14188 (N_14188,N_13368,N_12671);
nand U14189 (N_14189,N_13459,N_13639);
nand U14190 (N_14190,N_12058,N_13999);
and U14191 (N_14191,N_12746,N_12709);
or U14192 (N_14192,N_13436,N_12617);
and U14193 (N_14193,N_13975,N_13106);
nand U14194 (N_14194,N_12073,N_12777);
or U14195 (N_14195,N_13380,N_13460);
nor U14196 (N_14196,N_13945,N_13289);
or U14197 (N_14197,N_13749,N_13913);
nand U14198 (N_14198,N_12435,N_12349);
nand U14199 (N_14199,N_12291,N_13898);
xnor U14200 (N_14200,N_12012,N_12874);
or U14201 (N_14201,N_13113,N_13141);
and U14202 (N_14202,N_13120,N_13774);
or U14203 (N_14203,N_13710,N_12249);
and U14204 (N_14204,N_12861,N_12864);
nand U14205 (N_14205,N_13408,N_13832);
and U14206 (N_14206,N_13959,N_12845);
xor U14207 (N_14207,N_12001,N_12740);
nand U14208 (N_14208,N_12418,N_12547);
xnor U14209 (N_14209,N_13498,N_12620);
and U14210 (N_14210,N_12601,N_12426);
and U14211 (N_14211,N_12238,N_13463);
nand U14212 (N_14212,N_12916,N_13964);
nand U14213 (N_14213,N_13934,N_13199);
nor U14214 (N_14214,N_12137,N_13746);
nor U14215 (N_14215,N_12941,N_12191);
or U14216 (N_14216,N_13027,N_13932);
and U14217 (N_14217,N_13569,N_13627);
or U14218 (N_14218,N_13473,N_13874);
or U14219 (N_14219,N_12705,N_13202);
nor U14220 (N_14220,N_13139,N_12337);
and U14221 (N_14221,N_12190,N_12328);
xnor U14222 (N_14222,N_12917,N_12441);
nor U14223 (N_14223,N_13149,N_13503);
and U14224 (N_14224,N_12103,N_12391);
and U14225 (N_14225,N_12247,N_12380);
or U14226 (N_14226,N_12517,N_12896);
or U14227 (N_14227,N_13904,N_13672);
and U14228 (N_14228,N_13634,N_13900);
nor U14229 (N_14229,N_12665,N_13371);
xor U14230 (N_14230,N_13170,N_13418);
nor U14231 (N_14231,N_13303,N_13589);
nand U14232 (N_14232,N_12223,N_13329);
and U14233 (N_14233,N_12421,N_13482);
or U14234 (N_14234,N_13914,N_12723);
nand U14235 (N_14235,N_12248,N_13422);
and U14236 (N_14236,N_12141,N_13353);
or U14237 (N_14237,N_13159,N_13335);
nor U14238 (N_14238,N_12856,N_12759);
nor U14239 (N_14239,N_13584,N_12140);
nor U14240 (N_14240,N_12331,N_12100);
or U14241 (N_14241,N_13196,N_13491);
nor U14242 (N_14242,N_13475,N_12676);
nand U14243 (N_14243,N_13384,N_13485);
nor U14244 (N_14244,N_13192,N_12186);
and U14245 (N_14245,N_12781,N_12264);
xnor U14246 (N_14246,N_13080,N_13819);
nor U14247 (N_14247,N_13317,N_13127);
xor U14248 (N_14248,N_13903,N_13651);
nor U14249 (N_14249,N_13160,N_13519);
and U14250 (N_14250,N_12626,N_12134);
or U14251 (N_14251,N_12447,N_12733);
or U14252 (N_14252,N_13178,N_12675);
or U14253 (N_14253,N_13654,N_12586);
or U14254 (N_14254,N_12127,N_12108);
nor U14255 (N_14255,N_13146,N_13722);
nor U14256 (N_14256,N_13094,N_12000);
nand U14257 (N_14257,N_13545,N_12237);
xnor U14258 (N_14258,N_13441,N_12364);
and U14259 (N_14259,N_12553,N_13255);
nor U14260 (N_14260,N_12376,N_12884);
nor U14261 (N_14261,N_13064,N_13550);
nand U14262 (N_14262,N_12859,N_12123);
or U14263 (N_14263,N_13467,N_12167);
or U14264 (N_14264,N_12522,N_12498);
or U14265 (N_14265,N_12726,N_13111);
and U14266 (N_14266,N_13431,N_13417);
nor U14267 (N_14267,N_13708,N_13876);
and U14268 (N_14268,N_13624,N_12823);
nand U14269 (N_14269,N_13650,N_13065);
nand U14270 (N_14270,N_12126,N_12455);
xnor U14271 (N_14271,N_13133,N_12965);
nand U14272 (N_14272,N_12178,N_12151);
nor U14273 (N_14273,N_12198,N_13429);
nand U14274 (N_14274,N_13685,N_12589);
nor U14275 (N_14275,N_13849,N_13847);
or U14276 (N_14276,N_12868,N_13530);
nor U14277 (N_14277,N_13376,N_12422);
xnor U14278 (N_14278,N_13318,N_12728);
or U14279 (N_14279,N_12501,N_13177);
nor U14280 (N_14280,N_12483,N_13937);
and U14281 (N_14281,N_13164,N_13271);
nor U14282 (N_14282,N_12304,N_12575);
and U14283 (N_14283,N_12257,N_12336);
nand U14284 (N_14284,N_12900,N_13760);
nand U14285 (N_14285,N_13800,N_12101);
xor U14286 (N_14286,N_13674,N_13265);
nor U14287 (N_14287,N_13529,N_13712);
and U14288 (N_14288,N_12050,N_13750);
nor U14289 (N_14289,N_12510,N_12180);
and U14290 (N_14290,N_12912,N_12899);
nor U14291 (N_14291,N_12144,N_12914);
nand U14292 (N_14292,N_13899,N_13056);
or U14293 (N_14293,N_13062,N_12203);
or U14294 (N_14294,N_12593,N_12645);
xor U14295 (N_14295,N_12752,N_12226);
nor U14296 (N_14296,N_12524,N_12316);
nand U14297 (N_14297,N_12712,N_12775);
nor U14298 (N_14298,N_12890,N_13010);
nor U14299 (N_14299,N_12131,N_13152);
nor U14300 (N_14300,N_13481,N_13535);
xor U14301 (N_14301,N_12059,N_13872);
nand U14302 (N_14302,N_12982,N_12112);
or U14303 (N_14303,N_13968,N_13451);
and U14304 (N_14304,N_12536,N_13019);
nand U14305 (N_14305,N_13426,N_12189);
and U14306 (N_14306,N_13005,N_13327);
nand U14307 (N_14307,N_13308,N_13935);
nand U14308 (N_14308,N_12357,N_12082);
xor U14309 (N_14309,N_13777,N_12725);
and U14310 (N_14310,N_12672,N_12721);
nor U14311 (N_14311,N_13492,N_12323);
nand U14312 (N_14312,N_13824,N_13883);
nand U14313 (N_14313,N_12643,N_13140);
and U14314 (N_14314,N_13471,N_13676);
nor U14315 (N_14315,N_12678,N_13499);
nand U14316 (N_14316,N_13193,N_12756);
and U14317 (N_14317,N_12902,N_12305);
nand U14318 (N_14318,N_12596,N_12179);
nor U14319 (N_14319,N_13831,N_13740);
nor U14320 (N_14320,N_12898,N_13081);
nand U14321 (N_14321,N_12621,N_13727);
nand U14322 (N_14322,N_12734,N_13123);
or U14323 (N_14323,N_13424,N_13502);
nor U14324 (N_14324,N_12836,N_13973);
and U14325 (N_14325,N_12561,N_12296);
xnor U14326 (N_14326,N_13842,N_13373);
and U14327 (N_14327,N_12999,N_13294);
and U14328 (N_14328,N_13956,N_12019);
and U14329 (N_14329,N_13675,N_12843);
and U14330 (N_14330,N_12205,N_12919);
or U14331 (N_14331,N_13412,N_13362);
xnor U14332 (N_14332,N_12812,N_13958);
nor U14333 (N_14333,N_12708,N_13949);
or U14334 (N_14334,N_12468,N_12313);
or U14335 (N_14335,N_13806,N_13523);
xnor U14336 (N_14336,N_13761,N_13986);
nand U14337 (N_14337,N_12425,N_13948);
and U14338 (N_14338,N_13507,N_13602);
or U14339 (N_14339,N_13560,N_13835);
and U14340 (N_14340,N_12968,N_12437);
or U14341 (N_14341,N_12748,N_13379);
or U14342 (N_14342,N_13579,N_13447);
and U14343 (N_14343,N_12862,N_12372);
nand U14344 (N_14344,N_13423,N_12546);
or U14345 (N_14345,N_12322,N_12010);
nor U14346 (N_14346,N_12449,N_13566);
nand U14347 (N_14347,N_12765,N_13877);
or U14348 (N_14348,N_12005,N_12783);
nor U14349 (N_14349,N_13495,N_12953);
or U14350 (N_14350,N_13568,N_13009);
xor U14351 (N_14351,N_13328,N_13078);
or U14352 (N_14352,N_13000,N_12107);
and U14353 (N_14353,N_12217,N_12433);
or U14354 (N_14354,N_13076,N_13434);
or U14355 (N_14355,N_12551,N_13562);
and U14356 (N_14356,N_12817,N_12402);
and U14357 (N_14357,N_12996,N_12260);
or U14358 (N_14358,N_13930,N_13028);
nor U14359 (N_14359,N_12658,N_13580);
or U14360 (N_14360,N_13489,N_12630);
nand U14361 (N_14361,N_12766,N_13762);
nand U14362 (N_14362,N_12983,N_12910);
nor U14363 (N_14363,N_12527,N_12580);
xor U14364 (N_14364,N_13741,N_12950);
and U14365 (N_14365,N_12176,N_12928);
nand U14366 (N_14366,N_13858,N_12695);
nand U14367 (N_14367,N_13287,N_12029);
or U14368 (N_14368,N_12838,N_12473);
nor U14369 (N_14369,N_12306,N_13108);
and U14370 (N_14370,N_13609,N_12051);
nand U14371 (N_14371,N_12653,N_13637);
nand U14372 (N_14372,N_13635,N_13400);
nand U14373 (N_14373,N_12789,N_13506);
or U14374 (N_14374,N_12966,N_12930);
nand U14375 (N_14375,N_12085,N_13325);
and U14376 (N_14376,N_12771,N_13116);
nor U14377 (N_14377,N_13518,N_13739);
and U14378 (N_14378,N_13480,N_13047);
nor U14379 (N_14379,N_12410,N_13068);
nor U14380 (N_14380,N_12292,N_12432);
and U14381 (N_14381,N_13240,N_12246);
or U14382 (N_14382,N_12420,N_13403);
nor U14383 (N_14383,N_13378,N_12673);
nand U14384 (N_14384,N_12071,N_13604);
nor U14385 (N_14385,N_12025,N_12563);
nand U14386 (N_14386,N_13588,N_13861);
or U14387 (N_14387,N_12506,N_12924);
nand U14388 (N_14388,N_13033,N_13235);
and U14389 (N_14389,N_13521,N_12136);
nor U14390 (N_14390,N_12797,N_13500);
and U14391 (N_14391,N_13561,N_12714);
or U14392 (N_14392,N_12116,N_12936);
and U14393 (N_14393,N_12889,N_13001);
and U14394 (N_14394,N_13855,N_12737);
or U14395 (N_14395,N_12570,N_12346);
xnor U14396 (N_14396,N_12147,N_13401);
and U14397 (N_14397,N_13771,N_12476);
nor U14398 (N_14398,N_12955,N_12816);
or U14399 (N_14399,N_13246,N_12674);
nand U14400 (N_14400,N_13222,N_12104);
nand U14401 (N_14401,N_13462,N_13734);
or U14402 (N_14402,N_12744,N_12298);
nor U14403 (N_14403,N_13143,N_12367);
nand U14404 (N_14404,N_12474,N_12525);
nand U14405 (N_14405,N_12946,N_13184);
and U14406 (N_14406,N_12605,N_12267);
and U14407 (N_14407,N_12018,N_13244);
nand U14408 (N_14408,N_13640,N_13841);
and U14409 (N_14409,N_13388,N_12595);
and U14410 (N_14410,N_12780,N_13128);
nand U14411 (N_14411,N_12181,N_13103);
and U14412 (N_14412,N_13030,N_12371);
and U14413 (N_14413,N_12804,N_12622);
or U14414 (N_14414,N_12020,N_13767);
nor U14415 (N_14415,N_12963,N_12668);
and U14416 (N_14416,N_12951,N_12277);
nand U14417 (N_14417,N_12356,N_12979);
nand U14418 (N_14418,N_12314,N_12272);
or U14419 (N_14419,N_12288,N_12164);
nand U14420 (N_14420,N_12445,N_12387);
or U14421 (N_14421,N_12727,N_12096);
nor U14422 (N_14422,N_12087,N_13279);
xnor U14423 (N_14423,N_13314,N_13186);
nor U14424 (N_14424,N_12883,N_12332);
or U14425 (N_14425,N_13018,N_12039);
or U14426 (N_14426,N_12213,N_12600);
nor U14427 (N_14427,N_12826,N_13998);
nor U14428 (N_14428,N_12855,N_12651);
nand U14429 (N_14429,N_12344,N_13225);
nor U14430 (N_14430,N_13454,N_12379);
nor U14431 (N_14431,N_13752,N_12724);
nand U14432 (N_14432,N_13893,N_13117);
nand U14433 (N_14433,N_12374,N_13189);
nor U14434 (N_14434,N_12074,N_12276);
nor U14435 (N_14435,N_13210,N_12929);
and U14436 (N_14436,N_12193,N_12508);
nand U14437 (N_14437,N_12268,N_13970);
or U14438 (N_14438,N_13880,N_12345);
nor U14439 (N_14439,N_13364,N_13419);
and U14440 (N_14440,N_12688,N_13578);
and U14441 (N_14441,N_12614,N_13456);
nand U14442 (N_14442,N_12793,N_13098);
nor U14443 (N_14443,N_12698,N_12286);
nor U14444 (N_14444,N_12206,N_13779);
nor U14445 (N_14445,N_12485,N_13055);
nor U14446 (N_14446,N_13351,N_13668);
or U14447 (N_14447,N_13965,N_12088);
nand U14448 (N_14448,N_12573,N_12574);
nand U14449 (N_14449,N_12224,N_12048);
or U14450 (N_14450,N_13282,N_12528);
and U14451 (N_14451,N_12803,N_13438);
nor U14452 (N_14452,N_13176,N_12741);
and U14453 (N_14453,N_13439,N_12681);
nand U14454 (N_14454,N_13692,N_13788);
or U14455 (N_14455,N_13183,N_13286);
or U14456 (N_14456,N_13283,N_12062);
or U14457 (N_14457,N_12109,N_13190);
xor U14458 (N_14458,N_12256,N_12409);
or U14459 (N_14459,N_13795,N_13003);
and U14460 (N_14460,N_13660,N_12758);
nor U14461 (N_14461,N_13252,N_12294);
nand U14462 (N_14462,N_13590,N_13121);
and U14463 (N_14463,N_13690,N_13733);
or U14464 (N_14464,N_13864,N_13611);
and U14465 (N_14465,N_12407,N_13638);
and U14466 (N_14466,N_13525,N_13045);
xor U14467 (N_14467,N_13022,N_13472);
and U14468 (N_14468,N_12648,N_13758);
or U14469 (N_14469,N_12876,N_12458);
nand U14470 (N_14470,N_13340,N_13002);
nand U14471 (N_14471,N_12065,N_13486);
nand U14472 (N_14472,N_13916,N_12639);
nand U14473 (N_14473,N_12608,N_13667);
xnor U14474 (N_14474,N_12017,N_12948);
or U14475 (N_14475,N_12309,N_13277);
xnor U14476 (N_14476,N_12299,N_12977);
and U14477 (N_14477,N_13625,N_12791);
nor U14478 (N_14478,N_12399,N_13307);
xor U14479 (N_14479,N_12587,N_12138);
and U14480 (N_14480,N_12607,N_13729);
nand U14481 (N_14481,N_13334,N_13450);
nor U14482 (N_14482,N_13680,N_12453);
nor U14483 (N_14483,N_13509,N_13764);
xnor U14484 (N_14484,N_13599,N_13967);
nor U14485 (N_14485,N_12947,N_13886);
nand U14486 (N_14486,N_13154,N_12290);
and U14487 (N_14487,N_13306,N_13977);
or U14488 (N_14488,N_12208,N_12158);
xnor U14489 (N_14489,N_13406,N_12207);
nor U14490 (N_14490,N_12885,N_13790);
nor U14491 (N_14491,N_12319,N_12760);
nor U14492 (N_14492,N_12269,N_12106);
nor U14493 (N_14493,N_13345,N_13206);
and U14494 (N_14494,N_12110,N_12139);
nor U14495 (N_14495,N_12388,N_12556);
nand U14496 (N_14496,N_13032,N_12559);
or U14497 (N_14497,N_12550,N_13137);
nand U14498 (N_14498,N_12006,N_13086);
and U14499 (N_14499,N_13288,N_13856);
nor U14500 (N_14500,N_12685,N_13694);
nor U14501 (N_14501,N_12124,N_12013);
xnor U14502 (N_14502,N_12092,N_13822);
and U14503 (N_14503,N_12722,N_13781);
or U14504 (N_14504,N_13105,N_13698);
and U14505 (N_14505,N_13805,N_12117);
nand U14506 (N_14506,N_13553,N_12480);
nand U14507 (N_14507,N_13902,N_12199);
or U14508 (N_14508,N_13665,N_12219);
and U14509 (N_14509,N_12988,N_13347);
nor U14510 (N_14510,N_12068,N_12667);
nand U14511 (N_14511,N_13510,N_13875);
and U14512 (N_14512,N_12354,N_13751);
xor U14513 (N_14513,N_12800,N_12696);
nor U14514 (N_14514,N_12507,N_12706);
or U14515 (N_14515,N_13280,N_12537);
nand U14516 (N_14516,N_13229,N_13107);
and U14517 (N_14517,N_12584,N_12417);
nand U14518 (N_14518,N_13947,N_13520);
and U14519 (N_14519,N_13995,N_12778);
or U14520 (N_14520,N_12462,N_13405);
and U14521 (N_14521,N_12784,N_13702);
nand U14522 (N_14522,N_13382,N_13185);
nand U14523 (N_14523,N_12469,N_13505);
xnor U14524 (N_14524,N_12656,N_13697);
and U14525 (N_14525,N_12631,N_13274);
nand U14526 (N_14526,N_13082,N_13428);
nor U14527 (N_14527,N_13936,N_12482);
or U14528 (N_14528,N_13787,N_13704);
nor U14529 (N_14529,N_13333,N_13971);
nand U14530 (N_14530,N_13319,N_12962);
or U14531 (N_14531,N_12887,N_12512);
nor U14532 (N_14532,N_13158,N_13259);
and U14533 (N_14533,N_12054,N_13214);
xor U14534 (N_14534,N_12679,N_12976);
or U14535 (N_14535,N_13079,N_13596);
nand U14536 (N_14536,N_12429,N_13465);
and U14537 (N_14537,N_12704,N_13567);
or U14538 (N_14538,N_13386,N_13326);
and U14539 (N_14539,N_12670,N_13217);
nand U14540 (N_14540,N_12650,N_13536);
nor U14541 (N_14541,N_13248,N_13616);
nor U14542 (N_14542,N_13501,N_12275);
and U14543 (N_14543,N_13843,N_13955);
nor U14544 (N_14544,N_13060,N_13359);
or U14545 (N_14545,N_13444,N_13541);
or U14546 (N_14546,N_13039,N_13354);
nand U14547 (N_14547,N_12519,N_12129);
or U14548 (N_14548,N_12279,N_13866);
nor U14549 (N_14549,N_12931,N_13918);
and U14550 (N_14550,N_13458,N_13896);
and U14551 (N_14551,N_13349,N_13261);
nor U14552 (N_14552,N_12169,N_13791);
nand U14553 (N_14553,N_13850,N_13344);
or U14554 (N_14554,N_12035,N_12989);
nand U14555 (N_14555,N_12404,N_13961);
and U14556 (N_14556,N_12523,N_13034);
nor U14557 (N_14557,N_12022,N_12597);
and U14558 (N_14558,N_12099,N_12490);
or U14559 (N_14559,N_12080,N_12244);
nor U14560 (N_14560,N_12602,N_12278);
nand U14561 (N_14561,N_12629,N_13647);
and U14562 (N_14562,N_13910,N_12084);
nor U14563 (N_14563,N_13670,N_12097);
nor U14564 (N_14564,N_13468,N_13570);
nor U14565 (N_14565,N_12933,N_13093);
xor U14566 (N_14566,N_12647,N_12538);
nand U14567 (N_14567,N_13257,N_13960);
or U14568 (N_14568,N_12549,N_13072);
nor U14569 (N_14569,N_13134,N_12066);
xnor U14570 (N_14570,N_13731,N_13565);
nand U14571 (N_14571,N_12718,N_12870);
xor U14572 (N_14572,N_12424,N_12825);
or U14573 (N_14573,N_13024,N_13759);
and U14574 (N_14574,N_13928,N_13237);
and U14575 (N_14575,N_13621,N_12202);
nor U14576 (N_14576,N_12687,N_13693);
nand U14577 (N_14577,N_12452,N_12368);
xor U14578 (N_14578,N_12821,N_13617);
and U14579 (N_14579,N_13440,N_12369);
or U14580 (N_14580,N_12984,N_13049);
and U14581 (N_14581,N_13394,N_13011);
and U14582 (N_14582,N_13369,N_13919);
nor U14583 (N_14583,N_13784,N_12412);
and U14584 (N_14584,N_12324,N_12295);
xor U14585 (N_14585,N_13871,N_13194);
nor U14586 (N_14586,N_13743,N_12909);
nand U14587 (N_14587,N_13487,N_13276);
nor U14588 (N_14588,N_12959,N_13631);
and U14589 (N_14589,N_12616,N_13924);
and U14590 (N_14590,N_12534,N_12841);
and U14591 (N_14591,N_12911,N_13042);
or U14592 (N_14592,N_13413,N_12554);
nor U14593 (N_14593,N_13963,N_12310);
or U14594 (N_14594,N_12363,N_13564);
and U14595 (N_14595,N_13833,N_12502);
or U14596 (N_14596,N_12232,N_13104);
nor U14597 (N_14597,N_12083,N_12301);
and U14598 (N_14598,N_12133,N_13593);
nand U14599 (N_14599,N_13622,N_13138);
or U14600 (N_14600,N_13469,N_13054);
or U14601 (N_14601,N_13802,N_12079);
xnor U14602 (N_14602,N_12263,N_13031);
nor U14603 (N_14603,N_13008,N_13649);
and U14604 (N_14604,N_12153,N_13316);
xor U14605 (N_14605,N_13844,N_12044);
nor U14606 (N_14606,N_12794,N_12731);
and U14607 (N_14607,N_13182,N_12182);
nor U14608 (N_14608,N_13313,N_13171);
nand U14609 (N_14609,N_13768,N_13909);
nand U14610 (N_14610,N_13829,N_13224);
nor U14611 (N_14611,N_12053,N_13618);
or U14612 (N_14612,N_12183,N_12444);
nand U14613 (N_14613,N_13643,N_13013);
nor U14614 (N_14614,N_13264,N_12197);
nand U14615 (N_14615,N_13922,N_12567);
and U14616 (N_14616,N_12509,N_13360);
xnor U14617 (N_14617,N_13595,N_12231);
nand U14618 (N_14618,N_13298,N_12873);
nand U14619 (N_14619,N_12814,N_13448);
nor U14620 (N_14620,N_12343,N_13058);
or U14621 (N_14621,N_12613,N_13851);
nor U14622 (N_14622,N_12839,N_13552);
and U14623 (N_14623,N_13583,N_13052);
or U14624 (N_14624,N_12239,N_12847);
nor U14625 (N_14625,N_12768,N_12923);
nand U14626 (N_14626,N_12937,N_12666);
and U14627 (N_14627,N_13539,N_12353);
or U14628 (N_14628,N_12114,N_13641);
or U14629 (N_14629,N_12282,N_12822);
and U14630 (N_14630,N_12145,N_12633);
or U14631 (N_14631,N_13172,N_12878);
nand U14632 (N_14632,N_12581,N_12229);
nor U14633 (N_14633,N_13059,N_12382);
nand U14634 (N_14634,N_13012,N_12091);
or U14635 (N_14635,N_13040,N_13180);
nor U14636 (N_14636,N_12064,N_12960);
or U14637 (N_14637,N_12415,N_13988);
and U14638 (N_14638,N_13398,N_12918);
xor U14639 (N_14639,N_12949,N_13219);
nand U14640 (N_14640,N_13242,N_13483);
nor U14641 (N_14641,N_12590,N_12423);
nand U14642 (N_14642,N_13980,N_13695);
nor U14643 (N_14643,N_12265,N_12513);
or U14644 (N_14644,N_12395,N_12684);
nor U14645 (N_14645,N_12491,N_12786);
nand U14646 (N_14646,N_13852,N_12833);
nand U14647 (N_14647,N_13310,N_12618);
xnor U14648 (N_14648,N_13389,N_13839);
xor U14649 (N_14649,N_13091,N_12401);
nor U14650 (N_14650,N_12779,N_13470);
xor U14651 (N_14651,N_12466,N_12904);
nand U14652 (N_14652,N_12359,N_13278);
and U14653 (N_14653,N_13407,N_13575);
nand U14654 (N_14654,N_12893,N_13612);
nand U14655 (N_14655,N_12261,N_13437);
nand U14656 (N_14656,N_13952,N_13513);
or U14657 (N_14657,N_12063,N_12956);
or U14658 (N_14658,N_12735,N_12366);
nor U14659 (N_14659,N_12830,N_13321);
or U14660 (N_14660,N_12903,N_12118);
nor U14661 (N_14661,N_12488,N_12927);
and U14662 (N_14662,N_13410,N_12230);
or U14663 (N_14663,N_13531,N_12612);
and U14664 (N_14664,N_13073,N_13163);
nor U14665 (N_14665,N_12762,N_13757);
or U14666 (N_14666,N_12747,N_13381);
and U14667 (N_14667,N_12479,N_13925);
xor U14668 (N_14668,N_13773,N_13455);
xor U14669 (N_14669,N_12400,N_13110);
nand U14670 (N_14670,N_13017,N_13221);
and U14671 (N_14671,N_12188,N_13243);
and U14672 (N_14672,N_12348,N_13632);
and U14673 (N_14673,N_13785,N_13747);
nand U14674 (N_14674,N_13854,N_13923);
nand U14675 (N_14675,N_12763,N_12477);
or U14676 (N_14676,N_12055,N_12072);
xnor U14677 (N_14677,N_13304,N_12961);
nand U14678 (N_14678,N_12406,N_13067);
nand U14679 (N_14679,N_12090,N_13814);
or U14680 (N_14680,N_12545,N_12274);
and U14681 (N_14681,N_12964,N_12408);
nor U14682 (N_14682,N_12113,N_13608);
and U14683 (N_14683,N_12184,N_13338);
nor U14684 (N_14684,N_13126,N_12003);
nand U14685 (N_14685,N_13863,N_13320);
and U14686 (N_14686,N_13322,N_12732);
xor U14687 (N_14687,N_12555,N_13494);
and U14688 (N_14688,N_13581,N_12700);
or U14689 (N_14689,N_13869,N_13155);
or U14690 (N_14690,N_12243,N_12077);
and U14691 (N_14691,N_12935,N_13323);
and U14692 (N_14692,N_12287,N_12008);
and U14693 (N_14693,N_12460,N_12334);
or U14694 (N_14694,N_12635,N_13563);
nand U14695 (N_14695,N_12981,N_13859);
or U14696 (N_14696,N_12098,N_13912);
and U14697 (N_14697,N_12591,N_12450);
and U14698 (N_14698,N_12165,N_12592);
or U14699 (N_14699,N_13512,N_12266);
and U14700 (N_14700,N_12234,N_12598);
nor U14701 (N_14701,N_12854,N_13538);
nor U14702 (N_14702,N_12250,N_13356);
nand U14703 (N_14703,N_12236,N_12241);
or U14704 (N_14704,N_13397,N_13239);
or U14705 (N_14705,N_12338,N_12032);
and U14706 (N_14706,N_13051,N_13737);
or U14707 (N_14707,N_12398,N_13285);
or U14708 (N_14708,N_13387,N_13092);
nor U14709 (N_14709,N_12627,N_13476);
or U14710 (N_14710,N_13046,N_12649);
nor U14711 (N_14711,N_12558,N_12228);
and U14712 (N_14712,N_12835,N_13187);
or U14713 (N_14713,N_13195,N_13102);
and U14714 (N_14714,N_12975,N_12235);
and U14715 (N_14715,N_12428,N_12500);
and U14716 (N_14716,N_12659,N_13250);
or U14717 (N_14717,N_13921,N_12185);
nor U14718 (N_14718,N_13614,N_13534);
xor U14719 (N_14719,N_12143,N_12464);
nor U14720 (N_14720,N_12922,N_12457);
nor U14721 (N_14721,N_12467,N_12440);
nor U14722 (N_14722,N_12751,N_12403);
and U14723 (N_14723,N_13112,N_12216);
nand U14724 (N_14724,N_12505,N_13799);
xnor U14725 (N_14725,N_12720,N_12664);
xnor U14726 (N_14726,N_13522,N_12148);
nor U14727 (N_14727,N_12863,N_12703);
nor U14728 (N_14728,N_12451,N_13821);
or U14729 (N_14729,N_12162,N_13885);
nand U14730 (N_14730,N_13646,N_12283);
xnor U14731 (N_14731,N_12484,N_12443);
nand U14732 (N_14732,N_13157,N_12390);
nor U14733 (N_14733,N_13950,N_13894);
or U14734 (N_14734,N_13272,N_12220);
xnor U14735 (N_14735,N_12540,N_12105);
xnor U14736 (N_14736,N_12086,N_13148);
nand U14737 (N_14737,N_12945,N_12942);
nand U14738 (N_14738,N_13267,N_13097);
nand U14739 (N_14739,N_12102,N_12773);
and U14740 (N_14740,N_13393,N_13181);
or U14741 (N_14741,N_12394,N_13897);
or U14742 (N_14742,N_12308,N_13994);
or U14743 (N_14743,N_12757,N_12564);
nor U14744 (N_14744,N_12327,N_13305);
or U14745 (N_14745,N_12807,N_13857);
nor U14746 (N_14746,N_13556,N_13296);
nor U14747 (N_14747,N_13269,N_13301);
or U14748 (N_14748,N_12624,N_13477);
nor U14749 (N_14749,N_13220,N_12365);
nand U14750 (N_14750,N_13713,N_13586);
and U14751 (N_14751,N_12693,N_12532);
nand U14752 (N_14752,N_12669,N_12222);
nand U14753 (N_14753,N_12697,N_12971);
and U14754 (N_14754,N_12330,N_13830);
or U14755 (N_14755,N_13548,N_12307);
nand U14756 (N_14756,N_12713,N_12610);
nand U14757 (N_14757,N_12609,N_12252);
nand U14758 (N_14758,N_13263,N_12069);
or U14759 (N_14759,N_12761,N_12439);
nand U14760 (N_14760,N_12492,N_12386);
nand U14761 (N_14761,N_13908,N_12560);
xor U14762 (N_14762,N_13848,N_12599);
nand U14763 (N_14763,N_12520,N_12710);
xnor U14764 (N_14764,N_12037,N_12075);
or U14765 (N_14765,N_13236,N_12895);
and U14766 (N_14766,N_13197,N_13165);
nand U14767 (N_14767,N_12471,N_13946);
and U14768 (N_14768,N_12819,N_13636);
nor U14769 (N_14769,N_13130,N_12707);
xnor U14770 (N_14770,N_13873,N_12853);
xor U14771 (N_14771,N_13982,N_13457);
or U14772 (N_14772,N_13115,N_13006);
nor U14773 (N_14773,N_13628,N_12038);
or U14774 (N_14774,N_12827,N_12967);
and U14775 (N_14775,N_12259,N_12489);
nand U14776 (N_14776,N_12121,N_12729);
or U14777 (N_14777,N_13820,N_13816);
and U14778 (N_14778,N_13940,N_13275);
or U14779 (N_14779,N_13151,N_12475);
nor U14780 (N_14780,N_13358,N_12738);
nor U14781 (N_14781,N_12168,N_13655);
nor U14782 (N_14782,N_13544,N_12637);
nor U14783 (N_14783,N_13361,N_12691);
and U14784 (N_14784,N_12872,N_12041);
nor U14785 (N_14785,N_12795,N_13207);
nor U14786 (N_14786,N_13689,N_12015);
and U14787 (N_14787,N_12033,N_12504);
nor U14788 (N_14788,N_12745,N_12882);
nand U14789 (N_14789,N_13493,N_13057);
or U14790 (N_14790,N_12657,N_12993);
nand U14791 (N_14791,N_12515,N_12615);
nand U14792 (N_14792,N_12470,N_12312);
nor U14793 (N_14793,N_12195,N_12776);
xor U14794 (N_14794,N_12806,N_13496);
xor U14795 (N_14795,N_12588,N_13725);
or U14796 (N_14796,N_12413,N_13150);
nor U14797 (N_14797,N_13415,N_12297);
xnor U14798 (N_14798,N_12511,N_12694);
nand U14799 (N_14799,N_13085,N_12541);
nor U14800 (N_14800,N_12200,N_12769);
nand U14801 (N_14801,N_12049,N_13678);
nand U14802 (N_14802,N_13260,N_13656);
and U14803 (N_14803,N_12837,N_12682);
nor U14804 (N_14804,N_13336,N_12891);
or U14805 (N_14805,N_12970,N_12258);
nand U14806 (N_14806,N_12004,N_12844);
or U14807 (N_14807,N_12552,N_12201);
or U14808 (N_14808,N_13453,N_13377);
or U14809 (N_14809,N_12925,N_13089);
or U14810 (N_14810,N_13901,N_12991);
xor U14811 (N_14811,N_13063,N_12644);
nor U14812 (N_14812,N_12808,N_13430);
and U14813 (N_14813,N_12427,N_12585);
nor U14814 (N_14814,N_13987,N_12014);
or U14815 (N_14815,N_12430,N_13700);
or U14816 (N_14816,N_12915,N_12221);
nor U14817 (N_14817,N_13881,N_13597);
or U14818 (N_14818,N_12849,N_13783);
nor U14819 (N_14819,N_13173,N_12952);
xor U14820 (N_14820,N_13585,N_13041);
and U14821 (N_14821,N_12135,N_13490);
xnor U14822 (N_14822,N_12174,N_13684);
nor U14823 (N_14823,N_12892,N_13728);
nand U14824 (N_14824,N_12211,N_13029);
nor U14825 (N_14825,N_13391,N_13511);
nor U14826 (N_14826,N_13324,N_12373);
nor U14827 (N_14827,N_13865,N_12926);
nor U14828 (N_14828,N_12218,N_13592);
and U14829 (N_14829,N_13911,N_13129);
nand U14830 (N_14830,N_13302,N_12225);
nor U14831 (N_14831,N_12329,N_12802);
or U14832 (N_14832,N_13879,N_12254);
or U14833 (N_14833,N_13118,N_13792);
and U14834 (N_14834,N_12634,N_13542);
nand U14835 (N_14835,N_13125,N_12974);
or U14836 (N_14836,N_12998,N_13043);
and U14837 (N_14837,N_13915,N_13119);
or U14838 (N_14838,N_13686,N_13153);
nor U14839 (N_14839,N_13446,N_13755);
xor U14840 (N_14840,N_13218,N_13309);
nor U14841 (N_14841,N_13644,N_13984);
nand U14842 (N_14842,N_12533,N_13228);
nor U14843 (N_14843,N_12481,N_12743);
or U14844 (N_14844,N_13991,N_13109);
and U14845 (N_14845,N_13688,N_13605);
xnor U14846 (N_14846,N_13962,N_13794);
nand U14847 (N_14847,N_13840,N_12692);
and U14848 (N_14848,N_12846,N_12972);
or U14849 (N_14849,N_13633,N_13753);
and U14850 (N_14850,N_12156,N_12702);
nand U14851 (N_14851,N_12565,N_13142);
nand U14852 (N_14852,N_12699,N_13425);
or U14853 (N_14853,N_12204,N_12886);
nand U14854 (N_14854,N_12320,N_13549);
nor U14855 (N_14855,N_12809,N_13663);
or U14856 (N_14856,N_12340,N_13363);
xor U14857 (N_14857,N_13882,N_12535);
and U14858 (N_14858,N_12171,N_12603);
nand U14859 (N_14859,N_13537,N_13392);
and U14860 (N_14860,N_12973,N_13238);
and U14861 (N_14861,N_13432,N_13366);
and U14862 (N_14862,N_13020,N_12848);
nor U14863 (N_14863,N_12661,N_13135);
and U14864 (N_14864,N_13610,N_13895);
or U14865 (N_14865,N_12894,N_13920);
or U14866 (N_14866,N_13803,N_13778);
and U14867 (N_14867,N_13517,N_13868);
or U14868 (N_14868,N_12980,N_13527);
nand U14869 (N_14869,N_13048,N_13077);
nor U14870 (N_14870,N_12578,N_13719);
and U14871 (N_14871,N_12411,N_13433);
or U14872 (N_14872,N_13682,N_12568);
and U14873 (N_14873,N_12021,N_12719);
nor U14874 (N_14874,N_12146,N_12623);
and U14875 (N_14875,N_13209,N_13299);
nand U14876 (N_14876,N_12997,N_12940);
nor U14877 (N_14877,N_13348,N_13331);
xnor U14878 (N_14878,N_12377,N_13007);
nand U14879 (N_14879,N_13374,N_12920);
nand U14880 (N_14880,N_13071,N_13343);
or U14881 (N_14881,N_13466,N_12431);
nand U14882 (N_14882,N_12381,N_13657);
and U14883 (N_14883,N_13191,N_13951);
and U14884 (N_14884,N_13131,N_13083);
xor U14885 (N_14885,N_13074,N_13744);
nor U14886 (N_14886,N_13626,N_13642);
xnor U14887 (N_14887,N_13804,N_13297);
or U14888 (N_14888,N_12067,N_13101);
and U14889 (N_14889,N_12214,N_13488);
nand U14890 (N_14890,N_12499,N_13718);
and U14891 (N_14891,N_12378,N_13036);
nor U14892 (N_14892,N_12496,N_13979);
nor U14893 (N_14893,N_13607,N_12985);
and U14894 (N_14894,N_13526,N_13707);
and U14895 (N_14895,N_12251,N_12990);
and U14896 (N_14896,N_12212,N_13330);
nand U14897 (N_14897,N_12548,N_13095);
nor U14898 (N_14898,N_13615,N_13203);
or U14899 (N_14899,N_13156,N_12888);
and U14900 (N_14900,N_13367,N_13997);
nand U14901 (N_14901,N_13293,N_12240);
or U14902 (N_14902,N_12461,N_13825);
nor U14903 (N_14903,N_12161,N_12566);
nor U14904 (N_14904,N_13132,N_13846);
nor U14905 (N_14905,N_13122,N_13205);
xnor U14906 (N_14906,N_13603,N_13699);
nand U14907 (N_14907,N_12061,N_13766);
or U14908 (N_14908,N_12046,N_13669);
nor U14909 (N_14909,N_13720,N_12969);
nor U14910 (N_14910,N_13938,N_12271);
xnor U14911 (N_14911,N_12317,N_13927);
and U14912 (N_14912,N_12736,N_13715);
nand U14913 (N_14913,N_13053,N_13528);
xor U14914 (N_14914,N_12360,N_12370);
xnor U14915 (N_14915,N_13653,N_12384);
or U14916 (N_14916,N_13245,N_13888);
and U14917 (N_14917,N_12638,N_13917);
nand U14918 (N_14918,N_12253,N_13557);
or U14919 (N_14919,N_12155,N_13551);
xnor U14920 (N_14920,N_12043,N_12333);
or U14921 (N_14921,N_12215,N_13421);
nand U14922 (N_14922,N_13295,N_13717);
nor U14923 (N_14923,N_13989,N_12303);
and U14924 (N_14924,N_13478,N_12300);
nand U14925 (N_14925,N_13810,N_12810);
nand U14926 (N_14926,N_12361,N_12820);
nand U14927 (N_14927,N_12518,N_13372);
or U14928 (N_14928,N_13061,N_12824);
nor U14929 (N_14929,N_13342,N_13188);
nor U14930 (N_14930,N_13037,N_12571);
nand U14931 (N_14931,N_12834,N_13812);
xor U14932 (N_14932,N_12582,N_12871);
nand U14933 (N_14933,N_12289,N_12943);
and U14934 (N_14934,N_12787,N_12149);
or U14935 (N_14935,N_12739,N_13797);
and U14936 (N_14936,N_13981,N_13161);
and U14937 (N_14937,N_13445,N_13664);
nand U14938 (N_14938,N_13671,N_13147);
and U14939 (N_14939,N_13474,N_12865);
and U14940 (N_14940,N_13162,N_13714);
nor U14941 (N_14941,N_12057,N_13452);
nor U14942 (N_14942,N_13247,N_13204);
nand U14943 (N_14943,N_13166,N_12027);
or U14944 (N_14944,N_12355,N_12921);
xnor U14945 (N_14945,N_13944,N_13023);
xor U14946 (N_14946,N_12009,N_12790);
xnor U14947 (N_14947,N_13658,N_12095);
or U14948 (N_14948,N_13711,N_13281);
nor U14949 (N_14949,N_13290,N_13256);
nand U14950 (N_14950,N_12818,N_13514);
nor U14951 (N_14951,N_12392,N_13770);
nand U14952 (N_14952,N_13978,N_12529);
and U14953 (N_14953,N_13337,N_12583);
or U14954 (N_14954,N_12419,N_13853);
nand U14955 (N_14955,N_12715,N_13623);
nand U14956 (N_14956,N_12750,N_13620);
nand U14957 (N_14957,N_12414,N_13573);
nand U14958 (N_14958,N_13870,N_13396);
nor U14959 (N_14959,N_12245,N_13696);
nand U14960 (N_14960,N_13926,N_12662);
and U14961 (N_14961,N_12163,N_13929);
or U14962 (N_14962,N_12628,N_12242);
or U14963 (N_14963,N_12742,N_12152);
or U14964 (N_14964,N_12089,N_12111);
nand U14965 (N_14965,N_12562,N_13993);
or U14966 (N_14966,N_12641,N_12749);
nand U14967 (N_14967,N_13953,N_13026);
or U14968 (N_14968,N_12906,N_13996);
nor U14969 (N_14969,N_13227,N_13300);
or U14970 (N_14970,N_13701,N_12132);
nor U14971 (N_14971,N_12632,N_13088);
and U14972 (N_14972,N_13357,N_12939);
nor U14973 (N_14973,N_12858,N_13677);
and U14974 (N_14974,N_12572,N_13990);
nand U14975 (N_14975,N_12811,N_12389);
nand U14976 (N_14976,N_13273,N_12879);
or U14977 (N_14977,N_12636,N_12007);
xnor U14978 (N_14978,N_12717,N_13284);
xor U14979 (N_14979,N_12060,N_12175);
nor U14980 (N_14980,N_12857,N_12992);
and U14981 (N_14981,N_12683,N_12284);
xnor U14982 (N_14982,N_13629,N_12755);
and U14983 (N_14983,N_13532,N_12579);
and U14984 (N_14984,N_12128,N_13648);
nor U14985 (N_14985,N_13038,N_13014);
nor U14986 (N_14986,N_13726,N_12465);
and U14987 (N_14987,N_12028,N_12436);
xnor U14988 (N_14988,N_12619,N_12994);
and U14989 (N_14989,N_12442,N_12177);
nor U14990 (N_14990,N_13395,N_13817);
or U14991 (N_14991,N_12680,N_13793);
or U14992 (N_14992,N_12852,N_12150);
or U14993 (N_14993,N_13748,N_13826);
nand U14994 (N_14994,N_12026,N_12270);
nand U14995 (N_14995,N_12396,N_12434);
xor U14996 (N_14996,N_12342,N_12045);
and U14997 (N_14997,N_13907,N_13860);
nand U14998 (N_14998,N_13661,N_13390);
or U14999 (N_14999,N_12285,N_13765);
and U15000 (N_15000,N_12789,N_13638);
or U15001 (N_15001,N_12720,N_13306);
or U15002 (N_15002,N_13049,N_12145);
or U15003 (N_15003,N_13467,N_13349);
or U15004 (N_15004,N_13864,N_13170);
or U15005 (N_15005,N_12400,N_13129);
and U15006 (N_15006,N_13619,N_13875);
and U15007 (N_15007,N_13765,N_13391);
nand U15008 (N_15008,N_13979,N_12368);
or U15009 (N_15009,N_12092,N_12873);
nand U15010 (N_15010,N_13602,N_13942);
or U15011 (N_15011,N_13780,N_12912);
and U15012 (N_15012,N_12196,N_12209);
nand U15013 (N_15013,N_13022,N_12121);
or U15014 (N_15014,N_13667,N_13220);
nor U15015 (N_15015,N_12322,N_13673);
or U15016 (N_15016,N_13088,N_13164);
and U15017 (N_15017,N_13841,N_13520);
or U15018 (N_15018,N_12596,N_13010);
and U15019 (N_15019,N_12101,N_12423);
nor U15020 (N_15020,N_13772,N_13365);
or U15021 (N_15021,N_12526,N_13161);
xor U15022 (N_15022,N_13799,N_12013);
xnor U15023 (N_15023,N_13608,N_12178);
nor U15024 (N_15024,N_12743,N_12547);
nand U15025 (N_15025,N_13407,N_12440);
xor U15026 (N_15026,N_12291,N_12392);
nand U15027 (N_15027,N_13741,N_12852);
xnor U15028 (N_15028,N_13753,N_12833);
or U15029 (N_15029,N_12693,N_13750);
or U15030 (N_15030,N_13207,N_12911);
and U15031 (N_15031,N_12717,N_12722);
nor U15032 (N_15032,N_12924,N_13972);
nand U15033 (N_15033,N_12835,N_13050);
and U15034 (N_15034,N_13198,N_12235);
nor U15035 (N_15035,N_13055,N_12122);
and U15036 (N_15036,N_13414,N_12231);
and U15037 (N_15037,N_12377,N_13264);
nand U15038 (N_15038,N_12441,N_13218);
or U15039 (N_15039,N_12638,N_12549);
and U15040 (N_15040,N_13899,N_12723);
nor U15041 (N_15041,N_13407,N_12611);
xor U15042 (N_15042,N_12642,N_12529);
and U15043 (N_15043,N_12880,N_13564);
and U15044 (N_15044,N_12333,N_13745);
xor U15045 (N_15045,N_12592,N_12786);
xor U15046 (N_15046,N_12818,N_12779);
xor U15047 (N_15047,N_12035,N_12472);
and U15048 (N_15048,N_12238,N_13168);
or U15049 (N_15049,N_13211,N_13955);
nor U15050 (N_15050,N_12107,N_12283);
xnor U15051 (N_15051,N_13477,N_13784);
or U15052 (N_15052,N_12563,N_13008);
and U15053 (N_15053,N_13401,N_13901);
or U15054 (N_15054,N_13927,N_12251);
nand U15055 (N_15055,N_12605,N_12170);
or U15056 (N_15056,N_13069,N_12188);
and U15057 (N_15057,N_12978,N_13853);
and U15058 (N_15058,N_13013,N_12196);
and U15059 (N_15059,N_13701,N_13453);
nor U15060 (N_15060,N_12507,N_13151);
or U15061 (N_15061,N_12388,N_12810);
or U15062 (N_15062,N_12133,N_12607);
or U15063 (N_15063,N_13809,N_12809);
nor U15064 (N_15064,N_12220,N_13664);
and U15065 (N_15065,N_13646,N_13699);
nand U15066 (N_15066,N_12483,N_13635);
nand U15067 (N_15067,N_12413,N_13865);
nand U15068 (N_15068,N_13987,N_13430);
nor U15069 (N_15069,N_12480,N_12652);
nor U15070 (N_15070,N_13113,N_13957);
nand U15071 (N_15071,N_12600,N_12457);
xnor U15072 (N_15072,N_13804,N_12579);
or U15073 (N_15073,N_13538,N_12671);
nor U15074 (N_15074,N_13341,N_12918);
xnor U15075 (N_15075,N_13252,N_12374);
nor U15076 (N_15076,N_12093,N_12787);
and U15077 (N_15077,N_13691,N_12059);
or U15078 (N_15078,N_12568,N_12702);
nand U15079 (N_15079,N_13156,N_13549);
or U15080 (N_15080,N_12552,N_13576);
nor U15081 (N_15081,N_13750,N_12968);
or U15082 (N_15082,N_12681,N_12742);
nor U15083 (N_15083,N_12689,N_13595);
or U15084 (N_15084,N_13870,N_13399);
and U15085 (N_15085,N_12542,N_12407);
or U15086 (N_15086,N_13802,N_12517);
nand U15087 (N_15087,N_13287,N_12568);
xor U15088 (N_15088,N_13555,N_12105);
nor U15089 (N_15089,N_13375,N_13490);
nand U15090 (N_15090,N_12113,N_12712);
nor U15091 (N_15091,N_13485,N_13882);
or U15092 (N_15092,N_13715,N_12323);
nor U15093 (N_15093,N_13827,N_13179);
and U15094 (N_15094,N_12454,N_12331);
or U15095 (N_15095,N_12158,N_12303);
or U15096 (N_15096,N_13037,N_12195);
xnor U15097 (N_15097,N_12002,N_12371);
and U15098 (N_15098,N_12593,N_12038);
nor U15099 (N_15099,N_12081,N_13020);
and U15100 (N_15100,N_13039,N_12344);
nand U15101 (N_15101,N_12706,N_12205);
xor U15102 (N_15102,N_12063,N_13784);
or U15103 (N_15103,N_13974,N_13703);
and U15104 (N_15104,N_13615,N_13387);
or U15105 (N_15105,N_12226,N_13065);
or U15106 (N_15106,N_12467,N_12978);
nand U15107 (N_15107,N_12541,N_13786);
or U15108 (N_15108,N_12326,N_12916);
nand U15109 (N_15109,N_12274,N_13900);
or U15110 (N_15110,N_13391,N_13814);
and U15111 (N_15111,N_13307,N_12113);
or U15112 (N_15112,N_13296,N_13999);
nand U15113 (N_15113,N_12085,N_13102);
or U15114 (N_15114,N_13103,N_12775);
and U15115 (N_15115,N_13942,N_12390);
xnor U15116 (N_15116,N_12045,N_12575);
xor U15117 (N_15117,N_13065,N_12295);
nand U15118 (N_15118,N_13999,N_13297);
and U15119 (N_15119,N_13443,N_12448);
nand U15120 (N_15120,N_13225,N_13794);
nor U15121 (N_15121,N_12479,N_12946);
nor U15122 (N_15122,N_12793,N_12499);
and U15123 (N_15123,N_12997,N_13591);
and U15124 (N_15124,N_13991,N_13810);
or U15125 (N_15125,N_12401,N_12690);
nor U15126 (N_15126,N_13661,N_13270);
xnor U15127 (N_15127,N_13934,N_13013);
or U15128 (N_15128,N_13168,N_13190);
and U15129 (N_15129,N_13491,N_13086);
nand U15130 (N_15130,N_13619,N_13466);
or U15131 (N_15131,N_12033,N_12510);
and U15132 (N_15132,N_12677,N_13206);
and U15133 (N_15133,N_13732,N_12138);
nand U15134 (N_15134,N_12006,N_13420);
nand U15135 (N_15135,N_13102,N_12306);
xor U15136 (N_15136,N_13550,N_12660);
and U15137 (N_15137,N_12555,N_13190);
or U15138 (N_15138,N_12136,N_13427);
or U15139 (N_15139,N_12625,N_13404);
nand U15140 (N_15140,N_12914,N_13294);
nor U15141 (N_15141,N_13897,N_12332);
and U15142 (N_15142,N_12485,N_12107);
nor U15143 (N_15143,N_13542,N_13962);
xnor U15144 (N_15144,N_12216,N_12765);
nand U15145 (N_15145,N_13369,N_12679);
nand U15146 (N_15146,N_13583,N_13207);
nor U15147 (N_15147,N_12875,N_13732);
nor U15148 (N_15148,N_12573,N_13528);
and U15149 (N_15149,N_12652,N_13345);
nor U15150 (N_15150,N_13371,N_13288);
nor U15151 (N_15151,N_12137,N_12105);
nor U15152 (N_15152,N_13106,N_13435);
and U15153 (N_15153,N_12925,N_12821);
and U15154 (N_15154,N_13048,N_13938);
nor U15155 (N_15155,N_13948,N_12303);
nor U15156 (N_15156,N_12483,N_13602);
or U15157 (N_15157,N_12669,N_13272);
and U15158 (N_15158,N_12419,N_13263);
nor U15159 (N_15159,N_13429,N_12018);
and U15160 (N_15160,N_12861,N_13418);
nor U15161 (N_15161,N_12804,N_12302);
or U15162 (N_15162,N_12015,N_12116);
nor U15163 (N_15163,N_12549,N_13871);
and U15164 (N_15164,N_12230,N_13926);
and U15165 (N_15165,N_12454,N_12367);
nor U15166 (N_15166,N_13070,N_12593);
xor U15167 (N_15167,N_13760,N_12159);
nand U15168 (N_15168,N_12706,N_13142);
nor U15169 (N_15169,N_12050,N_12691);
nand U15170 (N_15170,N_13649,N_13582);
xor U15171 (N_15171,N_13087,N_13708);
or U15172 (N_15172,N_12578,N_13015);
or U15173 (N_15173,N_13927,N_12560);
and U15174 (N_15174,N_12265,N_13573);
nor U15175 (N_15175,N_13110,N_12429);
and U15176 (N_15176,N_13900,N_12940);
nor U15177 (N_15177,N_13349,N_12486);
or U15178 (N_15178,N_13812,N_12749);
and U15179 (N_15179,N_13071,N_13139);
nor U15180 (N_15180,N_13149,N_12187);
and U15181 (N_15181,N_12862,N_13036);
or U15182 (N_15182,N_12636,N_12956);
nand U15183 (N_15183,N_13806,N_13569);
nor U15184 (N_15184,N_13126,N_13083);
xnor U15185 (N_15185,N_13190,N_13715);
nand U15186 (N_15186,N_13920,N_12306);
nand U15187 (N_15187,N_12374,N_13038);
nor U15188 (N_15188,N_12018,N_12381);
nand U15189 (N_15189,N_12713,N_13643);
or U15190 (N_15190,N_13835,N_12019);
nand U15191 (N_15191,N_12176,N_13239);
xor U15192 (N_15192,N_13054,N_13401);
nor U15193 (N_15193,N_13901,N_13645);
nand U15194 (N_15194,N_12146,N_12010);
nor U15195 (N_15195,N_13813,N_12506);
and U15196 (N_15196,N_12645,N_12187);
nor U15197 (N_15197,N_13975,N_13272);
and U15198 (N_15198,N_12937,N_13163);
xor U15199 (N_15199,N_12828,N_13598);
nand U15200 (N_15200,N_13734,N_13892);
and U15201 (N_15201,N_12545,N_13505);
nor U15202 (N_15202,N_13241,N_13032);
nand U15203 (N_15203,N_12490,N_12332);
and U15204 (N_15204,N_13600,N_12172);
nor U15205 (N_15205,N_13207,N_12114);
or U15206 (N_15206,N_13425,N_12228);
or U15207 (N_15207,N_13833,N_13736);
nand U15208 (N_15208,N_13156,N_12392);
nor U15209 (N_15209,N_13143,N_12961);
or U15210 (N_15210,N_12839,N_13503);
nand U15211 (N_15211,N_12854,N_12949);
and U15212 (N_15212,N_13741,N_13087);
nor U15213 (N_15213,N_12908,N_13412);
nor U15214 (N_15214,N_13402,N_13311);
nor U15215 (N_15215,N_13735,N_12971);
and U15216 (N_15216,N_12896,N_13105);
nor U15217 (N_15217,N_12543,N_13161);
nand U15218 (N_15218,N_12732,N_12007);
or U15219 (N_15219,N_13842,N_13700);
or U15220 (N_15220,N_13280,N_12387);
or U15221 (N_15221,N_12029,N_12075);
nor U15222 (N_15222,N_12790,N_13418);
or U15223 (N_15223,N_12102,N_12754);
or U15224 (N_15224,N_12890,N_13500);
or U15225 (N_15225,N_12611,N_13283);
and U15226 (N_15226,N_13249,N_13569);
and U15227 (N_15227,N_12131,N_13079);
xor U15228 (N_15228,N_12457,N_13354);
or U15229 (N_15229,N_12146,N_12891);
nand U15230 (N_15230,N_13592,N_12063);
and U15231 (N_15231,N_12474,N_12769);
nand U15232 (N_15232,N_12399,N_13756);
nor U15233 (N_15233,N_12035,N_12604);
nand U15234 (N_15234,N_13448,N_12766);
nand U15235 (N_15235,N_12257,N_13884);
xnor U15236 (N_15236,N_13953,N_12645);
nand U15237 (N_15237,N_13734,N_12449);
nand U15238 (N_15238,N_12412,N_12070);
nor U15239 (N_15239,N_13008,N_13476);
nand U15240 (N_15240,N_13591,N_12874);
or U15241 (N_15241,N_12629,N_13697);
nand U15242 (N_15242,N_13027,N_13872);
nor U15243 (N_15243,N_12888,N_13240);
or U15244 (N_15244,N_12267,N_12148);
and U15245 (N_15245,N_12608,N_12007);
xor U15246 (N_15246,N_13704,N_13327);
nor U15247 (N_15247,N_13147,N_12060);
and U15248 (N_15248,N_13510,N_12316);
or U15249 (N_15249,N_12456,N_13908);
and U15250 (N_15250,N_13670,N_12910);
and U15251 (N_15251,N_12916,N_13737);
xor U15252 (N_15252,N_12135,N_13217);
or U15253 (N_15253,N_12589,N_13918);
nand U15254 (N_15254,N_13818,N_13425);
or U15255 (N_15255,N_12517,N_12119);
and U15256 (N_15256,N_13036,N_13527);
xnor U15257 (N_15257,N_12716,N_13089);
and U15258 (N_15258,N_13495,N_13686);
nand U15259 (N_15259,N_13444,N_12188);
or U15260 (N_15260,N_12101,N_13575);
or U15261 (N_15261,N_12909,N_13844);
and U15262 (N_15262,N_13983,N_13579);
xor U15263 (N_15263,N_13742,N_12971);
and U15264 (N_15264,N_13145,N_12453);
nand U15265 (N_15265,N_12794,N_13670);
nor U15266 (N_15266,N_13843,N_13535);
nor U15267 (N_15267,N_12475,N_12238);
nor U15268 (N_15268,N_13151,N_13669);
nand U15269 (N_15269,N_12680,N_12923);
and U15270 (N_15270,N_13403,N_13218);
nand U15271 (N_15271,N_13933,N_12361);
or U15272 (N_15272,N_12639,N_13665);
or U15273 (N_15273,N_12285,N_13531);
xor U15274 (N_15274,N_12335,N_12206);
nand U15275 (N_15275,N_12586,N_12021);
or U15276 (N_15276,N_13582,N_12708);
or U15277 (N_15277,N_12314,N_13495);
nand U15278 (N_15278,N_12675,N_12509);
nor U15279 (N_15279,N_12683,N_13329);
and U15280 (N_15280,N_13053,N_12111);
and U15281 (N_15281,N_12479,N_13361);
and U15282 (N_15282,N_12045,N_12563);
nor U15283 (N_15283,N_13238,N_12934);
nand U15284 (N_15284,N_12846,N_12814);
nor U15285 (N_15285,N_12097,N_13572);
nand U15286 (N_15286,N_13296,N_12718);
nand U15287 (N_15287,N_12716,N_13925);
nor U15288 (N_15288,N_13130,N_13310);
nor U15289 (N_15289,N_12462,N_12401);
nand U15290 (N_15290,N_12610,N_13634);
xor U15291 (N_15291,N_12467,N_12511);
nor U15292 (N_15292,N_13470,N_13025);
and U15293 (N_15293,N_13813,N_12333);
nor U15294 (N_15294,N_13956,N_13990);
nand U15295 (N_15295,N_12806,N_13355);
or U15296 (N_15296,N_12456,N_13381);
nor U15297 (N_15297,N_12608,N_13379);
nor U15298 (N_15298,N_12128,N_12293);
nand U15299 (N_15299,N_13741,N_12878);
and U15300 (N_15300,N_13150,N_12674);
or U15301 (N_15301,N_13988,N_13993);
or U15302 (N_15302,N_12911,N_12676);
xnor U15303 (N_15303,N_13673,N_12672);
and U15304 (N_15304,N_13238,N_13352);
or U15305 (N_15305,N_13333,N_12400);
and U15306 (N_15306,N_13491,N_12848);
nor U15307 (N_15307,N_13638,N_13239);
nand U15308 (N_15308,N_13121,N_13776);
and U15309 (N_15309,N_13491,N_12605);
xor U15310 (N_15310,N_13189,N_13907);
and U15311 (N_15311,N_13977,N_12678);
nor U15312 (N_15312,N_13730,N_12763);
or U15313 (N_15313,N_12648,N_12105);
and U15314 (N_15314,N_13105,N_12599);
or U15315 (N_15315,N_13587,N_12181);
or U15316 (N_15316,N_13364,N_12836);
nand U15317 (N_15317,N_13542,N_12674);
xor U15318 (N_15318,N_12887,N_12172);
and U15319 (N_15319,N_13369,N_12816);
nor U15320 (N_15320,N_13066,N_13284);
or U15321 (N_15321,N_12983,N_13189);
and U15322 (N_15322,N_12414,N_13633);
nand U15323 (N_15323,N_12034,N_12357);
xor U15324 (N_15324,N_12281,N_13821);
nand U15325 (N_15325,N_12430,N_12348);
or U15326 (N_15326,N_12022,N_12806);
nor U15327 (N_15327,N_12632,N_13098);
nor U15328 (N_15328,N_12462,N_12915);
nand U15329 (N_15329,N_13297,N_12713);
nor U15330 (N_15330,N_13470,N_12117);
or U15331 (N_15331,N_13605,N_13483);
nand U15332 (N_15332,N_12536,N_13592);
xnor U15333 (N_15333,N_13112,N_12230);
or U15334 (N_15334,N_13159,N_13077);
and U15335 (N_15335,N_13488,N_13953);
or U15336 (N_15336,N_13927,N_12697);
or U15337 (N_15337,N_12405,N_13895);
or U15338 (N_15338,N_13550,N_13692);
and U15339 (N_15339,N_12151,N_12866);
or U15340 (N_15340,N_13832,N_12531);
or U15341 (N_15341,N_12401,N_12614);
nand U15342 (N_15342,N_12671,N_12634);
nor U15343 (N_15343,N_13615,N_13205);
xor U15344 (N_15344,N_13256,N_13141);
nand U15345 (N_15345,N_13297,N_12363);
and U15346 (N_15346,N_12232,N_12489);
xor U15347 (N_15347,N_12400,N_12705);
nand U15348 (N_15348,N_12988,N_13109);
nand U15349 (N_15349,N_13947,N_13466);
or U15350 (N_15350,N_12140,N_13527);
xnor U15351 (N_15351,N_13981,N_12579);
or U15352 (N_15352,N_12837,N_13446);
nand U15353 (N_15353,N_13574,N_12199);
and U15354 (N_15354,N_12197,N_13239);
and U15355 (N_15355,N_13531,N_12682);
or U15356 (N_15356,N_13642,N_13952);
nand U15357 (N_15357,N_13981,N_13477);
nand U15358 (N_15358,N_13512,N_12593);
nand U15359 (N_15359,N_13955,N_12130);
nand U15360 (N_15360,N_12834,N_12658);
nor U15361 (N_15361,N_12008,N_12662);
nor U15362 (N_15362,N_12761,N_13366);
or U15363 (N_15363,N_12992,N_13794);
xor U15364 (N_15364,N_12677,N_12146);
and U15365 (N_15365,N_12677,N_12283);
nor U15366 (N_15366,N_12728,N_12048);
and U15367 (N_15367,N_13876,N_13321);
nor U15368 (N_15368,N_13927,N_12058);
and U15369 (N_15369,N_13593,N_12442);
or U15370 (N_15370,N_13626,N_12382);
nor U15371 (N_15371,N_12610,N_13056);
and U15372 (N_15372,N_12555,N_13719);
or U15373 (N_15373,N_13538,N_12836);
or U15374 (N_15374,N_12111,N_12687);
or U15375 (N_15375,N_12518,N_12845);
nand U15376 (N_15376,N_12122,N_12533);
or U15377 (N_15377,N_12260,N_12569);
nor U15378 (N_15378,N_12186,N_13158);
or U15379 (N_15379,N_13021,N_12974);
and U15380 (N_15380,N_13708,N_13200);
or U15381 (N_15381,N_13083,N_13477);
or U15382 (N_15382,N_12732,N_12806);
xnor U15383 (N_15383,N_13127,N_13333);
and U15384 (N_15384,N_13674,N_12431);
and U15385 (N_15385,N_13523,N_13292);
nor U15386 (N_15386,N_12542,N_13795);
nor U15387 (N_15387,N_13629,N_13986);
nor U15388 (N_15388,N_13710,N_12295);
nor U15389 (N_15389,N_13505,N_12832);
nor U15390 (N_15390,N_12522,N_12159);
and U15391 (N_15391,N_12353,N_13250);
nand U15392 (N_15392,N_13500,N_12156);
or U15393 (N_15393,N_13485,N_13969);
and U15394 (N_15394,N_12496,N_13075);
or U15395 (N_15395,N_13425,N_12974);
nand U15396 (N_15396,N_12895,N_12737);
nor U15397 (N_15397,N_12059,N_13405);
nor U15398 (N_15398,N_12108,N_13247);
xnor U15399 (N_15399,N_12607,N_12762);
and U15400 (N_15400,N_12660,N_13732);
nand U15401 (N_15401,N_12545,N_13495);
nand U15402 (N_15402,N_12804,N_12725);
and U15403 (N_15403,N_12419,N_12498);
nor U15404 (N_15404,N_13412,N_12938);
nand U15405 (N_15405,N_13841,N_13579);
nand U15406 (N_15406,N_12024,N_13552);
xnor U15407 (N_15407,N_12630,N_12461);
nor U15408 (N_15408,N_13657,N_13035);
and U15409 (N_15409,N_13189,N_12708);
nor U15410 (N_15410,N_13477,N_13294);
nor U15411 (N_15411,N_13167,N_12084);
xor U15412 (N_15412,N_12246,N_13713);
and U15413 (N_15413,N_13536,N_12998);
nand U15414 (N_15414,N_12002,N_12990);
nand U15415 (N_15415,N_12075,N_13377);
nand U15416 (N_15416,N_13430,N_12564);
or U15417 (N_15417,N_12028,N_13501);
nor U15418 (N_15418,N_12571,N_13835);
nor U15419 (N_15419,N_12377,N_12485);
and U15420 (N_15420,N_13020,N_12851);
nor U15421 (N_15421,N_13213,N_13300);
nor U15422 (N_15422,N_12982,N_13128);
and U15423 (N_15423,N_13488,N_13057);
or U15424 (N_15424,N_13732,N_13051);
or U15425 (N_15425,N_13702,N_13309);
nand U15426 (N_15426,N_12867,N_12651);
and U15427 (N_15427,N_12628,N_12223);
and U15428 (N_15428,N_12428,N_12006);
or U15429 (N_15429,N_13223,N_12856);
or U15430 (N_15430,N_12281,N_12469);
and U15431 (N_15431,N_12531,N_12902);
and U15432 (N_15432,N_12414,N_13647);
and U15433 (N_15433,N_12366,N_13869);
nor U15434 (N_15434,N_12184,N_12054);
xnor U15435 (N_15435,N_13649,N_12163);
nor U15436 (N_15436,N_13424,N_12861);
nor U15437 (N_15437,N_12412,N_12788);
and U15438 (N_15438,N_12016,N_12838);
nand U15439 (N_15439,N_12242,N_12603);
or U15440 (N_15440,N_12264,N_13130);
xnor U15441 (N_15441,N_13155,N_13834);
nand U15442 (N_15442,N_13024,N_13118);
and U15443 (N_15443,N_12130,N_13474);
and U15444 (N_15444,N_12238,N_12611);
or U15445 (N_15445,N_13759,N_12704);
xnor U15446 (N_15446,N_12807,N_12486);
and U15447 (N_15447,N_12810,N_12042);
or U15448 (N_15448,N_13451,N_13711);
nand U15449 (N_15449,N_12982,N_13635);
or U15450 (N_15450,N_12379,N_12323);
nand U15451 (N_15451,N_12179,N_12219);
or U15452 (N_15452,N_13876,N_12667);
nor U15453 (N_15453,N_13213,N_13585);
nor U15454 (N_15454,N_12442,N_12494);
nor U15455 (N_15455,N_12930,N_13572);
nand U15456 (N_15456,N_12332,N_12872);
and U15457 (N_15457,N_12931,N_12881);
nand U15458 (N_15458,N_12239,N_12215);
nor U15459 (N_15459,N_13665,N_13982);
nor U15460 (N_15460,N_12736,N_12517);
or U15461 (N_15461,N_13940,N_13088);
nor U15462 (N_15462,N_13289,N_13513);
nand U15463 (N_15463,N_13340,N_12619);
or U15464 (N_15464,N_12776,N_13141);
nor U15465 (N_15465,N_12925,N_12995);
nor U15466 (N_15466,N_12154,N_13054);
and U15467 (N_15467,N_12730,N_13339);
nand U15468 (N_15468,N_13260,N_12360);
or U15469 (N_15469,N_13993,N_12346);
and U15470 (N_15470,N_12017,N_12106);
and U15471 (N_15471,N_13925,N_13594);
or U15472 (N_15472,N_12491,N_13595);
xor U15473 (N_15473,N_12998,N_12945);
and U15474 (N_15474,N_13982,N_12126);
nand U15475 (N_15475,N_13545,N_13080);
nand U15476 (N_15476,N_13983,N_13573);
nor U15477 (N_15477,N_13695,N_12725);
or U15478 (N_15478,N_13287,N_13973);
and U15479 (N_15479,N_12314,N_13482);
and U15480 (N_15480,N_13771,N_12479);
nor U15481 (N_15481,N_12791,N_13093);
nor U15482 (N_15482,N_12903,N_13791);
or U15483 (N_15483,N_13828,N_12083);
and U15484 (N_15484,N_12451,N_13295);
xor U15485 (N_15485,N_12599,N_13083);
or U15486 (N_15486,N_12814,N_13636);
nor U15487 (N_15487,N_12270,N_12062);
nor U15488 (N_15488,N_13526,N_13199);
or U15489 (N_15489,N_12079,N_12796);
or U15490 (N_15490,N_13269,N_13575);
nor U15491 (N_15491,N_12451,N_12418);
and U15492 (N_15492,N_13827,N_12530);
nand U15493 (N_15493,N_13134,N_12064);
nand U15494 (N_15494,N_13979,N_13939);
nor U15495 (N_15495,N_13029,N_12284);
or U15496 (N_15496,N_12730,N_12920);
or U15497 (N_15497,N_12216,N_12289);
nand U15498 (N_15498,N_12925,N_12960);
or U15499 (N_15499,N_12870,N_12880);
and U15500 (N_15500,N_13137,N_13957);
nand U15501 (N_15501,N_12066,N_12889);
nor U15502 (N_15502,N_13369,N_13367);
or U15503 (N_15503,N_12180,N_13959);
or U15504 (N_15504,N_12264,N_13686);
xor U15505 (N_15505,N_13209,N_12791);
xnor U15506 (N_15506,N_13762,N_12467);
nor U15507 (N_15507,N_12279,N_13818);
xor U15508 (N_15508,N_13991,N_13770);
nor U15509 (N_15509,N_13877,N_12266);
or U15510 (N_15510,N_12548,N_13259);
or U15511 (N_15511,N_13658,N_13067);
and U15512 (N_15512,N_13158,N_13397);
and U15513 (N_15513,N_13503,N_12973);
nor U15514 (N_15514,N_13231,N_12826);
xnor U15515 (N_15515,N_13868,N_13555);
nor U15516 (N_15516,N_13100,N_13005);
and U15517 (N_15517,N_12112,N_13954);
and U15518 (N_15518,N_13541,N_12460);
and U15519 (N_15519,N_13325,N_12862);
nor U15520 (N_15520,N_12901,N_12509);
nand U15521 (N_15521,N_12740,N_13571);
nand U15522 (N_15522,N_12301,N_13318);
nor U15523 (N_15523,N_12195,N_12819);
xor U15524 (N_15524,N_13678,N_13066);
or U15525 (N_15525,N_13065,N_12091);
and U15526 (N_15526,N_12503,N_12939);
nand U15527 (N_15527,N_12516,N_13513);
nand U15528 (N_15528,N_12493,N_13407);
nor U15529 (N_15529,N_13281,N_13809);
nand U15530 (N_15530,N_12517,N_13108);
nor U15531 (N_15531,N_12842,N_13731);
nand U15532 (N_15532,N_13016,N_13702);
and U15533 (N_15533,N_13312,N_12757);
nand U15534 (N_15534,N_13012,N_12658);
or U15535 (N_15535,N_13800,N_12628);
or U15536 (N_15536,N_12653,N_13703);
nor U15537 (N_15537,N_13939,N_13728);
nand U15538 (N_15538,N_12313,N_12784);
nand U15539 (N_15539,N_12624,N_12406);
and U15540 (N_15540,N_13971,N_12987);
or U15541 (N_15541,N_13839,N_12741);
or U15542 (N_15542,N_12688,N_13715);
or U15543 (N_15543,N_12279,N_13876);
and U15544 (N_15544,N_13795,N_12744);
and U15545 (N_15545,N_13220,N_12085);
nand U15546 (N_15546,N_12184,N_13297);
and U15547 (N_15547,N_12711,N_12736);
and U15548 (N_15548,N_12389,N_12963);
or U15549 (N_15549,N_12594,N_12101);
or U15550 (N_15550,N_13804,N_12218);
nand U15551 (N_15551,N_13537,N_13511);
and U15552 (N_15552,N_12065,N_12005);
xnor U15553 (N_15553,N_13621,N_13450);
and U15554 (N_15554,N_12035,N_13396);
or U15555 (N_15555,N_13967,N_12302);
nor U15556 (N_15556,N_13415,N_13438);
nor U15557 (N_15557,N_12458,N_13969);
nor U15558 (N_15558,N_12811,N_12091);
or U15559 (N_15559,N_13814,N_12025);
xnor U15560 (N_15560,N_12269,N_13076);
nor U15561 (N_15561,N_13376,N_12821);
or U15562 (N_15562,N_13660,N_13115);
or U15563 (N_15563,N_12170,N_12539);
and U15564 (N_15564,N_12375,N_13623);
nor U15565 (N_15565,N_13359,N_13295);
or U15566 (N_15566,N_13980,N_12811);
nand U15567 (N_15567,N_13123,N_12760);
and U15568 (N_15568,N_13318,N_13537);
and U15569 (N_15569,N_12630,N_13369);
nor U15570 (N_15570,N_12858,N_13329);
xor U15571 (N_15571,N_12864,N_13325);
and U15572 (N_15572,N_12247,N_13089);
or U15573 (N_15573,N_13318,N_12628);
and U15574 (N_15574,N_13544,N_12869);
nand U15575 (N_15575,N_13487,N_13880);
nor U15576 (N_15576,N_13964,N_13643);
or U15577 (N_15577,N_13499,N_13245);
nor U15578 (N_15578,N_12639,N_13007);
nand U15579 (N_15579,N_12582,N_13788);
nand U15580 (N_15580,N_12158,N_12206);
nand U15581 (N_15581,N_13731,N_12197);
nor U15582 (N_15582,N_12739,N_13179);
nand U15583 (N_15583,N_13595,N_12247);
nor U15584 (N_15584,N_12334,N_12469);
or U15585 (N_15585,N_13723,N_13358);
nand U15586 (N_15586,N_13564,N_13661);
and U15587 (N_15587,N_12018,N_13562);
or U15588 (N_15588,N_13701,N_13952);
nand U15589 (N_15589,N_12401,N_13648);
xor U15590 (N_15590,N_12800,N_13080);
xor U15591 (N_15591,N_12467,N_12685);
nand U15592 (N_15592,N_12615,N_12156);
nor U15593 (N_15593,N_12876,N_13646);
and U15594 (N_15594,N_12674,N_12832);
nand U15595 (N_15595,N_13809,N_13986);
nand U15596 (N_15596,N_13990,N_13471);
nand U15597 (N_15597,N_12990,N_12198);
xor U15598 (N_15598,N_13105,N_12461);
or U15599 (N_15599,N_12853,N_12450);
xnor U15600 (N_15600,N_12693,N_12419);
nand U15601 (N_15601,N_13992,N_13710);
nand U15602 (N_15602,N_13015,N_13115);
nand U15603 (N_15603,N_13829,N_12017);
nand U15604 (N_15604,N_12401,N_13917);
or U15605 (N_15605,N_12018,N_12100);
or U15606 (N_15606,N_13130,N_13799);
nor U15607 (N_15607,N_12233,N_13425);
nand U15608 (N_15608,N_12280,N_13345);
nor U15609 (N_15609,N_13155,N_13408);
or U15610 (N_15610,N_12949,N_12557);
xnor U15611 (N_15611,N_13168,N_12355);
nand U15612 (N_15612,N_12710,N_13189);
nand U15613 (N_15613,N_12139,N_12633);
nand U15614 (N_15614,N_13724,N_12231);
nand U15615 (N_15615,N_13318,N_12928);
nor U15616 (N_15616,N_13181,N_12861);
nor U15617 (N_15617,N_12283,N_13316);
or U15618 (N_15618,N_12432,N_13685);
nor U15619 (N_15619,N_13249,N_13099);
and U15620 (N_15620,N_13058,N_12708);
or U15621 (N_15621,N_13365,N_13721);
nand U15622 (N_15622,N_13070,N_13912);
or U15623 (N_15623,N_12587,N_12506);
or U15624 (N_15624,N_12215,N_13204);
nand U15625 (N_15625,N_13856,N_12065);
and U15626 (N_15626,N_13824,N_12091);
nand U15627 (N_15627,N_12588,N_13960);
and U15628 (N_15628,N_13849,N_12761);
and U15629 (N_15629,N_13014,N_13507);
and U15630 (N_15630,N_13937,N_12637);
nor U15631 (N_15631,N_13124,N_13659);
nand U15632 (N_15632,N_12633,N_12556);
or U15633 (N_15633,N_13724,N_13995);
nor U15634 (N_15634,N_12044,N_13647);
or U15635 (N_15635,N_13490,N_12325);
nand U15636 (N_15636,N_13659,N_13886);
and U15637 (N_15637,N_12274,N_13088);
and U15638 (N_15638,N_12485,N_13804);
nor U15639 (N_15639,N_12096,N_12480);
and U15640 (N_15640,N_13736,N_13622);
nand U15641 (N_15641,N_13246,N_13755);
nor U15642 (N_15642,N_12706,N_13334);
nor U15643 (N_15643,N_12892,N_13331);
and U15644 (N_15644,N_13535,N_13280);
nor U15645 (N_15645,N_12425,N_12377);
nand U15646 (N_15646,N_12597,N_13667);
and U15647 (N_15647,N_13901,N_12161);
nand U15648 (N_15648,N_12587,N_12395);
and U15649 (N_15649,N_13711,N_12396);
nand U15650 (N_15650,N_12038,N_13976);
and U15651 (N_15651,N_12993,N_13725);
nand U15652 (N_15652,N_12146,N_13632);
nand U15653 (N_15653,N_12975,N_12452);
or U15654 (N_15654,N_12173,N_13571);
or U15655 (N_15655,N_12506,N_12000);
or U15656 (N_15656,N_13944,N_12081);
or U15657 (N_15657,N_12209,N_12225);
and U15658 (N_15658,N_12844,N_13289);
or U15659 (N_15659,N_13546,N_12485);
nor U15660 (N_15660,N_13783,N_12080);
nand U15661 (N_15661,N_12522,N_12421);
or U15662 (N_15662,N_13097,N_13273);
or U15663 (N_15663,N_13853,N_12165);
nor U15664 (N_15664,N_12932,N_13099);
xor U15665 (N_15665,N_13952,N_12777);
or U15666 (N_15666,N_13604,N_13112);
or U15667 (N_15667,N_13447,N_13811);
and U15668 (N_15668,N_12473,N_13534);
nor U15669 (N_15669,N_13880,N_12803);
nor U15670 (N_15670,N_12044,N_13618);
or U15671 (N_15671,N_12996,N_12623);
nand U15672 (N_15672,N_12371,N_12896);
nand U15673 (N_15673,N_13886,N_13290);
and U15674 (N_15674,N_13990,N_12082);
and U15675 (N_15675,N_12055,N_12570);
nand U15676 (N_15676,N_12855,N_13462);
or U15677 (N_15677,N_13265,N_13631);
nor U15678 (N_15678,N_12770,N_13440);
or U15679 (N_15679,N_12729,N_12720);
nor U15680 (N_15680,N_12558,N_13510);
and U15681 (N_15681,N_13140,N_13620);
and U15682 (N_15682,N_13121,N_12605);
xor U15683 (N_15683,N_12178,N_13486);
nor U15684 (N_15684,N_12115,N_12727);
nor U15685 (N_15685,N_12970,N_13385);
nor U15686 (N_15686,N_12113,N_12211);
nor U15687 (N_15687,N_12063,N_13759);
and U15688 (N_15688,N_13468,N_12725);
and U15689 (N_15689,N_13132,N_12834);
nand U15690 (N_15690,N_13118,N_13092);
or U15691 (N_15691,N_13694,N_13152);
nor U15692 (N_15692,N_13161,N_12904);
xnor U15693 (N_15693,N_13480,N_13972);
xor U15694 (N_15694,N_12210,N_13522);
nor U15695 (N_15695,N_12809,N_12462);
and U15696 (N_15696,N_13432,N_12698);
nand U15697 (N_15697,N_12826,N_12048);
or U15698 (N_15698,N_12969,N_12950);
and U15699 (N_15699,N_13729,N_13615);
or U15700 (N_15700,N_13768,N_13809);
xor U15701 (N_15701,N_12745,N_13666);
nor U15702 (N_15702,N_13532,N_13518);
or U15703 (N_15703,N_12130,N_12882);
and U15704 (N_15704,N_12650,N_13284);
nor U15705 (N_15705,N_13652,N_12033);
and U15706 (N_15706,N_13187,N_12602);
or U15707 (N_15707,N_12378,N_12132);
nand U15708 (N_15708,N_12454,N_12615);
nand U15709 (N_15709,N_12108,N_13716);
and U15710 (N_15710,N_12914,N_13760);
nor U15711 (N_15711,N_13371,N_13853);
or U15712 (N_15712,N_12524,N_13045);
and U15713 (N_15713,N_13076,N_13002);
or U15714 (N_15714,N_13707,N_12382);
nor U15715 (N_15715,N_12926,N_13031);
xnor U15716 (N_15716,N_13207,N_13047);
nand U15717 (N_15717,N_13285,N_13695);
or U15718 (N_15718,N_13792,N_12004);
nand U15719 (N_15719,N_13080,N_13048);
and U15720 (N_15720,N_12910,N_13744);
or U15721 (N_15721,N_12185,N_12626);
nand U15722 (N_15722,N_12011,N_13051);
or U15723 (N_15723,N_12166,N_12440);
nor U15724 (N_15724,N_12122,N_12151);
and U15725 (N_15725,N_13083,N_13616);
or U15726 (N_15726,N_12333,N_12556);
and U15727 (N_15727,N_13015,N_13996);
nor U15728 (N_15728,N_13007,N_12054);
nand U15729 (N_15729,N_12219,N_13592);
and U15730 (N_15730,N_13745,N_12099);
or U15731 (N_15731,N_13053,N_13157);
nand U15732 (N_15732,N_12173,N_12702);
and U15733 (N_15733,N_13418,N_12984);
nand U15734 (N_15734,N_12991,N_13042);
nand U15735 (N_15735,N_13787,N_12644);
or U15736 (N_15736,N_12427,N_13435);
xnor U15737 (N_15737,N_13036,N_12214);
nor U15738 (N_15738,N_13992,N_12322);
and U15739 (N_15739,N_13037,N_13254);
nand U15740 (N_15740,N_12927,N_13618);
nor U15741 (N_15741,N_12033,N_13455);
and U15742 (N_15742,N_13805,N_13979);
xnor U15743 (N_15743,N_12659,N_12742);
nand U15744 (N_15744,N_12448,N_13349);
and U15745 (N_15745,N_12262,N_12759);
and U15746 (N_15746,N_13143,N_13381);
nor U15747 (N_15747,N_12363,N_12034);
nor U15748 (N_15748,N_13943,N_13054);
nor U15749 (N_15749,N_12352,N_13130);
nand U15750 (N_15750,N_13903,N_13669);
nand U15751 (N_15751,N_12189,N_12290);
or U15752 (N_15752,N_12576,N_13936);
nor U15753 (N_15753,N_13645,N_13837);
nor U15754 (N_15754,N_13591,N_13237);
or U15755 (N_15755,N_12353,N_13128);
or U15756 (N_15756,N_13324,N_12772);
and U15757 (N_15757,N_12293,N_13400);
nor U15758 (N_15758,N_13980,N_13744);
nand U15759 (N_15759,N_12134,N_12028);
xor U15760 (N_15760,N_12503,N_13403);
nor U15761 (N_15761,N_12556,N_13697);
and U15762 (N_15762,N_12906,N_13274);
nand U15763 (N_15763,N_13247,N_13364);
nand U15764 (N_15764,N_13049,N_12027);
nor U15765 (N_15765,N_13613,N_12640);
or U15766 (N_15766,N_13776,N_12467);
nand U15767 (N_15767,N_12196,N_12374);
nor U15768 (N_15768,N_13557,N_12125);
nor U15769 (N_15769,N_13832,N_13919);
nor U15770 (N_15770,N_13637,N_12101);
or U15771 (N_15771,N_13534,N_12442);
xor U15772 (N_15772,N_13226,N_12762);
nor U15773 (N_15773,N_12436,N_13225);
or U15774 (N_15774,N_12537,N_13764);
and U15775 (N_15775,N_13711,N_12193);
nand U15776 (N_15776,N_12986,N_12341);
xnor U15777 (N_15777,N_12184,N_12250);
nand U15778 (N_15778,N_13514,N_13029);
or U15779 (N_15779,N_12205,N_12913);
nor U15780 (N_15780,N_12902,N_13282);
and U15781 (N_15781,N_12327,N_12457);
nand U15782 (N_15782,N_13395,N_12965);
and U15783 (N_15783,N_13686,N_12968);
nor U15784 (N_15784,N_12336,N_12041);
xnor U15785 (N_15785,N_13269,N_13468);
and U15786 (N_15786,N_13672,N_13645);
nor U15787 (N_15787,N_12966,N_12131);
or U15788 (N_15788,N_13128,N_12784);
nand U15789 (N_15789,N_12523,N_12875);
nor U15790 (N_15790,N_12946,N_12444);
and U15791 (N_15791,N_13906,N_13844);
and U15792 (N_15792,N_12142,N_12552);
or U15793 (N_15793,N_12305,N_12351);
nand U15794 (N_15794,N_13213,N_12869);
xnor U15795 (N_15795,N_13933,N_12769);
nand U15796 (N_15796,N_12928,N_12474);
xnor U15797 (N_15797,N_12075,N_12495);
nor U15798 (N_15798,N_13456,N_12275);
nor U15799 (N_15799,N_13115,N_12519);
or U15800 (N_15800,N_12878,N_12715);
or U15801 (N_15801,N_13912,N_13282);
nand U15802 (N_15802,N_13725,N_13026);
or U15803 (N_15803,N_13258,N_12083);
nor U15804 (N_15804,N_12489,N_13978);
nand U15805 (N_15805,N_12936,N_12738);
nor U15806 (N_15806,N_13406,N_13361);
or U15807 (N_15807,N_13006,N_13078);
or U15808 (N_15808,N_13357,N_12949);
nor U15809 (N_15809,N_12628,N_12447);
nand U15810 (N_15810,N_13134,N_12721);
and U15811 (N_15811,N_13336,N_13337);
nor U15812 (N_15812,N_13691,N_13171);
nor U15813 (N_15813,N_12989,N_12813);
nor U15814 (N_15814,N_13273,N_13619);
and U15815 (N_15815,N_12737,N_12696);
and U15816 (N_15816,N_12870,N_13111);
and U15817 (N_15817,N_12215,N_13829);
and U15818 (N_15818,N_12368,N_13405);
and U15819 (N_15819,N_13588,N_13271);
nor U15820 (N_15820,N_12477,N_13354);
and U15821 (N_15821,N_12542,N_13364);
nor U15822 (N_15822,N_12022,N_12740);
xnor U15823 (N_15823,N_12695,N_13239);
or U15824 (N_15824,N_12015,N_13220);
or U15825 (N_15825,N_12418,N_12540);
and U15826 (N_15826,N_12548,N_12814);
nand U15827 (N_15827,N_13678,N_13441);
nor U15828 (N_15828,N_13852,N_12973);
xor U15829 (N_15829,N_12749,N_13478);
nand U15830 (N_15830,N_13247,N_13722);
and U15831 (N_15831,N_13211,N_13623);
nor U15832 (N_15832,N_12374,N_12008);
nor U15833 (N_15833,N_12787,N_12193);
or U15834 (N_15834,N_13891,N_12530);
and U15835 (N_15835,N_12174,N_13520);
or U15836 (N_15836,N_13797,N_12957);
and U15837 (N_15837,N_13178,N_13755);
xor U15838 (N_15838,N_13610,N_13073);
and U15839 (N_15839,N_12530,N_13539);
xnor U15840 (N_15840,N_12452,N_13801);
or U15841 (N_15841,N_12618,N_12487);
and U15842 (N_15842,N_13598,N_12332);
and U15843 (N_15843,N_12040,N_12801);
nor U15844 (N_15844,N_13826,N_12664);
nand U15845 (N_15845,N_13048,N_12149);
or U15846 (N_15846,N_13202,N_12655);
nand U15847 (N_15847,N_13964,N_13591);
and U15848 (N_15848,N_12843,N_12570);
and U15849 (N_15849,N_12307,N_13845);
and U15850 (N_15850,N_13829,N_13061);
nand U15851 (N_15851,N_12014,N_13593);
or U15852 (N_15852,N_13974,N_13344);
xnor U15853 (N_15853,N_12979,N_12072);
and U15854 (N_15854,N_13453,N_12051);
and U15855 (N_15855,N_12098,N_13179);
and U15856 (N_15856,N_12728,N_12023);
nor U15857 (N_15857,N_13974,N_12939);
or U15858 (N_15858,N_13443,N_13854);
nor U15859 (N_15859,N_13272,N_12790);
nand U15860 (N_15860,N_12535,N_12904);
nor U15861 (N_15861,N_12807,N_12180);
nand U15862 (N_15862,N_13774,N_12947);
nor U15863 (N_15863,N_13707,N_13678);
nand U15864 (N_15864,N_12668,N_12482);
and U15865 (N_15865,N_12358,N_12285);
nor U15866 (N_15866,N_12996,N_13486);
or U15867 (N_15867,N_12000,N_12972);
nor U15868 (N_15868,N_13012,N_12872);
nor U15869 (N_15869,N_12048,N_13954);
or U15870 (N_15870,N_13219,N_13652);
nor U15871 (N_15871,N_13130,N_12052);
nor U15872 (N_15872,N_13446,N_12174);
and U15873 (N_15873,N_13724,N_13790);
and U15874 (N_15874,N_13167,N_13283);
or U15875 (N_15875,N_13237,N_13401);
xor U15876 (N_15876,N_13947,N_12869);
nand U15877 (N_15877,N_12263,N_13412);
nand U15878 (N_15878,N_13922,N_12900);
nor U15879 (N_15879,N_13243,N_13768);
xor U15880 (N_15880,N_12538,N_13329);
nor U15881 (N_15881,N_12294,N_12837);
or U15882 (N_15882,N_12672,N_13385);
and U15883 (N_15883,N_12762,N_13132);
and U15884 (N_15884,N_13878,N_13116);
and U15885 (N_15885,N_13559,N_13817);
nand U15886 (N_15886,N_13046,N_13751);
and U15887 (N_15887,N_13849,N_12463);
nor U15888 (N_15888,N_12267,N_13668);
nand U15889 (N_15889,N_13820,N_12138);
nand U15890 (N_15890,N_12200,N_12860);
or U15891 (N_15891,N_12445,N_13552);
xor U15892 (N_15892,N_13497,N_13128);
nor U15893 (N_15893,N_13305,N_12432);
and U15894 (N_15894,N_12296,N_12963);
nand U15895 (N_15895,N_12732,N_13930);
and U15896 (N_15896,N_12157,N_13974);
or U15897 (N_15897,N_13586,N_13819);
nand U15898 (N_15898,N_13624,N_12539);
nand U15899 (N_15899,N_12528,N_12006);
nand U15900 (N_15900,N_12766,N_12397);
nor U15901 (N_15901,N_12768,N_12822);
and U15902 (N_15902,N_13282,N_12860);
nor U15903 (N_15903,N_12207,N_12460);
or U15904 (N_15904,N_12669,N_13131);
nand U15905 (N_15905,N_13784,N_13821);
nor U15906 (N_15906,N_13164,N_12394);
nor U15907 (N_15907,N_13209,N_12268);
xor U15908 (N_15908,N_13164,N_13580);
and U15909 (N_15909,N_13450,N_12761);
xnor U15910 (N_15910,N_13871,N_13045);
and U15911 (N_15911,N_12316,N_12546);
nor U15912 (N_15912,N_12097,N_12795);
nor U15913 (N_15913,N_12659,N_13264);
xnor U15914 (N_15914,N_12510,N_13875);
xnor U15915 (N_15915,N_13143,N_13590);
nand U15916 (N_15916,N_13563,N_13367);
and U15917 (N_15917,N_12822,N_12903);
nor U15918 (N_15918,N_12377,N_13532);
and U15919 (N_15919,N_13063,N_12189);
or U15920 (N_15920,N_12501,N_12026);
or U15921 (N_15921,N_12981,N_13593);
and U15922 (N_15922,N_13839,N_13461);
xor U15923 (N_15923,N_13766,N_12118);
or U15924 (N_15924,N_12291,N_13883);
nor U15925 (N_15925,N_13230,N_13017);
xor U15926 (N_15926,N_12188,N_12618);
nor U15927 (N_15927,N_13245,N_12776);
and U15928 (N_15928,N_12391,N_12091);
nand U15929 (N_15929,N_12729,N_13872);
nor U15930 (N_15930,N_13137,N_13819);
and U15931 (N_15931,N_13124,N_12259);
nand U15932 (N_15932,N_12307,N_13667);
nand U15933 (N_15933,N_12700,N_13295);
and U15934 (N_15934,N_12794,N_12335);
and U15935 (N_15935,N_12230,N_12444);
nor U15936 (N_15936,N_12643,N_12290);
nor U15937 (N_15937,N_12265,N_12960);
and U15938 (N_15938,N_12471,N_13800);
nor U15939 (N_15939,N_12582,N_13322);
nor U15940 (N_15940,N_13129,N_12298);
or U15941 (N_15941,N_12735,N_12560);
nand U15942 (N_15942,N_12450,N_12978);
nor U15943 (N_15943,N_12832,N_12372);
nor U15944 (N_15944,N_13192,N_13416);
or U15945 (N_15945,N_13175,N_13514);
and U15946 (N_15946,N_12043,N_13447);
nand U15947 (N_15947,N_12726,N_13160);
or U15948 (N_15948,N_12580,N_13602);
and U15949 (N_15949,N_12186,N_12509);
nand U15950 (N_15950,N_13731,N_13342);
nand U15951 (N_15951,N_13011,N_12428);
nand U15952 (N_15952,N_12152,N_12271);
nor U15953 (N_15953,N_12364,N_13256);
nand U15954 (N_15954,N_13684,N_12606);
xor U15955 (N_15955,N_12794,N_13891);
nand U15956 (N_15956,N_13271,N_12689);
or U15957 (N_15957,N_12908,N_12638);
or U15958 (N_15958,N_13419,N_12000);
or U15959 (N_15959,N_13250,N_12113);
and U15960 (N_15960,N_12120,N_12867);
xnor U15961 (N_15961,N_12134,N_13630);
nor U15962 (N_15962,N_12958,N_13536);
nand U15963 (N_15963,N_12621,N_13333);
xor U15964 (N_15964,N_12183,N_12932);
or U15965 (N_15965,N_13550,N_12293);
nor U15966 (N_15966,N_12314,N_13585);
or U15967 (N_15967,N_13975,N_13884);
or U15968 (N_15968,N_12326,N_13621);
xor U15969 (N_15969,N_12413,N_12441);
nor U15970 (N_15970,N_12829,N_12401);
and U15971 (N_15971,N_13486,N_13524);
and U15972 (N_15972,N_13749,N_12747);
xor U15973 (N_15973,N_12957,N_13961);
and U15974 (N_15974,N_13885,N_13161);
and U15975 (N_15975,N_13402,N_12521);
or U15976 (N_15976,N_13911,N_12832);
and U15977 (N_15977,N_13277,N_12510);
xor U15978 (N_15978,N_13833,N_13309);
nor U15979 (N_15979,N_13993,N_13707);
xor U15980 (N_15980,N_13911,N_12138);
or U15981 (N_15981,N_12461,N_12211);
nand U15982 (N_15982,N_12622,N_12955);
and U15983 (N_15983,N_13311,N_12368);
nand U15984 (N_15984,N_13185,N_12484);
nand U15985 (N_15985,N_12766,N_12898);
and U15986 (N_15986,N_13324,N_12803);
or U15987 (N_15987,N_13700,N_13621);
and U15988 (N_15988,N_13295,N_13740);
or U15989 (N_15989,N_13944,N_13288);
and U15990 (N_15990,N_13975,N_13979);
or U15991 (N_15991,N_13985,N_13956);
or U15992 (N_15992,N_13497,N_12313);
nor U15993 (N_15993,N_13528,N_13066);
and U15994 (N_15994,N_12318,N_13144);
and U15995 (N_15995,N_12146,N_13142);
and U15996 (N_15996,N_12995,N_12096);
nor U15997 (N_15997,N_13252,N_12509);
xnor U15998 (N_15998,N_12547,N_12864);
or U15999 (N_15999,N_13234,N_12639);
or U16000 (N_16000,N_14322,N_14453);
xnor U16001 (N_16001,N_15658,N_15159);
nor U16002 (N_16002,N_14640,N_15085);
or U16003 (N_16003,N_15964,N_14288);
nor U16004 (N_16004,N_14589,N_14693);
nand U16005 (N_16005,N_14158,N_14708);
nand U16006 (N_16006,N_14414,N_14222);
nor U16007 (N_16007,N_15685,N_15565);
or U16008 (N_16008,N_14686,N_14817);
nand U16009 (N_16009,N_14723,N_15483);
nor U16010 (N_16010,N_15393,N_15370);
xor U16011 (N_16011,N_14378,N_14198);
nand U16012 (N_16012,N_15260,N_15618);
nand U16013 (N_16013,N_15637,N_15388);
or U16014 (N_16014,N_15094,N_15163);
or U16015 (N_16015,N_14568,N_15353);
nand U16016 (N_16016,N_14056,N_14417);
and U16017 (N_16017,N_14086,N_14891);
nor U16018 (N_16018,N_14267,N_14487);
xor U16019 (N_16019,N_15998,N_14060);
xnor U16020 (N_16020,N_14053,N_14984);
nor U16021 (N_16021,N_15671,N_14518);
and U16022 (N_16022,N_14889,N_14540);
or U16023 (N_16023,N_14863,N_14968);
or U16024 (N_16024,N_14124,N_15712);
or U16025 (N_16025,N_14527,N_14070);
nor U16026 (N_16026,N_14625,N_14818);
and U16027 (N_16027,N_14998,N_14459);
nand U16028 (N_16028,N_14659,N_15286);
nand U16029 (N_16029,N_15012,N_15013);
nand U16030 (N_16030,N_15317,N_14499);
or U16031 (N_16031,N_14711,N_14166);
and U16032 (N_16032,N_15421,N_14190);
nor U16033 (N_16033,N_14134,N_15843);
and U16034 (N_16034,N_15446,N_15066);
nand U16035 (N_16035,N_14989,N_15281);
nand U16036 (N_16036,N_15879,N_15303);
nand U16037 (N_16037,N_15238,N_14494);
nor U16038 (N_16038,N_15399,N_14358);
nand U16039 (N_16039,N_14421,N_14474);
nand U16040 (N_16040,N_14546,N_15220);
xnor U16041 (N_16041,N_15874,N_14795);
and U16042 (N_16042,N_15920,N_15691);
nor U16043 (N_16043,N_15102,N_15620);
nor U16044 (N_16044,N_14061,N_14464);
nor U16045 (N_16045,N_14851,N_15128);
xnor U16046 (N_16046,N_14553,N_14885);
nor U16047 (N_16047,N_15268,N_15850);
and U16048 (N_16048,N_14768,N_15975);
and U16049 (N_16049,N_14560,N_15166);
nor U16050 (N_16050,N_14620,N_15600);
and U16051 (N_16051,N_14974,N_14072);
or U16052 (N_16052,N_15398,N_14339);
and U16053 (N_16053,N_15563,N_15132);
nand U16054 (N_16054,N_15262,N_15787);
xor U16055 (N_16055,N_15913,N_15909);
nor U16056 (N_16056,N_14800,N_14558);
nand U16057 (N_16057,N_14763,N_14648);
or U16058 (N_16058,N_15289,N_14202);
nor U16059 (N_16059,N_14477,N_14674);
nor U16060 (N_16060,N_15251,N_15462);
xor U16061 (N_16061,N_15065,N_15616);
or U16062 (N_16062,N_14063,N_14455);
or U16063 (N_16063,N_14710,N_15481);
nand U16064 (N_16064,N_14450,N_14257);
and U16065 (N_16065,N_14367,N_14255);
and U16066 (N_16066,N_14581,N_14532);
nand U16067 (N_16067,N_14750,N_14058);
nor U16068 (N_16068,N_14254,N_14246);
nor U16069 (N_16069,N_15641,N_15117);
and U16070 (N_16070,N_15182,N_15177);
and U16071 (N_16071,N_15753,N_14442);
nand U16072 (N_16072,N_14767,N_15394);
nand U16073 (N_16073,N_15782,N_15922);
nor U16074 (N_16074,N_15836,N_14176);
or U16075 (N_16075,N_14836,N_14935);
nor U16076 (N_16076,N_14735,N_14361);
and U16077 (N_16077,N_15968,N_14893);
xor U16078 (N_16078,N_15125,N_14468);
or U16079 (N_16079,N_14566,N_15130);
and U16080 (N_16080,N_15871,N_14543);
nor U16081 (N_16081,N_15445,N_14724);
nor U16082 (N_16082,N_15041,N_14187);
nand U16083 (N_16083,N_15058,N_15672);
or U16084 (N_16084,N_14276,N_15164);
nor U16085 (N_16085,N_14503,N_14208);
xor U16086 (N_16086,N_15501,N_15716);
and U16087 (N_16087,N_15588,N_15544);
and U16088 (N_16088,N_14268,N_14656);
nand U16089 (N_16089,N_14122,N_14995);
or U16090 (N_16090,N_14856,N_15929);
and U16091 (N_16091,N_15143,N_15208);
nor U16092 (N_16092,N_14688,N_14346);
and U16093 (N_16093,N_15688,N_14316);
or U16094 (N_16094,N_14396,N_14399);
xor U16095 (N_16095,N_15257,N_14441);
and U16096 (N_16096,N_14824,N_14776);
xor U16097 (N_16097,N_14615,N_15005);
nand U16098 (N_16098,N_14846,N_14365);
nor U16099 (N_16099,N_14658,N_15504);
or U16100 (N_16100,N_14229,N_15571);
nand U16101 (N_16101,N_14606,N_14162);
nand U16102 (N_16102,N_14431,N_14928);
and U16103 (N_16103,N_14621,N_15342);
nand U16104 (N_16104,N_14895,N_15387);
nor U16105 (N_16105,N_14880,N_14142);
or U16106 (N_16106,N_14603,N_14547);
or U16107 (N_16107,N_14242,N_14508);
nor U16108 (N_16108,N_15271,N_14234);
xnor U16109 (N_16109,N_14952,N_14900);
nor U16110 (N_16110,N_15466,N_15146);
and U16111 (N_16111,N_15063,N_15852);
nor U16112 (N_16112,N_15966,N_15420);
nand U16113 (N_16113,N_14252,N_15527);
and U16114 (N_16114,N_14381,N_14784);
and U16115 (N_16115,N_14154,N_15924);
nor U16116 (N_16116,N_15232,N_14323);
or U16117 (N_16117,N_15280,N_15030);
nand U16118 (N_16118,N_14164,N_14296);
nand U16119 (N_16119,N_15261,N_15425);
and U16120 (N_16120,N_14579,N_15096);
nand U16121 (N_16121,N_14590,N_15773);
and U16122 (N_16122,N_15193,N_15677);
nor U16123 (N_16123,N_14028,N_14282);
nor U16124 (N_16124,N_15776,N_14835);
or U16125 (N_16125,N_15140,N_15845);
xor U16126 (N_16126,N_15956,N_14596);
or U16127 (N_16127,N_14264,N_15367);
xnor U16128 (N_16128,N_15898,N_15690);
nand U16129 (N_16129,N_15868,N_14614);
nor U16130 (N_16130,N_15026,N_15596);
and U16131 (N_16131,N_14838,N_15572);
or U16132 (N_16132,N_15792,N_14143);
nand U16133 (N_16133,N_14876,N_15722);
and U16134 (N_16134,N_15386,N_14423);
nand U16135 (N_16135,N_15650,N_15171);
or U16136 (N_16136,N_14217,N_15001);
nor U16137 (N_16137,N_14557,N_14864);
xnor U16138 (N_16138,N_15778,N_15983);
nand U16139 (N_16139,N_15918,N_14182);
xnor U16140 (N_16140,N_15475,N_15168);
or U16141 (N_16141,N_15478,N_15930);
and U16142 (N_16142,N_15101,N_15474);
nand U16143 (N_16143,N_15804,N_15380);
nand U16144 (N_16144,N_14313,N_14324);
nand U16145 (N_16145,N_14292,N_14087);
nor U16146 (N_16146,N_14754,N_15512);
or U16147 (N_16147,N_14329,N_15218);
and U16148 (N_16148,N_14703,N_15011);
and U16149 (N_16149,N_14663,N_14704);
xnor U16150 (N_16150,N_14847,N_14673);
and U16151 (N_16151,N_14940,N_15557);
nand U16152 (N_16152,N_15376,N_14751);
or U16153 (N_16153,N_15739,N_14115);
nor U16154 (N_16154,N_15862,N_14443);
and U16155 (N_16155,N_15578,N_15647);
nor U16156 (N_16156,N_14643,N_15599);
xor U16157 (N_16157,N_14395,N_15540);
nand U16158 (N_16158,N_14777,N_14602);
and U16159 (N_16159,N_15795,N_14130);
xor U16160 (N_16160,N_15495,N_15246);
nor U16161 (N_16161,N_14570,N_15138);
xor U16162 (N_16162,N_14571,N_14233);
nor U16163 (N_16163,N_14064,N_14251);
nor U16164 (N_16164,N_14669,N_14588);
nand U16165 (N_16165,N_14761,N_14966);
nand U16166 (N_16166,N_15666,N_14016);
nor U16167 (N_16167,N_15496,N_14528);
or U16168 (N_16168,N_15925,N_14375);
and U16169 (N_16169,N_14787,N_15332);
and U16170 (N_16170,N_14432,N_15884);
or U16171 (N_16171,N_15943,N_15176);
nor U16172 (N_16172,N_15839,N_15683);
nand U16173 (N_16173,N_15746,N_15907);
nand U16174 (N_16174,N_14644,N_15382);
and U16175 (N_16175,N_14728,N_14000);
or U16176 (N_16176,N_15927,N_14120);
and U16177 (N_16177,N_15695,N_15396);
nor U16178 (N_16178,N_14806,N_14752);
or U16179 (N_16179,N_15161,N_15076);
or U16180 (N_16180,N_14738,N_14116);
or U16181 (N_16181,N_14672,N_14213);
or U16182 (N_16182,N_14103,N_14489);
or U16183 (N_16183,N_15053,N_14456);
nand U16184 (N_16184,N_14383,N_15921);
nand U16185 (N_16185,N_15269,N_14266);
nor U16186 (N_16186,N_15427,N_15613);
and U16187 (N_16187,N_14287,N_14556);
and U16188 (N_16188,N_15025,N_15513);
nand U16189 (N_16189,N_14232,N_15562);
nor U16190 (N_16190,N_14597,N_14924);
or U16191 (N_16191,N_15331,N_15097);
and U16192 (N_16192,N_14145,N_14428);
nand U16193 (N_16193,N_14011,N_15978);
nand U16194 (N_16194,N_14567,N_15211);
and U16195 (N_16195,N_15379,N_14224);
nor U16196 (N_16196,N_14912,N_15510);
or U16197 (N_16197,N_15072,N_14054);
nand U16198 (N_16198,N_14194,N_14306);
nand U16199 (N_16199,N_15514,N_15633);
nor U16200 (N_16200,N_14920,N_15437);
nand U16201 (N_16201,N_15108,N_14493);
xor U16202 (N_16202,N_14852,N_14585);
nand U16203 (N_16203,N_15236,N_14963);
nand U16204 (N_16204,N_15465,N_15873);
xnor U16205 (N_16205,N_15299,N_14366);
nand U16206 (N_16206,N_14805,N_14107);
or U16207 (N_16207,N_15865,N_15904);
nor U16208 (N_16208,N_14015,N_14249);
nor U16209 (N_16209,N_14498,N_15917);
nand U16210 (N_16210,N_14867,N_15830);
and U16211 (N_16211,N_14328,N_14958);
nand U16212 (N_16212,N_15070,N_15590);
or U16213 (N_16213,N_14804,N_15890);
nor U16214 (N_16214,N_14985,N_15459);
and U16215 (N_16215,N_15078,N_14156);
nor U16216 (N_16216,N_14630,N_14183);
and U16217 (N_16217,N_14382,N_14564);
nand U16218 (N_16218,N_14170,N_15032);
nor U16219 (N_16219,N_15264,N_14744);
nand U16220 (N_16220,N_15700,N_14020);
or U16221 (N_16221,N_15018,N_15634);
or U16222 (N_16222,N_15003,N_14126);
nor U16223 (N_16223,N_15511,N_15574);
nand U16224 (N_16224,N_14512,N_14247);
or U16225 (N_16225,N_14253,N_15452);
and U16226 (N_16226,N_15363,N_15629);
nor U16227 (N_16227,N_15582,N_14894);
nand U16228 (N_16228,N_14331,N_15556);
or U16229 (N_16229,N_14879,N_15867);
nand U16230 (N_16230,N_15622,N_15110);
and U16231 (N_16231,N_15490,N_15015);
nor U16232 (N_16232,N_14429,N_14745);
xor U16233 (N_16233,N_15704,N_14841);
nand U16234 (N_16234,N_14539,N_14374);
xnor U16235 (N_16235,N_15186,N_15765);
xnor U16236 (N_16236,N_14839,N_14196);
nand U16237 (N_16237,N_14720,N_15508);
and U16238 (N_16238,N_15853,N_15876);
xnor U16239 (N_16239,N_15995,N_14362);
and U16240 (N_16240,N_15114,N_15219);
nor U16241 (N_16241,N_14731,N_15350);
nor U16242 (N_16242,N_15115,N_14529);
nor U16243 (N_16243,N_15384,N_14632);
nor U16244 (N_16244,N_14778,N_15049);
xor U16245 (N_16245,N_15713,N_14189);
nor U16246 (N_16246,N_14332,N_14363);
nand U16247 (N_16247,N_15999,N_15725);
and U16248 (N_16248,N_14259,N_15696);
or U16249 (N_16249,N_14823,N_14080);
and U16250 (N_16250,N_15347,N_15763);
xnor U16251 (N_16251,N_14269,N_15467);
nand U16252 (N_16252,N_14899,N_14733);
and U16253 (N_16253,N_15880,N_14144);
or U16254 (N_16254,N_14830,N_14681);
xor U16255 (N_16255,N_14992,N_15283);
and U16256 (N_16256,N_14572,N_15856);
and U16257 (N_16257,N_15042,N_14427);
xor U16258 (N_16258,N_14317,N_15893);
nand U16259 (N_16259,N_14480,N_15112);
or U16260 (N_16260,N_15638,N_14452);
nor U16261 (N_16261,N_14803,N_15560);
nor U16262 (N_16262,N_15265,N_14682);
nor U16263 (N_16263,N_15945,N_14609);
and U16264 (N_16264,N_15413,N_14272);
nand U16265 (N_16265,N_14436,N_14994);
or U16266 (N_16266,N_15073,N_14519);
or U16267 (N_16267,N_15373,N_14128);
nand U16268 (N_16268,N_14444,N_14779);
and U16269 (N_16269,N_15100,N_15301);
and U16270 (N_16270,N_14404,N_14280);
nand U16271 (N_16271,N_15858,N_15305);
or U16272 (N_16272,N_14454,N_15891);
or U16273 (N_16273,N_14790,N_15545);
nand U16274 (N_16274,N_15422,N_15412);
or U16275 (N_16275,N_14402,N_14598);
nand U16276 (N_16276,N_15121,N_15180);
nand U16277 (N_16277,N_15814,N_15083);
xor U16278 (N_16278,N_15566,N_14907);
nand U16279 (N_16279,N_15585,N_14069);
or U16280 (N_16280,N_15098,N_15418);
or U16281 (N_16281,N_15727,N_15962);
xor U16282 (N_16282,N_15986,N_15882);
nand U16283 (N_16283,N_15610,N_14769);
and U16284 (N_16284,N_14019,N_14814);
and U16285 (N_16285,N_14749,N_15549);
nand U16286 (N_16286,N_15266,N_14671);
nor U16287 (N_16287,N_14027,N_15229);
and U16288 (N_16288,N_14721,N_15223);
nor U16289 (N_16289,N_14353,N_14073);
or U16290 (N_16290,N_15506,N_15270);
nor U16291 (N_16291,N_14902,N_15675);
and U16292 (N_16292,N_15334,N_14099);
nor U16293 (N_16293,N_15938,N_14921);
nor U16294 (N_16294,N_15628,N_14179);
nand U16295 (N_16295,N_14380,N_14554);
nand U16296 (N_16296,N_14403,N_14228);
nand U16297 (N_16297,N_15067,N_15838);
nand U16298 (N_16298,N_14278,N_15181);
nor U16299 (N_16299,N_14742,N_15002);
nor U16300 (N_16300,N_14235,N_15916);
nor U16301 (N_16301,N_14368,N_14398);
xor U16302 (N_16302,N_15680,N_14067);
or U16303 (N_16303,N_15614,N_14949);
or U16304 (N_16304,N_15595,N_14506);
or U16305 (N_16305,N_14865,N_14076);
or U16306 (N_16306,N_14858,N_15768);
or U16307 (N_16307,N_14942,N_14953);
nand U16308 (N_16308,N_14369,N_14815);
and U16309 (N_16309,N_14138,N_15872);
nor U16310 (N_16310,N_15653,N_14033);
nand U16311 (N_16311,N_14133,N_15046);
nand U16312 (N_16312,N_15377,N_14679);
and U16313 (N_16313,N_14521,N_15451);
nand U16314 (N_16314,N_15592,N_14667);
and U16315 (N_16315,N_14757,N_14509);
xor U16316 (N_16316,N_14490,N_15227);
and U16317 (N_16317,N_15661,N_15894);
and U16318 (N_16318,N_15287,N_15607);
or U16319 (N_16319,N_14739,N_15939);
nand U16320 (N_16320,N_15199,N_15766);
or U16321 (N_16321,N_14938,N_15149);
nand U16322 (N_16322,N_14236,N_15756);
nand U16323 (N_16323,N_15365,N_15226);
xor U16324 (N_16324,N_15198,N_15554);
xor U16325 (N_16325,N_14100,N_15997);
nor U16326 (N_16326,N_15823,N_14660);
or U16327 (N_16327,N_15254,N_15312);
or U16328 (N_16328,N_15644,N_14351);
or U16329 (N_16329,N_14996,N_15436);
nor U16330 (N_16330,N_14001,N_14319);
nand U16331 (N_16331,N_15010,N_15136);
nor U16332 (N_16332,N_15252,N_15431);
nor U16333 (N_16333,N_15196,N_15908);
and U16334 (N_16334,N_15579,N_14798);
nand U16335 (N_16335,N_15656,N_15815);
or U16336 (N_16336,N_15390,N_15507);
nor U16337 (N_16337,N_15061,N_15423);
nand U16338 (N_16338,N_15558,N_14705);
nor U16339 (N_16339,N_15409,N_14916);
nand U16340 (N_16340,N_15749,N_14636);
or U16341 (N_16341,N_14623,N_15869);
and U16342 (N_16342,N_14003,N_14225);
xor U16343 (N_16343,N_14294,N_14783);
and U16344 (N_16344,N_15697,N_15471);
and U16345 (N_16345,N_15681,N_15155);
nor U16346 (N_16346,N_14796,N_14038);
nand U16347 (N_16347,N_14909,N_14822);
nor U16348 (N_16348,N_15528,N_14240);
nand U16349 (N_16349,N_14105,N_14277);
nor U16350 (N_16350,N_15439,N_15643);
xor U16351 (N_16351,N_14756,N_14786);
and U16352 (N_16352,N_15583,N_15952);
and U16353 (N_16353,N_14601,N_15256);
nand U16354 (N_16354,N_14511,N_15803);
or U16355 (N_16355,N_15400,N_15297);
nand U16356 (N_16356,N_15173,N_15044);
or U16357 (N_16357,N_15764,N_15516);
and U16358 (N_16358,N_15194,N_14775);
xnor U16359 (N_16359,N_14422,N_14821);
nand U16360 (N_16360,N_14675,N_14297);
and U16361 (N_16361,N_15676,N_14734);
and U16362 (N_16362,N_15936,N_14552);
or U16363 (N_16363,N_14025,N_15651);
xnor U16364 (N_16364,N_14258,N_14925);
nor U16365 (N_16365,N_14337,N_15974);
or U16366 (N_16366,N_14030,N_15313);
nand U16367 (N_16367,N_14286,N_15842);
xor U16368 (N_16368,N_15131,N_15428);
xor U16369 (N_16369,N_15686,N_14869);
xnor U16370 (N_16370,N_15861,N_14727);
nor U16371 (N_16371,N_15231,N_14523);
nand U16372 (N_16372,N_15796,N_14993);
or U16373 (N_16373,N_14241,N_15859);
nor U16374 (N_16374,N_14210,N_14849);
xnor U16375 (N_16375,N_15951,N_14868);
and U16376 (N_16376,N_15267,N_15961);
or U16377 (N_16377,N_14018,N_14031);
nand U16378 (N_16378,N_14906,N_14913);
and U16379 (N_16379,N_14608,N_15292);
xor U16380 (N_16380,N_15954,N_14997);
and U16381 (N_16381,N_14904,N_15037);
nor U16382 (N_16382,N_15253,N_14321);
nor U16383 (N_16383,N_15158,N_15649);
nand U16384 (N_16384,N_14678,N_15659);
and U16385 (N_16385,N_14825,N_14155);
and U16386 (N_16386,N_15296,N_15789);
nand U16387 (N_16387,N_15381,N_14212);
nand U16388 (N_16388,N_14092,N_14690);
xor U16389 (N_16389,N_14799,N_15214);
and U16390 (N_16390,N_15051,N_15914);
or U16391 (N_16391,N_14279,N_15461);
xnor U16392 (N_16392,N_15529,N_15447);
nand U16393 (N_16393,N_15819,N_14348);
nor U16394 (N_16394,N_14626,N_14026);
or U16395 (N_16395,N_14718,N_14457);
or U16396 (N_16396,N_15801,N_14012);
or U16397 (N_16397,N_15440,N_15576);
nand U16398 (N_16398,N_14075,N_14333);
and U16399 (N_16399,N_15417,N_15430);
xnor U16400 (N_16400,N_15981,N_15760);
nor U16401 (N_16401,N_15724,N_15017);
or U16402 (N_16402,N_14843,N_14094);
and U16403 (N_16403,N_14513,N_15802);
or U16404 (N_16404,N_15984,N_15240);
nand U16405 (N_16405,N_14483,N_14274);
nand U16406 (N_16406,N_14357,N_15550);
nor U16407 (N_16407,N_15547,N_15933);
xor U16408 (N_16408,N_15485,N_15000);
or U16409 (N_16409,N_15468,N_14981);
and U16410 (N_16410,N_15870,N_14438);
or U16411 (N_16411,N_15230,N_14541);
nor U16412 (N_16412,N_14409,N_14139);
or U16413 (N_16413,N_14413,N_14975);
nand U16414 (N_16414,N_15369,N_14447);
or U16415 (N_16415,N_14627,N_14782);
nand U16416 (N_16416,N_15406,N_14544);
xnor U16417 (N_16417,N_15769,N_15693);
nor U16418 (N_16418,N_15024,N_15328);
and U16419 (N_16419,N_14119,N_15008);
or U16420 (N_16420,N_15307,N_15120);
nand U16421 (N_16421,N_15284,N_15940);
and U16422 (N_16422,N_15355,N_15294);
xor U16423 (N_16423,N_15416,N_14460);
nand U16424 (N_16424,N_15323,N_14017);
xor U16425 (N_16425,N_14857,N_14551);
nand U16426 (N_16426,N_14200,N_14950);
and U16427 (N_16427,N_14842,N_14537);
or U16428 (N_16428,N_15004,N_15694);
xor U16429 (N_16429,N_15410,N_14021);
or U16430 (N_16430,N_15237,N_14978);
nand U16431 (N_16431,N_14536,N_14344);
nor U16432 (N_16432,N_15494,N_15738);
nor U16433 (N_16433,N_14157,N_15258);
or U16434 (N_16434,N_15729,N_14173);
xnor U16435 (N_16435,N_15318,N_14748);
or U16436 (N_16436,N_15705,N_15949);
nand U16437 (N_16437,N_15316,N_15732);
nor U16438 (N_16438,N_14495,N_15048);
nor U16439 (N_16439,N_14256,N_14408);
xor U16440 (N_16440,N_14582,N_14022);
and U16441 (N_16441,N_15503,N_15309);
and U16442 (N_16442,N_14077,N_14216);
nor U16443 (N_16443,N_15127,N_14081);
nand U16444 (N_16444,N_14376,N_14129);
and U16445 (N_16445,N_15277,N_15457);
and U16446 (N_16446,N_14986,N_15752);
nand U16447 (N_16447,N_15454,N_14741);
or U16448 (N_16448,N_14005,N_14922);
nand U16449 (N_16449,N_14855,N_15087);
and U16450 (N_16450,N_15426,N_15486);
nand U16451 (N_16451,N_14616,N_14476);
nor U16452 (N_16452,N_15487,N_15341);
or U16453 (N_16453,N_14044,N_14149);
xnor U16454 (N_16454,N_15126,N_14619);
nand U16455 (N_16455,N_14961,N_15805);
and U16456 (N_16456,N_15524,N_14976);
or U16457 (N_16457,N_14685,N_15960);
nor U16458 (N_16458,N_14036,N_15084);
or U16459 (N_16459,N_15818,N_14931);
and U16460 (N_16460,N_14041,N_15973);
and U16461 (N_16461,N_15747,N_14219);
or U16462 (N_16462,N_14238,N_15937);
nand U16463 (N_16463,N_15532,N_15142);
nor U16464 (N_16464,N_15119,N_15711);
nor U16465 (N_16465,N_15460,N_15631);
nor U16466 (N_16466,N_15109,N_14172);
nor U16467 (N_16467,N_14911,N_14774);
nand U16468 (N_16468,N_15179,N_15689);
or U16469 (N_16469,N_15709,N_15217);
and U16470 (N_16470,N_15090,N_15124);
nand U16471 (N_16471,N_14577,N_14684);
nor U16472 (N_16472,N_15188,N_15931);
nor U16473 (N_16473,N_15408,N_14500);
and U16474 (N_16474,N_15980,N_14325);
nor U16475 (N_16475,N_15152,N_14420);
nand U16476 (N_16476,N_14707,N_14914);
nor U16477 (N_16477,N_14725,N_15797);
or U16478 (N_16478,N_15175,N_14651);
or U16479 (N_16479,N_14930,N_14694);
and U16480 (N_16480,N_14957,N_15291);
and U16481 (N_16481,N_15151,N_14762);
nor U16482 (N_16482,N_14295,N_14765);
xor U16483 (N_16483,N_15245,N_15790);
and U16484 (N_16484,N_14697,N_14118);
and U16485 (N_16485,N_14770,N_15274);
nand U16486 (N_16486,N_14501,N_14426);
and U16487 (N_16487,N_15444,N_15941);
nor U16488 (N_16488,N_14591,N_15911);
or U16489 (N_16489,N_14009,N_15069);
and U16490 (N_16490,N_15847,N_15455);
or U16491 (N_16491,N_15584,N_14947);
or U16492 (N_16492,N_15885,N_14004);
and U16493 (N_16493,N_14927,N_15655);
nand U16494 (N_16494,N_14372,N_14665);
xor U16495 (N_16495,N_14214,N_15829);
or U16496 (N_16496,N_14184,N_14106);
nor U16497 (N_16497,N_15210,N_15033);
or U16498 (N_16498,N_14434,N_14151);
nor U16499 (N_16499,N_15555,N_14882);
nor U16500 (N_16500,N_15982,N_15021);
and U16501 (N_16501,N_14517,N_14310);
nand U16502 (N_16502,N_14792,N_15737);
nand U16503 (N_16503,N_14809,N_15023);
nor U16504 (N_16504,N_14781,N_15947);
nand U16505 (N_16505,N_15456,N_14013);
and U16506 (N_16506,N_15335,N_14112);
or U16507 (N_16507,N_15338,N_14700);
nor U16508 (N_16508,N_14275,N_14641);
or U16509 (N_16509,N_14638,N_14263);
or U16510 (N_16510,N_14309,N_14083);
xor U16511 (N_16511,N_14764,N_14874);
and U16512 (N_16512,N_14525,N_15903);
and U16513 (N_16513,N_15346,N_15889);
or U16514 (N_16514,N_14110,N_15139);
or U16515 (N_16515,N_15535,N_14545);
nor U16516 (N_16516,N_15187,N_14548);
and U16517 (N_16517,N_15178,N_15699);
nand U16518 (N_16518,N_15278,N_15162);
nand U16519 (N_16519,N_14612,N_15054);
nand U16520 (N_16520,N_14169,N_14967);
xor U16521 (N_16521,N_14698,N_15953);
or U16522 (N_16522,N_14469,N_15742);
nand U16523 (N_16523,N_15407,N_15537);
nand U16524 (N_16524,N_14834,N_15123);
and U16525 (N_16525,N_14416,N_14478);
nor U16526 (N_16526,N_14873,N_14390);
nand U16527 (N_16527,N_14095,N_15698);
nor U16528 (N_16528,N_14057,N_15133);
nor U16529 (N_16529,N_14034,N_14719);
and U16530 (N_16530,N_14937,N_15568);
and U16531 (N_16531,N_15344,N_14113);
and U16532 (N_16532,N_15811,N_14746);
nor U16533 (N_16533,N_14617,N_14929);
or U16534 (N_16534,N_14370,N_15714);
nand U16535 (N_16535,N_15905,N_14098);
or U16536 (N_16536,N_15591,N_14029);
or U16537 (N_16537,N_15987,N_15009);
or U16538 (N_16538,N_15300,N_14239);
and U16539 (N_16539,N_14446,N_15721);
nand U16540 (N_16540,N_15617,N_14604);
nand U16541 (N_16541,N_14023,N_15944);
or U16542 (N_16542,N_15640,N_15167);
nor U16543 (N_16543,N_14066,N_14607);
xnor U16544 (N_16544,N_15314,N_15403);
nand U16545 (N_16545,N_14530,N_15833);
nand U16546 (N_16546,N_15419,N_14618);
nor U16547 (N_16547,N_14482,N_15209);
nor U16548 (N_16548,N_15707,N_14091);
or U16549 (N_16549,N_14565,N_15472);
xor U16550 (N_16550,N_14097,N_15543);
nand U16551 (N_16551,N_15733,N_14624);
nand U16552 (N_16552,N_14167,N_14415);
xnor U16553 (N_16553,N_14007,N_15477);
and U16554 (N_16554,N_15014,N_15972);
and U16555 (N_16555,N_15881,N_15156);
and U16556 (N_16556,N_15348,N_14192);
xnor U16557 (N_16557,N_14969,N_15036);
and U16558 (N_16558,N_14772,N_15915);
nand U16559 (N_16559,N_15358,N_15969);
nor U16560 (N_16560,N_15104,N_15411);
or U16561 (N_16561,N_15895,N_15826);
or U16562 (N_16562,N_15957,N_14691);
xor U16563 (N_16563,N_15505,N_14440);
or U16564 (N_16564,N_15371,N_14584);
nand U16565 (N_16565,N_14722,N_14898);
or U16566 (N_16566,N_14141,N_14035);
nand U16567 (N_16567,N_15354,N_15095);
or U16568 (N_16568,N_15668,N_14227);
nand U16569 (N_16569,N_14605,N_15141);
or U16570 (N_16570,N_14435,N_15703);
nand U16571 (N_16571,N_14970,N_14524);
or U16572 (N_16572,N_14877,N_15664);
nor U16573 (N_16573,N_15539,N_14542);
or U16574 (N_16574,N_15988,N_14290);
nor U16575 (N_16575,N_14973,N_15731);
and U16576 (N_16576,N_14801,N_14813);
nand U16577 (N_16577,N_14265,N_14311);
nor U16578 (N_16578,N_15375,N_15172);
or U16579 (N_16579,N_15081,N_15575);
nor U16580 (N_16580,N_14730,N_14689);
or U16581 (N_16581,N_15212,N_14336);
or U16582 (N_16582,N_15684,N_15105);
nand U16583 (N_16583,N_14692,N_14109);
or U16584 (N_16584,N_14211,N_14244);
nand U16585 (N_16585,N_14231,N_14870);
nor U16586 (N_16586,N_15762,N_15285);
and U16587 (N_16587,N_15985,N_15831);
and U16588 (N_16588,N_14534,N_15405);
nor U16589 (N_16589,N_14962,N_14872);
nand U16590 (N_16590,N_14793,N_14104);
xor U16591 (N_16591,N_14785,N_14758);
nor U16592 (N_16592,N_15497,N_14954);
xor U16593 (N_16593,N_14260,N_14531);
and U16594 (N_16594,N_14737,N_14549);
nor U16595 (N_16595,N_15827,N_14479);
or U16596 (N_16596,N_15034,N_14289);
nand U16597 (N_16597,N_14043,N_15197);
xnor U16598 (N_16598,N_14533,N_15608);
nand U16599 (N_16599,N_14637,N_14117);
or U16600 (N_16600,N_14046,N_15234);
nor U16601 (N_16601,N_14298,N_14379);
nand U16602 (N_16602,N_15896,N_15016);
nand U16603 (N_16603,N_15745,N_14918);
or U16604 (N_16604,N_15639,N_15772);
or U16605 (N_16605,N_15470,N_15275);
and U16606 (N_16606,N_15662,N_14699);
nand U16607 (N_16607,N_15780,N_15148);
nor U16608 (N_16608,N_15429,N_14578);
nand U16609 (N_16609,N_15955,N_14203);
nand U16610 (N_16610,N_15785,N_15432);
and U16611 (N_16611,N_15934,N_14759);
nor U16612 (N_16612,N_15415,N_15816);
or U16613 (N_16613,N_14875,N_15337);
nor U16614 (N_16614,N_15099,N_14844);
and U16615 (N_16615,N_15910,N_15719);
nor U16616 (N_16616,N_14204,N_15356);
nand U16617 (N_16617,N_15499,N_14988);
nor U16618 (N_16618,N_14941,N_15160);
and U16619 (N_16619,N_14188,N_15674);
nor U16620 (N_16620,N_15604,N_14655);
nand U16621 (N_16621,N_15935,N_14024);
nor U16622 (N_16622,N_15646,N_15533);
and U16623 (N_16623,N_14394,N_14650);
and U16624 (N_16624,N_14791,N_15362);
and U16625 (N_16625,N_15809,N_14716);
and U16626 (N_16626,N_15720,N_14903);
xor U16627 (N_16627,N_15897,N_15625);
nor U16628 (N_16628,N_14635,N_15723);
xnor U16629 (N_16629,N_14049,N_15329);
nor U16630 (N_16630,N_15340,N_15755);
nor U16631 (N_16631,N_15476,N_15757);
nand U16632 (N_16632,N_14209,N_14859);
nand U16633 (N_16633,N_15701,N_14794);
nor U16634 (N_16634,N_15247,N_15089);
nand U16635 (N_16635,N_14657,N_15450);
nor U16636 (N_16636,N_15480,N_15068);
xnor U16637 (N_16637,N_14285,N_15311);
nor U16638 (N_16638,N_14051,N_14629);
nor U16639 (N_16639,N_14613,N_15056);
and U16640 (N_16640,N_15031,N_14896);
nand U16641 (N_16641,N_15990,N_15587);
nor U16642 (N_16642,N_14569,N_14068);
and U16643 (N_16643,N_15518,N_14833);
nand U16644 (N_16644,N_15530,N_15391);
or U16645 (N_16645,N_14812,N_14936);
nor U16646 (N_16646,N_15667,N_14713);
xor U16647 (N_16647,N_15434,N_14360);
or U16648 (N_16648,N_14850,N_14575);
or U16649 (N_16649,N_15228,N_14419);
xor U16650 (N_16650,N_15906,N_14195);
nand U16651 (N_16651,N_14347,N_14683);
and U16652 (N_16652,N_15129,N_14301);
or U16653 (N_16653,N_15221,N_15817);
and U16654 (N_16654,N_14327,N_15244);
nand U16655 (N_16655,N_15263,N_15551);
xnor U16656 (N_16656,N_15029,N_15788);
or U16657 (N_16657,N_15813,N_14861);
xor U16658 (N_16658,N_15484,N_15799);
and U16659 (N_16659,N_15824,N_14982);
or U16660 (N_16660,N_14163,N_14008);
or U16661 (N_16661,N_14304,N_15994);
nand U16662 (N_16662,N_15374,N_14649);
or U16663 (N_16663,N_15458,N_15402);
and U16664 (N_16664,N_15991,N_14300);
xnor U16665 (N_16665,N_15116,N_14504);
or U16666 (N_16666,N_15243,N_14886);
or U16667 (N_16667,N_15057,N_14808);
or U16668 (N_16668,N_14388,N_14526);
nor U16669 (N_16669,N_14411,N_15523);
nor U16670 (N_16670,N_14299,N_14965);
nor U16671 (N_16671,N_14883,N_14802);
and U16672 (N_16672,N_14520,N_14045);
or U16673 (N_16673,N_15453,N_14945);
xnor U16674 (N_16674,N_15154,N_15993);
nor U16675 (N_16675,N_15433,N_14826);
nand U16676 (N_16676,N_14747,N_14854);
nor U16677 (N_16677,N_14386,N_15624);
or U16678 (N_16678,N_14816,N_15071);
and U16679 (N_16679,N_14178,N_15621);
nor U16680 (N_16680,N_15153,N_14284);
nand U16681 (N_16681,N_14373,N_15215);
xor U16682 (N_16682,N_14473,N_15660);
and U16683 (N_16683,N_15635,N_14944);
or U16684 (N_16684,N_15665,N_15106);
or U16685 (N_16685,N_15007,N_14146);
nand U16686 (N_16686,N_15673,N_15092);
and U16687 (N_16687,N_14152,N_14771);
or U16688 (N_16688,N_15573,N_14377);
nand U16689 (N_16689,N_15047,N_14502);
nor U16690 (N_16690,N_15808,N_15103);
nor U16691 (N_16691,N_14654,N_15793);
and U16692 (N_16692,N_15259,N_15959);
and U16693 (N_16693,N_15233,N_15812);
and U16694 (N_16694,N_14159,N_15569);
and U16695 (N_16695,N_14150,N_15308);
nand U16696 (N_16696,N_15282,N_15754);
and U16697 (N_16697,N_15976,N_15327);
nand U16698 (N_16698,N_14320,N_15213);
or U16699 (N_16699,N_15627,N_14979);
and U16700 (N_16700,N_14471,N_15035);
nor U16701 (N_16701,N_15841,N_15404);
or U16702 (N_16702,N_14062,N_15840);
nand U16703 (N_16703,N_15606,N_14355);
nand U16704 (N_16704,N_15967,N_14934);
nand U16705 (N_16705,N_15603,N_14732);
and U16706 (N_16706,N_15948,N_15928);
nor U16707 (N_16707,N_15517,N_15538);
nand U16708 (N_16708,N_15692,N_15864);
and U16709 (N_16709,N_14191,N_14932);
nand U16710 (N_16710,N_14050,N_14407);
and U16711 (N_16711,N_15059,N_14342);
or U16712 (N_16712,N_15580,N_14451);
nand U16713 (N_16713,N_14350,N_15189);
and U16714 (N_16714,N_15239,N_15743);
xnor U16715 (N_16715,N_14881,N_15715);
nor U16716 (N_16716,N_15926,N_14645);
xnor U16717 (N_16717,N_14807,N_14127);
nand U16718 (N_16718,N_15279,N_15784);
nand U16719 (N_16719,N_14515,N_15204);
or U16720 (N_16720,N_15687,N_15088);
nor U16721 (N_16721,N_14039,N_15783);
or U16722 (N_16722,N_14283,N_14481);
nor U16723 (N_16723,N_14666,N_14470);
nand U16724 (N_16724,N_14014,N_15657);
xor U16725 (N_16725,N_15645,N_15570);
nor U16726 (N_16726,N_15310,N_14392);
or U16727 (N_16727,N_15325,N_14701);
or U16728 (N_16728,N_15855,N_14341);
xnor U16729 (N_16729,N_15542,N_15389);
nor U16730 (N_16730,N_14071,N_15806);
and U16731 (N_16731,N_15500,N_14079);
nand U16732 (N_16732,N_14797,N_15052);
nand U16733 (N_16733,N_15531,N_15849);
or U16734 (N_16734,N_15892,N_14334);
and U16735 (N_16735,N_14562,N_15702);
nand U16736 (N_16736,N_14201,N_14972);
or U16737 (N_16737,N_14218,N_15736);
nand U16738 (N_16738,N_15970,N_15050);
or U16739 (N_16739,N_15519,N_14884);
nor U16740 (N_16740,N_15932,N_15963);
and U16741 (N_16741,N_15134,N_15594);
or U16742 (N_16742,N_14354,N_15118);
and U16743 (N_16743,N_15383,N_15942);
nor U16744 (N_16744,N_15493,N_14599);
and U16745 (N_16745,N_15589,N_15598);
and U16746 (N_16746,N_14960,N_15272);
nor U16747 (N_16747,N_14461,N_15039);
nand U16748 (N_16748,N_14610,N_14174);
nor U16749 (N_16749,N_15632,N_15349);
or U16750 (N_16750,N_14631,N_15027);
nor U16751 (N_16751,N_15534,N_15441);
and U16752 (N_16752,N_15863,N_14135);
xor U16753 (N_16753,N_15888,N_15079);
or U16754 (N_16754,N_15900,N_14811);
and U16755 (N_16755,N_14303,N_14040);
nor U16756 (N_16756,N_15235,N_14010);
or U16757 (N_16757,N_14535,N_14510);
nor U16758 (N_16758,N_15740,N_15250);
nor U16759 (N_16759,N_14084,N_15878);
nor U16760 (N_16760,N_14687,N_14819);
nand U16761 (N_16761,N_15321,N_15750);
and U16762 (N_16762,N_14462,N_15734);
nand U16763 (N_16763,N_15679,N_14717);
and U16764 (N_16764,N_15877,N_14335);
nand U16765 (N_16765,N_15564,N_14491);
nor U16766 (N_16766,N_14753,N_14458);
or U16767 (N_16767,N_14497,N_15184);
nand U16768 (N_16768,N_14827,N_14832);
nor U16769 (N_16769,N_14848,N_14773);
nor U16770 (N_16770,N_15111,N_14291);
and U16771 (N_16771,N_14661,N_15759);
nor U16772 (N_16772,N_15887,N_14712);
and U16773 (N_16773,N_15190,N_14425);
xor U16774 (N_16774,N_14496,N_15726);
nor U16775 (N_16775,N_15216,N_15435);
or U16776 (N_16776,N_15392,N_15601);
nand U16777 (N_16777,N_14405,N_15170);
nor U16778 (N_16778,N_14860,N_14002);
and U16779 (N_16779,N_15043,N_15192);
nand U16780 (N_16780,N_14507,N_15611);
and U16781 (N_16781,N_15137,N_15045);
nor U16782 (N_16782,N_14977,N_14467);
xor U16783 (N_16783,N_15006,N_14516);
xor U16784 (N_16784,N_14177,N_15751);
and U16785 (N_16785,N_14611,N_14389);
nand U16786 (N_16786,N_14829,N_15255);
nor U16787 (N_16787,N_15979,N_14696);
nor U16788 (N_16788,N_14563,N_14393);
nand U16789 (N_16789,N_14262,N_14652);
xnor U16790 (N_16790,N_14538,N_14102);
nor U16791 (N_16791,N_15901,N_14006);
or U16792 (N_16792,N_14223,N_14114);
nand U16793 (N_16793,N_15361,N_14780);
or U16794 (N_16794,N_15781,N_14245);
and U16795 (N_16795,N_15364,N_15522);
nand U16796 (N_16796,N_14897,N_14397);
or U16797 (N_16797,N_14052,N_15359);
nand U16798 (N_16798,N_15761,N_14890);
nor U16799 (N_16799,N_14946,N_15019);
or U16800 (N_16800,N_14888,N_15336);
and U16801 (N_16801,N_15619,N_14715);
or U16802 (N_16802,N_15609,N_15249);
nor U16803 (N_16803,N_15851,N_15678);
nor U16804 (N_16804,N_14788,N_15304);
xnor U16805 (N_16805,N_15273,N_14237);
nand U16806 (N_16806,N_14161,N_15848);
nor U16807 (N_16807,N_15028,N_14055);
nand U16808 (N_16808,N_15357,N_14125);
and U16809 (N_16809,N_14919,N_15378);
nand U16810 (N_16810,N_15135,N_15810);
nor U16811 (N_16811,N_14905,N_14307);
or U16812 (N_16812,N_15958,N_15717);
xnor U16813 (N_16813,N_14653,N_14391);
and U16814 (N_16814,N_15372,N_14964);
or U16815 (N_16815,N_15022,N_15442);
or U16816 (N_16816,N_14132,N_15602);
or U16817 (N_16817,N_15735,N_15821);
or U16818 (N_16818,N_14089,N_15205);
xnor U16819 (N_16819,N_14831,N_14485);
nor U16820 (N_16820,N_14472,N_14197);
nand U16821 (N_16821,N_15536,N_14340);
nand U16822 (N_16822,N_15586,N_14199);
nor U16823 (N_16823,N_15515,N_14165);
nand U16824 (N_16824,N_15866,N_14093);
nor U16825 (N_16825,N_14948,N_14486);
nor U16826 (N_16826,N_14955,N_15469);
nor U16827 (N_16827,N_14078,N_14343);
nor U16828 (N_16828,N_15844,N_15902);
nor U16829 (N_16829,N_15395,N_15597);
nor U16830 (N_16830,N_14639,N_15195);
nor U16831 (N_16831,N_14600,N_14910);
nor U16832 (N_16832,N_15225,N_15082);
nand U16833 (N_16833,N_15552,N_15883);
xnor U16834 (N_16834,N_15315,N_14433);
nand U16835 (N_16835,N_14185,N_15038);
and U16836 (N_16836,N_15791,N_15401);
nand U16837 (N_16837,N_15174,N_15144);
nand U16838 (N_16838,N_14933,N_14308);
nor U16839 (N_16839,N_14315,N_15147);
or U16840 (N_16840,N_14622,N_14418);
or U16841 (N_16841,N_15203,N_15055);
and U16842 (N_16842,N_15971,N_14406);
and U16843 (N_16843,N_14633,N_14586);
nor U16844 (N_16844,N_14959,N_14345);
nor U16845 (N_16845,N_15488,N_14755);
and U16846 (N_16846,N_15464,N_15080);
nor U16847 (N_16847,N_15020,N_15912);
nand U16848 (N_16848,N_14646,N_15438);
nor U16849 (N_16849,N_14820,N_14048);
and U16850 (N_16850,N_15525,N_15145);
nand U16851 (N_16851,N_15886,N_15615);
nor U16852 (N_16852,N_15185,N_14153);
nor U16853 (N_16853,N_14991,N_15875);
nor U16854 (N_16854,N_14676,N_14248);
nand U16855 (N_16855,N_14261,N_14137);
or U16856 (N_16856,N_14449,N_14088);
xnor U16857 (N_16857,N_14168,N_15822);
nand U16858 (N_16858,N_14215,N_14983);
and U16859 (N_16859,N_15612,N_14160);
and U16860 (N_16860,N_15860,N_14463);
xor U16861 (N_16861,N_15553,N_15366);
or U16862 (N_16862,N_15091,N_15919);
nor U16863 (N_16863,N_15654,N_14059);
xor U16864 (N_16864,N_15541,N_14580);
or U16865 (N_16865,N_14475,N_14175);
nor U16866 (N_16866,N_14302,N_14559);
or U16867 (N_16867,N_14729,N_15837);
nor U16868 (N_16868,N_15165,N_15605);
and U16869 (N_16869,N_14845,N_15491);
nor U16870 (N_16870,N_15786,N_14042);
nor U16871 (N_16871,N_15248,N_14108);
nor U16872 (N_16872,N_15352,N_15333);
and U16873 (N_16873,N_15526,N_14140);
and U16874 (N_16874,N_15977,N_15950);
or U16875 (N_16875,N_14980,N_14484);
nand U16876 (N_16876,N_15385,N_14305);
or U16877 (N_16877,N_15169,N_14410);
or U16878 (N_16878,N_14573,N_14956);
and U16879 (N_16879,N_14492,N_15113);
nand U16880 (N_16880,N_15345,N_15498);
nand U16881 (N_16881,N_14271,N_15339);
nor U16882 (N_16882,N_15546,N_15157);
xor U16883 (N_16883,N_14592,N_14789);
and U16884 (N_16884,N_14628,N_15559);
and U16885 (N_16885,N_15730,N_15324);
nor U16886 (N_16886,N_15577,N_14917);
or U16887 (N_16887,N_15561,N_14837);
nor U16888 (N_16888,N_15899,N_14680);
or U16889 (N_16889,N_14205,N_14384);
and U16890 (N_16890,N_14047,N_14293);
nor U16891 (N_16891,N_15290,N_15448);
xnor U16892 (N_16892,N_15832,N_14677);
nand U16893 (N_16893,N_14206,N_14706);
nor U16894 (N_16894,N_14385,N_14437);
nor U16895 (N_16895,N_15319,N_15074);
and U16896 (N_16896,N_14576,N_15062);
nand U16897 (N_16897,N_14709,N_14193);
nor U16898 (N_16898,N_15183,N_15748);
nor U16899 (N_16899,N_14445,N_14111);
or U16900 (N_16900,N_15835,N_15150);
or U16901 (N_16901,N_15636,N_15191);
nor U16902 (N_16902,N_15306,N_15449);
nand U16903 (N_16903,N_14171,N_15276);
xnor U16904 (N_16904,N_14574,N_14090);
nor U16905 (N_16905,N_14522,N_15777);
and U16906 (N_16906,N_15798,N_14349);
and U16907 (N_16907,N_14439,N_14594);
and U16908 (N_16908,N_15682,N_15320);
and U16909 (N_16909,N_15800,N_15770);
xor U16910 (N_16910,N_15567,N_15708);
nand U16911 (N_16911,N_15923,N_15207);
nor U16912 (N_16912,N_14999,N_14695);
nor U16913 (N_16913,N_14273,N_14583);
nor U16914 (N_16914,N_14810,N_15623);
nor U16915 (N_16915,N_15086,N_15548);
nand U16916 (N_16916,N_15626,N_14740);
or U16917 (N_16917,N_14714,N_15846);
nor U16918 (N_16918,N_15581,N_15224);
nor U16919 (N_16919,N_15206,N_14862);
nor U16920 (N_16920,N_14082,N_14330);
nand U16921 (N_16921,N_14668,N_15509);
xor U16922 (N_16922,N_15718,N_14131);
nand U16923 (N_16923,N_15520,N_15200);
and U16924 (N_16924,N_14400,N_14338);
and U16925 (N_16925,N_14314,N_14951);
nor U16926 (N_16926,N_14352,N_15060);
nor U16927 (N_16927,N_14448,N_14121);
or U16928 (N_16928,N_15075,N_14878);
and U16929 (N_16929,N_14647,N_15741);
nand U16930 (N_16930,N_15322,N_14871);
and U16931 (N_16931,N_15648,N_14587);
xnor U16932 (N_16932,N_15854,N_14595);
nor U16933 (N_16933,N_14923,N_14181);
or U16934 (N_16934,N_15093,N_14514);
nor U16935 (N_16935,N_14726,N_15767);
or U16936 (N_16936,N_15992,N_15710);
nand U16937 (N_16937,N_15521,N_14736);
nand U16938 (N_16938,N_14908,N_14743);
nand U16939 (N_16939,N_14555,N_15242);
and U16940 (N_16940,N_15293,N_15758);
nor U16941 (N_16941,N_15779,N_15302);
or U16942 (N_16942,N_15774,N_14065);
and U16943 (N_16943,N_15397,N_15857);
xnor U16944 (N_16944,N_14186,N_15489);
and U16945 (N_16945,N_15473,N_14226);
and U16946 (N_16946,N_15965,N_14096);
nor U16947 (N_16947,N_15298,N_14561);
nand U16948 (N_16948,N_14642,N_14270);
and U16949 (N_16949,N_14828,N_15295);
and U16950 (N_16950,N_14866,N_14207);
or U16951 (N_16951,N_15064,N_14220);
and U16952 (N_16952,N_15663,N_15288);
and U16953 (N_16953,N_14032,N_14101);
nand U16954 (N_16954,N_15825,N_14243);
nand U16955 (N_16955,N_15834,N_14915);
nor U16956 (N_16956,N_14356,N_15326);
nor U16957 (N_16957,N_15122,N_15424);
nor U16958 (N_16958,N_15670,N_14180);
and U16959 (N_16959,N_14971,N_15744);
nor U16960 (N_16960,N_14593,N_14670);
nor U16961 (N_16961,N_14136,N_14887);
or U16962 (N_16962,N_14926,N_14359);
xnor U16963 (N_16963,N_15989,N_15728);
nor U16964 (N_16964,N_14990,N_14318);
and U16965 (N_16965,N_14664,N_15593);
nand U16966 (N_16966,N_14939,N_15502);
or U16967 (N_16967,N_15807,N_14505);
and U16968 (N_16968,N_15630,N_14550);
and U16969 (N_16969,N_14371,N_14326);
and U16970 (N_16970,N_14147,N_14085);
or U16971 (N_16971,N_15482,N_15479);
and U16972 (N_16972,N_15492,N_14943);
nor U16973 (N_16973,N_15775,N_15652);
xnor U16974 (N_16974,N_14430,N_14148);
or U16975 (N_16975,N_14424,N_15794);
nor U16976 (N_16976,N_15414,N_14853);
and U16977 (N_16977,N_15107,N_14702);
nor U16978 (N_16978,N_15642,N_15202);
xor U16979 (N_16979,N_14230,N_15443);
nor U16980 (N_16980,N_14987,N_14892);
or U16981 (N_16981,N_14250,N_15996);
nor U16982 (N_16982,N_14901,N_14401);
nor U16983 (N_16983,N_15368,N_14840);
or U16984 (N_16984,N_14364,N_15222);
nor U16985 (N_16985,N_15077,N_14037);
nand U16986 (N_16986,N_15946,N_14123);
nand U16987 (N_16987,N_14634,N_15828);
nand U16988 (N_16988,N_14387,N_15241);
and U16989 (N_16989,N_15820,N_15360);
nor U16990 (N_16990,N_15706,N_15771);
and U16991 (N_16991,N_14465,N_14662);
nor U16992 (N_16992,N_14760,N_14766);
nor U16993 (N_16993,N_15669,N_14466);
or U16994 (N_16994,N_14412,N_15343);
nor U16995 (N_16995,N_14221,N_15463);
nand U16996 (N_16996,N_15040,N_15351);
nor U16997 (N_16997,N_14281,N_14488);
and U16998 (N_16998,N_15201,N_14312);
nand U16999 (N_16999,N_14074,N_15330);
or U17000 (N_17000,N_15762,N_14762);
nor U17001 (N_17001,N_14614,N_14277);
nor U17002 (N_17002,N_15770,N_15748);
nor U17003 (N_17003,N_15747,N_14403);
nand U17004 (N_17004,N_14365,N_15973);
nor U17005 (N_17005,N_14851,N_14668);
or U17006 (N_17006,N_15720,N_14464);
and U17007 (N_17007,N_15320,N_14610);
nand U17008 (N_17008,N_14535,N_14316);
and U17009 (N_17009,N_15231,N_15114);
and U17010 (N_17010,N_14111,N_14733);
nand U17011 (N_17011,N_15994,N_14002);
nor U17012 (N_17012,N_15990,N_14835);
nand U17013 (N_17013,N_15868,N_15545);
nor U17014 (N_17014,N_14091,N_15441);
nand U17015 (N_17015,N_15368,N_15014);
or U17016 (N_17016,N_14065,N_14796);
or U17017 (N_17017,N_15382,N_15026);
and U17018 (N_17018,N_15025,N_14097);
xor U17019 (N_17019,N_14024,N_15808);
nand U17020 (N_17020,N_14484,N_15295);
nand U17021 (N_17021,N_15860,N_14486);
or U17022 (N_17022,N_14130,N_15644);
xor U17023 (N_17023,N_15837,N_15078);
nor U17024 (N_17024,N_14390,N_15977);
nand U17025 (N_17025,N_14755,N_14342);
and U17026 (N_17026,N_14185,N_14448);
and U17027 (N_17027,N_15372,N_15770);
or U17028 (N_17028,N_14201,N_15248);
xor U17029 (N_17029,N_15120,N_15188);
and U17030 (N_17030,N_15427,N_14751);
nand U17031 (N_17031,N_15072,N_14999);
or U17032 (N_17032,N_14464,N_14348);
xor U17033 (N_17033,N_15154,N_15251);
and U17034 (N_17034,N_14569,N_15034);
or U17035 (N_17035,N_15986,N_14477);
and U17036 (N_17036,N_14203,N_14164);
nor U17037 (N_17037,N_15423,N_14305);
nand U17038 (N_17038,N_15517,N_14097);
and U17039 (N_17039,N_14019,N_15736);
nand U17040 (N_17040,N_14498,N_15212);
or U17041 (N_17041,N_14399,N_14353);
or U17042 (N_17042,N_15267,N_15881);
nand U17043 (N_17043,N_15046,N_15197);
or U17044 (N_17044,N_14610,N_15627);
or U17045 (N_17045,N_15022,N_14051);
nor U17046 (N_17046,N_15697,N_14801);
xor U17047 (N_17047,N_14116,N_14012);
nand U17048 (N_17048,N_15763,N_15563);
and U17049 (N_17049,N_14352,N_15467);
nand U17050 (N_17050,N_15616,N_14485);
or U17051 (N_17051,N_15430,N_15348);
nor U17052 (N_17052,N_14109,N_15537);
nor U17053 (N_17053,N_15651,N_14652);
xnor U17054 (N_17054,N_14101,N_15791);
nand U17055 (N_17055,N_15023,N_15931);
nor U17056 (N_17056,N_15693,N_15023);
or U17057 (N_17057,N_15712,N_15557);
and U17058 (N_17058,N_15863,N_15493);
or U17059 (N_17059,N_15876,N_15200);
or U17060 (N_17060,N_14833,N_14768);
nand U17061 (N_17061,N_15381,N_15040);
nor U17062 (N_17062,N_14124,N_14529);
xnor U17063 (N_17063,N_14566,N_15182);
nand U17064 (N_17064,N_14885,N_15552);
or U17065 (N_17065,N_14440,N_14050);
or U17066 (N_17066,N_15834,N_14608);
or U17067 (N_17067,N_15483,N_14177);
nor U17068 (N_17068,N_15604,N_15885);
or U17069 (N_17069,N_15997,N_14505);
or U17070 (N_17070,N_15804,N_14424);
nor U17071 (N_17071,N_14673,N_15892);
and U17072 (N_17072,N_15598,N_15338);
nor U17073 (N_17073,N_14102,N_14068);
nand U17074 (N_17074,N_15160,N_15580);
nand U17075 (N_17075,N_14222,N_14748);
and U17076 (N_17076,N_14313,N_15545);
nand U17077 (N_17077,N_14904,N_14466);
or U17078 (N_17078,N_14639,N_15008);
and U17079 (N_17079,N_14691,N_15721);
nand U17080 (N_17080,N_15768,N_15009);
or U17081 (N_17081,N_15134,N_14129);
or U17082 (N_17082,N_14168,N_15921);
nor U17083 (N_17083,N_15572,N_14964);
nand U17084 (N_17084,N_14123,N_14087);
nand U17085 (N_17085,N_14142,N_14493);
or U17086 (N_17086,N_15984,N_14240);
nand U17087 (N_17087,N_14714,N_14153);
nand U17088 (N_17088,N_15046,N_15908);
nor U17089 (N_17089,N_14748,N_14794);
nand U17090 (N_17090,N_14637,N_14092);
nand U17091 (N_17091,N_14021,N_15398);
and U17092 (N_17092,N_15052,N_15840);
xnor U17093 (N_17093,N_15504,N_14734);
or U17094 (N_17094,N_15096,N_15715);
nor U17095 (N_17095,N_15376,N_14105);
and U17096 (N_17096,N_14147,N_14097);
nand U17097 (N_17097,N_14353,N_14237);
and U17098 (N_17098,N_14353,N_15764);
xor U17099 (N_17099,N_14376,N_14277);
or U17100 (N_17100,N_14491,N_15846);
and U17101 (N_17101,N_14174,N_14592);
nand U17102 (N_17102,N_15512,N_15238);
and U17103 (N_17103,N_15520,N_14743);
xor U17104 (N_17104,N_15250,N_15847);
xor U17105 (N_17105,N_15743,N_14271);
nand U17106 (N_17106,N_14232,N_15902);
and U17107 (N_17107,N_14502,N_15766);
nor U17108 (N_17108,N_15256,N_15525);
nor U17109 (N_17109,N_15211,N_15332);
nor U17110 (N_17110,N_15194,N_15164);
and U17111 (N_17111,N_14824,N_14791);
or U17112 (N_17112,N_15274,N_14941);
and U17113 (N_17113,N_14103,N_15252);
and U17114 (N_17114,N_14782,N_14669);
nor U17115 (N_17115,N_14173,N_14720);
nor U17116 (N_17116,N_14226,N_15472);
nand U17117 (N_17117,N_14876,N_15202);
nor U17118 (N_17118,N_14022,N_14365);
nand U17119 (N_17119,N_15881,N_14109);
nand U17120 (N_17120,N_15410,N_15924);
and U17121 (N_17121,N_14599,N_14093);
nor U17122 (N_17122,N_14622,N_14253);
or U17123 (N_17123,N_15220,N_15702);
and U17124 (N_17124,N_14833,N_14667);
and U17125 (N_17125,N_14204,N_15175);
nor U17126 (N_17126,N_14381,N_14500);
nor U17127 (N_17127,N_14344,N_15256);
xor U17128 (N_17128,N_14926,N_15459);
or U17129 (N_17129,N_15973,N_14816);
xor U17130 (N_17130,N_15669,N_15112);
or U17131 (N_17131,N_15078,N_14597);
and U17132 (N_17132,N_14167,N_15278);
xnor U17133 (N_17133,N_14049,N_14176);
nor U17134 (N_17134,N_14923,N_14914);
and U17135 (N_17135,N_15332,N_14808);
and U17136 (N_17136,N_15762,N_15931);
nand U17137 (N_17137,N_15638,N_14074);
and U17138 (N_17138,N_14688,N_14802);
and U17139 (N_17139,N_15142,N_15669);
xnor U17140 (N_17140,N_15556,N_15573);
and U17141 (N_17141,N_14396,N_15952);
nand U17142 (N_17142,N_15608,N_14084);
nor U17143 (N_17143,N_15844,N_14439);
nor U17144 (N_17144,N_14622,N_14533);
nor U17145 (N_17145,N_14761,N_14946);
and U17146 (N_17146,N_14911,N_14250);
or U17147 (N_17147,N_15085,N_14119);
or U17148 (N_17148,N_15899,N_14269);
or U17149 (N_17149,N_15949,N_15256);
or U17150 (N_17150,N_15282,N_14339);
nand U17151 (N_17151,N_15384,N_14457);
and U17152 (N_17152,N_15626,N_15453);
and U17153 (N_17153,N_14948,N_14089);
nor U17154 (N_17154,N_14520,N_14083);
xnor U17155 (N_17155,N_15228,N_15938);
nor U17156 (N_17156,N_14240,N_15723);
nor U17157 (N_17157,N_15715,N_15712);
nor U17158 (N_17158,N_15086,N_15869);
nor U17159 (N_17159,N_15323,N_14102);
and U17160 (N_17160,N_14851,N_14412);
nand U17161 (N_17161,N_14620,N_15570);
nand U17162 (N_17162,N_14816,N_15830);
xnor U17163 (N_17163,N_15058,N_15734);
xor U17164 (N_17164,N_15349,N_14759);
or U17165 (N_17165,N_15387,N_14027);
xor U17166 (N_17166,N_14829,N_14869);
and U17167 (N_17167,N_15218,N_15408);
nor U17168 (N_17168,N_14761,N_14256);
and U17169 (N_17169,N_14997,N_15885);
nand U17170 (N_17170,N_15153,N_15775);
xor U17171 (N_17171,N_15977,N_15648);
nand U17172 (N_17172,N_15306,N_15272);
or U17173 (N_17173,N_14313,N_14432);
xnor U17174 (N_17174,N_14982,N_15055);
or U17175 (N_17175,N_14222,N_15625);
xor U17176 (N_17176,N_14985,N_15695);
nor U17177 (N_17177,N_14734,N_14301);
and U17178 (N_17178,N_15368,N_14707);
nor U17179 (N_17179,N_15399,N_14114);
nor U17180 (N_17180,N_14295,N_15313);
and U17181 (N_17181,N_15005,N_15934);
or U17182 (N_17182,N_15745,N_14870);
or U17183 (N_17183,N_14818,N_15315);
and U17184 (N_17184,N_15544,N_14536);
or U17185 (N_17185,N_14261,N_14039);
nand U17186 (N_17186,N_15626,N_14446);
nand U17187 (N_17187,N_15431,N_15393);
nand U17188 (N_17188,N_15409,N_15098);
and U17189 (N_17189,N_15140,N_14507);
and U17190 (N_17190,N_14906,N_14195);
nand U17191 (N_17191,N_14153,N_14185);
and U17192 (N_17192,N_14163,N_15126);
and U17193 (N_17193,N_14872,N_15766);
nand U17194 (N_17194,N_15743,N_15510);
and U17195 (N_17195,N_14567,N_14471);
and U17196 (N_17196,N_15679,N_14227);
nor U17197 (N_17197,N_14163,N_14920);
and U17198 (N_17198,N_15766,N_15770);
and U17199 (N_17199,N_14726,N_14116);
or U17200 (N_17200,N_14332,N_14751);
and U17201 (N_17201,N_15414,N_15721);
nor U17202 (N_17202,N_15145,N_15270);
or U17203 (N_17203,N_14584,N_15461);
and U17204 (N_17204,N_14793,N_14150);
nand U17205 (N_17205,N_15698,N_14043);
nor U17206 (N_17206,N_14837,N_14377);
nand U17207 (N_17207,N_15217,N_14177);
and U17208 (N_17208,N_14511,N_15416);
or U17209 (N_17209,N_14850,N_15485);
nand U17210 (N_17210,N_15497,N_14278);
nor U17211 (N_17211,N_14476,N_15108);
nand U17212 (N_17212,N_14432,N_14090);
nor U17213 (N_17213,N_14435,N_14309);
or U17214 (N_17214,N_15108,N_14143);
xor U17215 (N_17215,N_15158,N_15397);
nor U17216 (N_17216,N_15242,N_15856);
or U17217 (N_17217,N_15813,N_15668);
nand U17218 (N_17218,N_14712,N_15236);
and U17219 (N_17219,N_14032,N_15611);
nand U17220 (N_17220,N_14458,N_14537);
or U17221 (N_17221,N_14936,N_15142);
nor U17222 (N_17222,N_14118,N_14780);
nand U17223 (N_17223,N_14663,N_14126);
or U17224 (N_17224,N_15312,N_15150);
nand U17225 (N_17225,N_15215,N_15957);
nand U17226 (N_17226,N_14972,N_14089);
or U17227 (N_17227,N_14127,N_14876);
nor U17228 (N_17228,N_15543,N_15051);
and U17229 (N_17229,N_14466,N_15435);
and U17230 (N_17230,N_14498,N_14951);
and U17231 (N_17231,N_15897,N_15628);
or U17232 (N_17232,N_14861,N_15861);
xor U17233 (N_17233,N_15693,N_15338);
nor U17234 (N_17234,N_15774,N_14996);
xor U17235 (N_17235,N_15943,N_14046);
and U17236 (N_17236,N_15835,N_15499);
and U17237 (N_17237,N_14139,N_15692);
xnor U17238 (N_17238,N_15862,N_15176);
nand U17239 (N_17239,N_15763,N_14330);
nor U17240 (N_17240,N_14907,N_15576);
and U17241 (N_17241,N_14770,N_15602);
or U17242 (N_17242,N_14733,N_15157);
xnor U17243 (N_17243,N_15677,N_14862);
and U17244 (N_17244,N_15740,N_14810);
nor U17245 (N_17245,N_14572,N_14367);
or U17246 (N_17246,N_14480,N_14262);
nor U17247 (N_17247,N_15658,N_14671);
nor U17248 (N_17248,N_14787,N_15688);
or U17249 (N_17249,N_15974,N_15819);
nor U17250 (N_17250,N_14902,N_15692);
nor U17251 (N_17251,N_14942,N_15103);
and U17252 (N_17252,N_15356,N_14351);
or U17253 (N_17253,N_14976,N_15978);
nand U17254 (N_17254,N_14265,N_15759);
nor U17255 (N_17255,N_14338,N_14814);
nor U17256 (N_17256,N_14317,N_15211);
nor U17257 (N_17257,N_14305,N_14740);
nand U17258 (N_17258,N_14582,N_15969);
nand U17259 (N_17259,N_15689,N_15366);
and U17260 (N_17260,N_14008,N_14220);
and U17261 (N_17261,N_14178,N_14805);
and U17262 (N_17262,N_14098,N_15269);
and U17263 (N_17263,N_15764,N_14682);
or U17264 (N_17264,N_14040,N_14280);
or U17265 (N_17265,N_15486,N_14652);
nor U17266 (N_17266,N_14018,N_15646);
or U17267 (N_17267,N_15304,N_15115);
and U17268 (N_17268,N_14883,N_14405);
nand U17269 (N_17269,N_15589,N_14160);
nand U17270 (N_17270,N_14352,N_15380);
nand U17271 (N_17271,N_14758,N_14262);
and U17272 (N_17272,N_14736,N_15224);
xor U17273 (N_17273,N_14268,N_14400);
or U17274 (N_17274,N_14080,N_14439);
nor U17275 (N_17275,N_14255,N_15001);
and U17276 (N_17276,N_15049,N_15016);
and U17277 (N_17277,N_15507,N_14710);
nand U17278 (N_17278,N_15299,N_15482);
xnor U17279 (N_17279,N_15158,N_15625);
nand U17280 (N_17280,N_14228,N_15661);
and U17281 (N_17281,N_15803,N_14671);
or U17282 (N_17282,N_15002,N_15746);
nand U17283 (N_17283,N_15248,N_15382);
or U17284 (N_17284,N_15396,N_15063);
or U17285 (N_17285,N_15332,N_15367);
nand U17286 (N_17286,N_15958,N_15404);
nor U17287 (N_17287,N_14123,N_14218);
nor U17288 (N_17288,N_15303,N_15486);
nor U17289 (N_17289,N_15013,N_14453);
nand U17290 (N_17290,N_14267,N_14133);
nand U17291 (N_17291,N_14804,N_14590);
nand U17292 (N_17292,N_14791,N_15572);
xor U17293 (N_17293,N_15066,N_15309);
nor U17294 (N_17294,N_14044,N_15574);
or U17295 (N_17295,N_15991,N_15850);
nor U17296 (N_17296,N_14541,N_15522);
or U17297 (N_17297,N_15190,N_15108);
nor U17298 (N_17298,N_15362,N_14280);
nor U17299 (N_17299,N_14777,N_15464);
nand U17300 (N_17300,N_15870,N_15999);
nor U17301 (N_17301,N_15844,N_15210);
nand U17302 (N_17302,N_15436,N_15743);
xor U17303 (N_17303,N_15020,N_15442);
and U17304 (N_17304,N_15188,N_15706);
and U17305 (N_17305,N_14041,N_15875);
or U17306 (N_17306,N_14864,N_15001);
nand U17307 (N_17307,N_15571,N_15256);
and U17308 (N_17308,N_14574,N_14882);
nor U17309 (N_17309,N_14559,N_14804);
nor U17310 (N_17310,N_14382,N_14433);
nor U17311 (N_17311,N_14105,N_14352);
or U17312 (N_17312,N_15151,N_15511);
xnor U17313 (N_17313,N_15094,N_15528);
or U17314 (N_17314,N_15028,N_14460);
nand U17315 (N_17315,N_15010,N_14540);
or U17316 (N_17316,N_15412,N_14503);
nor U17317 (N_17317,N_15729,N_15961);
and U17318 (N_17318,N_15705,N_14907);
or U17319 (N_17319,N_15966,N_15334);
xnor U17320 (N_17320,N_14533,N_14232);
or U17321 (N_17321,N_15058,N_14738);
and U17322 (N_17322,N_14914,N_15408);
nand U17323 (N_17323,N_14908,N_14247);
or U17324 (N_17324,N_15642,N_15342);
and U17325 (N_17325,N_14392,N_15206);
nor U17326 (N_17326,N_14051,N_15147);
nand U17327 (N_17327,N_15618,N_15395);
or U17328 (N_17328,N_15679,N_14517);
nand U17329 (N_17329,N_15487,N_15413);
nand U17330 (N_17330,N_14639,N_15730);
nor U17331 (N_17331,N_14219,N_14589);
or U17332 (N_17332,N_15132,N_15994);
nor U17333 (N_17333,N_15739,N_14076);
nand U17334 (N_17334,N_15033,N_14224);
and U17335 (N_17335,N_14485,N_15934);
nor U17336 (N_17336,N_15137,N_14882);
nand U17337 (N_17337,N_14753,N_15425);
nand U17338 (N_17338,N_15010,N_15823);
nand U17339 (N_17339,N_15641,N_15032);
or U17340 (N_17340,N_15034,N_14118);
nor U17341 (N_17341,N_15120,N_15369);
nand U17342 (N_17342,N_14244,N_14220);
xor U17343 (N_17343,N_14335,N_15609);
xor U17344 (N_17344,N_15244,N_15122);
nor U17345 (N_17345,N_15227,N_14528);
nor U17346 (N_17346,N_15248,N_14395);
nand U17347 (N_17347,N_15054,N_15216);
and U17348 (N_17348,N_14990,N_15586);
or U17349 (N_17349,N_14355,N_14766);
and U17350 (N_17350,N_15411,N_15345);
nor U17351 (N_17351,N_14467,N_15429);
xor U17352 (N_17352,N_15621,N_15123);
nor U17353 (N_17353,N_15420,N_14412);
nand U17354 (N_17354,N_14877,N_15476);
nor U17355 (N_17355,N_15664,N_15359);
xnor U17356 (N_17356,N_14698,N_15363);
nand U17357 (N_17357,N_14022,N_14756);
nand U17358 (N_17358,N_15675,N_15025);
nor U17359 (N_17359,N_15265,N_15402);
and U17360 (N_17360,N_14618,N_15140);
nor U17361 (N_17361,N_14737,N_14328);
and U17362 (N_17362,N_14433,N_14708);
and U17363 (N_17363,N_14480,N_14836);
or U17364 (N_17364,N_14762,N_15274);
nand U17365 (N_17365,N_14527,N_14627);
nand U17366 (N_17366,N_14537,N_14586);
nor U17367 (N_17367,N_15687,N_14803);
nor U17368 (N_17368,N_14917,N_15545);
nand U17369 (N_17369,N_15477,N_14679);
xnor U17370 (N_17370,N_15100,N_14970);
nor U17371 (N_17371,N_15022,N_14827);
nand U17372 (N_17372,N_15708,N_15799);
nor U17373 (N_17373,N_15257,N_15752);
and U17374 (N_17374,N_14050,N_15261);
and U17375 (N_17375,N_14780,N_14646);
and U17376 (N_17376,N_14793,N_14001);
or U17377 (N_17377,N_14840,N_14408);
or U17378 (N_17378,N_15994,N_14306);
nand U17379 (N_17379,N_14955,N_15824);
nand U17380 (N_17380,N_14112,N_14358);
and U17381 (N_17381,N_15004,N_15439);
xor U17382 (N_17382,N_14264,N_14014);
or U17383 (N_17383,N_14154,N_15682);
nand U17384 (N_17384,N_15476,N_14820);
nand U17385 (N_17385,N_14779,N_15362);
and U17386 (N_17386,N_15921,N_15002);
and U17387 (N_17387,N_15191,N_14478);
or U17388 (N_17388,N_15999,N_15891);
nor U17389 (N_17389,N_15722,N_15660);
nand U17390 (N_17390,N_14794,N_15416);
or U17391 (N_17391,N_14445,N_15973);
nor U17392 (N_17392,N_15539,N_14885);
or U17393 (N_17393,N_14999,N_14602);
nor U17394 (N_17394,N_15849,N_15032);
nand U17395 (N_17395,N_14240,N_15566);
and U17396 (N_17396,N_15438,N_15513);
nand U17397 (N_17397,N_14408,N_15981);
nor U17398 (N_17398,N_14526,N_15628);
nor U17399 (N_17399,N_15183,N_14017);
and U17400 (N_17400,N_15890,N_14764);
nor U17401 (N_17401,N_14438,N_15143);
and U17402 (N_17402,N_15546,N_14112);
nor U17403 (N_17403,N_14711,N_15094);
nor U17404 (N_17404,N_15954,N_14249);
or U17405 (N_17405,N_15050,N_14767);
or U17406 (N_17406,N_15158,N_14872);
nor U17407 (N_17407,N_14157,N_15690);
and U17408 (N_17408,N_14079,N_14761);
or U17409 (N_17409,N_14586,N_14764);
nand U17410 (N_17410,N_15470,N_15072);
nor U17411 (N_17411,N_15137,N_14737);
or U17412 (N_17412,N_15427,N_15513);
nand U17413 (N_17413,N_15075,N_15980);
nand U17414 (N_17414,N_15203,N_14429);
and U17415 (N_17415,N_14595,N_15407);
nor U17416 (N_17416,N_14829,N_15964);
xor U17417 (N_17417,N_14482,N_15353);
nor U17418 (N_17418,N_14395,N_14043);
or U17419 (N_17419,N_15117,N_14392);
nor U17420 (N_17420,N_14776,N_15176);
xnor U17421 (N_17421,N_15829,N_14430);
nor U17422 (N_17422,N_14537,N_14776);
nand U17423 (N_17423,N_15962,N_15984);
nand U17424 (N_17424,N_14315,N_14242);
and U17425 (N_17425,N_15441,N_15172);
nor U17426 (N_17426,N_14269,N_14095);
nand U17427 (N_17427,N_15839,N_14018);
nand U17428 (N_17428,N_14144,N_15979);
and U17429 (N_17429,N_14584,N_15049);
and U17430 (N_17430,N_15486,N_14476);
nand U17431 (N_17431,N_14208,N_14071);
xor U17432 (N_17432,N_14303,N_15060);
nor U17433 (N_17433,N_15988,N_14868);
or U17434 (N_17434,N_15251,N_15669);
and U17435 (N_17435,N_15207,N_14197);
and U17436 (N_17436,N_15050,N_14829);
xor U17437 (N_17437,N_14173,N_15605);
nor U17438 (N_17438,N_14596,N_15552);
nand U17439 (N_17439,N_14314,N_14351);
and U17440 (N_17440,N_15859,N_15940);
nor U17441 (N_17441,N_15257,N_14371);
xnor U17442 (N_17442,N_15784,N_15168);
or U17443 (N_17443,N_14815,N_15188);
or U17444 (N_17444,N_15858,N_15743);
or U17445 (N_17445,N_14445,N_15899);
nor U17446 (N_17446,N_15573,N_14100);
nor U17447 (N_17447,N_15091,N_14636);
or U17448 (N_17448,N_14104,N_15181);
or U17449 (N_17449,N_15294,N_15729);
or U17450 (N_17450,N_15517,N_15870);
nor U17451 (N_17451,N_15674,N_14761);
and U17452 (N_17452,N_15999,N_15516);
nand U17453 (N_17453,N_14861,N_15713);
nor U17454 (N_17454,N_14430,N_15553);
nor U17455 (N_17455,N_14895,N_14588);
or U17456 (N_17456,N_15986,N_14383);
and U17457 (N_17457,N_14339,N_15678);
and U17458 (N_17458,N_15745,N_14010);
or U17459 (N_17459,N_14803,N_15284);
nor U17460 (N_17460,N_14072,N_15729);
nor U17461 (N_17461,N_15590,N_14618);
or U17462 (N_17462,N_14409,N_15030);
nand U17463 (N_17463,N_14340,N_15820);
or U17464 (N_17464,N_15344,N_14413);
nand U17465 (N_17465,N_14449,N_15568);
nand U17466 (N_17466,N_14188,N_14003);
or U17467 (N_17467,N_14185,N_14776);
and U17468 (N_17468,N_14340,N_14811);
or U17469 (N_17469,N_14811,N_15812);
nand U17470 (N_17470,N_14478,N_15395);
nor U17471 (N_17471,N_15712,N_14783);
or U17472 (N_17472,N_15123,N_15780);
nor U17473 (N_17473,N_15713,N_14430);
nor U17474 (N_17474,N_15860,N_14681);
and U17475 (N_17475,N_14088,N_15505);
nor U17476 (N_17476,N_15954,N_15808);
or U17477 (N_17477,N_15130,N_14832);
nor U17478 (N_17478,N_15728,N_14450);
nor U17479 (N_17479,N_14098,N_15766);
or U17480 (N_17480,N_14048,N_14114);
nor U17481 (N_17481,N_15884,N_14280);
and U17482 (N_17482,N_14298,N_15764);
nand U17483 (N_17483,N_15177,N_15440);
nand U17484 (N_17484,N_14218,N_14530);
and U17485 (N_17485,N_14215,N_15946);
and U17486 (N_17486,N_15822,N_15837);
nor U17487 (N_17487,N_14746,N_15979);
or U17488 (N_17488,N_15592,N_14308);
nor U17489 (N_17489,N_14073,N_15042);
nand U17490 (N_17490,N_15925,N_15570);
nor U17491 (N_17491,N_15583,N_15718);
and U17492 (N_17492,N_15468,N_14136);
nand U17493 (N_17493,N_15065,N_15286);
nor U17494 (N_17494,N_15407,N_14089);
or U17495 (N_17495,N_14751,N_15614);
nand U17496 (N_17496,N_15116,N_15039);
nand U17497 (N_17497,N_14193,N_15572);
nor U17498 (N_17498,N_14541,N_14902);
or U17499 (N_17499,N_14606,N_14832);
or U17500 (N_17500,N_14852,N_14561);
nor U17501 (N_17501,N_15246,N_15582);
nand U17502 (N_17502,N_15823,N_15928);
or U17503 (N_17503,N_15480,N_14849);
nand U17504 (N_17504,N_14842,N_15922);
nor U17505 (N_17505,N_14790,N_15030);
and U17506 (N_17506,N_14552,N_15221);
and U17507 (N_17507,N_15924,N_15932);
nand U17508 (N_17508,N_14854,N_15444);
and U17509 (N_17509,N_14838,N_15313);
nor U17510 (N_17510,N_15669,N_14677);
nor U17511 (N_17511,N_14242,N_15718);
nand U17512 (N_17512,N_15045,N_14467);
xor U17513 (N_17513,N_14117,N_14477);
nand U17514 (N_17514,N_14440,N_14034);
xnor U17515 (N_17515,N_15044,N_14881);
or U17516 (N_17516,N_15245,N_14010);
and U17517 (N_17517,N_15099,N_15817);
or U17518 (N_17518,N_14125,N_15202);
xor U17519 (N_17519,N_15477,N_15113);
or U17520 (N_17520,N_15683,N_15666);
nand U17521 (N_17521,N_15013,N_15563);
and U17522 (N_17522,N_15335,N_15889);
and U17523 (N_17523,N_15819,N_14829);
nand U17524 (N_17524,N_15517,N_14860);
and U17525 (N_17525,N_15082,N_14315);
and U17526 (N_17526,N_14839,N_15138);
nand U17527 (N_17527,N_15904,N_15936);
or U17528 (N_17528,N_15947,N_14573);
and U17529 (N_17529,N_15756,N_14521);
and U17530 (N_17530,N_14571,N_15388);
nor U17531 (N_17531,N_14060,N_15454);
xnor U17532 (N_17532,N_14056,N_15259);
and U17533 (N_17533,N_14302,N_14927);
and U17534 (N_17534,N_15064,N_15498);
nor U17535 (N_17535,N_15891,N_15565);
and U17536 (N_17536,N_15432,N_14650);
or U17537 (N_17537,N_14039,N_14492);
nand U17538 (N_17538,N_14410,N_15928);
nor U17539 (N_17539,N_15992,N_14187);
or U17540 (N_17540,N_14933,N_14197);
nand U17541 (N_17541,N_14948,N_15866);
nor U17542 (N_17542,N_15018,N_14621);
nand U17543 (N_17543,N_15432,N_14514);
xnor U17544 (N_17544,N_15097,N_14343);
and U17545 (N_17545,N_14738,N_14675);
xor U17546 (N_17546,N_14209,N_14094);
nor U17547 (N_17547,N_15157,N_15489);
and U17548 (N_17548,N_14096,N_14004);
nor U17549 (N_17549,N_14865,N_15226);
nand U17550 (N_17550,N_15951,N_14286);
and U17551 (N_17551,N_15899,N_14950);
nor U17552 (N_17552,N_15948,N_14572);
nor U17553 (N_17553,N_15137,N_14045);
or U17554 (N_17554,N_14369,N_15068);
nor U17555 (N_17555,N_15708,N_15779);
nand U17556 (N_17556,N_14951,N_14980);
and U17557 (N_17557,N_14887,N_14680);
or U17558 (N_17558,N_15039,N_15609);
or U17559 (N_17559,N_14741,N_15913);
or U17560 (N_17560,N_14437,N_15792);
or U17561 (N_17561,N_15069,N_15950);
nand U17562 (N_17562,N_15647,N_15198);
or U17563 (N_17563,N_15625,N_15511);
nand U17564 (N_17564,N_15336,N_14317);
and U17565 (N_17565,N_15357,N_15770);
nor U17566 (N_17566,N_14056,N_14603);
and U17567 (N_17567,N_15423,N_14076);
nor U17568 (N_17568,N_14969,N_14205);
nand U17569 (N_17569,N_14417,N_15409);
nand U17570 (N_17570,N_14225,N_15121);
nand U17571 (N_17571,N_14991,N_14019);
and U17572 (N_17572,N_14565,N_14927);
or U17573 (N_17573,N_15087,N_14081);
nor U17574 (N_17574,N_15584,N_14713);
nand U17575 (N_17575,N_15863,N_15740);
and U17576 (N_17576,N_14965,N_14334);
and U17577 (N_17577,N_14551,N_15270);
or U17578 (N_17578,N_14295,N_15678);
nor U17579 (N_17579,N_15385,N_14931);
xnor U17580 (N_17580,N_15160,N_15688);
nor U17581 (N_17581,N_15893,N_14701);
and U17582 (N_17582,N_15259,N_14063);
or U17583 (N_17583,N_14688,N_14068);
and U17584 (N_17584,N_15858,N_14583);
and U17585 (N_17585,N_14530,N_14001);
or U17586 (N_17586,N_14547,N_15352);
nor U17587 (N_17587,N_15287,N_14386);
nor U17588 (N_17588,N_15423,N_15923);
xor U17589 (N_17589,N_14045,N_15129);
nor U17590 (N_17590,N_14408,N_14223);
nand U17591 (N_17591,N_14960,N_14891);
nand U17592 (N_17592,N_14171,N_15312);
and U17593 (N_17593,N_15463,N_15500);
and U17594 (N_17594,N_15601,N_15369);
or U17595 (N_17595,N_15510,N_14901);
or U17596 (N_17596,N_14229,N_15396);
nor U17597 (N_17597,N_15682,N_15464);
and U17598 (N_17598,N_15731,N_15711);
or U17599 (N_17599,N_14819,N_14390);
or U17600 (N_17600,N_14768,N_14516);
and U17601 (N_17601,N_14124,N_14643);
or U17602 (N_17602,N_15378,N_15732);
or U17603 (N_17603,N_15292,N_14939);
nor U17604 (N_17604,N_14348,N_15154);
and U17605 (N_17605,N_14439,N_15619);
nand U17606 (N_17606,N_15407,N_14869);
xnor U17607 (N_17607,N_15875,N_15905);
xnor U17608 (N_17608,N_14006,N_15283);
nand U17609 (N_17609,N_15711,N_15118);
and U17610 (N_17610,N_14880,N_14405);
nor U17611 (N_17611,N_15853,N_15380);
nor U17612 (N_17612,N_14425,N_15698);
xnor U17613 (N_17613,N_15266,N_14171);
xnor U17614 (N_17614,N_15441,N_14137);
nand U17615 (N_17615,N_14623,N_15847);
nor U17616 (N_17616,N_15372,N_14010);
and U17617 (N_17617,N_15273,N_14725);
and U17618 (N_17618,N_15274,N_15027);
and U17619 (N_17619,N_15848,N_14963);
nor U17620 (N_17620,N_15147,N_15881);
nand U17621 (N_17621,N_15443,N_14992);
and U17622 (N_17622,N_15821,N_15036);
nand U17623 (N_17623,N_14942,N_14844);
nor U17624 (N_17624,N_15441,N_15482);
and U17625 (N_17625,N_15188,N_14276);
and U17626 (N_17626,N_14053,N_14259);
nand U17627 (N_17627,N_14788,N_14833);
nor U17628 (N_17628,N_14651,N_15405);
nor U17629 (N_17629,N_14661,N_14608);
nor U17630 (N_17630,N_15200,N_15355);
or U17631 (N_17631,N_15302,N_15794);
or U17632 (N_17632,N_14915,N_15432);
nor U17633 (N_17633,N_14058,N_15642);
and U17634 (N_17634,N_14177,N_15912);
and U17635 (N_17635,N_15448,N_15392);
or U17636 (N_17636,N_15419,N_14481);
nand U17637 (N_17637,N_14859,N_14929);
and U17638 (N_17638,N_14679,N_15325);
nand U17639 (N_17639,N_15391,N_14828);
or U17640 (N_17640,N_14018,N_15549);
or U17641 (N_17641,N_14050,N_15595);
and U17642 (N_17642,N_14105,N_14074);
nand U17643 (N_17643,N_14051,N_15671);
xor U17644 (N_17644,N_15342,N_15645);
xor U17645 (N_17645,N_14781,N_15868);
nor U17646 (N_17646,N_15414,N_14729);
or U17647 (N_17647,N_15297,N_15825);
nand U17648 (N_17648,N_15477,N_14576);
nand U17649 (N_17649,N_14237,N_15468);
or U17650 (N_17650,N_14205,N_15744);
and U17651 (N_17651,N_15420,N_14306);
nor U17652 (N_17652,N_15736,N_15027);
xnor U17653 (N_17653,N_14245,N_14686);
or U17654 (N_17654,N_15777,N_14843);
nor U17655 (N_17655,N_15774,N_15578);
nand U17656 (N_17656,N_14325,N_15293);
nand U17657 (N_17657,N_15835,N_15915);
nand U17658 (N_17658,N_14418,N_14997);
nor U17659 (N_17659,N_14774,N_14682);
nor U17660 (N_17660,N_14250,N_14179);
nand U17661 (N_17661,N_15090,N_14616);
nor U17662 (N_17662,N_14882,N_15063);
and U17663 (N_17663,N_14631,N_14123);
nand U17664 (N_17664,N_15733,N_15049);
xnor U17665 (N_17665,N_14382,N_14747);
and U17666 (N_17666,N_14704,N_14745);
nand U17667 (N_17667,N_15531,N_15854);
or U17668 (N_17668,N_15013,N_15392);
nand U17669 (N_17669,N_14131,N_15228);
xor U17670 (N_17670,N_14542,N_14055);
xor U17671 (N_17671,N_15091,N_14198);
or U17672 (N_17672,N_14770,N_14718);
nor U17673 (N_17673,N_15514,N_15298);
nand U17674 (N_17674,N_15958,N_15941);
nor U17675 (N_17675,N_15757,N_15507);
and U17676 (N_17676,N_15447,N_14592);
nor U17677 (N_17677,N_15139,N_15244);
nand U17678 (N_17678,N_14020,N_14575);
and U17679 (N_17679,N_14771,N_14784);
nand U17680 (N_17680,N_14447,N_15831);
nand U17681 (N_17681,N_14027,N_14520);
nor U17682 (N_17682,N_14227,N_15683);
or U17683 (N_17683,N_15302,N_14926);
and U17684 (N_17684,N_15890,N_15587);
or U17685 (N_17685,N_14595,N_15944);
xor U17686 (N_17686,N_15946,N_14020);
nor U17687 (N_17687,N_15434,N_14000);
or U17688 (N_17688,N_15225,N_15845);
nor U17689 (N_17689,N_14156,N_14832);
and U17690 (N_17690,N_15988,N_15513);
nor U17691 (N_17691,N_15739,N_15246);
or U17692 (N_17692,N_14077,N_14751);
or U17693 (N_17693,N_15697,N_14824);
nor U17694 (N_17694,N_15518,N_14522);
nand U17695 (N_17695,N_14239,N_14700);
xnor U17696 (N_17696,N_15277,N_15147);
and U17697 (N_17697,N_15875,N_14502);
or U17698 (N_17698,N_15899,N_15887);
or U17699 (N_17699,N_15502,N_15622);
nand U17700 (N_17700,N_14223,N_14805);
and U17701 (N_17701,N_15885,N_15910);
or U17702 (N_17702,N_14150,N_15748);
nand U17703 (N_17703,N_14673,N_15721);
or U17704 (N_17704,N_15091,N_15998);
nand U17705 (N_17705,N_15546,N_15698);
nand U17706 (N_17706,N_15378,N_15362);
nand U17707 (N_17707,N_14678,N_15714);
nand U17708 (N_17708,N_15919,N_15177);
xor U17709 (N_17709,N_15629,N_15083);
xor U17710 (N_17710,N_15503,N_15341);
nor U17711 (N_17711,N_14414,N_15015);
and U17712 (N_17712,N_14190,N_14195);
and U17713 (N_17713,N_15795,N_15509);
nor U17714 (N_17714,N_15292,N_14128);
xnor U17715 (N_17715,N_15208,N_14715);
nor U17716 (N_17716,N_14601,N_15110);
nand U17717 (N_17717,N_15760,N_15913);
or U17718 (N_17718,N_15618,N_15164);
nand U17719 (N_17719,N_15821,N_14640);
nand U17720 (N_17720,N_14582,N_14058);
nor U17721 (N_17721,N_14371,N_14955);
xor U17722 (N_17722,N_15916,N_14482);
xnor U17723 (N_17723,N_14089,N_15751);
nand U17724 (N_17724,N_15990,N_15694);
xor U17725 (N_17725,N_14437,N_15617);
or U17726 (N_17726,N_15294,N_14025);
nor U17727 (N_17727,N_14430,N_14827);
or U17728 (N_17728,N_14048,N_15252);
xnor U17729 (N_17729,N_15412,N_14469);
nand U17730 (N_17730,N_15969,N_14416);
nor U17731 (N_17731,N_15524,N_14536);
nor U17732 (N_17732,N_15101,N_14971);
or U17733 (N_17733,N_14256,N_14679);
or U17734 (N_17734,N_15954,N_15113);
nand U17735 (N_17735,N_14528,N_14027);
nand U17736 (N_17736,N_15005,N_14814);
nand U17737 (N_17737,N_15445,N_15198);
nand U17738 (N_17738,N_14429,N_14389);
or U17739 (N_17739,N_15868,N_14273);
nand U17740 (N_17740,N_15939,N_14668);
nor U17741 (N_17741,N_14527,N_15788);
nor U17742 (N_17742,N_15801,N_15762);
or U17743 (N_17743,N_15377,N_14532);
nand U17744 (N_17744,N_14514,N_14171);
nand U17745 (N_17745,N_14642,N_15945);
or U17746 (N_17746,N_14213,N_14066);
nand U17747 (N_17747,N_14243,N_15585);
and U17748 (N_17748,N_15677,N_15942);
and U17749 (N_17749,N_15311,N_14571);
or U17750 (N_17750,N_15165,N_15992);
nor U17751 (N_17751,N_14258,N_15236);
nand U17752 (N_17752,N_14973,N_15070);
and U17753 (N_17753,N_15217,N_14445);
or U17754 (N_17754,N_14884,N_14481);
xor U17755 (N_17755,N_14081,N_15341);
xnor U17756 (N_17756,N_14650,N_15399);
and U17757 (N_17757,N_15915,N_14045);
and U17758 (N_17758,N_15950,N_15866);
xor U17759 (N_17759,N_14687,N_15152);
nor U17760 (N_17760,N_14604,N_15599);
nor U17761 (N_17761,N_14160,N_14964);
nand U17762 (N_17762,N_15371,N_15594);
nand U17763 (N_17763,N_15988,N_14469);
nor U17764 (N_17764,N_14316,N_15102);
nor U17765 (N_17765,N_14114,N_14035);
and U17766 (N_17766,N_15985,N_15350);
or U17767 (N_17767,N_14896,N_14814);
or U17768 (N_17768,N_15593,N_14969);
xnor U17769 (N_17769,N_14211,N_14048);
and U17770 (N_17770,N_14751,N_14604);
nand U17771 (N_17771,N_14723,N_14895);
nand U17772 (N_17772,N_15697,N_15630);
nand U17773 (N_17773,N_15962,N_15653);
nor U17774 (N_17774,N_15036,N_15928);
nor U17775 (N_17775,N_14916,N_15204);
nand U17776 (N_17776,N_14068,N_14712);
nor U17777 (N_17777,N_15923,N_15502);
nand U17778 (N_17778,N_15363,N_14554);
and U17779 (N_17779,N_15265,N_15009);
xor U17780 (N_17780,N_14583,N_15427);
or U17781 (N_17781,N_14545,N_14749);
xor U17782 (N_17782,N_14648,N_14088);
xnor U17783 (N_17783,N_14513,N_14664);
or U17784 (N_17784,N_15154,N_14147);
or U17785 (N_17785,N_14284,N_15078);
and U17786 (N_17786,N_14804,N_15226);
nor U17787 (N_17787,N_14303,N_15756);
xor U17788 (N_17788,N_15218,N_15883);
nand U17789 (N_17789,N_14504,N_15048);
and U17790 (N_17790,N_14308,N_15927);
nor U17791 (N_17791,N_14172,N_15750);
nor U17792 (N_17792,N_15700,N_15126);
nor U17793 (N_17793,N_15899,N_15838);
xnor U17794 (N_17794,N_15090,N_15709);
and U17795 (N_17795,N_15360,N_15839);
nand U17796 (N_17796,N_15955,N_15824);
nor U17797 (N_17797,N_14756,N_15449);
nor U17798 (N_17798,N_15721,N_14578);
and U17799 (N_17799,N_15739,N_15740);
nor U17800 (N_17800,N_15152,N_15084);
nor U17801 (N_17801,N_15567,N_14654);
nor U17802 (N_17802,N_14228,N_15785);
xor U17803 (N_17803,N_15551,N_14125);
nor U17804 (N_17804,N_15736,N_15236);
or U17805 (N_17805,N_15105,N_15771);
nand U17806 (N_17806,N_15090,N_15574);
xnor U17807 (N_17807,N_15090,N_15930);
and U17808 (N_17808,N_15738,N_14848);
or U17809 (N_17809,N_14426,N_15534);
and U17810 (N_17810,N_15712,N_15650);
and U17811 (N_17811,N_15208,N_15785);
nor U17812 (N_17812,N_15460,N_15652);
nor U17813 (N_17813,N_15466,N_14016);
nor U17814 (N_17814,N_14805,N_15379);
xnor U17815 (N_17815,N_14220,N_14793);
nand U17816 (N_17816,N_15978,N_14032);
nor U17817 (N_17817,N_14028,N_15709);
and U17818 (N_17818,N_15308,N_14577);
or U17819 (N_17819,N_14134,N_14356);
nand U17820 (N_17820,N_14207,N_14305);
or U17821 (N_17821,N_15728,N_14018);
and U17822 (N_17822,N_15840,N_15367);
or U17823 (N_17823,N_14878,N_14964);
nand U17824 (N_17824,N_14213,N_15444);
and U17825 (N_17825,N_14128,N_15995);
nor U17826 (N_17826,N_14047,N_14505);
and U17827 (N_17827,N_15887,N_14550);
nand U17828 (N_17828,N_14132,N_15451);
xor U17829 (N_17829,N_15684,N_14369);
or U17830 (N_17830,N_14499,N_15681);
nand U17831 (N_17831,N_14939,N_14891);
nand U17832 (N_17832,N_14668,N_15460);
xnor U17833 (N_17833,N_15980,N_14498);
and U17834 (N_17834,N_14188,N_14424);
and U17835 (N_17835,N_14545,N_15231);
nor U17836 (N_17836,N_15468,N_14289);
nor U17837 (N_17837,N_15321,N_14386);
nand U17838 (N_17838,N_14969,N_14362);
nor U17839 (N_17839,N_14860,N_14507);
nand U17840 (N_17840,N_15297,N_15464);
xnor U17841 (N_17841,N_15001,N_14893);
nand U17842 (N_17842,N_15843,N_15614);
nand U17843 (N_17843,N_15460,N_14717);
and U17844 (N_17844,N_15180,N_14295);
and U17845 (N_17845,N_14715,N_15610);
xnor U17846 (N_17846,N_14662,N_15088);
nand U17847 (N_17847,N_14176,N_15587);
and U17848 (N_17848,N_15920,N_15501);
nand U17849 (N_17849,N_14386,N_15657);
xnor U17850 (N_17850,N_14222,N_15741);
nor U17851 (N_17851,N_14596,N_15263);
nor U17852 (N_17852,N_15986,N_14115);
nor U17853 (N_17853,N_14045,N_14881);
nand U17854 (N_17854,N_15373,N_14431);
nor U17855 (N_17855,N_14631,N_15670);
nand U17856 (N_17856,N_15384,N_14730);
nor U17857 (N_17857,N_14361,N_14391);
nor U17858 (N_17858,N_15001,N_14687);
nand U17859 (N_17859,N_15928,N_15126);
nor U17860 (N_17860,N_15550,N_15942);
nand U17861 (N_17861,N_14616,N_15107);
or U17862 (N_17862,N_15621,N_14283);
or U17863 (N_17863,N_14502,N_15572);
and U17864 (N_17864,N_14658,N_15898);
xnor U17865 (N_17865,N_14269,N_14240);
nand U17866 (N_17866,N_15718,N_14537);
or U17867 (N_17867,N_14490,N_14023);
and U17868 (N_17868,N_14953,N_14056);
nand U17869 (N_17869,N_15179,N_15426);
or U17870 (N_17870,N_14225,N_14285);
and U17871 (N_17871,N_14273,N_15683);
nor U17872 (N_17872,N_14057,N_14812);
nor U17873 (N_17873,N_15781,N_15144);
xnor U17874 (N_17874,N_14384,N_15939);
and U17875 (N_17875,N_15497,N_15733);
and U17876 (N_17876,N_15812,N_15465);
or U17877 (N_17877,N_14400,N_15290);
and U17878 (N_17878,N_14459,N_15228);
nand U17879 (N_17879,N_14326,N_15862);
and U17880 (N_17880,N_15338,N_14087);
xnor U17881 (N_17881,N_15984,N_15333);
or U17882 (N_17882,N_14345,N_15858);
or U17883 (N_17883,N_15247,N_14420);
and U17884 (N_17884,N_15507,N_14517);
or U17885 (N_17885,N_14315,N_14873);
nand U17886 (N_17886,N_14505,N_14758);
or U17887 (N_17887,N_15096,N_14582);
or U17888 (N_17888,N_15527,N_15899);
or U17889 (N_17889,N_15411,N_15985);
xor U17890 (N_17890,N_14517,N_15688);
nand U17891 (N_17891,N_15307,N_14948);
nor U17892 (N_17892,N_15117,N_14811);
nor U17893 (N_17893,N_15286,N_15351);
nand U17894 (N_17894,N_14848,N_15548);
nand U17895 (N_17895,N_14027,N_15655);
or U17896 (N_17896,N_15827,N_15453);
and U17897 (N_17897,N_15333,N_14398);
nor U17898 (N_17898,N_14766,N_15495);
or U17899 (N_17899,N_14864,N_15780);
xnor U17900 (N_17900,N_15388,N_14222);
nor U17901 (N_17901,N_14241,N_14247);
and U17902 (N_17902,N_14561,N_14219);
or U17903 (N_17903,N_14151,N_14352);
nand U17904 (N_17904,N_14161,N_15576);
or U17905 (N_17905,N_14381,N_14595);
and U17906 (N_17906,N_14304,N_15158);
and U17907 (N_17907,N_14184,N_14933);
nand U17908 (N_17908,N_15344,N_15224);
or U17909 (N_17909,N_14318,N_15512);
nor U17910 (N_17910,N_15623,N_15358);
or U17911 (N_17911,N_15944,N_15965);
and U17912 (N_17912,N_15117,N_15669);
nor U17913 (N_17913,N_15030,N_15252);
or U17914 (N_17914,N_14878,N_15133);
or U17915 (N_17915,N_15463,N_15321);
and U17916 (N_17916,N_14904,N_15920);
nand U17917 (N_17917,N_14601,N_15884);
or U17918 (N_17918,N_15448,N_14880);
nor U17919 (N_17919,N_15708,N_14224);
nand U17920 (N_17920,N_15219,N_14634);
nand U17921 (N_17921,N_15423,N_15599);
nand U17922 (N_17922,N_14436,N_14328);
nor U17923 (N_17923,N_14909,N_15318);
or U17924 (N_17924,N_15237,N_14825);
nor U17925 (N_17925,N_14945,N_15401);
and U17926 (N_17926,N_15210,N_14807);
or U17927 (N_17927,N_15633,N_15483);
or U17928 (N_17928,N_14197,N_14593);
nor U17929 (N_17929,N_15768,N_14692);
xor U17930 (N_17930,N_15427,N_15108);
and U17931 (N_17931,N_14787,N_15892);
nor U17932 (N_17932,N_15502,N_15808);
and U17933 (N_17933,N_15113,N_14561);
nand U17934 (N_17934,N_15927,N_15027);
xnor U17935 (N_17935,N_14931,N_14878);
xnor U17936 (N_17936,N_15079,N_14765);
nor U17937 (N_17937,N_15114,N_14287);
nand U17938 (N_17938,N_14421,N_15950);
and U17939 (N_17939,N_14471,N_15108);
nand U17940 (N_17940,N_14501,N_14491);
nand U17941 (N_17941,N_15264,N_14591);
or U17942 (N_17942,N_14113,N_14567);
nor U17943 (N_17943,N_15729,N_14193);
nor U17944 (N_17944,N_14662,N_15007);
nand U17945 (N_17945,N_14498,N_15986);
nor U17946 (N_17946,N_14827,N_14376);
or U17947 (N_17947,N_15616,N_14567);
nor U17948 (N_17948,N_14428,N_15725);
nor U17949 (N_17949,N_15489,N_14111);
xnor U17950 (N_17950,N_15269,N_15183);
or U17951 (N_17951,N_15992,N_14567);
nand U17952 (N_17952,N_15214,N_14310);
nor U17953 (N_17953,N_14699,N_14357);
or U17954 (N_17954,N_15702,N_15736);
nand U17955 (N_17955,N_15409,N_15422);
and U17956 (N_17956,N_14577,N_15440);
and U17957 (N_17957,N_14725,N_15789);
and U17958 (N_17958,N_14447,N_14327);
and U17959 (N_17959,N_15699,N_14938);
nand U17960 (N_17960,N_14626,N_14262);
nand U17961 (N_17961,N_14916,N_15738);
or U17962 (N_17962,N_15793,N_14512);
nor U17963 (N_17963,N_14380,N_14114);
nor U17964 (N_17964,N_15550,N_14652);
or U17965 (N_17965,N_14931,N_15487);
or U17966 (N_17966,N_14595,N_14376);
and U17967 (N_17967,N_15123,N_15474);
xor U17968 (N_17968,N_14953,N_14315);
or U17969 (N_17969,N_15283,N_15104);
or U17970 (N_17970,N_14302,N_15287);
or U17971 (N_17971,N_15017,N_15359);
nand U17972 (N_17972,N_14878,N_14560);
nand U17973 (N_17973,N_15065,N_14668);
nand U17974 (N_17974,N_14291,N_14051);
or U17975 (N_17975,N_15097,N_14749);
or U17976 (N_17976,N_15751,N_14419);
nor U17977 (N_17977,N_15310,N_15739);
and U17978 (N_17978,N_14711,N_14034);
nor U17979 (N_17979,N_15077,N_14340);
nor U17980 (N_17980,N_14540,N_14222);
or U17981 (N_17981,N_14209,N_15798);
xnor U17982 (N_17982,N_14761,N_14329);
xnor U17983 (N_17983,N_14496,N_14987);
nand U17984 (N_17984,N_15645,N_15083);
nand U17985 (N_17985,N_15365,N_14643);
nor U17986 (N_17986,N_15014,N_14201);
nand U17987 (N_17987,N_14568,N_15138);
nand U17988 (N_17988,N_15681,N_15787);
nor U17989 (N_17989,N_15546,N_15815);
and U17990 (N_17990,N_14919,N_15025);
and U17991 (N_17991,N_14443,N_14598);
nor U17992 (N_17992,N_14470,N_15101);
and U17993 (N_17993,N_15709,N_15374);
nor U17994 (N_17994,N_15495,N_15852);
nor U17995 (N_17995,N_15739,N_14613);
nand U17996 (N_17996,N_15059,N_14913);
nand U17997 (N_17997,N_14804,N_14245);
nand U17998 (N_17998,N_15613,N_15516);
or U17999 (N_17999,N_14653,N_15070);
nor U18000 (N_18000,N_16112,N_17692);
or U18001 (N_18001,N_17919,N_16714);
and U18002 (N_18002,N_17854,N_16424);
nor U18003 (N_18003,N_16785,N_16365);
and U18004 (N_18004,N_17670,N_16308);
and U18005 (N_18005,N_17950,N_16091);
or U18006 (N_18006,N_16184,N_17767);
or U18007 (N_18007,N_17113,N_16322);
nand U18008 (N_18008,N_16875,N_16569);
nand U18009 (N_18009,N_16800,N_17313);
and U18010 (N_18010,N_17367,N_17247);
or U18011 (N_18011,N_17745,N_17957);
nor U18012 (N_18012,N_17798,N_17475);
nand U18013 (N_18013,N_16392,N_16903);
xnor U18014 (N_18014,N_16044,N_17938);
nand U18015 (N_18015,N_17254,N_16481);
nor U18016 (N_18016,N_16774,N_17080);
and U18017 (N_18017,N_16966,N_17599);
nand U18018 (N_18018,N_16218,N_17374);
xnor U18019 (N_18019,N_17872,N_17699);
nor U18020 (N_18020,N_16255,N_17473);
or U18021 (N_18021,N_16089,N_17811);
xnor U18022 (N_18022,N_16069,N_16414);
or U18023 (N_18023,N_17366,N_16085);
xnor U18024 (N_18024,N_16252,N_16137);
and U18025 (N_18025,N_17742,N_17657);
nor U18026 (N_18026,N_17708,N_17306);
xnor U18027 (N_18027,N_16542,N_16355);
nor U18028 (N_18028,N_16861,N_16822);
or U18029 (N_18029,N_16663,N_16843);
and U18030 (N_18030,N_17283,N_17329);
nand U18031 (N_18031,N_17216,N_17459);
nor U18032 (N_18032,N_16844,N_16659);
nand U18033 (N_18033,N_17842,N_16752);
nand U18034 (N_18034,N_17073,N_17969);
nor U18035 (N_18035,N_16307,N_16235);
and U18036 (N_18036,N_17922,N_17646);
or U18037 (N_18037,N_17365,N_17307);
nand U18038 (N_18038,N_17241,N_17725);
or U18039 (N_18039,N_16905,N_17397);
nand U18040 (N_18040,N_17839,N_17350);
or U18041 (N_18041,N_17300,N_17522);
nand U18042 (N_18042,N_16304,N_17487);
and U18043 (N_18043,N_17823,N_16129);
nor U18044 (N_18044,N_17163,N_17213);
or U18045 (N_18045,N_16500,N_16934);
and U18046 (N_18046,N_16581,N_17391);
nor U18047 (N_18047,N_16501,N_16380);
or U18048 (N_18048,N_17244,N_16865);
nor U18049 (N_18049,N_16601,N_17086);
nor U18050 (N_18050,N_17743,N_17735);
xnor U18051 (N_18051,N_16758,N_17311);
xor U18052 (N_18052,N_16283,N_16003);
or U18053 (N_18053,N_17220,N_17333);
nand U18054 (N_18054,N_17828,N_16570);
xnor U18055 (N_18055,N_17824,N_16797);
nor U18056 (N_18056,N_16909,N_16401);
or U18057 (N_18057,N_16121,N_16262);
nand U18058 (N_18058,N_16995,N_16383);
or U18059 (N_18059,N_17578,N_17211);
and U18060 (N_18060,N_16344,N_17291);
and U18061 (N_18061,N_16202,N_17998);
or U18062 (N_18062,N_16832,N_17382);
or U18063 (N_18063,N_17036,N_17643);
nand U18064 (N_18064,N_17664,N_16454);
and U18065 (N_18065,N_17790,N_17188);
nand U18066 (N_18066,N_17323,N_17848);
or U18067 (N_18067,N_16607,N_17486);
nor U18068 (N_18068,N_17056,N_16884);
and U18069 (N_18069,N_16827,N_17935);
xnor U18070 (N_18070,N_16437,N_17519);
xnor U18071 (N_18071,N_16866,N_16650);
and U18072 (N_18072,N_16075,N_17668);
nand U18073 (N_18073,N_17422,N_17704);
nor U18074 (N_18074,N_16559,N_16712);
xnor U18075 (N_18075,N_17035,N_16362);
and U18076 (N_18076,N_17444,N_16405);
or U18077 (N_18077,N_16166,N_16094);
nor U18078 (N_18078,N_17673,N_16889);
and U18079 (N_18079,N_17736,N_17066);
or U18080 (N_18080,N_17057,N_17165);
or U18081 (N_18081,N_16158,N_17024);
nand U18082 (N_18082,N_17787,N_16951);
nor U18083 (N_18083,N_16942,N_17625);
or U18084 (N_18084,N_16710,N_16703);
nor U18085 (N_18085,N_17503,N_17794);
nand U18086 (N_18086,N_17343,N_16653);
xnor U18087 (N_18087,N_17852,N_17504);
or U18088 (N_18088,N_16023,N_16916);
nor U18089 (N_18089,N_16492,N_17301);
or U18090 (N_18090,N_17455,N_17224);
or U18091 (N_18091,N_17807,N_16807);
nand U18092 (N_18092,N_17732,N_16212);
xor U18093 (N_18093,N_16289,N_17903);
nand U18094 (N_18094,N_17543,N_16810);
and U18095 (N_18095,N_17063,N_17602);
nor U18096 (N_18096,N_16791,N_16005);
nand U18097 (N_18097,N_16987,N_17078);
and U18098 (N_18098,N_16247,N_17218);
nor U18099 (N_18099,N_16118,N_16537);
nor U18100 (N_18100,N_17184,N_16461);
or U18101 (N_18101,N_16669,N_16136);
nand U18102 (N_18102,N_17143,N_17279);
nand U18103 (N_18103,N_16447,N_17123);
and U18104 (N_18104,N_16314,N_17262);
nor U18105 (N_18105,N_16275,N_17437);
nor U18106 (N_18106,N_17644,N_17114);
nand U18107 (N_18107,N_17014,N_16020);
nand U18108 (N_18108,N_17744,N_17820);
or U18109 (N_18109,N_16319,N_16972);
nand U18110 (N_18110,N_17288,N_16170);
and U18111 (N_18111,N_17714,N_16046);
nor U18112 (N_18112,N_17545,N_17172);
and U18113 (N_18113,N_16002,N_16572);
and U18114 (N_18114,N_17116,N_16346);
or U18115 (N_18115,N_16818,N_17492);
or U18116 (N_18116,N_16065,N_16610);
nand U18117 (N_18117,N_17517,N_16926);
nor U18118 (N_18118,N_17145,N_16169);
nor U18119 (N_18119,N_17941,N_17748);
nand U18120 (N_18120,N_16410,N_16468);
or U18121 (N_18121,N_16297,N_17430);
xor U18122 (N_18122,N_17840,N_17393);
and U18123 (N_18123,N_17337,N_17104);
nand U18124 (N_18124,N_16970,N_16193);
nor U18125 (N_18125,N_17128,N_16991);
or U18126 (N_18126,N_16755,N_16960);
and U18127 (N_18127,N_16302,N_16589);
nand U18128 (N_18128,N_16620,N_16736);
and U18129 (N_18129,N_16512,N_16498);
nand U18130 (N_18130,N_17701,N_17727);
nor U18131 (N_18131,N_16740,N_17565);
and U18132 (N_18132,N_17791,N_17821);
nand U18133 (N_18133,N_16667,N_17152);
nand U18134 (N_18134,N_17650,N_17419);
or U18135 (N_18135,N_16415,N_16210);
nand U18136 (N_18136,N_17574,N_17045);
or U18137 (N_18137,N_17896,N_16323);
and U18138 (N_18138,N_16338,N_16787);
nor U18139 (N_18139,N_16370,N_16382);
or U18140 (N_18140,N_17720,N_16681);
and U18141 (N_18141,N_17912,N_16716);
nand U18142 (N_18142,N_16938,N_17524);
or U18143 (N_18143,N_16575,N_17191);
nor U18144 (N_18144,N_17022,N_16566);
nor U18145 (N_18145,N_16761,N_17827);
nand U18146 (N_18146,N_16001,N_17619);
or U18147 (N_18147,N_17551,N_17906);
or U18148 (N_18148,N_16376,N_17067);
nand U18149 (N_18149,N_17582,N_17598);
and U18150 (N_18150,N_17434,N_16041);
xor U18151 (N_18151,N_16826,N_17411);
nand U18152 (N_18152,N_16749,N_17955);
or U18153 (N_18153,N_17031,N_17992);
or U18154 (N_18154,N_17554,N_17200);
and U18155 (N_18155,N_16604,N_17100);
nor U18156 (N_18156,N_17253,N_17869);
and U18157 (N_18157,N_16402,N_16428);
nor U18158 (N_18158,N_17189,N_16538);
or U18159 (N_18159,N_17069,N_17741);
nand U18160 (N_18160,N_17924,N_16475);
or U18161 (N_18161,N_17738,N_17389);
xnor U18162 (N_18162,N_17686,N_16494);
or U18163 (N_18163,N_16790,N_17449);
and U18164 (N_18164,N_16444,N_17198);
or U18165 (N_18165,N_16342,N_17181);
nor U18166 (N_18166,N_17385,N_16056);
nor U18167 (N_18167,N_17669,N_17401);
and U18168 (N_18168,N_16426,N_16352);
or U18169 (N_18169,N_16029,N_17226);
and U18170 (N_18170,N_17887,N_17860);
nand U18171 (N_18171,N_16326,N_16691);
nand U18172 (N_18172,N_16831,N_17883);
xnor U18173 (N_18173,N_17777,N_16778);
or U18174 (N_18174,N_16052,N_17196);
and U18175 (N_18175,N_17917,N_16239);
nor U18176 (N_18176,N_16812,N_16595);
and U18177 (N_18177,N_17325,N_17814);
nor U18178 (N_18178,N_16353,N_16014);
nor U18179 (N_18179,N_17150,N_17167);
xor U18180 (N_18180,N_16514,N_17918);
and U18181 (N_18181,N_17098,N_16408);
nor U18182 (N_18182,N_16798,N_17539);
or U18183 (N_18183,N_16312,N_16597);
xor U18184 (N_18184,N_16240,N_16278);
or U18185 (N_18185,N_16183,N_16162);
or U18186 (N_18186,N_16441,N_16140);
nor U18187 (N_18187,N_16568,N_17890);
nand U18188 (N_18188,N_16585,N_16694);
or U18189 (N_18189,N_16050,N_16175);
nand U18190 (N_18190,N_17785,N_17677);
nor U18191 (N_18191,N_17166,N_16871);
nand U18192 (N_18192,N_17858,N_17162);
nand U18193 (N_18193,N_16395,N_17529);
nor U18194 (N_18194,N_17460,N_17611);
or U18195 (N_18195,N_16033,N_16756);
nand U18196 (N_18196,N_17471,N_17608);
nor U18197 (N_18197,N_17292,N_16974);
nor U18198 (N_18198,N_17020,N_16745);
xnor U18199 (N_18199,N_17416,N_16801);
and U18200 (N_18200,N_17270,N_17691);
nand U18201 (N_18201,N_17804,N_16935);
nor U18202 (N_18202,N_17132,N_17654);
xor U18203 (N_18203,N_17157,N_17299);
nand U18204 (N_18204,N_16433,N_17206);
or U18205 (N_18205,N_16911,N_17579);
or U18206 (N_18206,N_17536,N_17707);
nand U18207 (N_18207,N_17494,N_16837);
and U18208 (N_18208,N_17671,N_16562);
xnor U18209 (N_18209,N_16068,N_16896);
nand U18210 (N_18210,N_16161,N_16186);
and U18211 (N_18211,N_16484,N_17496);
nand U18212 (N_18212,N_17454,N_17258);
and U18213 (N_18213,N_17874,N_16195);
nand U18214 (N_18214,N_16693,N_16878);
nand U18215 (N_18215,N_17141,N_17015);
or U18216 (N_18216,N_16423,N_17390);
or U18217 (N_18217,N_16351,N_17921);
xnor U18218 (N_18218,N_16086,N_17420);
and U18219 (N_18219,N_16508,N_16808);
nor U18220 (N_18220,N_16900,N_17174);
nand U18221 (N_18221,N_16036,N_17518);
and U18222 (N_18222,N_16469,N_16549);
nor U18223 (N_18223,N_16630,N_17263);
nand U18224 (N_18224,N_16567,N_17055);
xor U18225 (N_18225,N_17928,N_17812);
or U18226 (N_18226,N_17029,N_16332);
nor U18227 (N_18227,N_16173,N_16457);
and U18228 (N_18228,N_17068,N_16211);
nand U18229 (N_18229,N_16404,N_16833);
xor U18230 (N_18230,N_17511,N_17415);
or U18231 (N_18231,N_16250,N_16389);
and U18232 (N_18232,N_17010,N_16254);
nand U18233 (N_18233,N_17974,N_16301);
or U18234 (N_18234,N_17542,N_16083);
xor U18235 (N_18235,N_17376,N_16919);
and U18236 (N_18236,N_16430,N_17287);
and U18237 (N_18237,N_16178,N_17515);
xor U18238 (N_18238,N_17610,N_17688);
nand U18239 (N_18239,N_16750,N_17980);
xor U18240 (N_18240,N_17910,N_17058);
nor U18241 (N_18241,N_16409,N_16399);
and U18242 (N_18242,N_16368,N_17975);
nor U18243 (N_18243,N_16596,N_17514);
nor U18244 (N_18244,N_17559,N_16217);
or U18245 (N_18245,N_17596,N_17477);
nor U18246 (N_18246,N_16286,N_17395);
nor U18247 (N_18247,N_17937,N_16510);
nand U18248 (N_18248,N_17318,N_17796);
nor U18249 (N_18249,N_16760,N_16340);
nand U18250 (N_18250,N_17825,N_16113);
nand U18251 (N_18251,N_17908,N_16325);
nand U18252 (N_18252,N_17583,N_17694);
nand U18253 (N_18253,N_17886,N_16413);
nand U18254 (N_18254,N_17427,N_16460);
and U18255 (N_18255,N_16486,N_17070);
or U18256 (N_18256,N_17655,N_16147);
nor U18257 (N_18257,N_16683,N_16298);
nand U18258 (N_18258,N_16770,N_16135);
nand U18259 (N_18259,N_17750,N_17038);
nor U18260 (N_18260,N_17914,N_17926);
nor U18261 (N_18261,N_16040,N_17392);
and U18262 (N_18262,N_17558,N_17109);
nor U18263 (N_18263,N_16443,N_16379);
nand U18264 (N_18264,N_16906,N_17408);
nand U18265 (N_18265,N_16391,N_16529);
nor U18266 (N_18266,N_17607,N_16261);
nor U18267 (N_18267,N_17567,N_17101);
and U18268 (N_18268,N_17665,N_17990);
xnor U18269 (N_18269,N_16964,N_17818);
nor U18270 (N_18270,N_17676,N_17880);
nor U18271 (N_18271,N_17954,N_17647);
or U18272 (N_18272,N_17594,N_17698);
nand U18273 (N_18273,N_17468,N_16257);
and U18274 (N_18274,N_16780,N_17281);
nor U18275 (N_18275,N_16682,N_16598);
nor U18276 (N_18276,N_17194,N_16015);
and U18277 (N_18277,N_16841,N_17195);
and U18278 (N_18278,N_17185,N_16759);
nand U18279 (N_18279,N_17484,N_16613);
nor U18280 (N_18280,N_17381,N_16556);
and U18281 (N_18281,N_16393,N_17943);
xor U18282 (N_18282,N_17277,N_16335);
nor U18283 (N_18283,N_17981,N_17850);
nor U18284 (N_18284,N_17330,N_16796);
nor U18285 (N_18285,N_17899,N_16997);
nand U18286 (N_18286,N_17799,N_17276);
and U18287 (N_18287,N_17465,N_17480);
or U18288 (N_18288,N_16544,N_16127);
and U18289 (N_18289,N_17341,N_16729);
and U18290 (N_18290,N_16006,N_16678);
and U18291 (N_18291,N_17043,N_17873);
xnor U18292 (N_18292,N_16983,N_17351);
nand U18293 (N_18293,N_17803,N_16267);
nor U18294 (N_18294,N_17637,N_17144);
xor U18295 (N_18295,N_16825,N_16064);
nor U18296 (N_18296,N_16107,N_17105);
and U18297 (N_18297,N_16248,N_16638);
nor U18298 (N_18298,N_17965,N_16609);
xor U18299 (N_18299,N_17636,N_16488);
nor U18300 (N_18300,N_17147,N_17032);
nand U18301 (N_18301,N_16773,N_16489);
nand U18302 (N_18302,N_16366,N_17103);
nand U18303 (N_18303,N_16132,N_17316);
nand U18304 (N_18304,N_17305,N_16509);
and U18305 (N_18305,N_16855,N_17988);
and U18306 (N_18306,N_17019,N_16159);
nor U18307 (N_18307,N_16615,N_17479);
or U18308 (N_18308,N_16846,N_17793);
xor U18309 (N_18309,N_16821,N_16584);
and U18310 (N_18310,N_17091,N_16655);
and U18311 (N_18311,N_16245,N_16450);
or U18312 (N_18312,N_17778,N_16677);
nand U18313 (N_18313,N_17161,N_17005);
nand U18314 (N_18314,N_17176,N_17356);
nand U18315 (N_18315,N_16000,N_16493);
or U18316 (N_18316,N_17342,N_16626);
and U18317 (N_18317,N_16842,N_16114);
nand U18318 (N_18318,N_17119,N_17417);
and U18319 (N_18319,N_16309,N_17936);
nand U18320 (N_18320,N_17940,N_17526);
and U18321 (N_18321,N_16658,N_16894);
or U18322 (N_18322,N_16098,N_17441);
nand U18323 (N_18323,N_17553,N_17754);
nor U18324 (N_18324,N_16232,N_17451);
or U18325 (N_18325,N_17958,N_16434);
or U18326 (N_18326,N_16743,N_16851);
and U18327 (N_18327,N_17040,N_16406);
nand U18328 (N_18328,N_16198,N_16466);
nor U18329 (N_18329,N_17203,N_17425);
nand U18330 (N_18330,N_16910,N_16647);
or U18331 (N_18331,N_17264,N_17630);
nand U18332 (N_18332,N_17978,N_17964);
or U18333 (N_18333,N_17979,N_16372);
xor U18334 (N_18334,N_17800,N_17640);
nand U18335 (N_18335,N_17813,N_16057);
nand U18336 (N_18336,N_16367,N_17659);
nand U18337 (N_18337,N_16009,N_16885);
or U18338 (N_18338,N_16704,N_17272);
and U18339 (N_18339,N_17186,N_16446);
nand U18340 (N_18340,N_17107,N_16281);
nand U18341 (N_18341,N_17483,N_17359);
nand U18342 (N_18342,N_16273,N_16013);
nor U18343 (N_18343,N_17829,N_17047);
nand U18344 (N_18344,N_16981,N_17809);
and U18345 (N_18345,N_16662,N_16521);
and U18346 (N_18346,N_17817,N_17159);
nor U18347 (N_18347,N_17112,N_17490);
and U18348 (N_18348,N_17645,N_16686);
nor U18349 (N_18349,N_16214,N_17457);
nor U18350 (N_18350,N_16194,N_17617);
or U18351 (N_18351,N_16251,N_17331);
nor U18352 (N_18352,N_16937,N_17094);
nor U18353 (N_18353,N_16285,N_17642);
xor U18354 (N_18354,N_17871,N_16676);
and U18355 (N_18355,N_17801,N_17830);
and U18356 (N_18356,N_16673,N_16892);
xnor U18357 (N_18357,N_16421,N_17945);
or U18358 (N_18358,N_16950,N_16226);
or U18359 (N_18359,N_17927,N_17095);
or U18360 (N_18360,N_16109,N_17773);
or U18361 (N_18361,N_16035,N_16329);
xnor U18362 (N_18362,N_17153,N_17905);
and U18363 (N_18363,N_17445,N_16788);
and U18364 (N_18364,N_17054,N_16181);
nor U18365 (N_18365,N_17168,N_16016);
and U18366 (N_18366,N_17207,N_16185);
and U18367 (N_18367,N_16071,N_16576);
and U18368 (N_18368,N_17233,N_17960);
nor U18369 (N_18369,N_17440,N_17901);
nand U18370 (N_18370,N_17633,N_16699);
xnor U18371 (N_18371,N_17530,N_16397);
nand U18372 (N_18372,N_17952,N_17011);
nor U18373 (N_18373,N_16836,N_16633);
or U18374 (N_18374,N_16848,N_17013);
nand U18375 (N_18375,N_16102,N_16820);
xnor U18376 (N_18376,N_16560,N_17808);
and U18377 (N_18377,N_16386,N_16429);
and U18378 (N_18378,N_17865,N_16923);
or U18379 (N_18379,N_17716,N_16961);
or U18380 (N_18380,N_17705,N_16028);
xor U18381 (N_18381,N_17328,N_17509);
nand U18382 (N_18382,N_16266,N_17672);
xnor U18383 (N_18383,N_16333,N_16438);
xor U18384 (N_18384,N_17148,N_17982);
nor U18385 (N_18385,N_17448,N_16725);
nand U18386 (N_18386,N_16915,N_16188);
and U18387 (N_18387,N_17177,N_16364);
and U18388 (N_18388,N_17002,N_16838);
nand U18389 (N_18389,N_16828,N_16721);
nand U18390 (N_18390,N_16225,N_17232);
or U18391 (N_18391,N_17626,N_16814);
and U18392 (N_18392,N_16546,N_17834);
or U18393 (N_18393,N_17278,N_16943);
or U18394 (N_18394,N_16119,N_16641);
or U18395 (N_18395,N_16599,N_16465);
and U18396 (N_18396,N_16403,N_17183);
or U18397 (N_18397,N_17718,N_16152);
nand U18398 (N_18398,N_16458,N_16640);
or U18399 (N_18399,N_16809,N_16886);
xor U18400 (N_18400,N_17606,N_16241);
and U18401 (N_18401,N_17648,N_17600);
and U18402 (N_18402,N_16737,N_16455);
nand U18403 (N_18403,N_17837,N_16835);
nand U18404 (N_18404,N_16299,N_16696);
and U18405 (N_18405,N_17139,N_16369);
or U18406 (N_18406,N_17347,N_16203);
xor U18407 (N_18407,N_17436,N_16929);
nand U18408 (N_18408,N_16144,N_17740);
and U18409 (N_18409,N_16092,N_17134);
xnor U18410 (N_18410,N_16702,N_16898);
nand U18411 (N_18411,N_16977,N_17271);
and U18412 (N_18412,N_16313,N_16928);
nor U18413 (N_18413,N_16573,N_16687);
nand U18414 (N_18414,N_17568,N_17863);
or U18415 (N_18415,N_16872,N_16347);
and U18416 (N_18416,N_17133,N_17780);
nand U18417 (N_18417,N_17911,N_17797);
nand U18418 (N_18418,N_17418,N_16477);
nand U18419 (N_18419,N_17488,N_17324);
or U18420 (N_18420,N_16793,N_16503);
and U18421 (N_18421,N_16887,N_16116);
xor U18422 (N_18422,N_17495,N_16555);
nand U18423 (N_18423,N_16047,N_16427);
or U18424 (N_18424,N_16296,N_17731);
nand U18425 (N_18425,N_17321,N_16327);
xor U18426 (N_18426,N_17396,N_17763);
nand U18427 (N_18427,N_16764,N_16249);
and U18428 (N_18428,N_17052,N_16051);
nor U18429 (N_18429,N_16482,N_16551);
nor U18430 (N_18430,N_17370,N_17726);
and U18431 (N_18431,N_16505,N_17085);
and U18432 (N_18432,N_17893,N_16839);
nand U18433 (N_18433,N_17360,N_17171);
or U18434 (N_18434,N_17154,N_16076);
nor U18435 (N_18435,N_17151,N_17339);
xnor U18436 (N_18436,N_17575,N_17219);
nor U18437 (N_18437,N_17160,N_17566);
or U18438 (N_18438,N_17939,N_17589);
or U18439 (N_18439,N_17228,N_17970);
and U18440 (N_18440,N_17994,N_16614);
or U18441 (N_18441,N_17348,N_16087);
and U18442 (N_18442,N_16027,N_17756);
xnor U18443 (N_18443,N_16473,N_16907);
or U18444 (N_18444,N_17076,N_17866);
or U18445 (N_18445,N_16079,N_16968);
nand U18446 (N_18446,N_17618,N_16624);
nand U18447 (N_18447,N_16583,N_17028);
and U18448 (N_18448,N_17653,N_17967);
nor U18449 (N_18449,N_17050,N_16010);
nor U18450 (N_18450,N_17007,N_16746);
and U18451 (N_18451,N_17931,N_16605);
or U18452 (N_18452,N_16328,N_16933);
or U18453 (N_18453,N_16108,N_16293);
or U18454 (N_18454,N_16927,N_16862);
and U18455 (N_18455,N_17953,N_17208);
or U18456 (N_18456,N_16709,N_16625);
nand U18457 (N_18457,N_17025,N_17312);
nor U18458 (N_18458,N_16622,N_17547);
nand U18459 (N_18459,N_17489,N_16830);
nor U18460 (N_18460,N_16253,N_16497);
or U18461 (N_18461,N_16303,N_17512);
nor U18462 (N_18462,N_17009,N_17158);
and U18463 (N_18463,N_16715,N_16619);
xnor U18464 (N_18464,N_17846,N_17771);
nand U18465 (N_18465,N_17164,N_16062);
or U18466 (N_18466,N_16361,N_17469);
nand U18467 (N_18467,N_17776,N_16600);
nand U18468 (N_18468,N_16661,N_17806);
nor U18469 (N_18469,N_16782,N_17661);
and U18470 (N_18470,N_16097,N_16767);
or U18471 (N_18471,N_16706,N_16204);
xnor U18472 (N_18472,N_16411,N_17675);
nand U18473 (N_18473,N_16897,N_16018);
nand U18474 (N_18474,N_16776,N_17711);
xor U18475 (N_18475,N_17792,N_17319);
nor U18476 (N_18476,N_17383,N_16072);
and U18477 (N_18477,N_17930,N_16282);
xor U18478 (N_18478,N_17421,N_16845);
or U18479 (N_18479,N_17257,N_17616);
nand U18480 (N_18480,N_17838,N_16148);
or U18481 (N_18481,N_16772,N_16805);
nand U18482 (N_18482,N_16025,N_17450);
xor U18483 (N_18483,N_16516,N_17538);
nand U18484 (N_18484,N_17248,N_16863);
and U18485 (N_18485,N_17977,N_17983);
nor U18486 (N_18486,N_16345,N_17667);
nand U18487 (N_18487,N_17130,N_17963);
and U18488 (N_18488,N_17217,N_16513);
nor U18489 (N_18489,N_16490,N_16485);
nor U18490 (N_18490,N_16969,N_17146);
nand U18491 (N_18491,N_16462,N_16646);
and U18492 (N_18492,N_16244,N_16577);
and U18493 (N_18493,N_16973,N_16967);
nand U18494 (N_18494,N_16506,N_16277);
or U18495 (N_18495,N_16873,N_16823);
and U18496 (N_18496,N_17096,N_17681);
or U18497 (N_18497,N_16634,N_17071);
nor U18498 (N_18498,N_17946,N_17576);
or U18499 (N_18499,N_17989,N_16698);
nor U18500 (N_18500,N_17971,N_16744);
nor U18501 (N_18501,N_16168,N_16418);
nand U18502 (N_18502,N_17326,N_16034);
or U18503 (N_18503,N_17406,N_17082);
nor U18504 (N_18504,N_17259,N_16270);
nor U18505 (N_18505,N_16123,N_17894);
nor U18506 (N_18506,N_17344,N_16978);
nand U18507 (N_18507,N_16483,N_17180);
nor U18508 (N_18508,N_16648,N_17414);
or U18509 (N_18509,N_17631,N_16111);
and U18510 (N_18510,N_17861,N_17588);
or U18511 (N_18511,N_17550,N_16877);
xnor U18512 (N_18512,N_17853,N_16753);
nor U18513 (N_18513,N_16701,N_16067);
and U18514 (N_18514,N_16627,N_17557);
or U18515 (N_18515,N_17273,N_16090);
and U18516 (N_18516,N_16936,N_16290);
or U18517 (N_18517,N_16074,N_17250);
xnor U18518 (N_18518,N_16789,N_16670);
or U18519 (N_18519,N_17634,N_16199);
or U18520 (N_18520,N_16138,N_17845);
nor U18521 (N_18521,N_17915,N_17739);
or U18522 (N_18522,N_16331,N_17991);
nor U18523 (N_18523,N_16571,N_16049);
and U18524 (N_18524,N_17230,N_17693);
xor U18525 (N_18525,N_17289,N_16017);
xor U18526 (N_18526,N_16007,N_17507);
or U18527 (N_18527,N_16157,N_17012);
and U18528 (N_18528,N_16420,N_17377);
xnor U18529 (N_18529,N_16958,N_16197);
nor U18530 (N_18530,N_16586,N_16311);
and U18531 (N_18531,N_16754,N_17296);
nand U18532 (N_18532,N_16563,N_16784);
nand U18533 (N_18533,N_16671,N_17265);
nand U18534 (N_18534,N_17290,N_16984);
and U18535 (N_18535,N_17238,N_16233);
nand U18536 (N_18536,N_17214,N_17870);
nand U18537 (N_18537,N_16478,N_17268);
and U18538 (N_18538,N_16895,N_16775);
nand U18539 (N_18539,N_16274,N_16176);
nand U18540 (N_18540,N_17709,N_16354);
and U18541 (N_18541,N_16602,N_17556);
and U18542 (N_18542,N_16305,N_16612);
and U18543 (N_18543,N_16971,N_16644);
and U18544 (N_18544,N_16317,N_16817);
nand U18545 (N_18545,N_16081,N_17682);
or U18546 (N_18546,N_17759,N_17084);
nor U18547 (N_18547,N_16957,N_16223);
and U18548 (N_18548,N_16642,N_17916);
or U18549 (N_18549,N_17280,N_17593);
and U18550 (N_18550,N_16463,N_17127);
or U18551 (N_18551,N_16026,N_16230);
and U18552 (N_18552,N_16105,N_17537);
nand U18553 (N_18553,N_16870,N_17004);
nor U18554 (N_18554,N_16914,N_16449);
and U18555 (N_18555,N_17947,N_17572);
xor U18556 (N_18556,N_17948,N_17765);
nand U18557 (N_18557,N_16799,N_16859);
xnor U18558 (N_18558,N_16227,N_17255);
or U18559 (N_18559,N_16918,N_17540);
nor U18560 (N_18560,N_17587,N_17609);
or U18561 (N_18561,N_16852,N_17284);
nor U18562 (N_18562,N_16982,N_16315);
or U18563 (N_18563,N_17156,N_17192);
or U18564 (N_18564,N_16629,N_16187);
nand U18565 (N_18565,N_16792,N_17628);
nor U18566 (N_18566,N_17571,N_17815);
xnor U18567 (N_18567,N_17678,N_17816);
nand U18568 (N_18568,N_16592,N_17135);
and U18569 (N_18569,N_16019,N_17913);
or U18570 (N_18570,N_17972,N_16398);
and U18571 (N_18571,N_17703,N_16762);
nand U18572 (N_18572,N_17826,N_17384);
nor U18573 (N_18573,N_16024,N_16539);
nand U18574 (N_18574,N_16747,N_16356);
nand U18575 (N_18575,N_17037,N_16816);
and U18576 (N_18576,N_17229,N_16189);
nor U18577 (N_18577,N_17612,N_17400);
xor U18578 (N_18578,N_17555,N_17223);
xor U18579 (N_18579,N_17199,N_16786);
nor U18580 (N_18580,N_16499,N_17762);
nor U18581 (N_18581,N_16130,N_17266);
and U18582 (N_18582,N_16436,N_17231);
or U18583 (N_18583,N_17752,N_17702);
xnor U18584 (N_18584,N_17864,N_16022);
or U18585 (N_18585,N_17929,N_17569);
nor U18586 (N_18586,N_16912,N_17126);
nand U18587 (N_18587,N_16700,N_16238);
nand U18588 (N_18588,N_17170,N_17336);
nor U18589 (N_18589,N_16153,N_16860);
and U18590 (N_18590,N_17959,N_17320);
nor U18591 (N_18591,N_17993,N_17293);
nand U18592 (N_18592,N_17822,N_17721);
nand U18593 (N_18593,N_17267,N_16946);
and U18594 (N_18594,N_16739,N_17197);
nand U18595 (N_18595,N_17629,N_16495);
nor U18596 (N_18596,N_16515,N_17680);
and U18597 (N_18597,N_16679,N_16947);
xor U18598 (N_18598,N_17746,N_17835);
nor U18599 (N_18599,N_16470,N_17895);
xor U18600 (N_18600,N_17755,N_17493);
nand U18601 (N_18601,N_16280,N_16526);
xnor U18602 (N_18602,N_17833,N_17573);
nand U18603 (N_18603,N_16265,N_17660);
or U18604 (N_18604,N_17561,N_17674);
nand U18605 (N_18605,N_16868,N_17624);
nor U18606 (N_18606,N_16588,N_16660);
or U18607 (N_18607,N_16357,N_17527);
or U18608 (N_18608,N_17995,N_16668);
xnor U18609 (N_18609,N_16234,N_17689);
nand U18610 (N_18610,N_17039,N_17137);
or U18611 (N_18611,N_17102,N_16949);
and U18612 (N_18612,N_17563,N_16996);
or U18613 (N_18613,N_16680,N_16396);
nand U18614 (N_18614,N_17666,N_17513);
nand U18615 (N_18615,N_17605,N_16557);
nand U18616 (N_18616,N_16779,N_16246);
nor U18617 (N_18617,N_16766,N_16664);
or U18618 (N_18618,N_16456,N_17018);
xnor U18619 (N_18619,N_16922,N_17093);
nor U18620 (N_18620,N_16374,N_17081);
and U18621 (N_18621,N_16435,N_17889);
nand U18622 (N_18622,N_17892,N_17729);
and U18623 (N_18623,N_16561,N_17205);
and U18624 (N_18624,N_17603,N_16442);
nor U18625 (N_18625,N_16858,N_16882);
nor U18626 (N_18626,N_17274,N_17239);
or U18627 (N_18627,N_17065,N_17783);
or U18628 (N_18628,N_16224,N_16216);
or U18629 (N_18629,N_17876,N_16416);
and U18630 (N_18630,N_17467,N_17046);
and U18631 (N_18631,N_17549,N_17240);
nor U18632 (N_18632,N_16623,N_17499);
and U18633 (N_18633,N_16713,N_16259);
nand U18634 (N_18634,N_17169,N_16139);
nand U18635 (N_18635,N_17841,N_16547);
or U18636 (N_18636,N_17388,N_16388);
nand U18637 (N_18637,N_16688,N_17684);
nor U18638 (N_18638,N_17369,N_17016);
and U18639 (N_18639,N_16209,N_17875);
and U18640 (N_18640,N_16502,N_16045);
nor U18641 (N_18641,N_17831,N_16066);
nand U18642 (N_18642,N_16594,N_17173);
xor U18643 (N_18643,N_16643,N_16854);
and U18644 (N_18644,N_16213,N_16011);
and U18645 (N_18645,N_16431,N_16552);
and U18646 (N_18646,N_16120,N_17003);
nor U18647 (N_18647,N_17961,N_17110);
nor U18648 (N_18648,N_17482,N_17877);
nor U18649 (N_18649,N_16048,N_16628);
xnor U18650 (N_18650,N_16084,N_16707);
nand U18651 (N_18651,N_17552,N_17786);
nor U18652 (N_18652,N_16394,N_17844);
xor U18653 (N_18653,N_17562,N_17802);
and U18654 (N_18654,N_17544,N_17663);
nor U18655 (N_18655,N_17304,N_17111);
nand U18656 (N_18656,N_16545,N_17059);
and U18657 (N_18657,N_17710,N_17027);
and U18658 (N_18658,N_17592,N_17261);
nor U18659 (N_18659,N_16891,N_17443);
nor U18660 (N_18660,N_16260,N_16932);
nor U18661 (N_18661,N_17749,N_17502);
nand U18662 (N_18662,N_16337,N_17017);
nand U18663 (N_18663,N_16864,N_17190);
nor U18664 (N_18664,N_17862,N_17256);
and U18665 (N_18665,N_16054,N_16794);
or U18666 (N_18666,N_16038,N_16453);
and U18667 (N_18667,N_17026,N_16077);
or U18668 (N_18668,N_17362,N_16192);
nand U18669 (N_18669,N_16522,N_16004);
nor U18670 (N_18670,N_17788,N_16452);
and U18671 (N_18671,N_16930,N_16264);
or U18672 (N_18672,N_17884,N_17857);
or U18673 (N_18673,N_17394,N_17730);
nor U18674 (N_18674,N_17500,N_17781);
and U18675 (N_18675,N_17380,N_17079);
nor U18676 (N_18676,N_17021,N_16705);
nor U18677 (N_18677,N_16881,N_17438);
nand U18678 (N_18678,N_16985,N_17000);
or U18679 (N_18679,N_16580,N_16272);
nor U18680 (N_18680,N_16652,N_17193);
nand U18681 (N_18681,N_17202,N_17413);
nand U18682 (N_18682,N_16917,N_16491);
or U18683 (N_18683,N_16876,N_17622);
or U18684 (N_18684,N_16829,N_17523);
xnor U18685 (N_18685,N_17008,N_17124);
nand U18686 (N_18686,N_17706,N_16989);
nand U18687 (N_18687,N_16030,N_17782);
nor U18688 (N_18688,N_16531,N_16904);
or U18689 (N_18689,N_17632,N_16840);
nand U18690 (N_18690,N_17237,N_16292);
nor U18691 (N_18691,N_17108,N_17368);
nor U18692 (N_18692,N_16813,N_17658);
nand U18693 (N_18693,N_16955,N_16334);
nand U18694 (N_18694,N_17049,N_16165);
nand U18695 (N_18695,N_17345,N_16530);
nand U18696 (N_18696,N_17696,N_17424);
and U18697 (N_18697,N_17712,N_17428);
nor U18698 (N_18698,N_16564,N_17620);
xnor U18699 (N_18699,N_17361,N_16608);
nand U18700 (N_18700,N_17878,N_16474);
xor U18701 (N_18701,N_16321,N_16341);
nor U18702 (N_18702,N_16467,N_17053);
nor U18703 (N_18703,N_16088,N_16400);
xor U18704 (N_18704,N_17309,N_16543);
nor U18705 (N_18705,N_16815,N_16952);
nand U18706 (N_18706,N_17332,N_17322);
or U18707 (N_18707,N_17528,N_16110);
and U18708 (N_18708,N_16371,N_16459);
nor U18709 (N_18709,N_16205,N_16856);
nand U18710 (N_18710,N_17303,N_16925);
or U18711 (N_18711,N_17508,N_17560);
nor U18712 (N_18712,N_17179,N_16039);
and U18713 (N_18713,N_17976,N_17187);
or U18714 (N_18714,N_17364,N_17387);
or U18715 (N_18715,N_16201,N_16310);
or U18716 (N_18716,N_17590,N_16155);
or U18717 (N_18717,N_16358,N_17532);
and U18718 (N_18718,N_16279,N_17760);
nor U18719 (N_18719,N_16536,N_16732);
nand U18720 (N_18720,N_16288,N_17106);
and U18721 (N_18721,N_16432,N_17357);
nor U18722 (N_18722,N_17138,N_16748);
or U18723 (N_18723,N_17683,N_16617);
nand U18724 (N_18724,N_16043,N_17118);
nand U18725 (N_18725,N_17456,N_17472);
and U18726 (N_18726,N_17464,N_16061);
or U18727 (N_18727,N_17904,N_17757);
and U18728 (N_18728,N_16349,N_17849);
nand U18729 (N_18729,N_17249,N_17120);
nor U18730 (N_18730,N_17805,N_17985);
nand U18731 (N_18731,N_16636,N_16963);
and U18732 (N_18732,N_17235,N_16385);
or U18733 (N_18733,N_16196,N_16666);
or U18734 (N_18734,N_16154,N_16728);
xnor U18735 (N_18735,N_16219,N_16541);
xor U18736 (N_18736,N_17882,N_17064);
nor U18737 (N_18737,N_16853,N_16795);
or U18738 (N_18738,N_17354,N_16979);
xnor U18739 (N_18739,N_17879,N_16164);
and U18740 (N_18740,N_17591,N_16377);
and U18741 (N_18741,N_17627,N_16783);
nand U18742 (N_18742,N_17178,N_16101);
nor U18743 (N_18743,N_16172,N_16824);
nand U18744 (N_18744,N_16975,N_16726);
nand U18745 (N_18745,N_16206,N_17090);
xor U18746 (N_18746,N_17564,N_17949);
and U18747 (N_18747,N_17294,N_16674);
nand U18748 (N_18748,N_16222,N_17097);
or U18749 (N_18749,N_17251,N_17819);
nor U18750 (N_18750,N_17491,N_16180);
nand U18751 (N_18751,N_16032,N_16174);
xnor U18752 (N_18752,N_17234,N_16554);
and U18753 (N_18753,N_17072,N_16781);
nand U18754 (N_18754,N_17030,N_16291);
xnor U18755 (N_18755,N_16339,N_16986);
or U18756 (N_18756,N_16632,N_16735);
or U18757 (N_18757,N_17652,N_16220);
or U18758 (N_18758,N_17753,N_17900);
nand U18759 (N_18759,N_16284,N_16060);
nand U18760 (N_18760,N_17402,N_16236);
nor U18761 (N_18761,N_17298,N_16651);
nand U18762 (N_18762,N_16381,N_16080);
and U18763 (N_18763,N_16931,N_16359);
or U18764 (N_18764,N_17088,N_17136);
nand U18765 (N_18765,N_17649,N_17353);
nand U18766 (N_18766,N_17403,N_16944);
nor U18767 (N_18767,N_17584,N_17581);
nor U18768 (N_18768,N_17868,N_17212);
and U18769 (N_18769,N_16734,N_16765);
and U18770 (N_18770,N_16685,N_17121);
nand U18771 (N_18771,N_17117,N_17966);
or U18772 (N_18772,N_16672,N_16558);
nand U18773 (N_18773,N_16330,N_16718);
nand U18774 (N_18774,N_17719,N_17236);
nor U18775 (N_18775,N_16124,N_17764);
nor U18776 (N_18776,N_16373,N_16417);
and U18777 (N_18777,N_17851,N_17613);
and U18778 (N_18778,N_17386,N_16511);
nand U18779 (N_18779,N_16603,N_17795);
and U18780 (N_18780,N_16143,N_17131);
and U18781 (N_18781,N_17201,N_17315);
nand U18782 (N_18782,N_17433,N_16221);
nor U18783 (N_18783,N_16684,N_17621);
xnor U18784 (N_18784,N_17286,N_17378);
and U18785 (N_18785,N_16976,N_17246);
and U18786 (N_18786,N_17586,N_16318);
or U18787 (N_18787,N_17074,N_17984);
or U18788 (N_18788,N_16920,N_17713);
nor U18789 (N_18789,N_17516,N_17439);
and U18790 (N_18790,N_17363,N_16507);
or U18791 (N_18791,N_17060,N_17447);
nor U18792 (N_18792,N_16128,N_17779);
and U18793 (N_18793,N_17282,N_17225);
nand U18794 (N_18794,N_16711,N_16998);
and U18795 (N_18795,N_16115,N_16869);
nor U18796 (N_18796,N_17129,N_16407);
or U18797 (N_18797,N_16142,N_17182);
nor U18798 (N_18798,N_17044,N_16390);
or U18799 (N_18799,N_17310,N_16874);
nand U18800 (N_18800,N_17083,N_16095);
nand U18801 (N_18801,N_17968,N_16723);
nor U18802 (N_18802,N_17245,N_16579);
xor U18803 (N_18803,N_17662,N_17275);
or U18804 (N_18804,N_17685,N_17925);
nand U18805 (N_18805,N_17897,N_16208);
nor U18806 (N_18806,N_16901,N_17252);
nor U18807 (N_18807,N_16122,N_17923);
nand U18808 (N_18808,N_17881,N_17615);
xor U18809 (N_18809,N_17453,N_17373);
and U18810 (N_18810,N_17867,N_17920);
nor U18811 (N_18811,N_16665,N_16419);
nand U18812 (N_18812,N_16591,N_17601);
or U18813 (N_18813,N_16548,N_16363);
nand U18814 (N_18814,N_16271,N_17335);
or U18815 (N_18815,N_17372,N_16611);
and U18816 (N_18816,N_16237,N_16179);
or U18817 (N_18817,N_16738,N_17243);
nand U18818 (N_18818,N_17352,N_16908);
nor U18819 (N_18819,N_16962,N_17215);
or U18820 (N_18820,N_16847,N_16519);
and U18821 (N_18821,N_16888,N_16472);
and U18822 (N_18822,N_17122,N_16439);
xor U18823 (N_18823,N_16993,N_17476);
nand U18824 (N_18824,N_17533,N_16771);
nand U18825 (N_18825,N_16635,N_16287);
and U18826 (N_18826,N_17379,N_17986);
nand U18827 (N_18827,N_16524,N_17210);
nand U18828 (N_18828,N_16445,N_16582);
nand U18829 (N_18829,N_16990,N_17944);
or U18830 (N_18830,N_16804,N_16448);
nor U18831 (N_18831,N_17635,N_16941);
nand U18832 (N_18832,N_17962,N_17077);
xnor U18833 (N_18833,N_16731,N_17404);
nor U18834 (N_18834,N_17768,N_17885);
nor U18835 (N_18835,N_17656,N_16689);
and U18836 (N_18836,N_16899,N_16879);
or U18837 (N_18837,N_16145,N_16733);
xnor U18838 (N_18838,N_17463,N_17733);
and U18839 (N_18839,N_16637,N_17051);
or U18840 (N_18840,N_17535,N_17260);
nand U18841 (N_18841,N_17766,N_16520);
nand U18842 (N_18842,N_16867,N_17435);
or U18843 (N_18843,N_16806,N_16757);
or U18844 (N_18844,N_17774,N_17570);
nor U18845 (N_18845,N_16645,N_16200);
nand U18846 (N_18846,N_17042,N_16742);
or U18847 (N_18847,N_17204,N_16104);
nor U18848 (N_18848,N_16378,N_16811);
nor U18849 (N_18849,N_16343,N_17614);
xnor U18850 (N_18850,N_17155,N_16082);
nor U18851 (N_18851,N_17717,N_16012);
or U18852 (N_18852,N_17751,N_17506);
or U18853 (N_18853,N_17638,N_17534);
nand U18854 (N_18854,N_17548,N_16992);
and U18855 (N_18855,N_17089,N_16058);
or U18856 (N_18856,N_17149,N_17898);
xor U18857 (N_18857,N_17942,N_17934);
nor U18858 (N_18858,N_17856,N_16523);
nor U18859 (N_18859,N_17399,N_17700);
nand U18860 (N_18860,N_17902,N_17832);
and U18861 (N_18861,N_16117,N_17891);
and U18862 (N_18862,N_16163,N_16242);
or U18863 (N_18863,N_17317,N_16695);
nor U18864 (N_18864,N_17023,N_16550);
or U18865 (N_18865,N_16125,N_16649);
and U18866 (N_18866,N_17327,N_17478);
and U18867 (N_18867,N_16021,N_16857);
xnor U18868 (N_18868,N_16587,N_17909);
or U18869 (N_18869,N_17474,N_16151);
and U18870 (N_18870,N_16300,N_16763);
and U18871 (N_18871,N_17520,N_16850);
and U18872 (N_18872,N_16535,N_16959);
xor U18873 (N_18873,N_17222,N_16675);
and U18874 (N_18874,N_16708,N_16565);
nor U18875 (N_18875,N_17001,N_16063);
or U18876 (N_18876,N_17996,N_17932);
or U18877 (N_18877,N_17349,N_16103);
nor U18878 (N_18878,N_16913,N_16167);
nand U18879 (N_18879,N_16031,N_17346);
and U18880 (N_18880,N_16883,N_16141);
nand U18881 (N_18881,N_16008,N_16803);
nor U18882 (N_18882,N_16945,N_16618);
nand U18883 (N_18883,N_17722,N_16384);
nor U18884 (N_18884,N_16360,N_17446);
or U18885 (N_18885,N_16504,N_16053);
nor U18886 (N_18886,N_17623,N_17431);
nor U18887 (N_18887,N_16953,N_16834);
and U18888 (N_18888,N_16268,N_16893);
nor U18889 (N_18889,N_17412,N_16156);
nand U18890 (N_18890,N_16073,N_17933);
xnor U18891 (N_18891,N_17041,N_16348);
and U18892 (N_18892,N_17597,N_16940);
and U18893 (N_18893,N_16777,N_17987);
and U18894 (N_18894,N_17531,N_16131);
xor U18895 (N_18895,N_16621,N_16480);
and U18896 (N_18896,N_16533,N_16527);
nor U18897 (N_18897,N_17697,N_16730);
nand U18898 (N_18898,N_16055,N_16106);
and U18899 (N_18899,N_16191,N_17295);
or U18900 (N_18900,N_16517,N_17075);
nand U18901 (N_18901,N_17595,N_17761);
or U18902 (N_18902,N_16999,N_16939);
or U18903 (N_18903,N_17142,N_17724);
nor U18904 (N_18904,N_17308,N_17175);
and U18905 (N_18905,N_17715,N_17639);
nand U18906 (N_18906,N_16496,N_17006);
nand U18907 (N_18907,N_16070,N_17099);
and U18908 (N_18908,N_16751,N_16954);
nor U18909 (N_18909,N_17442,N_17580);
xnor U18910 (N_18910,N_16692,N_17302);
nand U18911 (N_18911,N_17227,N_16890);
nor U18912 (N_18912,N_17772,N_16518);
and U18913 (N_18913,N_16190,N_17747);
or U18914 (N_18914,N_17843,N_17405);
nor U18915 (N_18915,N_16590,N_16231);
and U18916 (N_18916,N_17371,N_16654);
and U18917 (N_18917,N_17997,N_16534);
nor U18918 (N_18918,N_17242,N_17859);
or U18919 (N_18919,N_17546,N_17789);
and U18920 (N_18920,N_16697,N_16126);
and U18921 (N_18921,N_16375,N_17375);
and U18922 (N_18922,N_16965,N_16819);
nand U18923 (N_18923,N_16464,N_17470);
and U18924 (N_18924,N_17956,N_16948);
or U18925 (N_18925,N_17125,N_16171);
and U18926 (N_18926,N_16956,N_16724);
xor U18927 (N_18927,N_17775,N_16320);
and U18928 (N_18928,N_16306,N_16387);
nor U18929 (N_18929,N_16440,N_17462);
or U18930 (N_18930,N_16578,N_17338);
and U18931 (N_18931,N_16422,N_16078);
nand U18932 (N_18932,N_16769,N_16720);
and U18933 (N_18933,N_17510,N_16924);
xor U18934 (N_18934,N_16880,N_17758);
or U18935 (N_18935,N_17409,N_16258);
and U18936 (N_18936,N_17521,N_17285);
nor U18937 (N_18937,N_17687,N_16525);
nand U18938 (N_18938,N_16606,N_17466);
and U18939 (N_18939,N_17737,N_16412);
nand U18940 (N_18940,N_16902,N_16100);
and U18941 (N_18941,N_17485,N_17734);
xnor U18942 (N_18942,N_16528,N_16476);
and U18943 (N_18943,N_16256,N_16593);
and U18944 (N_18944,N_16574,N_16263);
or U18945 (N_18945,N_17062,N_17269);
nor U18946 (N_18946,N_17398,N_17498);
and U18947 (N_18947,N_17541,N_17297);
and U18948 (N_18948,N_17501,N_17784);
nor U18949 (N_18949,N_17525,N_17723);
and U18950 (N_18950,N_17641,N_16207);
or U18951 (N_18951,N_17115,N_16802);
nor U18952 (N_18952,N_16425,N_16093);
nor U18953 (N_18953,N_17690,N_16243);
and U18954 (N_18954,N_16146,N_16134);
nand U18955 (N_18955,N_17973,N_16324);
nor U18956 (N_18956,N_16228,N_16096);
xnor U18957 (N_18957,N_16980,N_16657);
and U18958 (N_18958,N_16768,N_16553);
nor U18959 (N_18959,N_16350,N_17651);
or U18960 (N_18960,N_17209,N_17907);
nand U18961 (N_18961,N_16727,N_16182);
nand U18962 (N_18962,N_17999,N_17770);
and U18963 (N_18963,N_17888,N_16042);
nand U18964 (N_18964,N_17087,N_17505);
nor U18965 (N_18965,N_16269,N_17061);
or U18966 (N_18966,N_16631,N_16471);
xor U18967 (N_18967,N_16921,N_16849);
or U18968 (N_18968,N_16451,N_17355);
nor U18969 (N_18969,N_16059,N_16616);
xor U18970 (N_18970,N_16532,N_17314);
or U18971 (N_18971,N_17951,N_17855);
and U18972 (N_18972,N_16690,N_16149);
and U18973 (N_18973,N_17728,N_17847);
nor U18974 (N_18974,N_16540,N_17092);
nor U18975 (N_18975,N_16722,N_17340);
nor U18976 (N_18976,N_16276,N_17461);
nand U18977 (N_18977,N_16295,N_17221);
and U18978 (N_18978,N_16037,N_17140);
and U18979 (N_18979,N_16336,N_17426);
xor U18980 (N_18980,N_16988,N_17358);
or U18981 (N_18981,N_16717,N_16316);
nand U18982 (N_18982,N_16639,N_16099);
nor U18983 (N_18983,N_17452,N_16177);
and U18984 (N_18984,N_16656,N_17407);
nand U18985 (N_18985,N_16487,N_17769);
xnor U18986 (N_18986,N_17033,N_17481);
xor U18987 (N_18987,N_17458,N_17048);
nand U18988 (N_18988,N_16719,N_17497);
or U18989 (N_18989,N_17604,N_16133);
nand U18990 (N_18990,N_17810,N_17334);
nor U18991 (N_18991,N_16994,N_17577);
or U18992 (N_18992,N_17423,N_17432);
nand U18993 (N_18993,N_16294,N_17410);
and U18994 (N_18994,N_16741,N_17585);
nand U18995 (N_18995,N_17695,N_16229);
or U18996 (N_18996,N_17679,N_16160);
nand U18997 (N_18997,N_17429,N_17836);
or U18998 (N_18998,N_16150,N_16479);
or U18999 (N_18999,N_17034,N_16215);
and U19000 (N_19000,N_16634,N_16561);
and U19001 (N_19001,N_16178,N_16063);
nor U19002 (N_19002,N_16412,N_17798);
and U19003 (N_19003,N_17055,N_17842);
nor U19004 (N_19004,N_16074,N_17893);
nor U19005 (N_19005,N_16025,N_17110);
or U19006 (N_19006,N_16489,N_17596);
and U19007 (N_19007,N_17809,N_17997);
or U19008 (N_19008,N_16730,N_17195);
or U19009 (N_19009,N_16673,N_17344);
or U19010 (N_19010,N_17592,N_17978);
nand U19011 (N_19011,N_17924,N_17575);
nand U19012 (N_19012,N_17733,N_17664);
and U19013 (N_19013,N_17021,N_16224);
nor U19014 (N_19014,N_17395,N_16491);
or U19015 (N_19015,N_16219,N_16150);
or U19016 (N_19016,N_17391,N_16750);
nor U19017 (N_19017,N_17638,N_17777);
and U19018 (N_19018,N_17415,N_16901);
nor U19019 (N_19019,N_16094,N_16030);
nor U19020 (N_19020,N_16387,N_17407);
xnor U19021 (N_19021,N_17045,N_17219);
or U19022 (N_19022,N_16521,N_17023);
nand U19023 (N_19023,N_16225,N_16321);
nor U19024 (N_19024,N_17026,N_16643);
and U19025 (N_19025,N_16677,N_16164);
and U19026 (N_19026,N_16309,N_17668);
xor U19027 (N_19027,N_16145,N_16910);
nor U19028 (N_19028,N_17327,N_16699);
nor U19029 (N_19029,N_17606,N_16397);
nand U19030 (N_19030,N_17272,N_16203);
or U19031 (N_19031,N_17538,N_17688);
and U19032 (N_19032,N_17023,N_17197);
nand U19033 (N_19033,N_16938,N_16310);
and U19034 (N_19034,N_17257,N_16261);
and U19035 (N_19035,N_17488,N_17543);
or U19036 (N_19036,N_16493,N_17577);
and U19037 (N_19037,N_16431,N_17677);
xor U19038 (N_19038,N_17543,N_17331);
nor U19039 (N_19039,N_16899,N_16425);
or U19040 (N_19040,N_16543,N_16626);
nor U19041 (N_19041,N_17093,N_17175);
and U19042 (N_19042,N_17247,N_16474);
xnor U19043 (N_19043,N_16027,N_16329);
nand U19044 (N_19044,N_16640,N_16859);
and U19045 (N_19045,N_16083,N_17915);
and U19046 (N_19046,N_17917,N_16706);
nand U19047 (N_19047,N_17561,N_16404);
xnor U19048 (N_19048,N_17270,N_16243);
xor U19049 (N_19049,N_17177,N_17116);
xnor U19050 (N_19050,N_17569,N_17303);
nand U19051 (N_19051,N_17683,N_16518);
and U19052 (N_19052,N_17714,N_16609);
or U19053 (N_19053,N_16091,N_16610);
and U19054 (N_19054,N_17783,N_16125);
nor U19055 (N_19055,N_16224,N_16137);
xor U19056 (N_19056,N_17135,N_16955);
and U19057 (N_19057,N_16626,N_16826);
nand U19058 (N_19058,N_16365,N_17901);
and U19059 (N_19059,N_17476,N_16106);
and U19060 (N_19060,N_16150,N_17535);
nor U19061 (N_19061,N_16602,N_17668);
or U19062 (N_19062,N_16747,N_17024);
and U19063 (N_19063,N_16009,N_16947);
and U19064 (N_19064,N_16229,N_16355);
nand U19065 (N_19065,N_17352,N_17643);
nor U19066 (N_19066,N_17082,N_17835);
nand U19067 (N_19067,N_17146,N_17347);
nand U19068 (N_19068,N_17833,N_17676);
or U19069 (N_19069,N_16463,N_16787);
or U19070 (N_19070,N_16150,N_17445);
and U19071 (N_19071,N_16900,N_17846);
nand U19072 (N_19072,N_16165,N_16464);
nor U19073 (N_19073,N_17347,N_16422);
or U19074 (N_19074,N_16611,N_17368);
and U19075 (N_19075,N_16500,N_16159);
nor U19076 (N_19076,N_17827,N_17000);
nand U19077 (N_19077,N_17006,N_16330);
and U19078 (N_19078,N_16613,N_16302);
and U19079 (N_19079,N_16205,N_17386);
xnor U19080 (N_19080,N_16575,N_16789);
or U19081 (N_19081,N_16783,N_17511);
and U19082 (N_19082,N_16833,N_17985);
or U19083 (N_19083,N_17773,N_17800);
and U19084 (N_19084,N_17126,N_17289);
or U19085 (N_19085,N_16977,N_17518);
or U19086 (N_19086,N_17536,N_17315);
and U19087 (N_19087,N_16940,N_17865);
xor U19088 (N_19088,N_17791,N_16143);
or U19089 (N_19089,N_17388,N_17177);
nor U19090 (N_19090,N_16874,N_17421);
or U19091 (N_19091,N_17482,N_17936);
xnor U19092 (N_19092,N_17328,N_17988);
nand U19093 (N_19093,N_17450,N_17101);
or U19094 (N_19094,N_17351,N_17633);
and U19095 (N_19095,N_17725,N_16182);
or U19096 (N_19096,N_17584,N_16603);
nor U19097 (N_19097,N_16732,N_17947);
xnor U19098 (N_19098,N_17180,N_17944);
and U19099 (N_19099,N_17041,N_16661);
and U19100 (N_19100,N_17103,N_16297);
and U19101 (N_19101,N_16859,N_16386);
nand U19102 (N_19102,N_17031,N_17614);
or U19103 (N_19103,N_16245,N_17731);
or U19104 (N_19104,N_17414,N_17016);
xor U19105 (N_19105,N_16934,N_17429);
or U19106 (N_19106,N_17142,N_17651);
or U19107 (N_19107,N_17646,N_16780);
nand U19108 (N_19108,N_17008,N_16460);
nand U19109 (N_19109,N_17231,N_16408);
nor U19110 (N_19110,N_16489,N_16669);
nor U19111 (N_19111,N_16494,N_16162);
or U19112 (N_19112,N_17402,N_17781);
nor U19113 (N_19113,N_16182,N_16862);
nand U19114 (N_19114,N_16135,N_17125);
nor U19115 (N_19115,N_16356,N_17562);
nor U19116 (N_19116,N_17642,N_16890);
xnor U19117 (N_19117,N_16764,N_17700);
nand U19118 (N_19118,N_16348,N_16954);
nand U19119 (N_19119,N_17172,N_17039);
or U19120 (N_19120,N_16801,N_17073);
or U19121 (N_19121,N_17481,N_16656);
and U19122 (N_19122,N_16578,N_16129);
nand U19123 (N_19123,N_16619,N_16486);
xnor U19124 (N_19124,N_16284,N_17706);
nor U19125 (N_19125,N_16518,N_17997);
nand U19126 (N_19126,N_16284,N_17769);
xnor U19127 (N_19127,N_16051,N_16607);
and U19128 (N_19128,N_17547,N_17016);
nor U19129 (N_19129,N_16704,N_17823);
or U19130 (N_19130,N_16200,N_17247);
and U19131 (N_19131,N_17007,N_16834);
or U19132 (N_19132,N_16501,N_17938);
xnor U19133 (N_19133,N_16447,N_17301);
nand U19134 (N_19134,N_17720,N_16801);
nor U19135 (N_19135,N_17732,N_17103);
or U19136 (N_19136,N_16079,N_16061);
xnor U19137 (N_19137,N_16799,N_16344);
nand U19138 (N_19138,N_17715,N_16618);
nor U19139 (N_19139,N_16719,N_17580);
and U19140 (N_19140,N_17634,N_17565);
or U19141 (N_19141,N_16766,N_16760);
xnor U19142 (N_19142,N_17827,N_17924);
nor U19143 (N_19143,N_17058,N_17447);
nand U19144 (N_19144,N_16579,N_17171);
xor U19145 (N_19145,N_16584,N_17920);
or U19146 (N_19146,N_16227,N_16035);
xnor U19147 (N_19147,N_17586,N_17132);
and U19148 (N_19148,N_16113,N_17596);
nor U19149 (N_19149,N_16300,N_17029);
nor U19150 (N_19150,N_16978,N_16168);
nand U19151 (N_19151,N_17376,N_17659);
and U19152 (N_19152,N_16164,N_17735);
and U19153 (N_19153,N_17630,N_16790);
nor U19154 (N_19154,N_17535,N_17656);
nand U19155 (N_19155,N_16952,N_17494);
nand U19156 (N_19156,N_17504,N_16679);
xor U19157 (N_19157,N_17649,N_17829);
and U19158 (N_19158,N_16271,N_16910);
nor U19159 (N_19159,N_17852,N_17492);
and U19160 (N_19160,N_16300,N_16257);
and U19161 (N_19161,N_16802,N_16901);
or U19162 (N_19162,N_17700,N_17032);
nand U19163 (N_19163,N_16166,N_16223);
or U19164 (N_19164,N_17195,N_17169);
or U19165 (N_19165,N_17679,N_16274);
and U19166 (N_19166,N_17551,N_16175);
and U19167 (N_19167,N_16588,N_16744);
nor U19168 (N_19168,N_17016,N_17572);
nand U19169 (N_19169,N_16507,N_16609);
or U19170 (N_19170,N_17019,N_16315);
or U19171 (N_19171,N_17593,N_17358);
nor U19172 (N_19172,N_17638,N_16898);
or U19173 (N_19173,N_16518,N_17927);
nor U19174 (N_19174,N_16023,N_16006);
or U19175 (N_19175,N_16108,N_17322);
nor U19176 (N_19176,N_16954,N_16505);
xor U19177 (N_19177,N_17167,N_17968);
nor U19178 (N_19178,N_16838,N_17263);
nand U19179 (N_19179,N_17460,N_16842);
xor U19180 (N_19180,N_17218,N_16122);
nand U19181 (N_19181,N_17782,N_16052);
nand U19182 (N_19182,N_17396,N_17969);
or U19183 (N_19183,N_17448,N_16846);
nand U19184 (N_19184,N_16364,N_16959);
and U19185 (N_19185,N_16947,N_16448);
or U19186 (N_19186,N_17614,N_16212);
or U19187 (N_19187,N_17691,N_16973);
or U19188 (N_19188,N_17899,N_17510);
nor U19189 (N_19189,N_17077,N_17755);
or U19190 (N_19190,N_16797,N_17135);
or U19191 (N_19191,N_17155,N_17012);
or U19192 (N_19192,N_16617,N_17509);
nor U19193 (N_19193,N_17352,N_16343);
or U19194 (N_19194,N_17357,N_17817);
and U19195 (N_19195,N_16720,N_17449);
nand U19196 (N_19196,N_17049,N_16001);
nand U19197 (N_19197,N_16950,N_17394);
xnor U19198 (N_19198,N_17509,N_17925);
or U19199 (N_19199,N_16410,N_17177);
and U19200 (N_19200,N_17593,N_16794);
nand U19201 (N_19201,N_16844,N_16038);
nand U19202 (N_19202,N_16906,N_17710);
nor U19203 (N_19203,N_17651,N_16716);
nand U19204 (N_19204,N_16108,N_16459);
or U19205 (N_19205,N_16202,N_16881);
or U19206 (N_19206,N_17106,N_16778);
nand U19207 (N_19207,N_16157,N_17589);
xnor U19208 (N_19208,N_16704,N_16879);
and U19209 (N_19209,N_17953,N_16092);
nand U19210 (N_19210,N_16372,N_16092);
nand U19211 (N_19211,N_16546,N_17987);
or U19212 (N_19212,N_17591,N_16426);
nor U19213 (N_19213,N_16919,N_17358);
or U19214 (N_19214,N_16421,N_17164);
nor U19215 (N_19215,N_17291,N_16632);
or U19216 (N_19216,N_16656,N_16649);
nand U19217 (N_19217,N_17155,N_17341);
or U19218 (N_19218,N_16868,N_16387);
xor U19219 (N_19219,N_16301,N_16180);
nand U19220 (N_19220,N_16504,N_17204);
nand U19221 (N_19221,N_16954,N_17329);
and U19222 (N_19222,N_17231,N_16011);
xor U19223 (N_19223,N_17183,N_16436);
nand U19224 (N_19224,N_17016,N_17266);
xnor U19225 (N_19225,N_17661,N_16361);
and U19226 (N_19226,N_17743,N_17217);
xnor U19227 (N_19227,N_17895,N_16983);
or U19228 (N_19228,N_17151,N_16648);
or U19229 (N_19229,N_17550,N_17765);
and U19230 (N_19230,N_16791,N_16767);
or U19231 (N_19231,N_17323,N_17633);
xnor U19232 (N_19232,N_17988,N_17802);
nand U19233 (N_19233,N_17339,N_17871);
nand U19234 (N_19234,N_17043,N_17885);
nor U19235 (N_19235,N_16619,N_16326);
nand U19236 (N_19236,N_16872,N_17210);
nor U19237 (N_19237,N_16455,N_17060);
xor U19238 (N_19238,N_17567,N_16351);
nand U19239 (N_19239,N_16596,N_16591);
and U19240 (N_19240,N_16382,N_16828);
nand U19241 (N_19241,N_17455,N_17756);
and U19242 (N_19242,N_17850,N_16285);
and U19243 (N_19243,N_16186,N_16543);
nor U19244 (N_19244,N_17890,N_17864);
nor U19245 (N_19245,N_16658,N_17247);
nand U19246 (N_19246,N_16253,N_17120);
and U19247 (N_19247,N_17224,N_17879);
nor U19248 (N_19248,N_17883,N_17663);
or U19249 (N_19249,N_16862,N_17992);
and U19250 (N_19250,N_16551,N_17754);
nor U19251 (N_19251,N_16782,N_17156);
and U19252 (N_19252,N_16137,N_16768);
nor U19253 (N_19253,N_16455,N_16678);
nor U19254 (N_19254,N_16805,N_17043);
or U19255 (N_19255,N_16788,N_16388);
nand U19256 (N_19256,N_17389,N_17207);
or U19257 (N_19257,N_16056,N_16306);
and U19258 (N_19258,N_16993,N_17609);
xor U19259 (N_19259,N_16919,N_16206);
nand U19260 (N_19260,N_17284,N_17960);
nor U19261 (N_19261,N_17059,N_16947);
and U19262 (N_19262,N_16702,N_17700);
or U19263 (N_19263,N_16593,N_17944);
and U19264 (N_19264,N_17742,N_16027);
and U19265 (N_19265,N_16388,N_17777);
or U19266 (N_19266,N_17208,N_17216);
nor U19267 (N_19267,N_17611,N_16612);
and U19268 (N_19268,N_16840,N_16681);
nand U19269 (N_19269,N_17795,N_16557);
nand U19270 (N_19270,N_16966,N_17872);
and U19271 (N_19271,N_16981,N_17876);
nand U19272 (N_19272,N_17816,N_16972);
nor U19273 (N_19273,N_16989,N_17255);
and U19274 (N_19274,N_17928,N_17509);
nand U19275 (N_19275,N_17154,N_16404);
and U19276 (N_19276,N_16822,N_16794);
nand U19277 (N_19277,N_16542,N_16739);
xor U19278 (N_19278,N_17441,N_17339);
nand U19279 (N_19279,N_17649,N_17257);
and U19280 (N_19280,N_16082,N_16129);
nor U19281 (N_19281,N_16337,N_17471);
nand U19282 (N_19282,N_16510,N_16657);
nand U19283 (N_19283,N_16605,N_16976);
nor U19284 (N_19284,N_17057,N_16476);
xnor U19285 (N_19285,N_17617,N_16388);
and U19286 (N_19286,N_16123,N_16365);
and U19287 (N_19287,N_16353,N_17526);
or U19288 (N_19288,N_16589,N_17828);
nor U19289 (N_19289,N_17361,N_16117);
nand U19290 (N_19290,N_16383,N_17290);
or U19291 (N_19291,N_16503,N_16850);
nand U19292 (N_19292,N_16413,N_16428);
and U19293 (N_19293,N_16084,N_17072);
nand U19294 (N_19294,N_17087,N_16271);
xor U19295 (N_19295,N_17674,N_16184);
and U19296 (N_19296,N_16515,N_16716);
nor U19297 (N_19297,N_17806,N_17354);
or U19298 (N_19298,N_17339,N_16401);
xnor U19299 (N_19299,N_16290,N_17007);
or U19300 (N_19300,N_16381,N_17757);
or U19301 (N_19301,N_17006,N_17453);
or U19302 (N_19302,N_16287,N_17925);
or U19303 (N_19303,N_16243,N_16735);
xnor U19304 (N_19304,N_16761,N_16675);
or U19305 (N_19305,N_16695,N_16819);
and U19306 (N_19306,N_16306,N_17727);
nand U19307 (N_19307,N_17106,N_16416);
and U19308 (N_19308,N_17530,N_17652);
or U19309 (N_19309,N_17876,N_17314);
and U19310 (N_19310,N_17500,N_16903);
nor U19311 (N_19311,N_17882,N_17488);
or U19312 (N_19312,N_17920,N_17560);
or U19313 (N_19313,N_16563,N_16103);
and U19314 (N_19314,N_17357,N_16066);
and U19315 (N_19315,N_17267,N_16672);
or U19316 (N_19316,N_16335,N_16665);
and U19317 (N_19317,N_16098,N_16125);
or U19318 (N_19318,N_16714,N_16783);
nor U19319 (N_19319,N_16287,N_16040);
nand U19320 (N_19320,N_17807,N_17314);
or U19321 (N_19321,N_17981,N_16837);
or U19322 (N_19322,N_17457,N_17304);
xor U19323 (N_19323,N_17561,N_16748);
nor U19324 (N_19324,N_16592,N_16661);
or U19325 (N_19325,N_16304,N_16003);
xnor U19326 (N_19326,N_17627,N_16479);
nor U19327 (N_19327,N_17264,N_17139);
xnor U19328 (N_19328,N_16609,N_17725);
nand U19329 (N_19329,N_17407,N_17155);
nand U19330 (N_19330,N_17063,N_16031);
and U19331 (N_19331,N_17569,N_17099);
xor U19332 (N_19332,N_16220,N_16092);
or U19333 (N_19333,N_17903,N_17632);
and U19334 (N_19334,N_17628,N_17197);
xnor U19335 (N_19335,N_17347,N_17548);
and U19336 (N_19336,N_17054,N_17832);
or U19337 (N_19337,N_16249,N_17055);
nand U19338 (N_19338,N_16841,N_16190);
or U19339 (N_19339,N_17564,N_17618);
or U19340 (N_19340,N_16704,N_17797);
or U19341 (N_19341,N_16720,N_17115);
and U19342 (N_19342,N_17230,N_16395);
nand U19343 (N_19343,N_16796,N_17857);
or U19344 (N_19344,N_17654,N_16326);
and U19345 (N_19345,N_17816,N_17863);
and U19346 (N_19346,N_17534,N_17330);
and U19347 (N_19347,N_17719,N_16972);
or U19348 (N_19348,N_17180,N_16865);
nor U19349 (N_19349,N_16806,N_17391);
or U19350 (N_19350,N_16143,N_17519);
nor U19351 (N_19351,N_17414,N_17509);
or U19352 (N_19352,N_17668,N_17194);
and U19353 (N_19353,N_16619,N_17095);
or U19354 (N_19354,N_16481,N_16498);
or U19355 (N_19355,N_16173,N_17396);
nand U19356 (N_19356,N_16156,N_17480);
or U19357 (N_19357,N_16756,N_17481);
nor U19358 (N_19358,N_17215,N_16746);
nand U19359 (N_19359,N_17371,N_17279);
or U19360 (N_19360,N_17691,N_17806);
and U19361 (N_19361,N_17196,N_16659);
and U19362 (N_19362,N_16068,N_16576);
xnor U19363 (N_19363,N_17094,N_17935);
nand U19364 (N_19364,N_16001,N_17598);
or U19365 (N_19365,N_17382,N_16730);
nor U19366 (N_19366,N_16725,N_16081);
and U19367 (N_19367,N_16708,N_16110);
nand U19368 (N_19368,N_17162,N_16471);
and U19369 (N_19369,N_17539,N_17257);
or U19370 (N_19370,N_17099,N_16938);
or U19371 (N_19371,N_17051,N_17615);
nand U19372 (N_19372,N_16619,N_17311);
xnor U19373 (N_19373,N_16664,N_17973);
nand U19374 (N_19374,N_17382,N_17250);
nor U19375 (N_19375,N_17929,N_16597);
and U19376 (N_19376,N_17140,N_17555);
or U19377 (N_19377,N_17377,N_17425);
and U19378 (N_19378,N_16737,N_17732);
nor U19379 (N_19379,N_17063,N_17994);
and U19380 (N_19380,N_16073,N_16968);
xor U19381 (N_19381,N_17342,N_17453);
and U19382 (N_19382,N_16875,N_17178);
or U19383 (N_19383,N_17997,N_16089);
nor U19384 (N_19384,N_17483,N_16018);
nand U19385 (N_19385,N_17735,N_17842);
and U19386 (N_19386,N_17365,N_16200);
and U19387 (N_19387,N_16441,N_17989);
xnor U19388 (N_19388,N_17906,N_16156);
nand U19389 (N_19389,N_16197,N_16684);
or U19390 (N_19390,N_16002,N_16537);
or U19391 (N_19391,N_17862,N_17786);
nor U19392 (N_19392,N_16895,N_16703);
and U19393 (N_19393,N_17799,N_17873);
nand U19394 (N_19394,N_16785,N_16131);
nor U19395 (N_19395,N_17840,N_16831);
nor U19396 (N_19396,N_17401,N_16785);
nor U19397 (N_19397,N_17790,N_16600);
nor U19398 (N_19398,N_17791,N_17814);
xor U19399 (N_19399,N_16560,N_17960);
nor U19400 (N_19400,N_17518,N_16854);
nand U19401 (N_19401,N_17254,N_16497);
nand U19402 (N_19402,N_17569,N_16378);
or U19403 (N_19403,N_16892,N_16408);
nor U19404 (N_19404,N_17255,N_16463);
nor U19405 (N_19405,N_17077,N_17513);
nand U19406 (N_19406,N_16721,N_17060);
and U19407 (N_19407,N_16499,N_16996);
nor U19408 (N_19408,N_17297,N_16784);
and U19409 (N_19409,N_16418,N_17474);
nor U19410 (N_19410,N_16557,N_16341);
nor U19411 (N_19411,N_16051,N_16923);
nand U19412 (N_19412,N_17589,N_17218);
nor U19413 (N_19413,N_17701,N_16033);
or U19414 (N_19414,N_17080,N_17526);
nor U19415 (N_19415,N_17926,N_16952);
nand U19416 (N_19416,N_17402,N_16300);
nor U19417 (N_19417,N_17760,N_16101);
and U19418 (N_19418,N_16292,N_17898);
nand U19419 (N_19419,N_16422,N_17339);
nand U19420 (N_19420,N_17191,N_16218);
nor U19421 (N_19421,N_16172,N_16367);
nor U19422 (N_19422,N_16347,N_17573);
nor U19423 (N_19423,N_17022,N_17231);
nor U19424 (N_19424,N_17084,N_16117);
and U19425 (N_19425,N_17016,N_16645);
or U19426 (N_19426,N_17314,N_17999);
or U19427 (N_19427,N_17286,N_17447);
nand U19428 (N_19428,N_17406,N_17211);
nor U19429 (N_19429,N_16806,N_17059);
nor U19430 (N_19430,N_17839,N_17077);
xnor U19431 (N_19431,N_17163,N_17886);
xor U19432 (N_19432,N_17080,N_16825);
nand U19433 (N_19433,N_16315,N_16029);
and U19434 (N_19434,N_16834,N_16216);
and U19435 (N_19435,N_17363,N_17074);
or U19436 (N_19436,N_17186,N_16922);
or U19437 (N_19437,N_16629,N_17537);
nor U19438 (N_19438,N_16378,N_17956);
and U19439 (N_19439,N_17207,N_17074);
or U19440 (N_19440,N_17125,N_16269);
or U19441 (N_19441,N_16841,N_17484);
nand U19442 (N_19442,N_17264,N_16338);
or U19443 (N_19443,N_17583,N_17606);
nand U19444 (N_19444,N_16508,N_17331);
nor U19445 (N_19445,N_16458,N_17493);
and U19446 (N_19446,N_17550,N_17990);
nand U19447 (N_19447,N_16598,N_16159);
and U19448 (N_19448,N_16200,N_17368);
or U19449 (N_19449,N_17664,N_16152);
nor U19450 (N_19450,N_16879,N_17861);
or U19451 (N_19451,N_17358,N_17836);
or U19452 (N_19452,N_16903,N_16916);
xnor U19453 (N_19453,N_16745,N_17797);
nor U19454 (N_19454,N_17287,N_16860);
or U19455 (N_19455,N_17098,N_17432);
or U19456 (N_19456,N_17751,N_17852);
xor U19457 (N_19457,N_17891,N_16487);
or U19458 (N_19458,N_17722,N_16289);
nor U19459 (N_19459,N_16655,N_16615);
or U19460 (N_19460,N_17657,N_17609);
nor U19461 (N_19461,N_16026,N_16842);
and U19462 (N_19462,N_17995,N_16643);
and U19463 (N_19463,N_16504,N_17413);
and U19464 (N_19464,N_16658,N_16748);
nand U19465 (N_19465,N_17726,N_16087);
nor U19466 (N_19466,N_17459,N_16563);
and U19467 (N_19467,N_17937,N_17795);
and U19468 (N_19468,N_16697,N_17122);
nand U19469 (N_19469,N_17896,N_16627);
and U19470 (N_19470,N_17269,N_17974);
nand U19471 (N_19471,N_16210,N_17092);
and U19472 (N_19472,N_16060,N_17414);
or U19473 (N_19473,N_17922,N_16205);
xnor U19474 (N_19474,N_16048,N_16044);
xnor U19475 (N_19475,N_17432,N_17868);
or U19476 (N_19476,N_16095,N_16805);
nand U19477 (N_19477,N_16811,N_16161);
or U19478 (N_19478,N_17102,N_17854);
and U19479 (N_19479,N_16649,N_17862);
nand U19480 (N_19480,N_17052,N_17562);
nand U19481 (N_19481,N_16571,N_16791);
xor U19482 (N_19482,N_17161,N_17246);
nand U19483 (N_19483,N_16085,N_16406);
and U19484 (N_19484,N_16980,N_17899);
nand U19485 (N_19485,N_16137,N_17189);
nand U19486 (N_19486,N_16244,N_17988);
nor U19487 (N_19487,N_16013,N_16762);
and U19488 (N_19488,N_16894,N_17200);
or U19489 (N_19489,N_17516,N_17894);
xnor U19490 (N_19490,N_17071,N_17334);
nand U19491 (N_19491,N_16128,N_16722);
nand U19492 (N_19492,N_17373,N_16906);
and U19493 (N_19493,N_17086,N_17435);
nor U19494 (N_19494,N_17815,N_17303);
and U19495 (N_19495,N_16893,N_16465);
nand U19496 (N_19496,N_17280,N_17881);
or U19497 (N_19497,N_16511,N_16809);
nand U19498 (N_19498,N_16104,N_16675);
or U19499 (N_19499,N_16684,N_17528);
nor U19500 (N_19500,N_16736,N_17677);
or U19501 (N_19501,N_17860,N_16807);
and U19502 (N_19502,N_17103,N_17507);
and U19503 (N_19503,N_16448,N_16517);
nor U19504 (N_19504,N_16071,N_17991);
xnor U19505 (N_19505,N_16256,N_17753);
or U19506 (N_19506,N_17446,N_17912);
nand U19507 (N_19507,N_16459,N_17876);
xor U19508 (N_19508,N_16888,N_16320);
nand U19509 (N_19509,N_17367,N_16996);
or U19510 (N_19510,N_16898,N_16283);
and U19511 (N_19511,N_16683,N_17107);
nor U19512 (N_19512,N_17598,N_16558);
nand U19513 (N_19513,N_16225,N_17118);
nand U19514 (N_19514,N_17374,N_16182);
nand U19515 (N_19515,N_17169,N_17697);
and U19516 (N_19516,N_17569,N_17738);
or U19517 (N_19517,N_17507,N_17935);
nand U19518 (N_19518,N_16256,N_17017);
or U19519 (N_19519,N_16231,N_17595);
nand U19520 (N_19520,N_17161,N_17618);
or U19521 (N_19521,N_16603,N_16249);
nand U19522 (N_19522,N_16905,N_17551);
xnor U19523 (N_19523,N_16224,N_17123);
nor U19524 (N_19524,N_17251,N_17693);
or U19525 (N_19525,N_17257,N_17085);
xnor U19526 (N_19526,N_16881,N_17526);
nor U19527 (N_19527,N_16613,N_16625);
xor U19528 (N_19528,N_17985,N_17321);
xnor U19529 (N_19529,N_16053,N_17030);
nand U19530 (N_19530,N_16748,N_17369);
or U19531 (N_19531,N_16615,N_17347);
or U19532 (N_19532,N_17288,N_17870);
nand U19533 (N_19533,N_16742,N_17238);
or U19534 (N_19534,N_17506,N_17013);
nand U19535 (N_19535,N_16974,N_17134);
and U19536 (N_19536,N_16270,N_16196);
and U19537 (N_19537,N_16670,N_16975);
xnor U19538 (N_19538,N_16115,N_17638);
or U19539 (N_19539,N_16328,N_16900);
or U19540 (N_19540,N_16996,N_17727);
or U19541 (N_19541,N_16090,N_17431);
or U19542 (N_19542,N_16792,N_17542);
or U19543 (N_19543,N_16163,N_16316);
nor U19544 (N_19544,N_16055,N_17866);
nand U19545 (N_19545,N_16301,N_16065);
or U19546 (N_19546,N_17529,N_16140);
nand U19547 (N_19547,N_17858,N_16258);
or U19548 (N_19548,N_16530,N_17115);
or U19549 (N_19549,N_17619,N_17759);
nand U19550 (N_19550,N_17919,N_16138);
nand U19551 (N_19551,N_16659,N_17240);
or U19552 (N_19552,N_16832,N_16654);
nand U19553 (N_19553,N_17828,N_17149);
or U19554 (N_19554,N_17131,N_17874);
or U19555 (N_19555,N_17577,N_16195);
nand U19556 (N_19556,N_17448,N_16194);
or U19557 (N_19557,N_17250,N_16761);
nor U19558 (N_19558,N_16432,N_17132);
nand U19559 (N_19559,N_17969,N_17324);
nor U19560 (N_19560,N_16531,N_17392);
or U19561 (N_19561,N_16284,N_17863);
nor U19562 (N_19562,N_16015,N_16442);
or U19563 (N_19563,N_16100,N_16361);
nor U19564 (N_19564,N_17485,N_16680);
nand U19565 (N_19565,N_17348,N_16688);
nand U19566 (N_19566,N_17240,N_17100);
or U19567 (N_19567,N_16022,N_16766);
or U19568 (N_19568,N_17979,N_17740);
nor U19569 (N_19569,N_16992,N_16176);
xor U19570 (N_19570,N_17408,N_17727);
and U19571 (N_19571,N_17975,N_17032);
and U19572 (N_19572,N_17272,N_16868);
nor U19573 (N_19573,N_16739,N_17788);
and U19574 (N_19574,N_16174,N_17557);
nand U19575 (N_19575,N_16612,N_16101);
and U19576 (N_19576,N_16200,N_17446);
nand U19577 (N_19577,N_16931,N_17287);
nor U19578 (N_19578,N_16378,N_17118);
nand U19579 (N_19579,N_16720,N_17827);
nor U19580 (N_19580,N_16293,N_17477);
and U19581 (N_19581,N_16538,N_16833);
nand U19582 (N_19582,N_16429,N_16236);
nor U19583 (N_19583,N_16377,N_16663);
or U19584 (N_19584,N_16130,N_16584);
and U19585 (N_19585,N_16486,N_16684);
and U19586 (N_19586,N_16710,N_16249);
nor U19587 (N_19587,N_16971,N_16043);
xor U19588 (N_19588,N_16552,N_17623);
and U19589 (N_19589,N_17587,N_16575);
and U19590 (N_19590,N_17284,N_17454);
and U19591 (N_19591,N_17725,N_16757);
or U19592 (N_19592,N_17393,N_17049);
nand U19593 (N_19593,N_16694,N_17109);
and U19594 (N_19594,N_17137,N_17686);
nor U19595 (N_19595,N_17086,N_17967);
nor U19596 (N_19596,N_16874,N_16041);
nor U19597 (N_19597,N_17292,N_16647);
nor U19598 (N_19598,N_16186,N_17625);
and U19599 (N_19599,N_17128,N_17173);
xor U19600 (N_19600,N_16137,N_17451);
and U19601 (N_19601,N_17442,N_16796);
nor U19602 (N_19602,N_16987,N_16143);
nor U19603 (N_19603,N_16391,N_16671);
nor U19604 (N_19604,N_16473,N_17129);
or U19605 (N_19605,N_16196,N_16894);
xor U19606 (N_19606,N_17451,N_17236);
nor U19607 (N_19607,N_17843,N_17406);
nor U19608 (N_19608,N_17256,N_17200);
nand U19609 (N_19609,N_17339,N_16331);
and U19610 (N_19610,N_16809,N_16490);
or U19611 (N_19611,N_16406,N_16171);
and U19612 (N_19612,N_17178,N_16881);
nor U19613 (N_19613,N_16048,N_17013);
nor U19614 (N_19614,N_16431,N_17288);
xnor U19615 (N_19615,N_16829,N_16007);
nand U19616 (N_19616,N_16064,N_17962);
nand U19617 (N_19617,N_16715,N_16487);
nand U19618 (N_19618,N_16747,N_16782);
nand U19619 (N_19619,N_17295,N_16820);
or U19620 (N_19620,N_16042,N_16138);
or U19621 (N_19621,N_17169,N_17617);
and U19622 (N_19622,N_16288,N_16009);
nand U19623 (N_19623,N_16025,N_16892);
or U19624 (N_19624,N_17507,N_17066);
nand U19625 (N_19625,N_17384,N_17491);
nand U19626 (N_19626,N_16100,N_16893);
or U19627 (N_19627,N_17670,N_17240);
nand U19628 (N_19628,N_17375,N_17324);
nand U19629 (N_19629,N_17272,N_16708);
nor U19630 (N_19630,N_17336,N_17353);
nor U19631 (N_19631,N_17578,N_17735);
nor U19632 (N_19632,N_17323,N_17085);
and U19633 (N_19633,N_16317,N_16154);
nand U19634 (N_19634,N_17593,N_17534);
nor U19635 (N_19635,N_17270,N_16690);
and U19636 (N_19636,N_16917,N_17269);
nor U19637 (N_19637,N_16583,N_17318);
or U19638 (N_19638,N_17078,N_16700);
nand U19639 (N_19639,N_17647,N_16133);
nor U19640 (N_19640,N_17971,N_17738);
xnor U19641 (N_19641,N_17528,N_16091);
nor U19642 (N_19642,N_17541,N_16208);
xor U19643 (N_19643,N_16485,N_17604);
or U19644 (N_19644,N_17985,N_17263);
and U19645 (N_19645,N_16815,N_17880);
xor U19646 (N_19646,N_17732,N_16590);
nor U19647 (N_19647,N_16314,N_16893);
nor U19648 (N_19648,N_16992,N_16846);
or U19649 (N_19649,N_17175,N_17059);
nor U19650 (N_19650,N_16907,N_17092);
nor U19651 (N_19651,N_17117,N_17626);
or U19652 (N_19652,N_17612,N_17801);
xor U19653 (N_19653,N_17017,N_16572);
nor U19654 (N_19654,N_17394,N_17002);
and U19655 (N_19655,N_16331,N_16954);
and U19656 (N_19656,N_17425,N_16800);
nor U19657 (N_19657,N_16112,N_17752);
and U19658 (N_19658,N_17556,N_17340);
nor U19659 (N_19659,N_16180,N_17214);
and U19660 (N_19660,N_16671,N_16706);
nand U19661 (N_19661,N_16960,N_16571);
and U19662 (N_19662,N_17607,N_16354);
or U19663 (N_19663,N_16448,N_17959);
or U19664 (N_19664,N_16280,N_17101);
or U19665 (N_19665,N_17724,N_16366);
and U19666 (N_19666,N_17315,N_17507);
xor U19667 (N_19667,N_17797,N_17107);
and U19668 (N_19668,N_16638,N_17122);
nand U19669 (N_19669,N_16221,N_17719);
nor U19670 (N_19670,N_16245,N_17733);
nor U19671 (N_19671,N_17272,N_16500);
or U19672 (N_19672,N_17679,N_17758);
xnor U19673 (N_19673,N_17442,N_17171);
or U19674 (N_19674,N_16160,N_16028);
nor U19675 (N_19675,N_17182,N_16326);
nand U19676 (N_19676,N_16803,N_16744);
nand U19677 (N_19677,N_17110,N_17202);
nor U19678 (N_19678,N_17419,N_16785);
or U19679 (N_19679,N_17864,N_16324);
nand U19680 (N_19680,N_17492,N_16342);
xnor U19681 (N_19681,N_16006,N_17191);
nor U19682 (N_19682,N_16945,N_17173);
nand U19683 (N_19683,N_16915,N_16585);
nand U19684 (N_19684,N_16996,N_16373);
and U19685 (N_19685,N_17529,N_16832);
nand U19686 (N_19686,N_16839,N_17708);
or U19687 (N_19687,N_16940,N_17641);
nand U19688 (N_19688,N_17260,N_16837);
and U19689 (N_19689,N_17014,N_16899);
or U19690 (N_19690,N_16689,N_16208);
nor U19691 (N_19691,N_16201,N_16939);
xnor U19692 (N_19692,N_16162,N_17742);
nor U19693 (N_19693,N_17168,N_16820);
nand U19694 (N_19694,N_17940,N_16339);
or U19695 (N_19695,N_16347,N_17577);
or U19696 (N_19696,N_17114,N_17361);
nand U19697 (N_19697,N_16592,N_17528);
nor U19698 (N_19698,N_16219,N_16091);
or U19699 (N_19699,N_17408,N_16435);
nand U19700 (N_19700,N_17357,N_16624);
and U19701 (N_19701,N_16190,N_16724);
nand U19702 (N_19702,N_17467,N_17975);
xnor U19703 (N_19703,N_17399,N_17627);
and U19704 (N_19704,N_17410,N_16138);
nor U19705 (N_19705,N_17858,N_17022);
and U19706 (N_19706,N_16926,N_16940);
nand U19707 (N_19707,N_17235,N_17419);
xor U19708 (N_19708,N_16686,N_16963);
nand U19709 (N_19709,N_17174,N_16253);
nor U19710 (N_19710,N_17687,N_17342);
and U19711 (N_19711,N_16900,N_17936);
and U19712 (N_19712,N_16558,N_16122);
or U19713 (N_19713,N_16234,N_16280);
xor U19714 (N_19714,N_17191,N_17771);
or U19715 (N_19715,N_16767,N_17998);
and U19716 (N_19716,N_16977,N_17050);
nand U19717 (N_19717,N_17229,N_16138);
and U19718 (N_19718,N_16037,N_16481);
xor U19719 (N_19719,N_16012,N_16898);
xnor U19720 (N_19720,N_16267,N_16412);
and U19721 (N_19721,N_16094,N_16224);
and U19722 (N_19722,N_16216,N_16981);
or U19723 (N_19723,N_16547,N_16545);
nand U19724 (N_19724,N_16748,N_17415);
nor U19725 (N_19725,N_17546,N_17182);
nor U19726 (N_19726,N_17149,N_17351);
or U19727 (N_19727,N_16680,N_16430);
or U19728 (N_19728,N_16708,N_16566);
or U19729 (N_19729,N_16821,N_16766);
or U19730 (N_19730,N_16612,N_16168);
xor U19731 (N_19731,N_16930,N_17562);
nor U19732 (N_19732,N_17615,N_16345);
and U19733 (N_19733,N_16513,N_17729);
nor U19734 (N_19734,N_16542,N_16290);
nor U19735 (N_19735,N_17229,N_17026);
xor U19736 (N_19736,N_16931,N_16930);
nor U19737 (N_19737,N_17098,N_17655);
or U19738 (N_19738,N_17035,N_17471);
nor U19739 (N_19739,N_16500,N_17199);
or U19740 (N_19740,N_16765,N_17058);
or U19741 (N_19741,N_16333,N_16513);
or U19742 (N_19742,N_16705,N_17510);
nor U19743 (N_19743,N_17753,N_17583);
nor U19744 (N_19744,N_17845,N_16117);
nand U19745 (N_19745,N_16646,N_17908);
or U19746 (N_19746,N_17607,N_17706);
nor U19747 (N_19747,N_16598,N_17059);
nand U19748 (N_19748,N_17832,N_16989);
and U19749 (N_19749,N_17492,N_16441);
nand U19750 (N_19750,N_17306,N_17177);
and U19751 (N_19751,N_17077,N_16760);
or U19752 (N_19752,N_17619,N_16018);
nand U19753 (N_19753,N_17828,N_16161);
and U19754 (N_19754,N_17934,N_16460);
nand U19755 (N_19755,N_17509,N_16534);
and U19756 (N_19756,N_17617,N_16441);
xnor U19757 (N_19757,N_17474,N_16586);
nor U19758 (N_19758,N_16203,N_16111);
or U19759 (N_19759,N_17323,N_17677);
or U19760 (N_19760,N_16779,N_17226);
nor U19761 (N_19761,N_16656,N_17066);
and U19762 (N_19762,N_16217,N_17855);
nor U19763 (N_19763,N_17043,N_16926);
or U19764 (N_19764,N_17318,N_16252);
and U19765 (N_19765,N_16133,N_16834);
and U19766 (N_19766,N_17674,N_16646);
nor U19767 (N_19767,N_17874,N_16609);
nor U19768 (N_19768,N_17343,N_16865);
nor U19769 (N_19769,N_16129,N_16764);
nand U19770 (N_19770,N_17002,N_16009);
nand U19771 (N_19771,N_17657,N_16689);
or U19772 (N_19772,N_16799,N_17440);
nor U19773 (N_19773,N_17662,N_16840);
nand U19774 (N_19774,N_17005,N_17749);
nand U19775 (N_19775,N_17175,N_17288);
and U19776 (N_19776,N_17098,N_17975);
nor U19777 (N_19777,N_16130,N_16219);
nand U19778 (N_19778,N_17414,N_16382);
and U19779 (N_19779,N_16681,N_16511);
and U19780 (N_19780,N_17168,N_16531);
nor U19781 (N_19781,N_17855,N_17422);
nor U19782 (N_19782,N_16435,N_16434);
nor U19783 (N_19783,N_16638,N_16724);
and U19784 (N_19784,N_17889,N_16192);
nor U19785 (N_19785,N_17256,N_16177);
or U19786 (N_19786,N_16155,N_16382);
nor U19787 (N_19787,N_16495,N_16857);
or U19788 (N_19788,N_16638,N_16169);
and U19789 (N_19789,N_16348,N_16973);
nand U19790 (N_19790,N_16662,N_16710);
nand U19791 (N_19791,N_17421,N_17694);
xnor U19792 (N_19792,N_16582,N_16641);
nor U19793 (N_19793,N_16845,N_16736);
xnor U19794 (N_19794,N_16766,N_17967);
and U19795 (N_19795,N_16669,N_17181);
or U19796 (N_19796,N_16238,N_16453);
nor U19797 (N_19797,N_16281,N_17732);
nor U19798 (N_19798,N_17016,N_16611);
nand U19799 (N_19799,N_17021,N_16192);
nor U19800 (N_19800,N_16917,N_16282);
or U19801 (N_19801,N_16158,N_17472);
nor U19802 (N_19802,N_16984,N_16836);
nor U19803 (N_19803,N_17777,N_17048);
nor U19804 (N_19804,N_16801,N_17335);
and U19805 (N_19805,N_17633,N_17500);
nand U19806 (N_19806,N_16918,N_17954);
nor U19807 (N_19807,N_16815,N_17393);
nand U19808 (N_19808,N_17917,N_16804);
nor U19809 (N_19809,N_17684,N_17251);
nor U19810 (N_19810,N_16629,N_17719);
and U19811 (N_19811,N_16314,N_16814);
nor U19812 (N_19812,N_17416,N_16172);
nand U19813 (N_19813,N_17234,N_16676);
nand U19814 (N_19814,N_17320,N_16759);
and U19815 (N_19815,N_17377,N_17035);
or U19816 (N_19816,N_16756,N_16472);
nor U19817 (N_19817,N_17602,N_16136);
nor U19818 (N_19818,N_16012,N_16926);
nand U19819 (N_19819,N_16541,N_17233);
xnor U19820 (N_19820,N_16986,N_16193);
and U19821 (N_19821,N_17088,N_17680);
or U19822 (N_19822,N_17496,N_16845);
nand U19823 (N_19823,N_17161,N_16901);
xor U19824 (N_19824,N_17088,N_17129);
or U19825 (N_19825,N_16077,N_16517);
nor U19826 (N_19826,N_17123,N_17623);
or U19827 (N_19827,N_17894,N_17992);
and U19828 (N_19828,N_16361,N_17523);
nand U19829 (N_19829,N_17385,N_17991);
nand U19830 (N_19830,N_17838,N_16226);
xor U19831 (N_19831,N_16787,N_17081);
or U19832 (N_19832,N_17518,N_16268);
and U19833 (N_19833,N_16865,N_16985);
nor U19834 (N_19834,N_17993,N_16317);
xnor U19835 (N_19835,N_16598,N_17175);
nor U19836 (N_19836,N_16485,N_16687);
and U19837 (N_19837,N_17523,N_16407);
and U19838 (N_19838,N_16803,N_17775);
nand U19839 (N_19839,N_17296,N_16572);
or U19840 (N_19840,N_16861,N_16063);
or U19841 (N_19841,N_16054,N_16382);
nor U19842 (N_19842,N_17296,N_16879);
and U19843 (N_19843,N_16565,N_16377);
nand U19844 (N_19844,N_16778,N_16672);
and U19845 (N_19845,N_17812,N_17328);
or U19846 (N_19846,N_16895,N_16747);
nor U19847 (N_19847,N_16601,N_17719);
or U19848 (N_19848,N_16889,N_17589);
nor U19849 (N_19849,N_16313,N_16665);
or U19850 (N_19850,N_16083,N_17772);
nand U19851 (N_19851,N_17373,N_16501);
or U19852 (N_19852,N_17694,N_17412);
xor U19853 (N_19853,N_16115,N_16175);
and U19854 (N_19854,N_17964,N_16068);
and U19855 (N_19855,N_16224,N_17395);
xor U19856 (N_19856,N_16789,N_17393);
nor U19857 (N_19857,N_17576,N_17707);
nand U19858 (N_19858,N_16953,N_17527);
or U19859 (N_19859,N_16082,N_16899);
or U19860 (N_19860,N_16270,N_17508);
or U19861 (N_19861,N_17413,N_17914);
or U19862 (N_19862,N_17276,N_17264);
nor U19863 (N_19863,N_17141,N_17256);
or U19864 (N_19864,N_17325,N_17774);
nor U19865 (N_19865,N_17758,N_16821);
xor U19866 (N_19866,N_17723,N_16819);
and U19867 (N_19867,N_17723,N_17227);
xor U19868 (N_19868,N_17697,N_17640);
xnor U19869 (N_19869,N_16605,N_16673);
nand U19870 (N_19870,N_16511,N_16623);
nand U19871 (N_19871,N_17565,N_16584);
nand U19872 (N_19872,N_17669,N_17472);
and U19873 (N_19873,N_17002,N_16852);
and U19874 (N_19874,N_17348,N_17614);
xor U19875 (N_19875,N_16640,N_16748);
nor U19876 (N_19876,N_17888,N_17562);
xor U19877 (N_19877,N_16356,N_17780);
and U19878 (N_19878,N_17249,N_16666);
nor U19879 (N_19879,N_17620,N_16541);
nand U19880 (N_19880,N_17687,N_17576);
and U19881 (N_19881,N_17895,N_16956);
and U19882 (N_19882,N_17917,N_17001);
and U19883 (N_19883,N_17269,N_17608);
nand U19884 (N_19884,N_16792,N_17675);
nor U19885 (N_19885,N_16942,N_17447);
xnor U19886 (N_19886,N_17788,N_16181);
nor U19887 (N_19887,N_17679,N_16860);
or U19888 (N_19888,N_17740,N_16307);
nand U19889 (N_19889,N_16699,N_16692);
or U19890 (N_19890,N_17008,N_16336);
nor U19891 (N_19891,N_17488,N_17408);
and U19892 (N_19892,N_17555,N_16218);
nor U19893 (N_19893,N_17817,N_16206);
xor U19894 (N_19894,N_16796,N_16757);
nand U19895 (N_19895,N_17081,N_17715);
nand U19896 (N_19896,N_17352,N_16669);
nand U19897 (N_19897,N_17562,N_16595);
and U19898 (N_19898,N_17060,N_16020);
or U19899 (N_19899,N_16295,N_16357);
or U19900 (N_19900,N_17817,N_16440);
nand U19901 (N_19901,N_16344,N_16185);
or U19902 (N_19902,N_17746,N_16872);
nor U19903 (N_19903,N_16160,N_17566);
and U19904 (N_19904,N_17047,N_16640);
or U19905 (N_19905,N_16220,N_16824);
nor U19906 (N_19906,N_16210,N_16357);
nor U19907 (N_19907,N_17545,N_17977);
or U19908 (N_19908,N_17774,N_16982);
and U19909 (N_19909,N_17711,N_17284);
and U19910 (N_19910,N_17111,N_16401);
and U19911 (N_19911,N_17459,N_17672);
and U19912 (N_19912,N_16166,N_17177);
or U19913 (N_19913,N_16453,N_17468);
or U19914 (N_19914,N_17474,N_17649);
nor U19915 (N_19915,N_17276,N_16691);
or U19916 (N_19916,N_16529,N_16816);
xor U19917 (N_19917,N_17266,N_17764);
nor U19918 (N_19918,N_16488,N_17863);
and U19919 (N_19919,N_16696,N_17794);
or U19920 (N_19920,N_17530,N_17671);
xor U19921 (N_19921,N_17057,N_17715);
nor U19922 (N_19922,N_16061,N_16239);
xnor U19923 (N_19923,N_16031,N_16829);
nand U19924 (N_19924,N_17373,N_17040);
nand U19925 (N_19925,N_16195,N_17025);
nor U19926 (N_19926,N_16980,N_17406);
or U19927 (N_19927,N_17024,N_16724);
xor U19928 (N_19928,N_16513,N_17097);
or U19929 (N_19929,N_17501,N_17082);
and U19930 (N_19930,N_16162,N_16544);
or U19931 (N_19931,N_16631,N_16464);
or U19932 (N_19932,N_17124,N_17194);
nor U19933 (N_19933,N_17335,N_17640);
nand U19934 (N_19934,N_16227,N_17363);
nand U19935 (N_19935,N_16705,N_16771);
nand U19936 (N_19936,N_17811,N_16074);
and U19937 (N_19937,N_17502,N_17252);
and U19938 (N_19938,N_17697,N_16771);
nand U19939 (N_19939,N_17646,N_16996);
nor U19940 (N_19940,N_17247,N_16490);
or U19941 (N_19941,N_16728,N_16846);
nor U19942 (N_19942,N_17508,N_16844);
or U19943 (N_19943,N_16768,N_17393);
nor U19944 (N_19944,N_17157,N_17763);
nand U19945 (N_19945,N_17925,N_16391);
nand U19946 (N_19946,N_16707,N_16290);
nand U19947 (N_19947,N_17559,N_17258);
nor U19948 (N_19948,N_17588,N_17879);
or U19949 (N_19949,N_17048,N_16866);
or U19950 (N_19950,N_16262,N_17065);
nor U19951 (N_19951,N_16370,N_17959);
and U19952 (N_19952,N_16082,N_16242);
xor U19953 (N_19953,N_17652,N_17297);
nor U19954 (N_19954,N_17129,N_16180);
nor U19955 (N_19955,N_16251,N_16666);
nor U19956 (N_19956,N_17218,N_16591);
and U19957 (N_19957,N_16585,N_17383);
or U19958 (N_19958,N_16697,N_16981);
and U19959 (N_19959,N_17024,N_16524);
nand U19960 (N_19960,N_17438,N_17895);
nor U19961 (N_19961,N_17325,N_16804);
and U19962 (N_19962,N_17869,N_17574);
and U19963 (N_19963,N_16013,N_16080);
or U19964 (N_19964,N_17720,N_16637);
or U19965 (N_19965,N_17983,N_17686);
and U19966 (N_19966,N_16446,N_17710);
or U19967 (N_19967,N_17095,N_16790);
and U19968 (N_19968,N_17426,N_17696);
and U19969 (N_19969,N_16099,N_16402);
nand U19970 (N_19970,N_17220,N_16290);
and U19971 (N_19971,N_17445,N_17295);
nand U19972 (N_19972,N_16467,N_16095);
or U19973 (N_19973,N_17285,N_16636);
nand U19974 (N_19974,N_16427,N_16395);
xnor U19975 (N_19975,N_17570,N_17005);
or U19976 (N_19976,N_17332,N_17693);
or U19977 (N_19977,N_17098,N_16746);
xor U19978 (N_19978,N_16627,N_17626);
and U19979 (N_19979,N_16876,N_17105);
and U19980 (N_19980,N_16179,N_16059);
or U19981 (N_19981,N_16385,N_17015);
or U19982 (N_19982,N_16538,N_16596);
nand U19983 (N_19983,N_17835,N_17688);
xnor U19984 (N_19984,N_17736,N_16065);
or U19985 (N_19985,N_17240,N_16360);
xnor U19986 (N_19986,N_17864,N_16192);
and U19987 (N_19987,N_16690,N_17985);
and U19988 (N_19988,N_16445,N_16909);
nor U19989 (N_19989,N_16577,N_16292);
xor U19990 (N_19990,N_17048,N_17662);
or U19991 (N_19991,N_17906,N_17536);
xnor U19992 (N_19992,N_17673,N_17039);
xor U19993 (N_19993,N_17489,N_16542);
and U19994 (N_19994,N_17555,N_16925);
or U19995 (N_19995,N_17949,N_17921);
and U19996 (N_19996,N_16694,N_16059);
nand U19997 (N_19997,N_16766,N_16515);
nand U19998 (N_19998,N_17014,N_16998);
nand U19999 (N_19999,N_16936,N_16665);
xor UO_0 (O_0,N_18134,N_18122);
nand UO_1 (O_1,N_18376,N_18042);
or UO_2 (O_2,N_18989,N_19021);
nand UO_3 (O_3,N_19428,N_18637);
xnor UO_4 (O_4,N_18858,N_19531);
xor UO_5 (O_5,N_18770,N_18589);
or UO_6 (O_6,N_19905,N_19857);
nand UO_7 (O_7,N_19980,N_18699);
and UO_8 (O_8,N_18564,N_18548);
nor UO_9 (O_9,N_19459,N_19227);
or UO_10 (O_10,N_18790,N_19489);
nor UO_11 (O_11,N_18505,N_18166);
and UO_12 (O_12,N_18050,N_19627);
and UO_13 (O_13,N_18774,N_18557);
nand UO_14 (O_14,N_19875,N_19977);
nand UO_15 (O_15,N_19701,N_18150);
nor UO_16 (O_16,N_19307,N_18411);
nor UO_17 (O_17,N_18162,N_18644);
and UO_18 (O_18,N_18247,N_19322);
or UO_19 (O_19,N_19380,N_19207);
nand UO_20 (O_20,N_19062,N_18563);
nor UO_21 (O_21,N_18343,N_19024);
nand UO_22 (O_22,N_19815,N_18843);
xnor UO_23 (O_23,N_18863,N_19522);
nand UO_24 (O_24,N_18213,N_19827);
nand UO_25 (O_25,N_19549,N_18091);
nor UO_26 (O_26,N_19669,N_19259);
or UO_27 (O_27,N_18633,N_19440);
nand UO_28 (O_28,N_18119,N_19639);
xnor UO_29 (O_29,N_19230,N_18340);
and UO_30 (O_30,N_18609,N_18757);
or UO_31 (O_31,N_18573,N_18281);
or UO_32 (O_32,N_18468,N_19364);
nand UO_33 (O_33,N_18691,N_18788);
nor UO_34 (O_34,N_18201,N_19610);
nand UO_35 (O_35,N_18590,N_18897);
nand UO_36 (O_36,N_19724,N_18437);
nor UO_37 (O_37,N_18246,N_19298);
nand UO_38 (O_38,N_19861,N_19629);
nor UO_39 (O_39,N_18995,N_18344);
xnor UO_40 (O_40,N_19763,N_19025);
nand UO_41 (O_41,N_18527,N_19251);
nor UO_42 (O_42,N_18908,N_19819);
and UO_43 (O_43,N_18158,N_18671);
and UO_44 (O_44,N_19390,N_18605);
nor UO_45 (O_45,N_19926,N_18192);
or UO_46 (O_46,N_19608,N_19636);
or UO_47 (O_47,N_19013,N_19743);
and UO_48 (O_48,N_18335,N_18891);
nor UO_49 (O_49,N_18276,N_18057);
and UO_50 (O_50,N_18345,N_18580);
nor UO_51 (O_51,N_18566,N_19809);
and UO_52 (O_52,N_18215,N_18888);
or UO_53 (O_53,N_18405,N_18726);
xor UO_54 (O_54,N_19456,N_18591);
nand UO_55 (O_55,N_19165,N_19734);
and UO_56 (O_56,N_19474,N_19874);
and UO_57 (O_57,N_18502,N_19195);
xnor UO_58 (O_58,N_19029,N_19341);
nor UO_59 (O_59,N_19732,N_19694);
and UO_60 (O_60,N_18689,N_19904);
and UO_61 (O_61,N_18872,N_19889);
or UO_62 (O_62,N_19956,N_19598);
and UO_63 (O_63,N_18098,N_19289);
and UO_64 (O_64,N_18945,N_18903);
nor UO_65 (O_65,N_19087,N_19234);
nand UO_66 (O_66,N_19587,N_18386);
nor UO_67 (O_67,N_18728,N_19236);
and UO_68 (O_68,N_18075,N_18499);
and UO_69 (O_69,N_18270,N_18883);
or UO_70 (O_70,N_18277,N_19678);
nand UO_71 (O_71,N_18651,N_18873);
and UO_72 (O_72,N_18646,N_19134);
or UO_73 (O_73,N_18598,N_18640);
or UO_74 (O_74,N_18526,N_18224);
or UO_75 (O_75,N_18205,N_19148);
nand UO_76 (O_76,N_18771,N_19737);
xor UO_77 (O_77,N_18353,N_19839);
or UO_78 (O_78,N_18009,N_18756);
nor UO_79 (O_79,N_18413,N_18919);
nand UO_80 (O_80,N_19880,N_18341);
nand UO_81 (O_81,N_19617,N_18541);
and UO_82 (O_82,N_18538,N_18494);
or UO_83 (O_83,N_18967,N_19156);
xor UO_84 (O_84,N_18832,N_19504);
nand UO_85 (O_85,N_18769,N_18078);
nand UO_86 (O_86,N_19922,N_18798);
and UO_87 (O_87,N_19334,N_19276);
or UO_88 (O_88,N_18680,N_18635);
and UO_89 (O_89,N_19699,N_18801);
xor UO_90 (O_90,N_19785,N_19347);
or UO_91 (O_91,N_18307,N_19125);
or UO_92 (O_92,N_18375,N_19594);
and UO_93 (O_93,N_18463,N_19797);
and UO_94 (O_94,N_18177,N_18156);
or UO_95 (O_95,N_19937,N_19019);
and UO_96 (O_96,N_19780,N_18773);
and UO_97 (O_97,N_19717,N_18423);
and UO_98 (O_98,N_19064,N_18944);
and UO_99 (O_99,N_18339,N_18806);
nor UO_100 (O_100,N_19108,N_19589);
or UO_101 (O_101,N_19993,N_19909);
and UO_102 (O_102,N_19676,N_18550);
or UO_103 (O_103,N_19677,N_18358);
nor UO_104 (O_104,N_18868,N_18291);
nor UO_105 (O_105,N_18731,N_18327);
nand UO_106 (O_106,N_18441,N_19103);
and UO_107 (O_107,N_19661,N_19398);
nand UO_108 (O_108,N_19620,N_18128);
and UO_109 (O_109,N_19917,N_18090);
nor UO_110 (O_110,N_19246,N_19060);
nor UO_111 (O_111,N_19487,N_19686);
and UO_112 (O_112,N_19329,N_19052);
nand UO_113 (O_113,N_18831,N_18673);
xor UO_114 (O_114,N_19213,N_19615);
nand UO_115 (O_115,N_19419,N_19853);
and UO_116 (O_116,N_19054,N_18647);
or UO_117 (O_117,N_18300,N_18244);
xor UO_118 (O_118,N_18565,N_19953);
xnor UO_119 (O_119,N_18927,N_19229);
or UO_120 (O_120,N_18266,N_18661);
and UO_121 (O_121,N_19557,N_19176);
and UO_122 (O_122,N_19050,N_18792);
xor UO_123 (O_123,N_18684,N_19936);
xor UO_124 (O_124,N_19547,N_19477);
or UO_125 (O_125,N_18223,N_19545);
nand UO_126 (O_126,N_18280,N_18132);
nor UO_127 (O_127,N_18096,N_19525);
nand UO_128 (O_128,N_19071,N_19957);
nand UO_129 (O_129,N_18429,N_19462);
xnor UO_130 (O_130,N_19619,N_19360);
nor UO_131 (O_131,N_18137,N_19911);
nand UO_132 (O_132,N_18398,N_19680);
or UO_133 (O_133,N_19458,N_19408);
or UO_134 (O_134,N_19974,N_18665);
xnor UO_135 (O_135,N_19424,N_19884);
or UO_136 (O_136,N_19015,N_18292);
nand UO_137 (O_137,N_19812,N_18937);
and UO_138 (O_138,N_18759,N_19327);
xnor UO_139 (O_139,N_18182,N_19973);
and UO_140 (O_140,N_19515,N_19215);
and UO_141 (O_141,N_19362,N_19662);
or UO_142 (O_142,N_19350,N_19453);
and UO_143 (O_143,N_18762,N_19344);
and UO_144 (O_144,N_18023,N_18392);
and UO_145 (O_145,N_18772,N_19443);
xnor UO_146 (O_146,N_19252,N_18662);
nand UO_147 (O_147,N_18072,N_18282);
and UO_148 (O_148,N_18139,N_19388);
nand UO_149 (O_149,N_18302,N_19495);
nor UO_150 (O_150,N_19172,N_18030);
or UO_151 (O_151,N_19208,N_19927);
and UO_152 (O_152,N_19439,N_19521);
nor UO_153 (O_153,N_18886,N_18370);
nand UO_154 (O_154,N_18459,N_18200);
nand UO_155 (O_155,N_18231,N_18932);
xnor UO_156 (O_156,N_19745,N_19243);
or UO_157 (O_157,N_18093,N_19469);
nor UO_158 (O_158,N_19817,N_18273);
or UO_159 (O_159,N_18059,N_19285);
or UO_160 (O_160,N_19028,N_19203);
and UO_161 (O_161,N_19121,N_19754);
or UO_162 (O_162,N_18606,N_18679);
nand UO_163 (O_163,N_18663,N_19828);
nand UO_164 (O_164,N_19850,N_19290);
xor UO_165 (O_165,N_19317,N_19033);
and UO_166 (O_166,N_19391,N_19591);
nand UO_167 (O_167,N_19007,N_18636);
nor UO_168 (O_168,N_19095,N_19012);
nand UO_169 (O_169,N_19444,N_18620);
and UO_170 (O_170,N_18439,N_19830);
and UO_171 (O_171,N_19561,N_18961);
or UO_172 (O_172,N_18087,N_19363);
nor UO_173 (O_173,N_18626,N_18144);
nor UO_174 (O_174,N_18037,N_18734);
and UO_175 (O_175,N_18109,N_19672);
and UO_176 (O_176,N_19768,N_19170);
and UO_177 (O_177,N_18498,N_19635);
nor UO_178 (O_178,N_18138,N_19090);
nand UO_179 (O_179,N_18904,N_19761);
xnor UO_180 (O_180,N_19325,N_18632);
xnor UO_181 (O_181,N_19590,N_19593);
nor UO_182 (O_182,N_19559,N_19681);
nand UO_183 (O_183,N_19175,N_19302);
xnor UO_184 (O_184,N_19653,N_19069);
or UO_185 (O_185,N_18417,N_18524);
nand UO_186 (O_186,N_18104,N_19178);
or UO_187 (O_187,N_19951,N_19253);
nand UO_188 (O_188,N_18004,N_19731);
xor UO_189 (O_189,N_18354,N_19145);
xor UO_190 (O_190,N_19383,N_18776);
nand UO_191 (O_191,N_19415,N_18333);
and UO_192 (O_192,N_18992,N_18403);
nand UO_193 (O_193,N_19571,N_19222);
nand UO_194 (O_194,N_19537,N_18296);
nand UO_195 (O_195,N_18553,N_18536);
nor UO_196 (O_196,N_19413,N_18763);
nand UO_197 (O_197,N_18672,N_18781);
and UO_198 (O_198,N_18739,N_18055);
or UO_199 (O_199,N_19088,N_19738);
or UO_200 (O_200,N_18986,N_19539);
or UO_201 (O_201,N_18245,N_18268);
nand UO_202 (O_202,N_19275,N_18416);
nand UO_203 (O_203,N_18603,N_18653);
or UO_204 (O_204,N_19824,N_18228);
nor UO_205 (O_205,N_19255,N_19356);
or UO_206 (O_206,N_18188,N_19393);
nand UO_207 (O_207,N_18551,N_19942);
and UO_208 (O_208,N_19368,N_19045);
nor UO_209 (O_209,N_19124,N_19755);
and UO_210 (O_210,N_19729,N_18926);
or UO_211 (O_211,N_19642,N_19741);
and UO_212 (O_212,N_19001,N_18033);
nor UO_213 (O_213,N_18758,N_19258);
or UO_214 (O_214,N_18859,N_19133);
or UO_215 (O_215,N_18220,N_18024);
and UO_216 (O_216,N_19727,N_19697);
nand UO_217 (O_217,N_18532,N_19074);
nand UO_218 (O_218,N_19336,N_19011);
or UO_219 (O_219,N_18575,N_18619);
nor UO_220 (O_220,N_18402,N_19529);
nor UO_221 (O_221,N_18373,N_18325);
or UO_222 (O_222,N_19041,N_18222);
and UO_223 (O_223,N_18153,N_19881);
nor UO_224 (O_224,N_18780,N_18737);
or UO_225 (O_225,N_18460,N_18053);
xnor UO_226 (O_226,N_18624,N_18847);
and UO_227 (O_227,N_18794,N_19656);
or UO_228 (O_228,N_19212,N_19059);
nor UO_229 (O_229,N_19540,N_19420);
nor UO_230 (O_230,N_18289,N_19712);
xnor UO_231 (O_231,N_19180,N_18625);
or UO_232 (O_232,N_19384,N_19422);
and UO_233 (O_233,N_19114,N_19882);
nand UO_234 (O_234,N_18933,N_19379);
nor UO_235 (O_235,N_19550,N_18185);
nor UO_236 (O_236,N_19655,N_18559);
nand UO_237 (O_237,N_18400,N_19784);
or UO_238 (O_238,N_19099,N_19193);
nand UO_239 (O_239,N_19284,N_19127);
xor UO_240 (O_240,N_18425,N_19139);
nor UO_241 (O_241,N_19442,N_18800);
xnor UO_242 (O_242,N_19473,N_19721);
or UO_243 (O_243,N_19106,N_19475);
and UO_244 (O_244,N_18943,N_18555);
nand UO_245 (O_245,N_19171,N_19032);
nor UO_246 (O_246,N_18510,N_19719);
or UO_247 (O_247,N_19497,N_19692);
nor UO_248 (O_248,N_19000,N_18131);
and UO_249 (O_249,N_19135,N_19866);
nand UO_250 (O_250,N_19138,N_19447);
or UO_251 (O_251,N_19119,N_18218);
and UO_252 (O_252,N_19781,N_19204);
and UO_253 (O_253,N_19810,N_18852);
or UO_254 (O_254,N_19343,N_18076);
and UO_255 (O_255,N_19894,N_18286);
and UO_256 (O_256,N_18730,N_18212);
and UO_257 (O_257,N_19989,N_19392);
nand UO_258 (O_258,N_19599,N_19657);
or UO_259 (O_259,N_19611,N_19425);
and UO_260 (O_260,N_19026,N_18766);
and UO_261 (O_261,N_19630,N_18649);
nand UO_262 (O_262,N_19143,N_18151);
and UO_263 (O_263,N_19022,N_18399);
nor UO_264 (O_264,N_18815,N_18741);
nor UO_265 (O_265,N_18881,N_19995);
nor UO_266 (O_266,N_19759,N_18818);
or UO_267 (O_267,N_19378,N_18261);
nand UO_268 (O_268,N_19962,N_18991);
nand UO_269 (O_269,N_18216,N_18235);
or UO_270 (O_270,N_18946,N_18043);
nand UO_271 (O_271,N_19693,N_18918);
nand UO_272 (O_272,N_19405,N_19696);
or UO_273 (O_273,N_19769,N_18178);
or UO_274 (O_274,N_18810,N_19563);
nor UO_275 (O_275,N_18172,N_18196);
and UO_276 (O_276,N_19199,N_19756);
or UO_277 (O_277,N_19313,N_18346);
or UO_278 (O_278,N_18194,N_19862);
nor UO_279 (O_279,N_18045,N_18948);
or UO_280 (O_280,N_18560,N_18383);
nor UO_281 (O_281,N_19932,N_18720);
xor UO_282 (O_282,N_18044,N_19018);
or UO_283 (O_283,N_18490,N_18260);
nand UO_284 (O_284,N_19441,N_18458);
nand UO_285 (O_285,N_19132,N_19645);
nand UO_286 (O_286,N_19247,N_19073);
and UO_287 (O_287,N_18319,N_19154);
or UO_288 (O_288,N_19128,N_19554);
nand UO_289 (O_289,N_19454,N_18539);
and UO_290 (O_290,N_18449,N_19934);
nor UO_291 (O_291,N_18389,N_19748);
xnor UO_292 (O_292,N_19113,N_18935);
or UO_293 (O_293,N_18784,N_18543);
and UO_294 (O_294,N_19533,N_19566);
and UO_295 (O_295,N_19924,N_18028);
and UO_296 (O_296,N_19793,N_19897);
and UO_297 (O_297,N_19933,N_18256);
or UO_298 (O_298,N_19968,N_18467);
nor UO_299 (O_299,N_19403,N_18914);
and UO_300 (O_300,N_19353,N_19847);
nor UO_301 (O_301,N_19842,N_18191);
or UO_302 (O_302,N_18176,N_18824);
nor UO_303 (O_303,N_19845,N_19164);
xnor UO_304 (O_304,N_19876,N_18225);
or UO_305 (O_305,N_19463,N_18743);
and UO_306 (O_306,N_19971,N_19218);
nor UO_307 (O_307,N_18595,N_19051);
nor UO_308 (O_308,N_19990,N_19049);
and UO_309 (O_309,N_19799,N_19264);
nor UO_310 (O_310,N_19492,N_18203);
nand UO_311 (O_311,N_19198,N_18356);
or UO_312 (O_312,N_19725,N_18645);
nand UO_313 (O_313,N_19899,N_18310);
nor UO_314 (O_314,N_19764,N_19270);
and UO_315 (O_315,N_19237,N_19902);
or UO_316 (O_316,N_18368,N_19580);
or UO_317 (O_317,N_18727,N_18793);
xor UO_318 (O_318,N_18929,N_18707);
or UO_319 (O_319,N_18685,N_18052);
nand UO_320 (O_320,N_19372,N_19448);
nor UO_321 (O_321,N_18157,N_18303);
or UO_322 (O_322,N_18917,N_19840);
nor UO_323 (O_323,N_19036,N_18114);
or UO_324 (O_324,N_19981,N_18288);
or UO_325 (O_325,N_19283,N_19584);
xnor UO_326 (O_326,N_18799,N_19790);
nor UO_327 (O_327,N_19151,N_19401);
nor UO_328 (O_328,N_18262,N_19010);
nand UO_329 (O_329,N_18775,N_18630);
nor UO_330 (O_330,N_19931,N_18081);
nand UO_331 (O_331,N_19109,N_19885);
nor UO_332 (O_332,N_18767,N_18495);
nand UO_333 (O_333,N_18819,N_18317);
xor UO_334 (O_334,N_18407,N_18849);
nand UO_335 (O_335,N_18953,N_19137);
and UO_336 (O_336,N_19192,N_18905);
or UO_337 (O_337,N_18982,N_19558);
nand UO_338 (O_338,N_19144,N_19216);
nor UO_339 (O_339,N_19233,N_19742);
nand UO_340 (O_340,N_19146,N_18294);
and UO_341 (O_341,N_18406,N_18657);
nand UO_342 (O_342,N_19958,N_19708);
nand UO_343 (O_343,N_19081,N_18071);
or UO_344 (O_344,N_18825,N_19573);
xor UO_345 (O_345,N_19245,N_19337);
xor UO_346 (O_346,N_19063,N_19295);
or UO_347 (O_347,N_19483,N_19939);
and UO_348 (O_348,N_19925,N_19838);
or UO_349 (O_349,N_18877,N_19169);
xor UO_350 (O_350,N_18058,N_18121);
nor UO_351 (O_351,N_19600,N_18522);
or UO_352 (O_352,N_19837,N_18841);
nor UO_353 (O_353,N_18126,N_19466);
and UO_354 (O_354,N_19299,N_18866);
nor UO_355 (O_355,N_19841,N_18264);
and UO_356 (O_356,N_18814,N_19798);
or UO_357 (O_357,N_18099,N_19345);
nand UO_358 (O_358,N_19339,N_19228);
or UO_359 (O_359,N_19574,N_18136);
and UO_360 (O_360,N_19888,N_18390);
nand UO_361 (O_361,N_19244,N_19324);
and UO_362 (O_362,N_18913,N_18086);
xnor UO_363 (O_363,N_19775,N_18934);
nor UO_364 (O_364,N_19659,N_18263);
and UO_365 (O_365,N_19994,N_18230);
xor UO_366 (O_366,N_18738,N_18979);
nor UO_367 (O_367,N_18796,N_18896);
nand UO_368 (O_368,N_19978,N_19512);
and UO_369 (O_369,N_18702,N_19895);
and UO_370 (O_370,N_18718,N_19271);
nor UO_371 (O_371,N_19648,N_19315);
xor UO_372 (O_372,N_19879,N_19886);
and UO_373 (O_373,N_19538,N_18387);
nand UO_374 (O_374,N_19631,N_19647);
or UO_375 (O_375,N_19498,N_19224);
nor UO_376 (O_376,N_18186,N_19367);
or UO_377 (O_377,N_18623,N_18311);
and UO_378 (O_378,N_19358,N_18457);
or UO_379 (O_379,N_18880,N_18778);
xor UO_380 (O_380,N_19825,N_19078);
nand UO_381 (O_381,N_18298,N_19832);
nor UO_382 (O_382,N_18805,N_18010);
or UO_383 (O_383,N_18285,N_19773);
nor UO_384 (O_384,N_18820,N_19072);
nor UO_385 (O_385,N_18654,N_19223);
nor UO_386 (O_386,N_18549,N_18688);
nand UO_387 (O_387,N_19188,N_18535);
nor UO_388 (O_388,N_19201,N_19433);
or UO_389 (O_389,N_18088,N_19831);
nand UO_390 (O_390,N_18427,N_18827);
nor UO_391 (O_391,N_18326,N_18503);
or UO_392 (O_392,N_18062,N_18195);
and UO_393 (O_393,N_19516,N_19700);
and UO_394 (O_394,N_18474,N_18314);
xor UO_395 (O_395,N_19189,N_19919);
nand UO_396 (O_396,N_18258,N_19250);
or UO_397 (O_397,N_18374,N_18960);
and UO_398 (O_398,N_18864,N_19804);
or UO_399 (O_399,N_18572,N_19122);
nand UO_400 (O_400,N_19575,N_18855);
and UO_401 (O_401,N_18110,N_19377);
nor UO_402 (O_402,N_19640,N_18723);
nor UO_403 (O_403,N_19003,N_19520);
nor UO_404 (O_404,N_19287,N_19646);
or UO_405 (O_405,N_18711,N_19753);
nor UO_406 (O_406,N_19046,N_19411);
nor UO_407 (O_407,N_18789,N_19998);
nand UO_408 (O_408,N_19077,N_18764);
or UO_409 (O_409,N_19963,N_18372);
xnor UO_410 (O_410,N_18909,N_19568);
or UO_411 (O_411,N_18716,N_19555);
or UO_412 (O_412,N_19084,N_18330);
and UO_413 (O_413,N_18011,N_19791);
xor UO_414 (O_414,N_18808,N_19310);
nand UO_415 (O_415,N_18838,N_18939);
or UO_416 (O_416,N_19546,N_19543);
nor UO_417 (O_417,N_18152,N_19726);
and UO_418 (O_418,N_18391,N_18027);
nor UO_419 (O_419,N_19965,N_18475);
nor UO_420 (O_420,N_19265,N_19382);
nand UO_421 (O_421,N_19964,N_19843);
or UO_422 (O_422,N_18695,N_18208);
and UO_423 (O_423,N_18629,N_19907);
or UO_424 (O_424,N_18471,N_18976);
or UO_425 (O_425,N_18969,N_19955);
or UO_426 (O_426,N_18890,N_18677);
or UO_427 (O_427,N_19565,N_18284);
or UO_428 (O_428,N_18751,N_18574);
xnor UO_429 (O_429,N_18893,N_19110);
nand UO_430 (O_430,N_19262,N_18385);
nor UO_431 (O_431,N_19163,N_18250);
nor UO_432 (O_432,N_18394,N_19733);
and UO_433 (O_433,N_18921,N_19588);
nor UO_434 (O_434,N_18545,N_18438);
or UO_435 (O_435,N_18660,N_19969);
and UO_436 (O_436,N_18513,N_18287);
and UO_437 (O_437,N_19535,N_19055);
nand UO_438 (O_438,N_18493,N_18065);
or UO_439 (O_439,N_19507,N_18032);
or UO_440 (O_440,N_19788,N_19746);
nand UO_441 (O_441,N_19455,N_19065);
or UO_442 (O_442,N_19848,N_18925);
or UO_443 (O_443,N_18962,N_18113);
nand UO_444 (O_444,N_19622,N_19960);
or UO_445 (O_445,N_18811,N_19159);
and UO_446 (O_446,N_18802,N_18997);
and UO_447 (O_447,N_19979,N_18204);
nor UO_448 (O_448,N_18401,N_19098);
and UO_449 (O_449,N_18981,N_18382);
and UO_450 (O_450,N_18430,N_18051);
nor UO_451 (O_451,N_18269,N_19235);
nand UO_452 (O_452,N_19174,N_19518);
nand UO_453 (O_453,N_19852,N_19654);
and UO_454 (O_454,N_19705,N_19190);
or UO_455 (O_455,N_18643,N_18462);
nand UO_456 (O_456,N_19490,N_18583);
nor UO_457 (O_457,N_18301,N_18608);
nor UO_458 (O_458,N_19846,N_19519);
nor UO_459 (O_459,N_18469,N_18111);
nor UO_460 (O_460,N_18304,N_18275);
or UO_461 (O_461,N_19038,N_19319);
nand UO_462 (O_462,N_19429,N_19682);
nor UO_463 (O_463,N_19445,N_19166);
or UO_464 (O_464,N_19140,N_18478);
or UO_465 (O_465,N_19883,N_19266);
nor UO_466 (O_466,N_18085,N_18082);
nor UO_467 (O_467,N_19306,N_19034);
and UO_468 (O_468,N_19102,N_19637);
or UO_469 (O_469,N_18988,N_18129);
or UO_470 (O_470,N_19461,N_18938);
or UO_471 (O_471,N_18607,N_19805);
or UO_472 (O_472,N_19966,N_18517);
or UO_473 (O_473,N_18352,N_19783);
and UO_474 (O_474,N_18243,N_19226);
or UO_475 (O_475,N_18145,N_18159);
nor UO_476 (O_476,N_19460,N_19735);
nor UO_477 (O_477,N_19118,N_18466);
nor UO_478 (O_478,N_19027,N_18839);
xnor UO_479 (O_479,N_19670,N_18323);
nand UO_480 (O_480,N_19056,N_19351);
nor UO_481 (O_481,N_19320,N_18117);
or UO_482 (O_482,N_18013,N_18334);
xor UO_483 (O_483,N_18002,N_19323);
and UO_484 (O_484,N_18958,N_18487);
or UO_485 (O_485,N_19663,N_18199);
nor UO_486 (O_486,N_19945,N_18163);
nand UO_487 (O_487,N_18005,N_19503);
and UO_488 (O_488,N_19017,N_18602);
xor UO_489 (O_489,N_19913,N_19120);
xor UO_490 (O_490,N_19569,N_18508);
nor UO_491 (O_491,N_19972,N_18489);
nor UO_492 (O_492,N_19822,N_18854);
and UO_493 (O_493,N_19153,N_19914);
nand UO_494 (O_494,N_18577,N_18106);
or UO_495 (O_495,N_19567,N_18167);
nor UO_496 (O_496,N_18928,N_19665);
nand UO_497 (O_497,N_18480,N_19892);
nand UO_498 (O_498,N_19016,N_18049);
nand UO_499 (O_499,N_18491,N_19173);
and UO_500 (O_500,N_19597,N_19954);
xnor UO_501 (O_501,N_18069,N_19157);
nor UO_502 (O_502,N_18857,N_18713);
nand UO_503 (O_503,N_19760,N_18377);
nand UO_504 (O_504,N_19623,N_18950);
nor UO_505 (O_505,N_18381,N_18107);
or UO_506 (O_506,N_18975,N_18347);
nor UO_507 (O_507,N_18529,N_18123);
or UO_508 (O_508,N_19186,N_18357);
or UO_509 (O_509,N_18994,N_19387);
and UO_510 (O_510,N_19147,N_19787);
nand UO_511 (O_511,N_18485,N_18056);
or UO_512 (O_512,N_19418,N_18419);
or UO_513 (O_513,N_19116,N_18492);
and UO_514 (O_514,N_18745,N_19395);
and UO_515 (O_515,N_18020,N_18744);
and UO_516 (O_516,N_19999,N_19005);
xor UO_517 (O_517,N_18740,N_19435);
nor UO_518 (O_518,N_18008,N_19097);
nor UO_519 (O_519,N_18848,N_18483);
nor UO_520 (O_520,N_18443,N_19710);
nand UO_521 (O_521,N_19814,N_18274);
and UO_522 (O_522,N_19111,N_18628);
or UO_523 (O_523,N_19472,N_19684);
and UO_524 (O_524,N_19404,N_19161);
xnor UO_525 (O_525,N_18965,N_18434);
or UO_526 (O_526,N_18320,N_18100);
and UO_527 (O_527,N_19349,N_18414);
xor UO_528 (O_528,N_18901,N_18143);
nand UO_529 (O_529,N_19844,N_19855);
xor UO_530 (O_530,N_18388,N_18064);
nor UO_531 (O_531,N_18754,N_19355);
xor UO_532 (O_532,N_18618,N_18812);
nand UO_533 (O_533,N_19040,N_19916);
and UO_534 (O_534,N_19004,N_19863);
or UO_535 (O_535,N_19946,N_18108);
nand UO_536 (O_536,N_18622,N_19471);
and UO_537 (O_537,N_18959,N_19241);
nand UO_538 (O_538,N_19796,N_19887);
nand UO_539 (O_539,N_19332,N_19465);
xor UO_540 (O_540,N_18936,N_18889);
nand UO_541 (O_541,N_19758,N_19261);
nor UO_542 (O_542,N_18063,N_19723);
or UO_543 (O_543,N_19083,N_19777);
and UO_544 (O_544,N_19976,N_18830);
nand UO_545 (O_545,N_19695,N_18253);
and UO_546 (O_546,N_18599,N_19718);
and UO_547 (O_547,N_19282,N_18765);
nor UO_548 (O_548,N_19514,N_18362);
nand UO_549 (O_549,N_19008,N_19603);
nor UO_550 (O_550,N_18931,N_18278);
or UO_551 (O_551,N_19660,N_19286);
nor UO_552 (O_552,N_18442,N_19606);
and UO_553 (O_553,N_18234,N_18729);
or UO_554 (O_554,N_19373,N_19691);
nor UO_555 (O_555,N_19365,N_18360);
and UO_556 (O_556,N_18160,N_19702);
nor UO_557 (O_557,N_19196,N_19058);
and UO_558 (O_558,N_18338,N_18512);
nor UO_559 (O_559,N_19864,N_19536);
xnor UO_560 (O_560,N_18174,N_18125);
and UO_561 (O_561,N_19576,N_19988);
and UO_562 (O_562,N_19249,N_18379);
and UO_563 (O_563,N_18714,N_18783);
or UO_564 (O_564,N_18650,N_18748);
or UO_565 (O_565,N_18676,N_19851);
and UO_566 (O_566,N_18898,N_19903);
or UO_567 (O_567,N_19479,N_18656);
nor UO_568 (O_568,N_18837,N_18217);
and UO_569 (O_569,N_18973,N_18433);
or UO_570 (O_570,N_18242,N_19427);
nand UO_571 (O_571,N_19912,N_18116);
nand UO_572 (O_572,N_18558,N_18755);
and UO_573 (O_573,N_18428,N_18501);
nand UO_574 (O_574,N_19406,N_19294);
and UO_575 (O_575,N_18206,N_19898);
nand UO_576 (O_576,N_18641,N_19184);
or UO_577 (O_577,N_19187,N_18435);
and UO_578 (O_578,N_18828,N_18687);
and UO_579 (O_579,N_19101,N_18506);
xnor UO_580 (O_580,N_18639,N_19480);
nand UO_581 (O_581,N_19744,N_19452);
or UO_582 (O_582,N_18180,N_18530);
or UO_583 (O_583,N_19602,N_18080);
nor UO_584 (O_584,N_19308,N_19944);
and UO_585 (O_585,N_18514,N_19200);
nor UO_586 (O_586,N_19240,N_18232);
and UO_587 (O_587,N_18970,N_18804);
xnor UO_588 (O_588,N_19205,N_18418);
xor UO_589 (O_589,N_18615,N_19493);
nor UO_590 (O_590,N_18257,N_18681);
and UO_591 (O_591,N_18604,N_18998);
and UO_592 (O_592,N_18709,N_19047);
or UO_593 (O_593,N_19220,N_18722);
or UO_594 (O_594,N_18885,N_19486);
or UO_595 (O_595,N_18207,N_19767);
and UO_596 (O_596,N_18568,N_18486);
nor UO_597 (O_597,N_18021,N_18170);
and UO_598 (O_598,N_19348,N_18464);
and UO_599 (O_599,N_19002,N_19321);
xnor UO_600 (O_600,N_19381,N_19407);
nand UO_601 (O_601,N_18272,N_18012);
xnor UO_602 (O_602,N_18912,N_18279);
nand UO_603 (O_603,N_18141,N_19750);
nand UO_604 (O_604,N_19984,N_19836);
nor UO_605 (O_605,N_18952,N_18440);
and UO_606 (O_606,N_18964,N_18614);
and UO_607 (O_607,N_19181,N_19312);
xnor UO_608 (O_608,N_19311,N_19873);
or UO_609 (O_609,N_18850,N_19947);
nor UO_610 (O_610,N_18534,N_18299);
and UO_611 (O_611,N_19160,N_19556);
xnor UO_612 (O_612,N_18924,N_19679);
and UO_613 (O_613,N_19191,N_18397);
nor UO_614 (O_614,N_18426,N_19079);
or UO_615 (O_615,N_19162,N_19779);
nand UO_616 (O_616,N_18408,N_18833);
nand UO_617 (O_617,N_18923,N_19397);
or UO_618 (O_618,N_18697,N_19009);
nand UO_619 (O_619,N_18198,N_19532);
xnor UO_620 (O_620,N_19214,N_18972);
nand UO_621 (O_621,N_18456,N_19553);
and UO_622 (O_622,N_18586,N_19961);
or UO_623 (O_623,N_19437,N_18875);
or UO_624 (O_624,N_18576,N_19506);
or UO_625 (O_625,N_18251,N_19096);
nand UO_626 (O_626,N_18101,N_18856);
nand UO_627 (O_627,N_18365,N_19436);
nor UO_628 (O_628,N_19410,N_19105);
or UO_629 (O_629,N_18942,N_18597);
and UO_630 (O_630,N_18957,N_19375);
nand UO_631 (O_631,N_19149,N_18105);
and UO_632 (O_632,N_19053,N_18211);
or UO_633 (O_633,N_18733,N_19130);
nor UO_634 (O_634,N_18951,N_18761);
or UO_635 (O_635,N_18694,N_18963);
or UO_636 (O_636,N_19714,N_19835);
and UO_637 (O_637,N_18581,N_19782);
nor UO_638 (O_638,N_18290,N_18306);
nor UO_639 (O_639,N_18692,N_18878);
nor UO_640 (O_640,N_19751,N_19970);
nor UO_641 (O_641,N_18627,N_18331);
xnor UO_642 (O_642,N_18017,N_18562);
or UO_643 (O_643,N_19687,N_19856);
nor UO_644 (O_644,N_19430,N_18149);
and UO_645 (O_645,N_19982,N_19509);
or UO_646 (O_646,N_18861,N_19707);
xnor UO_647 (O_647,N_19526,N_18659);
xnor UO_648 (O_648,N_18384,N_19006);
nand UO_649 (O_649,N_19068,N_18083);
nor UO_650 (O_650,N_18705,N_19478);
or UO_651 (O_651,N_18787,N_18034);
xnor UO_652 (O_652,N_18750,N_19578);
nor UO_653 (O_653,N_18834,N_18911);
nand UO_654 (O_654,N_18717,N_18473);
or UO_655 (O_655,N_19280,N_18454);
nand UO_656 (O_656,N_19100,N_18915);
nor UO_657 (O_657,N_19115,N_19820);
and UO_658 (O_658,N_19414,N_18060);
and UO_659 (O_659,N_19949,N_19941);
nor UO_660 (O_660,N_18415,N_19182);
or UO_661 (O_661,N_19818,N_18822);
and UO_662 (O_662,N_18040,N_18700);
nor UO_663 (O_663,N_19168,N_18666);
or UO_664 (O_664,N_19614,N_19385);
or UO_665 (O_665,N_19357,N_18404);
nand UO_666 (O_666,N_18351,N_18183);
nand UO_667 (O_667,N_18785,N_19551);
nand UO_668 (O_668,N_18461,N_18297);
xnor UO_669 (O_669,N_18588,N_19316);
and UO_670 (O_670,N_19938,N_18871);
or UO_671 (O_671,N_19354,N_18321);
nor UO_672 (O_672,N_19671,N_19242);
or UO_673 (O_673,N_18715,N_19142);
xor UO_674 (O_674,N_18987,N_19044);
or UO_675 (O_675,N_19394,N_18521);
nor UO_676 (O_676,N_19564,N_19470);
nor UO_677 (O_677,N_19915,N_18840);
xnor UO_678 (O_678,N_19595,N_19039);
nand UO_679 (O_679,N_18768,N_19829);
nand UO_680 (O_680,N_19803,N_18318);
or UO_681 (O_681,N_19030,N_19366);
and UO_682 (O_682,N_18118,N_19906);
nand UO_683 (O_683,N_19878,N_19293);
and UO_684 (O_684,N_18706,N_18436);
nor UO_685 (O_685,N_19952,N_19239);
and UO_686 (O_686,N_18900,N_19527);
and UO_687 (O_687,N_18255,N_18696);
and UO_688 (O_688,N_19967,N_18520);
and UO_689 (O_689,N_18315,N_19274);
or UO_690 (O_690,N_18993,N_18444);
and UO_691 (O_691,N_18252,N_19291);
nor UO_692 (O_692,N_18862,N_18197);
or UO_693 (O_693,N_18844,N_19632);
xor UO_694 (O_694,N_18148,N_19789);
or UO_695 (O_695,N_18999,N_19314);
or UO_696 (O_696,N_19624,N_18749);
nand UO_697 (O_697,N_18479,N_18124);
and UO_698 (O_698,N_19633,N_18214);
xnor UO_699 (O_699,N_18668,N_18966);
nor UO_700 (O_700,N_19890,N_18171);
xor UO_701 (O_701,N_18616,N_18983);
or UO_702 (O_702,N_19269,N_18316);
or UO_703 (O_703,N_18779,N_19296);
and UO_704 (O_704,N_19389,N_18359);
nand UO_705 (O_705,N_18329,N_18447);
nor UO_706 (O_706,N_18519,N_19080);
or UO_707 (O_707,N_19720,N_18821);
nor UO_708 (O_708,N_19991,N_18161);
or UO_709 (O_709,N_18350,N_19402);
nand UO_710 (O_710,N_18210,N_19093);
nor UO_711 (O_711,N_18669,N_18894);
or UO_712 (O_712,N_19300,N_18092);
nand UO_713 (O_713,N_18638,N_19112);
nor UO_714 (O_714,N_18348,N_18396);
and UO_715 (O_715,N_19075,N_18712);
or UO_716 (O_716,N_18974,N_18531);
nand UO_717 (O_717,N_19158,N_18001);
xor UO_718 (O_718,N_19704,N_19683);
and UO_719 (O_719,N_18016,N_19901);
and UO_720 (O_720,N_19409,N_19482);
xnor UO_721 (O_721,N_18876,N_19983);
and UO_722 (O_722,N_19524,N_19548);
xor UO_723 (O_723,N_19802,N_19202);
and UO_724 (O_724,N_18596,N_19658);
and UO_725 (O_725,N_18693,N_19674);
and UO_726 (O_726,N_18556,N_19807);
nand UO_727 (O_727,N_19500,N_19468);
and UO_728 (O_728,N_18410,N_19359);
nor UO_729 (O_729,N_19612,N_18613);
nor UO_730 (O_730,N_19736,N_18860);
or UO_731 (O_731,N_19728,N_19675);
xor UO_732 (O_732,N_19986,N_18146);
nor UO_733 (O_733,N_19155,N_19342);
or UO_734 (O_734,N_18190,N_19668);
and UO_735 (O_735,N_18193,N_18544);
nand UO_736 (O_736,N_18455,N_18546);
nor UO_737 (O_737,N_18807,N_19501);
nor UO_738 (O_738,N_18309,N_19221);
or UO_739 (O_739,N_18561,N_19638);
and UO_740 (O_740,N_19685,N_19197);
and UO_741 (O_741,N_18634,N_19872);
nand UO_742 (O_742,N_18658,N_18899);
nor UO_743 (O_743,N_19061,N_19371);
nand UO_744 (O_744,N_19066,N_19238);
nand UO_745 (O_745,N_19309,N_19910);
and UO_746 (O_746,N_18511,N_18642);
nor UO_747 (O_747,N_19908,N_19950);
xor UO_748 (O_748,N_19396,N_19369);
and UO_749 (O_749,N_18393,N_18584);
xnor UO_750 (O_750,N_18593,N_19667);
and UO_751 (O_751,N_18324,N_18378);
nand UO_752 (O_752,N_19057,N_19281);
or UO_753 (O_753,N_18732,N_18431);
and UO_754 (O_754,N_19476,N_19303);
nand UO_755 (O_755,N_18910,N_19335);
and UO_756 (O_756,N_19352,N_19167);
xnor UO_757 (O_757,N_18240,N_19801);
nand UO_758 (O_758,N_19921,N_19698);
or UO_759 (O_759,N_19399,N_18978);
or UO_760 (O_760,N_18571,N_19254);
nand UO_761 (O_761,N_18254,N_19975);
or UO_762 (O_762,N_18366,N_19330);
and UO_763 (O_763,N_18842,N_19706);
or UO_764 (O_764,N_18184,N_19628);
nor UO_765 (O_765,N_18984,N_18704);
and UO_766 (O_766,N_18022,N_18031);
nor UO_767 (O_767,N_18036,N_19859);
nand UO_768 (O_768,N_19771,N_18238);
or UO_769 (O_769,N_18267,N_18147);
nor UO_770 (O_770,N_19666,N_19257);
nand UO_771 (O_771,N_18355,N_18537);
or UO_772 (O_772,N_18578,N_19530);
nand UO_773 (O_773,N_18237,N_19834);
and UO_774 (O_774,N_18579,N_19256);
or UO_775 (O_775,N_18470,N_18686);
and UO_776 (O_776,N_19450,N_19792);
and UO_777 (O_777,N_19929,N_18569);
or UO_778 (O_778,N_18019,N_18481);
or UO_779 (O_779,N_19601,N_19037);
or UO_780 (O_780,N_18179,N_19940);
and UO_781 (O_781,N_18465,N_19997);
xor UO_782 (O_782,N_19092,N_18797);
or UO_783 (O_783,N_18585,N_18523);
nor UO_784 (O_784,N_18610,N_18648);
xnor UO_785 (O_785,N_18221,N_19816);
and UO_786 (O_786,N_19117,N_18189);
and UO_787 (O_787,N_18209,N_18533);
and UO_788 (O_788,N_19585,N_18054);
and UO_789 (O_789,N_18155,N_19304);
xor UO_790 (O_790,N_19141,N_18496);
and UO_791 (O_791,N_18173,N_19778);
or UO_792 (O_792,N_18867,N_19485);
or UO_793 (O_793,N_18753,N_19935);
nand UO_794 (O_794,N_19896,N_19690);
nor UO_795 (O_795,N_18484,N_19740);
or UO_796 (O_796,N_18865,N_18742);
or UO_797 (O_797,N_18026,N_18835);
nor UO_798 (O_798,N_18795,N_19776);
nand UO_799 (O_799,N_19517,N_18380);
and UO_800 (O_800,N_19094,N_19625);
nor UO_801 (O_801,N_18061,N_19481);
nor UO_802 (O_802,N_19930,N_19338);
nor UO_803 (O_803,N_19877,N_18922);
nand UO_804 (O_804,N_18412,N_18169);
and UO_805 (O_805,N_18500,N_19326);
or UO_806 (O_806,N_18369,N_19673);
nand UO_807 (O_807,N_19278,N_19715);
nand UO_808 (O_808,N_18236,N_18594);
or UO_809 (O_809,N_18295,N_18652);
or UO_810 (O_810,N_19206,N_18809);
or UO_811 (O_811,N_18869,N_18332);
and UO_812 (O_812,N_19082,N_18003);
nor UO_813 (O_813,N_19772,N_19579);
or UO_814 (O_814,N_19035,N_18168);
nand UO_815 (O_815,N_19664,N_19795);
nand UO_816 (O_816,N_18611,N_18451);
nand UO_817 (O_817,N_18229,N_19277);
and UO_818 (O_818,N_19340,N_19502);
or UO_819 (O_819,N_18187,N_19031);
and UO_820 (O_820,N_18670,N_19826);
nand UO_821 (O_821,N_19652,N_18079);
xnor UO_822 (O_822,N_19297,N_19757);
and UO_823 (O_823,N_18786,N_18617);
nor UO_824 (O_824,N_18095,N_19985);
nor UO_825 (O_825,N_18902,N_19749);
nand UO_826 (O_826,N_18736,N_18906);
nor UO_827 (O_827,N_19607,N_19431);
nand UO_828 (O_828,N_18476,N_19386);
and UO_829 (O_829,N_18308,N_19451);
xor UO_830 (O_830,N_18074,N_19494);
nor UO_831 (O_831,N_19528,N_19722);
and UO_832 (O_832,N_19273,N_19959);
nand UO_833 (O_833,N_18018,N_18971);
nor UO_834 (O_834,N_18895,N_18006);
and UO_835 (O_835,N_19703,N_19544);
and UO_836 (O_836,N_19689,N_19618);
nor UO_837 (O_837,N_19849,N_19987);
xnor UO_838 (O_838,N_19421,N_18046);
nand UO_839 (O_839,N_19869,N_19376);
or UO_840 (O_840,N_19918,N_18882);
and UO_841 (O_841,N_18698,N_19152);
nor UO_842 (O_842,N_19020,N_18477);
nor UO_843 (O_843,N_19806,N_19484);
nor UO_844 (O_844,N_18293,N_18202);
nor UO_845 (O_845,N_19823,N_18259);
nor UO_846 (O_846,N_18029,N_18395);
and UO_847 (O_847,N_18039,N_19713);
nor UO_848 (O_848,N_19609,N_19219);
nor UO_849 (O_849,N_18683,N_18248);
nand UO_850 (O_850,N_18916,N_19513);
or UO_851 (O_851,N_19794,N_18233);
nand UO_852 (O_852,N_18453,N_18164);
and UO_853 (O_853,N_19488,N_19496);
nor UO_854 (O_854,N_19412,N_19577);
nor UO_855 (O_855,N_18482,N_18515);
or UO_856 (O_856,N_19752,N_19267);
and UO_857 (O_857,N_19209,N_19217);
or UO_858 (O_858,N_18949,N_19562);
or UO_859 (O_859,N_18552,N_19508);
nor UO_860 (O_860,N_18181,N_19762);
or UO_861 (O_861,N_18853,N_19511);
nand UO_862 (O_862,N_18265,N_19541);
nand UO_863 (O_863,N_19651,N_18823);
nor UO_864 (O_864,N_18874,N_19457);
or UO_865 (O_865,N_18525,N_18542);
or UO_866 (O_866,N_18540,N_19583);
xor UO_867 (O_867,N_18879,N_19331);
nor UO_868 (O_868,N_19616,N_18884);
nor UO_869 (O_869,N_18990,N_19268);
nand UO_870 (O_870,N_19688,N_18226);
or UO_871 (O_871,N_19604,N_18089);
nand UO_872 (O_872,N_19260,N_18612);
and UO_873 (O_873,N_19833,N_18836);
xor UO_874 (O_874,N_19570,N_19318);
nor UO_875 (O_875,N_19333,N_18422);
nor UO_876 (O_876,N_19107,N_18655);
nand UO_877 (O_877,N_19811,N_19649);
or UO_878 (O_878,N_18664,N_19592);
nor UO_879 (O_879,N_18175,N_19210);
and UO_880 (O_880,N_18283,N_18239);
and UO_881 (O_881,N_18342,N_18445);
xor UO_882 (O_882,N_19076,N_18708);
nand UO_883 (O_883,N_18115,N_18135);
and UO_884 (O_884,N_19370,N_18000);
nand UO_885 (O_885,N_18725,N_18112);
nor UO_886 (O_886,N_18133,N_19943);
or UO_887 (O_887,N_18941,N_19770);
nor UO_888 (O_888,N_19716,N_18746);
and UO_889 (O_889,N_19423,N_18361);
nand UO_890 (O_890,N_19301,N_19417);
and UO_891 (O_891,N_19765,N_18829);
and UO_892 (O_892,N_18041,N_19867);
nand UO_893 (O_893,N_19305,N_19126);
nor UO_894 (O_894,N_18920,N_18219);
and UO_895 (O_895,N_19043,N_18448);
nor UO_896 (O_896,N_19865,N_19272);
nor UO_897 (O_897,N_18724,N_18621);
nor UO_898 (O_898,N_18084,N_18507);
nor UO_899 (O_899,N_19854,N_19085);
nor UO_900 (O_900,N_19179,N_18227);
xor UO_901 (O_901,N_18587,N_18504);
or UO_902 (O_902,N_18420,N_19542);
nor UO_903 (O_903,N_19534,N_19650);
and UO_904 (O_904,N_18068,N_19786);
and UO_905 (O_905,N_18048,N_18826);
nor UO_906 (O_906,N_19288,N_18582);
xor UO_907 (O_907,N_18547,N_18488);
nor UO_908 (O_908,N_18450,N_18947);
nor UO_909 (O_909,N_18241,N_18047);
or UO_910 (O_910,N_19123,N_19928);
nand UO_911 (O_911,N_18703,N_19996);
or UO_912 (O_912,N_19086,N_19070);
and UO_913 (O_913,N_18782,N_18592);
nand UO_914 (O_914,N_19023,N_18846);
or UO_915 (O_915,N_18432,N_18701);
or UO_916 (O_916,N_19858,N_18038);
nand UO_917 (O_917,N_18025,N_18363);
nor UO_918 (O_918,N_18120,N_18472);
nand UO_919 (O_919,N_19596,N_18719);
nand UO_920 (O_920,N_18336,N_18570);
or UO_921 (O_921,N_18305,N_19813);
or UO_922 (O_922,N_19432,N_18600);
or UO_923 (O_923,N_19870,N_19346);
nand UO_924 (O_924,N_18142,N_19136);
or UO_925 (O_925,N_18015,N_19893);
nand UO_926 (O_926,N_19709,N_18509);
and UO_927 (O_927,N_18271,N_18154);
nand UO_928 (O_928,N_18127,N_19467);
or UO_929 (O_929,N_19711,N_18674);
nand UO_930 (O_930,N_19582,N_19621);
nor UO_931 (O_931,N_19871,N_18968);
nand UO_932 (O_932,N_18328,N_18985);
nand UO_933 (O_933,N_19211,N_19948);
nor UO_934 (O_934,N_18077,N_18337);
and UO_935 (O_935,N_19185,N_18816);
nor UO_936 (O_936,N_18813,N_18955);
xnor UO_937 (O_937,N_18518,N_19891);
and UO_938 (O_938,N_19434,N_19499);
and UO_939 (O_939,N_18312,N_19292);
or UO_940 (O_940,N_18014,N_19232);
nor UO_941 (O_941,N_19605,N_18516);
and UO_942 (O_942,N_18940,N_18682);
and UO_943 (O_943,N_19613,N_19505);
and UO_944 (O_944,N_19523,N_18364);
or UO_945 (O_945,N_19446,N_18892);
nand UO_946 (O_946,N_18777,N_18791);
nor UO_947 (O_947,N_18845,N_18094);
nand UO_948 (O_948,N_18747,N_19374);
nor UO_949 (O_949,N_19586,N_19634);
and UO_950 (O_950,N_18678,N_19491);
and UO_951 (O_951,N_18721,N_19730);
nor UO_952 (O_952,N_18710,N_19808);
and UO_953 (O_953,N_19279,N_19920);
and UO_954 (O_954,N_19042,N_18249);
xnor UO_955 (O_955,N_19014,N_19900);
and UO_956 (O_956,N_19572,N_18130);
and UO_957 (O_957,N_18980,N_19510);
xnor UO_958 (O_958,N_19048,N_18102);
and UO_959 (O_959,N_18371,N_18887);
nor UO_960 (O_960,N_18035,N_18554);
nor UO_961 (O_961,N_18165,N_18070);
nor UO_962 (O_962,N_19992,N_18424);
xnor UO_963 (O_963,N_19416,N_19923);
and UO_964 (O_964,N_18760,N_18140);
nand UO_965 (O_965,N_18446,N_18313);
or UO_966 (O_966,N_19774,N_19449);
and UO_967 (O_967,N_19104,N_18996);
or UO_968 (O_968,N_19868,N_18367);
nand UO_969 (O_969,N_19552,N_18067);
nand UO_970 (O_970,N_19177,N_18567);
or UO_971 (O_971,N_19438,N_19091);
nand UO_972 (O_972,N_19581,N_19194);
nor UO_973 (O_973,N_19560,N_19231);
nand UO_974 (O_974,N_18421,N_18954);
nor UO_975 (O_975,N_19800,N_19821);
and UO_976 (O_976,N_19263,N_19426);
nand UO_977 (O_977,N_18956,N_19626);
and UO_978 (O_978,N_19641,N_18735);
and UO_979 (O_979,N_18601,N_18930);
nor UO_980 (O_980,N_18690,N_19150);
nor UO_981 (O_981,N_18073,N_18007);
or UO_982 (O_982,N_19739,N_19067);
nor UO_983 (O_983,N_19225,N_18497);
nor UO_984 (O_984,N_19464,N_18409);
nand UO_985 (O_985,N_18977,N_18103);
nor UO_986 (O_986,N_18752,N_19644);
nor UO_987 (O_987,N_19766,N_19183);
or UO_988 (O_988,N_19860,N_18667);
and UO_989 (O_989,N_19361,N_18803);
nor UO_990 (O_990,N_19400,N_18851);
xnor UO_991 (O_991,N_18870,N_18631);
nor UO_992 (O_992,N_18907,N_18675);
nand UO_993 (O_993,N_18817,N_19248);
or UO_994 (O_994,N_18066,N_19643);
and UO_995 (O_995,N_19328,N_18452);
nor UO_996 (O_996,N_18528,N_18349);
nor UO_997 (O_997,N_19089,N_19747);
or UO_998 (O_998,N_18322,N_19129);
xnor UO_999 (O_999,N_18097,N_19131);
nand UO_1000 (O_1000,N_18045,N_18137);
and UO_1001 (O_1001,N_19635,N_18944);
and UO_1002 (O_1002,N_19986,N_18175);
and UO_1003 (O_1003,N_18702,N_19660);
nand UO_1004 (O_1004,N_18707,N_18419);
or UO_1005 (O_1005,N_18920,N_19255);
or UO_1006 (O_1006,N_19272,N_18297);
and UO_1007 (O_1007,N_19151,N_19149);
and UO_1008 (O_1008,N_19346,N_19839);
or UO_1009 (O_1009,N_18072,N_18576);
nor UO_1010 (O_1010,N_18118,N_18629);
nor UO_1011 (O_1011,N_19080,N_18189);
xnor UO_1012 (O_1012,N_18336,N_19780);
xnor UO_1013 (O_1013,N_18397,N_18678);
nand UO_1014 (O_1014,N_19666,N_18541);
nand UO_1015 (O_1015,N_19951,N_19793);
nand UO_1016 (O_1016,N_18149,N_19539);
nand UO_1017 (O_1017,N_18622,N_18964);
xnor UO_1018 (O_1018,N_18578,N_19558);
or UO_1019 (O_1019,N_18345,N_18595);
nand UO_1020 (O_1020,N_19493,N_19249);
and UO_1021 (O_1021,N_18931,N_19509);
nand UO_1022 (O_1022,N_18633,N_18419);
nor UO_1023 (O_1023,N_19112,N_19991);
nand UO_1024 (O_1024,N_18733,N_18351);
xnor UO_1025 (O_1025,N_18332,N_19301);
nand UO_1026 (O_1026,N_18604,N_18178);
or UO_1027 (O_1027,N_19427,N_18101);
or UO_1028 (O_1028,N_19611,N_18490);
or UO_1029 (O_1029,N_19353,N_19193);
nand UO_1030 (O_1030,N_18885,N_19368);
nand UO_1031 (O_1031,N_19255,N_18446);
nand UO_1032 (O_1032,N_19594,N_18883);
nor UO_1033 (O_1033,N_18928,N_18794);
nand UO_1034 (O_1034,N_19036,N_19552);
nand UO_1035 (O_1035,N_18952,N_18411);
and UO_1036 (O_1036,N_19323,N_19322);
or UO_1037 (O_1037,N_19531,N_19944);
nor UO_1038 (O_1038,N_18223,N_19911);
xnor UO_1039 (O_1039,N_18291,N_18321);
or UO_1040 (O_1040,N_18099,N_18119);
and UO_1041 (O_1041,N_19490,N_19458);
or UO_1042 (O_1042,N_18022,N_19666);
xnor UO_1043 (O_1043,N_18180,N_18062);
and UO_1044 (O_1044,N_18217,N_19076);
xor UO_1045 (O_1045,N_18805,N_19347);
or UO_1046 (O_1046,N_19942,N_19884);
or UO_1047 (O_1047,N_18338,N_18162);
xnor UO_1048 (O_1048,N_19367,N_19937);
and UO_1049 (O_1049,N_19474,N_19233);
and UO_1050 (O_1050,N_19694,N_18141);
nand UO_1051 (O_1051,N_18099,N_19248);
nand UO_1052 (O_1052,N_18501,N_18656);
or UO_1053 (O_1053,N_19140,N_18680);
and UO_1054 (O_1054,N_19773,N_19264);
and UO_1055 (O_1055,N_18164,N_18607);
xnor UO_1056 (O_1056,N_18097,N_18697);
nor UO_1057 (O_1057,N_18109,N_18552);
and UO_1058 (O_1058,N_18296,N_18007);
or UO_1059 (O_1059,N_19410,N_19535);
xnor UO_1060 (O_1060,N_18574,N_19150);
nor UO_1061 (O_1061,N_19977,N_18242);
nand UO_1062 (O_1062,N_18531,N_19205);
or UO_1063 (O_1063,N_19622,N_19567);
nand UO_1064 (O_1064,N_18259,N_18645);
nor UO_1065 (O_1065,N_18019,N_18075);
nand UO_1066 (O_1066,N_18166,N_19002);
or UO_1067 (O_1067,N_18079,N_18070);
or UO_1068 (O_1068,N_19923,N_19842);
or UO_1069 (O_1069,N_18485,N_18857);
nor UO_1070 (O_1070,N_19529,N_18138);
nor UO_1071 (O_1071,N_18318,N_18153);
nor UO_1072 (O_1072,N_19317,N_19788);
nor UO_1073 (O_1073,N_18991,N_18231);
or UO_1074 (O_1074,N_18482,N_19171);
nor UO_1075 (O_1075,N_18284,N_19731);
nand UO_1076 (O_1076,N_19307,N_18266);
nand UO_1077 (O_1077,N_19619,N_19313);
nor UO_1078 (O_1078,N_18981,N_19684);
and UO_1079 (O_1079,N_19946,N_18837);
or UO_1080 (O_1080,N_19625,N_19758);
nor UO_1081 (O_1081,N_19960,N_19186);
nand UO_1082 (O_1082,N_18188,N_18012);
and UO_1083 (O_1083,N_19111,N_19767);
or UO_1084 (O_1084,N_19424,N_19131);
xor UO_1085 (O_1085,N_19602,N_19428);
and UO_1086 (O_1086,N_19812,N_18319);
and UO_1087 (O_1087,N_18197,N_18799);
or UO_1088 (O_1088,N_18029,N_18028);
nand UO_1089 (O_1089,N_19054,N_19474);
and UO_1090 (O_1090,N_18799,N_18901);
or UO_1091 (O_1091,N_18851,N_18166);
nand UO_1092 (O_1092,N_18733,N_19684);
nor UO_1093 (O_1093,N_19873,N_18205);
nor UO_1094 (O_1094,N_18850,N_19629);
or UO_1095 (O_1095,N_19780,N_18599);
and UO_1096 (O_1096,N_19706,N_19107);
nand UO_1097 (O_1097,N_18305,N_19533);
xor UO_1098 (O_1098,N_18928,N_19660);
and UO_1099 (O_1099,N_18365,N_18771);
nand UO_1100 (O_1100,N_19513,N_18175);
and UO_1101 (O_1101,N_18605,N_19820);
or UO_1102 (O_1102,N_19346,N_19619);
nand UO_1103 (O_1103,N_18470,N_18715);
nor UO_1104 (O_1104,N_19994,N_19869);
nor UO_1105 (O_1105,N_19034,N_18267);
nand UO_1106 (O_1106,N_19871,N_18330);
and UO_1107 (O_1107,N_19980,N_19103);
nand UO_1108 (O_1108,N_19763,N_19102);
xor UO_1109 (O_1109,N_18265,N_19349);
xnor UO_1110 (O_1110,N_19078,N_18250);
nand UO_1111 (O_1111,N_18967,N_19699);
and UO_1112 (O_1112,N_19515,N_19966);
xor UO_1113 (O_1113,N_18387,N_18469);
or UO_1114 (O_1114,N_19209,N_18214);
xor UO_1115 (O_1115,N_18953,N_18378);
or UO_1116 (O_1116,N_18666,N_18677);
or UO_1117 (O_1117,N_18390,N_18393);
xnor UO_1118 (O_1118,N_19734,N_18894);
and UO_1119 (O_1119,N_18104,N_18850);
nand UO_1120 (O_1120,N_19746,N_19643);
or UO_1121 (O_1121,N_18569,N_18855);
or UO_1122 (O_1122,N_19207,N_19595);
nor UO_1123 (O_1123,N_18554,N_19924);
or UO_1124 (O_1124,N_18653,N_19889);
nand UO_1125 (O_1125,N_19057,N_18811);
nor UO_1126 (O_1126,N_18262,N_18782);
and UO_1127 (O_1127,N_19303,N_19771);
and UO_1128 (O_1128,N_19610,N_19264);
and UO_1129 (O_1129,N_18331,N_18471);
and UO_1130 (O_1130,N_19847,N_18506);
and UO_1131 (O_1131,N_19683,N_19409);
nand UO_1132 (O_1132,N_19126,N_18347);
nand UO_1133 (O_1133,N_18874,N_19835);
nor UO_1134 (O_1134,N_18152,N_18206);
nand UO_1135 (O_1135,N_18096,N_19078);
nor UO_1136 (O_1136,N_19450,N_19281);
xor UO_1137 (O_1137,N_19935,N_18784);
nand UO_1138 (O_1138,N_18696,N_18148);
xnor UO_1139 (O_1139,N_19410,N_18291);
xnor UO_1140 (O_1140,N_19197,N_19104);
nor UO_1141 (O_1141,N_18163,N_18898);
or UO_1142 (O_1142,N_19011,N_19319);
nand UO_1143 (O_1143,N_18588,N_19091);
nand UO_1144 (O_1144,N_19309,N_19217);
or UO_1145 (O_1145,N_18077,N_18762);
or UO_1146 (O_1146,N_19154,N_19406);
or UO_1147 (O_1147,N_18621,N_18709);
nor UO_1148 (O_1148,N_19055,N_19737);
nor UO_1149 (O_1149,N_18426,N_18336);
and UO_1150 (O_1150,N_19543,N_18769);
nand UO_1151 (O_1151,N_18127,N_19925);
and UO_1152 (O_1152,N_19054,N_18450);
and UO_1153 (O_1153,N_18562,N_19624);
nand UO_1154 (O_1154,N_19271,N_19357);
nand UO_1155 (O_1155,N_18359,N_18015);
nand UO_1156 (O_1156,N_19038,N_18703);
nand UO_1157 (O_1157,N_18155,N_18003);
xor UO_1158 (O_1158,N_19388,N_19598);
and UO_1159 (O_1159,N_19256,N_19559);
nor UO_1160 (O_1160,N_18683,N_18206);
and UO_1161 (O_1161,N_19528,N_19355);
and UO_1162 (O_1162,N_19210,N_19979);
nand UO_1163 (O_1163,N_19128,N_18092);
nor UO_1164 (O_1164,N_18066,N_19993);
nand UO_1165 (O_1165,N_19393,N_18528);
nand UO_1166 (O_1166,N_19699,N_19881);
and UO_1167 (O_1167,N_18898,N_19909);
nand UO_1168 (O_1168,N_19704,N_19031);
or UO_1169 (O_1169,N_18315,N_19487);
xor UO_1170 (O_1170,N_19933,N_19337);
nor UO_1171 (O_1171,N_18781,N_18694);
xnor UO_1172 (O_1172,N_19592,N_18803);
nor UO_1173 (O_1173,N_18083,N_19405);
or UO_1174 (O_1174,N_19027,N_19569);
nand UO_1175 (O_1175,N_19223,N_19579);
nor UO_1176 (O_1176,N_19053,N_18679);
or UO_1177 (O_1177,N_18316,N_19284);
or UO_1178 (O_1178,N_18555,N_18860);
xor UO_1179 (O_1179,N_19506,N_19075);
and UO_1180 (O_1180,N_19973,N_18798);
nand UO_1181 (O_1181,N_18360,N_18996);
xor UO_1182 (O_1182,N_19263,N_19816);
or UO_1183 (O_1183,N_18551,N_18427);
nor UO_1184 (O_1184,N_19941,N_19602);
or UO_1185 (O_1185,N_19011,N_19417);
nand UO_1186 (O_1186,N_19932,N_18266);
nand UO_1187 (O_1187,N_18073,N_19565);
nand UO_1188 (O_1188,N_18186,N_19265);
xnor UO_1189 (O_1189,N_19671,N_19206);
nand UO_1190 (O_1190,N_18123,N_19523);
and UO_1191 (O_1191,N_19014,N_19243);
and UO_1192 (O_1192,N_18547,N_19974);
nor UO_1193 (O_1193,N_18583,N_18440);
nand UO_1194 (O_1194,N_18819,N_18607);
nand UO_1195 (O_1195,N_19643,N_19499);
nand UO_1196 (O_1196,N_18322,N_18306);
and UO_1197 (O_1197,N_19955,N_18114);
and UO_1198 (O_1198,N_19145,N_19299);
nor UO_1199 (O_1199,N_18159,N_19137);
and UO_1200 (O_1200,N_19404,N_19687);
or UO_1201 (O_1201,N_18552,N_19221);
nor UO_1202 (O_1202,N_18716,N_19450);
nor UO_1203 (O_1203,N_18759,N_19412);
nor UO_1204 (O_1204,N_18316,N_18989);
nand UO_1205 (O_1205,N_19302,N_18342);
and UO_1206 (O_1206,N_19045,N_18087);
nor UO_1207 (O_1207,N_18481,N_18354);
nand UO_1208 (O_1208,N_19582,N_19847);
nor UO_1209 (O_1209,N_18485,N_18558);
nor UO_1210 (O_1210,N_18606,N_18295);
and UO_1211 (O_1211,N_19702,N_19151);
and UO_1212 (O_1212,N_18170,N_19584);
xnor UO_1213 (O_1213,N_18425,N_18903);
and UO_1214 (O_1214,N_19621,N_18944);
xor UO_1215 (O_1215,N_18146,N_18675);
xnor UO_1216 (O_1216,N_18769,N_18613);
nor UO_1217 (O_1217,N_19785,N_19985);
xnor UO_1218 (O_1218,N_18427,N_18167);
or UO_1219 (O_1219,N_18901,N_18953);
or UO_1220 (O_1220,N_18301,N_19248);
or UO_1221 (O_1221,N_18742,N_19823);
nand UO_1222 (O_1222,N_19405,N_18084);
and UO_1223 (O_1223,N_19221,N_19749);
or UO_1224 (O_1224,N_18647,N_18944);
xnor UO_1225 (O_1225,N_19224,N_19303);
xnor UO_1226 (O_1226,N_19951,N_19338);
nor UO_1227 (O_1227,N_18716,N_19530);
nor UO_1228 (O_1228,N_19843,N_18165);
or UO_1229 (O_1229,N_18461,N_19760);
and UO_1230 (O_1230,N_19113,N_19562);
or UO_1231 (O_1231,N_18675,N_18919);
nor UO_1232 (O_1232,N_18413,N_18676);
nor UO_1233 (O_1233,N_18226,N_18337);
and UO_1234 (O_1234,N_18782,N_18557);
nand UO_1235 (O_1235,N_18447,N_19531);
nor UO_1236 (O_1236,N_19590,N_19824);
xor UO_1237 (O_1237,N_18963,N_18446);
nor UO_1238 (O_1238,N_19615,N_18411);
and UO_1239 (O_1239,N_18762,N_19134);
nand UO_1240 (O_1240,N_19943,N_19951);
nand UO_1241 (O_1241,N_18402,N_19046);
xnor UO_1242 (O_1242,N_18439,N_18500);
nor UO_1243 (O_1243,N_18196,N_19485);
and UO_1244 (O_1244,N_18071,N_19194);
or UO_1245 (O_1245,N_18452,N_19381);
nand UO_1246 (O_1246,N_19253,N_19525);
and UO_1247 (O_1247,N_19346,N_18225);
or UO_1248 (O_1248,N_19504,N_19505);
and UO_1249 (O_1249,N_18795,N_18428);
or UO_1250 (O_1250,N_18215,N_18521);
nand UO_1251 (O_1251,N_18736,N_19576);
xnor UO_1252 (O_1252,N_18311,N_19865);
nand UO_1253 (O_1253,N_19659,N_19796);
nor UO_1254 (O_1254,N_19966,N_18351);
and UO_1255 (O_1255,N_19986,N_19824);
nor UO_1256 (O_1256,N_18011,N_18498);
and UO_1257 (O_1257,N_18274,N_18600);
and UO_1258 (O_1258,N_19554,N_18967);
nand UO_1259 (O_1259,N_18110,N_18609);
nand UO_1260 (O_1260,N_18491,N_18467);
nand UO_1261 (O_1261,N_19260,N_19592);
and UO_1262 (O_1262,N_19786,N_18415);
and UO_1263 (O_1263,N_18818,N_19374);
nor UO_1264 (O_1264,N_18832,N_18036);
nor UO_1265 (O_1265,N_19673,N_19427);
xnor UO_1266 (O_1266,N_19348,N_18083);
xnor UO_1267 (O_1267,N_18222,N_18314);
nand UO_1268 (O_1268,N_18890,N_19369);
nand UO_1269 (O_1269,N_18219,N_19504);
nor UO_1270 (O_1270,N_19330,N_18828);
nand UO_1271 (O_1271,N_19988,N_18759);
xnor UO_1272 (O_1272,N_19722,N_19306);
and UO_1273 (O_1273,N_18427,N_18235);
nand UO_1274 (O_1274,N_18913,N_18833);
nor UO_1275 (O_1275,N_18511,N_18711);
nand UO_1276 (O_1276,N_18102,N_18490);
nand UO_1277 (O_1277,N_19357,N_18715);
xor UO_1278 (O_1278,N_19534,N_19474);
nand UO_1279 (O_1279,N_19313,N_19429);
xor UO_1280 (O_1280,N_18628,N_18791);
and UO_1281 (O_1281,N_19449,N_19167);
xnor UO_1282 (O_1282,N_19386,N_19999);
and UO_1283 (O_1283,N_19521,N_19520);
or UO_1284 (O_1284,N_19496,N_19808);
or UO_1285 (O_1285,N_19954,N_18414);
xor UO_1286 (O_1286,N_18348,N_18604);
or UO_1287 (O_1287,N_18827,N_19466);
xnor UO_1288 (O_1288,N_19036,N_18982);
or UO_1289 (O_1289,N_18272,N_18866);
xor UO_1290 (O_1290,N_19229,N_18598);
and UO_1291 (O_1291,N_18555,N_18319);
nor UO_1292 (O_1292,N_18778,N_18756);
nand UO_1293 (O_1293,N_18235,N_19853);
and UO_1294 (O_1294,N_18043,N_19915);
and UO_1295 (O_1295,N_18663,N_18497);
nand UO_1296 (O_1296,N_18668,N_19635);
nor UO_1297 (O_1297,N_19949,N_18378);
nand UO_1298 (O_1298,N_18301,N_19588);
and UO_1299 (O_1299,N_19188,N_19768);
nand UO_1300 (O_1300,N_19349,N_19252);
nor UO_1301 (O_1301,N_18487,N_18671);
or UO_1302 (O_1302,N_19975,N_19619);
nor UO_1303 (O_1303,N_18396,N_19183);
or UO_1304 (O_1304,N_19911,N_18861);
and UO_1305 (O_1305,N_19285,N_18029);
nor UO_1306 (O_1306,N_19672,N_19309);
or UO_1307 (O_1307,N_18902,N_18339);
nand UO_1308 (O_1308,N_19067,N_18757);
nor UO_1309 (O_1309,N_19039,N_19684);
nand UO_1310 (O_1310,N_19303,N_19380);
nor UO_1311 (O_1311,N_19861,N_18847);
nand UO_1312 (O_1312,N_19601,N_19279);
nand UO_1313 (O_1313,N_18715,N_19361);
or UO_1314 (O_1314,N_18727,N_18290);
nand UO_1315 (O_1315,N_18309,N_19443);
or UO_1316 (O_1316,N_19526,N_18512);
and UO_1317 (O_1317,N_19874,N_19201);
xnor UO_1318 (O_1318,N_18991,N_18571);
nor UO_1319 (O_1319,N_18230,N_18897);
or UO_1320 (O_1320,N_18637,N_19919);
xnor UO_1321 (O_1321,N_19689,N_19966);
nor UO_1322 (O_1322,N_19082,N_18925);
xnor UO_1323 (O_1323,N_19594,N_19190);
or UO_1324 (O_1324,N_19363,N_19046);
nand UO_1325 (O_1325,N_19802,N_19534);
nand UO_1326 (O_1326,N_18421,N_19111);
nor UO_1327 (O_1327,N_18288,N_19940);
and UO_1328 (O_1328,N_19165,N_19487);
xnor UO_1329 (O_1329,N_19496,N_19453);
nor UO_1330 (O_1330,N_19106,N_18018);
nor UO_1331 (O_1331,N_19689,N_18178);
and UO_1332 (O_1332,N_18943,N_19444);
nand UO_1333 (O_1333,N_18387,N_18560);
nor UO_1334 (O_1334,N_18498,N_19727);
nor UO_1335 (O_1335,N_18028,N_18094);
or UO_1336 (O_1336,N_18834,N_19905);
and UO_1337 (O_1337,N_18528,N_19960);
nand UO_1338 (O_1338,N_18525,N_18822);
nor UO_1339 (O_1339,N_19465,N_19041);
xnor UO_1340 (O_1340,N_18517,N_19455);
xnor UO_1341 (O_1341,N_18402,N_18643);
and UO_1342 (O_1342,N_19312,N_19389);
xor UO_1343 (O_1343,N_19798,N_18056);
xnor UO_1344 (O_1344,N_18561,N_19828);
and UO_1345 (O_1345,N_18775,N_18213);
xnor UO_1346 (O_1346,N_18754,N_19274);
and UO_1347 (O_1347,N_19433,N_18607);
xnor UO_1348 (O_1348,N_19753,N_18085);
xnor UO_1349 (O_1349,N_18206,N_19142);
xnor UO_1350 (O_1350,N_18881,N_18852);
and UO_1351 (O_1351,N_18872,N_18143);
nor UO_1352 (O_1352,N_19792,N_19790);
or UO_1353 (O_1353,N_19334,N_19695);
and UO_1354 (O_1354,N_18210,N_18324);
nor UO_1355 (O_1355,N_19248,N_18833);
nor UO_1356 (O_1356,N_19679,N_19975);
or UO_1357 (O_1357,N_19427,N_19496);
nand UO_1358 (O_1358,N_19732,N_19234);
nor UO_1359 (O_1359,N_18702,N_19248);
nor UO_1360 (O_1360,N_19490,N_18304);
and UO_1361 (O_1361,N_19775,N_18465);
or UO_1362 (O_1362,N_18529,N_18160);
nand UO_1363 (O_1363,N_18748,N_18283);
or UO_1364 (O_1364,N_18189,N_19859);
nand UO_1365 (O_1365,N_18652,N_18267);
xnor UO_1366 (O_1366,N_18649,N_18395);
nand UO_1367 (O_1367,N_18030,N_19965);
nand UO_1368 (O_1368,N_19604,N_19111);
or UO_1369 (O_1369,N_19741,N_19847);
nor UO_1370 (O_1370,N_19591,N_18906);
or UO_1371 (O_1371,N_18774,N_19317);
and UO_1372 (O_1372,N_18595,N_18909);
nand UO_1373 (O_1373,N_19994,N_18769);
or UO_1374 (O_1374,N_18094,N_18595);
and UO_1375 (O_1375,N_18273,N_19918);
nor UO_1376 (O_1376,N_19025,N_18079);
nor UO_1377 (O_1377,N_18318,N_19476);
and UO_1378 (O_1378,N_19064,N_19606);
or UO_1379 (O_1379,N_18323,N_19372);
nor UO_1380 (O_1380,N_19762,N_18843);
nand UO_1381 (O_1381,N_18763,N_18994);
nor UO_1382 (O_1382,N_19361,N_19098);
nand UO_1383 (O_1383,N_19197,N_18716);
or UO_1384 (O_1384,N_19553,N_18544);
or UO_1385 (O_1385,N_19268,N_19991);
and UO_1386 (O_1386,N_19380,N_18207);
nand UO_1387 (O_1387,N_18351,N_18190);
nor UO_1388 (O_1388,N_18317,N_19818);
and UO_1389 (O_1389,N_19963,N_19750);
or UO_1390 (O_1390,N_18635,N_19439);
nor UO_1391 (O_1391,N_18371,N_18701);
xnor UO_1392 (O_1392,N_18626,N_18715);
nor UO_1393 (O_1393,N_18675,N_18318);
nand UO_1394 (O_1394,N_19359,N_19387);
nor UO_1395 (O_1395,N_19626,N_18783);
nand UO_1396 (O_1396,N_18525,N_19506);
nor UO_1397 (O_1397,N_19737,N_18456);
nand UO_1398 (O_1398,N_18343,N_18761);
or UO_1399 (O_1399,N_19782,N_19899);
and UO_1400 (O_1400,N_19717,N_19345);
or UO_1401 (O_1401,N_18196,N_19129);
xnor UO_1402 (O_1402,N_19775,N_18229);
and UO_1403 (O_1403,N_18936,N_19505);
or UO_1404 (O_1404,N_18374,N_18175);
or UO_1405 (O_1405,N_19473,N_18449);
nor UO_1406 (O_1406,N_19571,N_18756);
or UO_1407 (O_1407,N_18798,N_18170);
or UO_1408 (O_1408,N_19448,N_18666);
or UO_1409 (O_1409,N_18028,N_19964);
nand UO_1410 (O_1410,N_18064,N_18427);
nand UO_1411 (O_1411,N_19082,N_18574);
nand UO_1412 (O_1412,N_18532,N_19304);
or UO_1413 (O_1413,N_18149,N_19682);
or UO_1414 (O_1414,N_19696,N_19477);
or UO_1415 (O_1415,N_19544,N_19903);
nand UO_1416 (O_1416,N_18388,N_19231);
nand UO_1417 (O_1417,N_19856,N_19280);
xor UO_1418 (O_1418,N_18627,N_19585);
nand UO_1419 (O_1419,N_18113,N_18790);
nor UO_1420 (O_1420,N_19217,N_19551);
or UO_1421 (O_1421,N_19093,N_19292);
nand UO_1422 (O_1422,N_18045,N_18386);
and UO_1423 (O_1423,N_18707,N_19484);
or UO_1424 (O_1424,N_19440,N_18672);
nor UO_1425 (O_1425,N_19235,N_19666);
nor UO_1426 (O_1426,N_18781,N_19119);
nor UO_1427 (O_1427,N_18498,N_19545);
xor UO_1428 (O_1428,N_19684,N_18264);
nor UO_1429 (O_1429,N_19103,N_18591);
nor UO_1430 (O_1430,N_18340,N_18886);
or UO_1431 (O_1431,N_19418,N_18929);
nor UO_1432 (O_1432,N_18016,N_19357);
nand UO_1433 (O_1433,N_18942,N_18137);
and UO_1434 (O_1434,N_19274,N_18640);
and UO_1435 (O_1435,N_19785,N_19892);
nor UO_1436 (O_1436,N_19724,N_18624);
or UO_1437 (O_1437,N_18174,N_18759);
or UO_1438 (O_1438,N_18511,N_19061);
and UO_1439 (O_1439,N_18538,N_18490);
and UO_1440 (O_1440,N_18794,N_19616);
or UO_1441 (O_1441,N_19468,N_19224);
or UO_1442 (O_1442,N_19355,N_19786);
or UO_1443 (O_1443,N_19013,N_19277);
and UO_1444 (O_1444,N_18047,N_18843);
nand UO_1445 (O_1445,N_19192,N_19525);
and UO_1446 (O_1446,N_19920,N_18051);
nand UO_1447 (O_1447,N_19079,N_19774);
or UO_1448 (O_1448,N_18754,N_18316);
or UO_1449 (O_1449,N_18519,N_18039);
and UO_1450 (O_1450,N_18441,N_19316);
or UO_1451 (O_1451,N_18160,N_19435);
nand UO_1452 (O_1452,N_19279,N_19026);
or UO_1453 (O_1453,N_19185,N_19043);
xnor UO_1454 (O_1454,N_18698,N_19077);
and UO_1455 (O_1455,N_19421,N_18015);
nor UO_1456 (O_1456,N_18497,N_18077);
or UO_1457 (O_1457,N_19908,N_18531);
nand UO_1458 (O_1458,N_19266,N_19209);
nand UO_1459 (O_1459,N_19736,N_19789);
and UO_1460 (O_1460,N_19037,N_18240);
and UO_1461 (O_1461,N_18615,N_19037);
or UO_1462 (O_1462,N_19538,N_18243);
xnor UO_1463 (O_1463,N_18515,N_19162);
nor UO_1464 (O_1464,N_19410,N_18608);
xnor UO_1465 (O_1465,N_19135,N_18347);
nor UO_1466 (O_1466,N_18247,N_19716);
xor UO_1467 (O_1467,N_18499,N_19843);
or UO_1468 (O_1468,N_19989,N_19039);
nor UO_1469 (O_1469,N_18381,N_19855);
or UO_1470 (O_1470,N_19131,N_19733);
or UO_1471 (O_1471,N_18544,N_19410);
and UO_1472 (O_1472,N_19484,N_18052);
or UO_1473 (O_1473,N_18456,N_18988);
and UO_1474 (O_1474,N_19066,N_19059);
xor UO_1475 (O_1475,N_18211,N_19760);
nand UO_1476 (O_1476,N_18741,N_19731);
nor UO_1477 (O_1477,N_18492,N_18335);
nand UO_1478 (O_1478,N_19319,N_19779);
and UO_1479 (O_1479,N_19954,N_18667);
and UO_1480 (O_1480,N_18613,N_19492);
nor UO_1481 (O_1481,N_18560,N_18723);
xnor UO_1482 (O_1482,N_18630,N_19994);
xnor UO_1483 (O_1483,N_18547,N_18361);
nand UO_1484 (O_1484,N_18673,N_18227);
nand UO_1485 (O_1485,N_18456,N_18529);
nand UO_1486 (O_1486,N_18811,N_18863);
nand UO_1487 (O_1487,N_19486,N_19161);
nand UO_1488 (O_1488,N_19957,N_18155);
or UO_1489 (O_1489,N_19053,N_19372);
and UO_1490 (O_1490,N_18895,N_18401);
nand UO_1491 (O_1491,N_19180,N_19595);
or UO_1492 (O_1492,N_18142,N_19385);
and UO_1493 (O_1493,N_19607,N_18913);
nand UO_1494 (O_1494,N_19183,N_19093);
or UO_1495 (O_1495,N_19300,N_18974);
or UO_1496 (O_1496,N_18836,N_19184);
nand UO_1497 (O_1497,N_19857,N_19286);
xnor UO_1498 (O_1498,N_19439,N_19586);
and UO_1499 (O_1499,N_19900,N_19757);
nor UO_1500 (O_1500,N_19168,N_19238);
nor UO_1501 (O_1501,N_19345,N_18766);
or UO_1502 (O_1502,N_19329,N_18053);
nor UO_1503 (O_1503,N_18868,N_19108);
and UO_1504 (O_1504,N_19472,N_18886);
nor UO_1505 (O_1505,N_18958,N_19166);
nand UO_1506 (O_1506,N_18964,N_19588);
nand UO_1507 (O_1507,N_18904,N_19037);
nor UO_1508 (O_1508,N_19035,N_18830);
and UO_1509 (O_1509,N_18718,N_19386);
nor UO_1510 (O_1510,N_19991,N_19194);
nor UO_1511 (O_1511,N_18577,N_19913);
nand UO_1512 (O_1512,N_18766,N_19120);
or UO_1513 (O_1513,N_18555,N_19342);
or UO_1514 (O_1514,N_18786,N_19985);
or UO_1515 (O_1515,N_18044,N_19005);
nand UO_1516 (O_1516,N_19999,N_18943);
or UO_1517 (O_1517,N_18717,N_19177);
nand UO_1518 (O_1518,N_19880,N_18858);
nor UO_1519 (O_1519,N_18975,N_18638);
nand UO_1520 (O_1520,N_18115,N_18930);
nand UO_1521 (O_1521,N_19430,N_18047);
and UO_1522 (O_1522,N_18942,N_19085);
nor UO_1523 (O_1523,N_18618,N_18983);
and UO_1524 (O_1524,N_19626,N_19943);
xnor UO_1525 (O_1525,N_18157,N_18938);
and UO_1526 (O_1526,N_18513,N_18427);
xor UO_1527 (O_1527,N_18779,N_19077);
or UO_1528 (O_1528,N_19325,N_19704);
xor UO_1529 (O_1529,N_18140,N_19275);
nand UO_1530 (O_1530,N_18407,N_18848);
xor UO_1531 (O_1531,N_19854,N_18502);
xor UO_1532 (O_1532,N_19710,N_18018);
nand UO_1533 (O_1533,N_18760,N_18721);
and UO_1534 (O_1534,N_18168,N_18427);
or UO_1535 (O_1535,N_19268,N_19409);
nand UO_1536 (O_1536,N_18742,N_19230);
or UO_1537 (O_1537,N_19784,N_18277);
or UO_1538 (O_1538,N_18116,N_18995);
nor UO_1539 (O_1539,N_19768,N_19936);
xnor UO_1540 (O_1540,N_18986,N_19608);
nor UO_1541 (O_1541,N_18979,N_19602);
nand UO_1542 (O_1542,N_18607,N_18003);
nand UO_1543 (O_1543,N_19090,N_18044);
xnor UO_1544 (O_1544,N_19929,N_19832);
or UO_1545 (O_1545,N_19029,N_18614);
nand UO_1546 (O_1546,N_18738,N_18840);
nand UO_1547 (O_1547,N_18204,N_18441);
or UO_1548 (O_1548,N_19705,N_18993);
or UO_1549 (O_1549,N_19663,N_18966);
and UO_1550 (O_1550,N_18802,N_19118);
or UO_1551 (O_1551,N_19716,N_19189);
and UO_1552 (O_1552,N_19967,N_19400);
nor UO_1553 (O_1553,N_19719,N_18499);
nand UO_1554 (O_1554,N_18248,N_18986);
and UO_1555 (O_1555,N_19681,N_18839);
nor UO_1556 (O_1556,N_18708,N_19179);
nor UO_1557 (O_1557,N_18025,N_19329);
nand UO_1558 (O_1558,N_19783,N_18952);
and UO_1559 (O_1559,N_18609,N_19398);
nor UO_1560 (O_1560,N_19754,N_19029);
and UO_1561 (O_1561,N_19071,N_18834);
or UO_1562 (O_1562,N_18589,N_19960);
nand UO_1563 (O_1563,N_19933,N_19228);
or UO_1564 (O_1564,N_18907,N_19968);
nand UO_1565 (O_1565,N_18663,N_19869);
xor UO_1566 (O_1566,N_18760,N_18467);
nor UO_1567 (O_1567,N_19110,N_18869);
nand UO_1568 (O_1568,N_19237,N_19368);
or UO_1569 (O_1569,N_19604,N_19531);
nor UO_1570 (O_1570,N_19324,N_19787);
or UO_1571 (O_1571,N_18946,N_19447);
and UO_1572 (O_1572,N_19768,N_19013);
xor UO_1573 (O_1573,N_19688,N_18356);
nand UO_1574 (O_1574,N_19024,N_18016);
xor UO_1575 (O_1575,N_19177,N_18533);
and UO_1576 (O_1576,N_18268,N_19956);
and UO_1577 (O_1577,N_19693,N_18133);
and UO_1578 (O_1578,N_19204,N_18025);
and UO_1579 (O_1579,N_18566,N_19380);
or UO_1580 (O_1580,N_19273,N_18526);
nand UO_1581 (O_1581,N_18041,N_18286);
nor UO_1582 (O_1582,N_18444,N_19681);
nor UO_1583 (O_1583,N_18138,N_19958);
nor UO_1584 (O_1584,N_18696,N_19728);
nand UO_1585 (O_1585,N_18366,N_18718);
nor UO_1586 (O_1586,N_19526,N_18570);
or UO_1587 (O_1587,N_18082,N_19767);
nor UO_1588 (O_1588,N_18097,N_18545);
or UO_1589 (O_1589,N_18663,N_18479);
nor UO_1590 (O_1590,N_19052,N_19331);
xor UO_1591 (O_1591,N_18947,N_19629);
or UO_1592 (O_1592,N_18970,N_19307);
and UO_1593 (O_1593,N_18258,N_19470);
or UO_1594 (O_1594,N_19756,N_18315);
or UO_1595 (O_1595,N_18373,N_19017);
or UO_1596 (O_1596,N_18717,N_19593);
or UO_1597 (O_1597,N_19618,N_18097);
xor UO_1598 (O_1598,N_18192,N_18739);
or UO_1599 (O_1599,N_19644,N_18568);
nand UO_1600 (O_1600,N_19104,N_19458);
nor UO_1601 (O_1601,N_19582,N_19577);
nor UO_1602 (O_1602,N_18755,N_18126);
nor UO_1603 (O_1603,N_18821,N_18931);
nor UO_1604 (O_1604,N_18518,N_18926);
nor UO_1605 (O_1605,N_19794,N_18283);
xor UO_1606 (O_1606,N_18542,N_18923);
and UO_1607 (O_1607,N_19695,N_19826);
nor UO_1608 (O_1608,N_18249,N_18763);
nand UO_1609 (O_1609,N_19049,N_19475);
or UO_1610 (O_1610,N_18528,N_19818);
nor UO_1611 (O_1611,N_19349,N_18954);
and UO_1612 (O_1612,N_19056,N_19625);
and UO_1613 (O_1613,N_18757,N_19035);
nand UO_1614 (O_1614,N_18039,N_18055);
nor UO_1615 (O_1615,N_19799,N_18889);
nor UO_1616 (O_1616,N_18640,N_18094);
or UO_1617 (O_1617,N_19227,N_19912);
nand UO_1618 (O_1618,N_18141,N_18491);
nand UO_1619 (O_1619,N_19548,N_19014);
and UO_1620 (O_1620,N_19824,N_18564);
or UO_1621 (O_1621,N_18406,N_18270);
nor UO_1622 (O_1622,N_19587,N_18879);
nor UO_1623 (O_1623,N_19236,N_19238);
xor UO_1624 (O_1624,N_19362,N_19333);
or UO_1625 (O_1625,N_18750,N_19958);
xor UO_1626 (O_1626,N_18054,N_19932);
or UO_1627 (O_1627,N_19242,N_18773);
or UO_1628 (O_1628,N_19003,N_18564);
or UO_1629 (O_1629,N_18508,N_19816);
nand UO_1630 (O_1630,N_18261,N_18326);
nor UO_1631 (O_1631,N_18099,N_19340);
xor UO_1632 (O_1632,N_19881,N_19629);
nand UO_1633 (O_1633,N_19702,N_19509);
xnor UO_1634 (O_1634,N_19364,N_18201);
nand UO_1635 (O_1635,N_18451,N_18099);
and UO_1636 (O_1636,N_19217,N_19937);
or UO_1637 (O_1637,N_19805,N_19149);
nand UO_1638 (O_1638,N_18556,N_19123);
nand UO_1639 (O_1639,N_19276,N_19704);
nor UO_1640 (O_1640,N_18358,N_18397);
or UO_1641 (O_1641,N_18768,N_18089);
and UO_1642 (O_1642,N_19603,N_19856);
nand UO_1643 (O_1643,N_19649,N_19905);
and UO_1644 (O_1644,N_18020,N_18178);
or UO_1645 (O_1645,N_18487,N_19074);
nor UO_1646 (O_1646,N_19089,N_19891);
nand UO_1647 (O_1647,N_19840,N_18199);
or UO_1648 (O_1648,N_18343,N_18739);
and UO_1649 (O_1649,N_18506,N_18008);
nor UO_1650 (O_1650,N_19973,N_19269);
and UO_1651 (O_1651,N_18997,N_18072);
nand UO_1652 (O_1652,N_19375,N_19918);
or UO_1653 (O_1653,N_18910,N_18328);
nor UO_1654 (O_1654,N_19757,N_18901);
and UO_1655 (O_1655,N_19247,N_19302);
xnor UO_1656 (O_1656,N_18302,N_19202);
nor UO_1657 (O_1657,N_19651,N_18633);
xor UO_1658 (O_1658,N_19998,N_19101);
and UO_1659 (O_1659,N_18821,N_19148);
or UO_1660 (O_1660,N_19084,N_19788);
nor UO_1661 (O_1661,N_18598,N_18344);
or UO_1662 (O_1662,N_19714,N_18020);
nor UO_1663 (O_1663,N_19049,N_18012);
nand UO_1664 (O_1664,N_19930,N_18126);
xor UO_1665 (O_1665,N_18809,N_19698);
or UO_1666 (O_1666,N_19437,N_19924);
and UO_1667 (O_1667,N_18210,N_19660);
or UO_1668 (O_1668,N_18899,N_19980);
nor UO_1669 (O_1669,N_19755,N_18821);
or UO_1670 (O_1670,N_19551,N_19320);
xnor UO_1671 (O_1671,N_18342,N_19479);
nand UO_1672 (O_1672,N_19499,N_19186);
nor UO_1673 (O_1673,N_19470,N_18801);
or UO_1674 (O_1674,N_19933,N_18928);
nand UO_1675 (O_1675,N_18090,N_19527);
nor UO_1676 (O_1676,N_18681,N_18861);
or UO_1677 (O_1677,N_18017,N_19759);
or UO_1678 (O_1678,N_19130,N_19785);
or UO_1679 (O_1679,N_18487,N_18995);
or UO_1680 (O_1680,N_18248,N_18669);
xnor UO_1681 (O_1681,N_19966,N_19096);
nor UO_1682 (O_1682,N_19728,N_18863);
nor UO_1683 (O_1683,N_19304,N_19302);
xnor UO_1684 (O_1684,N_19363,N_18413);
nor UO_1685 (O_1685,N_19327,N_18599);
xnor UO_1686 (O_1686,N_18512,N_18358);
or UO_1687 (O_1687,N_19959,N_19836);
nor UO_1688 (O_1688,N_18269,N_18416);
nand UO_1689 (O_1689,N_19031,N_19746);
nor UO_1690 (O_1690,N_18254,N_19268);
or UO_1691 (O_1691,N_19603,N_19612);
or UO_1692 (O_1692,N_18577,N_19453);
or UO_1693 (O_1693,N_19381,N_19939);
nand UO_1694 (O_1694,N_18277,N_18269);
nor UO_1695 (O_1695,N_19197,N_18583);
xnor UO_1696 (O_1696,N_18128,N_18200);
nor UO_1697 (O_1697,N_18440,N_19200);
nor UO_1698 (O_1698,N_18174,N_19993);
and UO_1699 (O_1699,N_18484,N_18603);
nand UO_1700 (O_1700,N_19040,N_18054);
nand UO_1701 (O_1701,N_18674,N_18036);
and UO_1702 (O_1702,N_18831,N_19207);
or UO_1703 (O_1703,N_18503,N_18022);
nand UO_1704 (O_1704,N_19849,N_18872);
nand UO_1705 (O_1705,N_19083,N_18990);
nor UO_1706 (O_1706,N_18342,N_18605);
nor UO_1707 (O_1707,N_19027,N_18435);
and UO_1708 (O_1708,N_19207,N_19571);
nand UO_1709 (O_1709,N_18403,N_19028);
nand UO_1710 (O_1710,N_18233,N_19985);
nor UO_1711 (O_1711,N_19384,N_19474);
or UO_1712 (O_1712,N_19990,N_19202);
or UO_1713 (O_1713,N_19488,N_19641);
or UO_1714 (O_1714,N_18059,N_18950);
nor UO_1715 (O_1715,N_19069,N_19972);
nand UO_1716 (O_1716,N_18229,N_19991);
nand UO_1717 (O_1717,N_19526,N_19384);
nor UO_1718 (O_1718,N_18558,N_19914);
and UO_1719 (O_1719,N_19751,N_18804);
nand UO_1720 (O_1720,N_19146,N_18657);
or UO_1721 (O_1721,N_19158,N_19830);
nand UO_1722 (O_1722,N_19915,N_18684);
xor UO_1723 (O_1723,N_18420,N_18035);
and UO_1724 (O_1724,N_19353,N_19407);
and UO_1725 (O_1725,N_19617,N_19546);
and UO_1726 (O_1726,N_18945,N_19040);
xnor UO_1727 (O_1727,N_19716,N_19656);
nor UO_1728 (O_1728,N_19925,N_18126);
nor UO_1729 (O_1729,N_18977,N_18141);
or UO_1730 (O_1730,N_19084,N_18069);
or UO_1731 (O_1731,N_19810,N_19602);
nand UO_1732 (O_1732,N_18512,N_19990);
nor UO_1733 (O_1733,N_19626,N_18492);
and UO_1734 (O_1734,N_19221,N_19240);
and UO_1735 (O_1735,N_18813,N_19740);
or UO_1736 (O_1736,N_18739,N_18783);
or UO_1737 (O_1737,N_18578,N_18265);
nand UO_1738 (O_1738,N_19692,N_19770);
nand UO_1739 (O_1739,N_18242,N_18804);
or UO_1740 (O_1740,N_19704,N_18047);
and UO_1741 (O_1741,N_19139,N_18027);
nor UO_1742 (O_1742,N_18504,N_18138);
nor UO_1743 (O_1743,N_19611,N_19618);
nor UO_1744 (O_1744,N_19047,N_18938);
or UO_1745 (O_1745,N_18672,N_18425);
nor UO_1746 (O_1746,N_18186,N_19481);
and UO_1747 (O_1747,N_18996,N_18159);
nor UO_1748 (O_1748,N_18108,N_18078);
nor UO_1749 (O_1749,N_19017,N_18368);
nor UO_1750 (O_1750,N_19344,N_18124);
and UO_1751 (O_1751,N_18342,N_18299);
xor UO_1752 (O_1752,N_18521,N_19388);
and UO_1753 (O_1753,N_19931,N_19476);
nor UO_1754 (O_1754,N_19485,N_18478);
xnor UO_1755 (O_1755,N_19191,N_18846);
or UO_1756 (O_1756,N_18427,N_19929);
xor UO_1757 (O_1757,N_19415,N_19047);
or UO_1758 (O_1758,N_18279,N_19959);
or UO_1759 (O_1759,N_19373,N_18181);
nand UO_1760 (O_1760,N_19215,N_18870);
nor UO_1761 (O_1761,N_18580,N_18005);
nand UO_1762 (O_1762,N_18800,N_18723);
nor UO_1763 (O_1763,N_18716,N_19736);
nor UO_1764 (O_1764,N_19537,N_18383);
nor UO_1765 (O_1765,N_18152,N_19096);
and UO_1766 (O_1766,N_19049,N_18449);
or UO_1767 (O_1767,N_19876,N_18349);
or UO_1768 (O_1768,N_18861,N_19659);
nand UO_1769 (O_1769,N_19235,N_18517);
nor UO_1770 (O_1770,N_18916,N_19076);
nand UO_1771 (O_1771,N_18964,N_19484);
nand UO_1772 (O_1772,N_18603,N_18379);
nor UO_1773 (O_1773,N_18121,N_18995);
nor UO_1774 (O_1774,N_18912,N_18880);
nand UO_1775 (O_1775,N_19671,N_18400);
and UO_1776 (O_1776,N_19825,N_19856);
or UO_1777 (O_1777,N_18390,N_18344);
or UO_1778 (O_1778,N_19472,N_19346);
or UO_1779 (O_1779,N_19388,N_19614);
and UO_1780 (O_1780,N_19175,N_18932);
nand UO_1781 (O_1781,N_18693,N_18035);
nor UO_1782 (O_1782,N_18474,N_18241);
and UO_1783 (O_1783,N_18650,N_18972);
or UO_1784 (O_1784,N_19404,N_18997);
xor UO_1785 (O_1785,N_18096,N_19537);
nor UO_1786 (O_1786,N_19595,N_18880);
nor UO_1787 (O_1787,N_18145,N_18769);
and UO_1788 (O_1788,N_18069,N_19463);
nand UO_1789 (O_1789,N_18352,N_18894);
or UO_1790 (O_1790,N_19450,N_18061);
xnor UO_1791 (O_1791,N_18009,N_18149);
and UO_1792 (O_1792,N_18870,N_18177);
and UO_1793 (O_1793,N_18939,N_19152);
nor UO_1794 (O_1794,N_18989,N_18041);
nand UO_1795 (O_1795,N_18999,N_19101);
nand UO_1796 (O_1796,N_19542,N_18543);
and UO_1797 (O_1797,N_19700,N_19623);
nand UO_1798 (O_1798,N_19300,N_19433);
and UO_1799 (O_1799,N_18432,N_18307);
and UO_1800 (O_1800,N_18924,N_18073);
nor UO_1801 (O_1801,N_19023,N_19065);
or UO_1802 (O_1802,N_18286,N_19530);
nand UO_1803 (O_1803,N_18785,N_18919);
nor UO_1804 (O_1804,N_18029,N_19002);
and UO_1805 (O_1805,N_19508,N_18607);
nor UO_1806 (O_1806,N_19156,N_18046);
nand UO_1807 (O_1807,N_18718,N_18922);
and UO_1808 (O_1808,N_19333,N_19830);
nor UO_1809 (O_1809,N_19359,N_18695);
and UO_1810 (O_1810,N_19816,N_19171);
or UO_1811 (O_1811,N_19559,N_19052);
xnor UO_1812 (O_1812,N_19799,N_18836);
nor UO_1813 (O_1813,N_19216,N_19547);
and UO_1814 (O_1814,N_19791,N_18442);
and UO_1815 (O_1815,N_19268,N_18498);
nand UO_1816 (O_1816,N_18608,N_18896);
nand UO_1817 (O_1817,N_18788,N_18726);
nand UO_1818 (O_1818,N_19632,N_19852);
or UO_1819 (O_1819,N_19433,N_18690);
nor UO_1820 (O_1820,N_19873,N_19399);
and UO_1821 (O_1821,N_18971,N_19019);
nand UO_1822 (O_1822,N_18269,N_19107);
and UO_1823 (O_1823,N_18063,N_19119);
nand UO_1824 (O_1824,N_19054,N_18739);
and UO_1825 (O_1825,N_19969,N_19222);
nand UO_1826 (O_1826,N_19459,N_19302);
and UO_1827 (O_1827,N_18193,N_18043);
and UO_1828 (O_1828,N_19658,N_18042);
and UO_1829 (O_1829,N_18924,N_19249);
nand UO_1830 (O_1830,N_19336,N_18116);
nor UO_1831 (O_1831,N_19212,N_19134);
and UO_1832 (O_1832,N_18155,N_18273);
and UO_1833 (O_1833,N_19972,N_18614);
nand UO_1834 (O_1834,N_19719,N_18804);
nand UO_1835 (O_1835,N_19653,N_19466);
and UO_1836 (O_1836,N_19062,N_18203);
or UO_1837 (O_1837,N_18239,N_19347);
nand UO_1838 (O_1838,N_19500,N_18242);
nand UO_1839 (O_1839,N_19727,N_19157);
nand UO_1840 (O_1840,N_19297,N_19651);
nor UO_1841 (O_1841,N_19365,N_19449);
nand UO_1842 (O_1842,N_19135,N_18863);
or UO_1843 (O_1843,N_19359,N_19919);
or UO_1844 (O_1844,N_19517,N_18135);
and UO_1845 (O_1845,N_18843,N_19848);
nor UO_1846 (O_1846,N_18451,N_19985);
and UO_1847 (O_1847,N_18951,N_18738);
and UO_1848 (O_1848,N_19167,N_19110);
nand UO_1849 (O_1849,N_18435,N_18280);
or UO_1850 (O_1850,N_18077,N_18529);
and UO_1851 (O_1851,N_19306,N_19186);
or UO_1852 (O_1852,N_18729,N_18906);
and UO_1853 (O_1853,N_18115,N_19957);
xor UO_1854 (O_1854,N_18058,N_19681);
and UO_1855 (O_1855,N_19037,N_18144);
or UO_1856 (O_1856,N_19854,N_18875);
and UO_1857 (O_1857,N_19805,N_18538);
nand UO_1858 (O_1858,N_19841,N_18196);
xor UO_1859 (O_1859,N_19274,N_18523);
nor UO_1860 (O_1860,N_19172,N_19882);
and UO_1861 (O_1861,N_18046,N_18186);
or UO_1862 (O_1862,N_18321,N_18519);
and UO_1863 (O_1863,N_19219,N_19533);
or UO_1864 (O_1864,N_18830,N_18146);
or UO_1865 (O_1865,N_18760,N_18435);
nand UO_1866 (O_1866,N_19324,N_18360);
or UO_1867 (O_1867,N_19381,N_19635);
or UO_1868 (O_1868,N_18336,N_19010);
nand UO_1869 (O_1869,N_18602,N_18473);
nor UO_1870 (O_1870,N_19768,N_18704);
nand UO_1871 (O_1871,N_18650,N_19622);
nor UO_1872 (O_1872,N_18675,N_18691);
and UO_1873 (O_1873,N_19254,N_18364);
nor UO_1874 (O_1874,N_19110,N_19613);
and UO_1875 (O_1875,N_19960,N_18223);
or UO_1876 (O_1876,N_19697,N_19200);
or UO_1877 (O_1877,N_18005,N_19786);
or UO_1878 (O_1878,N_18325,N_18203);
and UO_1879 (O_1879,N_18720,N_19306);
or UO_1880 (O_1880,N_19136,N_19215);
and UO_1881 (O_1881,N_19925,N_18470);
nand UO_1882 (O_1882,N_19679,N_18173);
xor UO_1883 (O_1883,N_18758,N_18502);
xnor UO_1884 (O_1884,N_19095,N_18047);
nand UO_1885 (O_1885,N_19830,N_19858);
nand UO_1886 (O_1886,N_18291,N_19895);
and UO_1887 (O_1887,N_18619,N_18709);
nand UO_1888 (O_1888,N_19208,N_18927);
nor UO_1889 (O_1889,N_18264,N_19060);
and UO_1890 (O_1890,N_19131,N_18161);
nand UO_1891 (O_1891,N_18483,N_19368);
and UO_1892 (O_1892,N_19005,N_19523);
and UO_1893 (O_1893,N_19519,N_19629);
or UO_1894 (O_1894,N_19904,N_19082);
nand UO_1895 (O_1895,N_19128,N_18529);
and UO_1896 (O_1896,N_19791,N_18600);
and UO_1897 (O_1897,N_18043,N_19008);
nand UO_1898 (O_1898,N_18224,N_19544);
and UO_1899 (O_1899,N_18712,N_19587);
and UO_1900 (O_1900,N_18190,N_18615);
nor UO_1901 (O_1901,N_19744,N_19700);
xnor UO_1902 (O_1902,N_19339,N_19124);
nor UO_1903 (O_1903,N_19275,N_19460);
nand UO_1904 (O_1904,N_18371,N_18494);
or UO_1905 (O_1905,N_18122,N_18534);
nor UO_1906 (O_1906,N_19514,N_19414);
nand UO_1907 (O_1907,N_18826,N_18314);
nor UO_1908 (O_1908,N_18217,N_19929);
and UO_1909 (O_1909,N_18878,N_19944);
and UO_1910 (O_1910,N_18864,N_18339);
and UO_1911 (O_1911,N_19350,N_18337);
and UO_1912 (O_1912,N_19766,N_19702);
or UO_1913 (O_1913,N_19071,N_18460);
or UO_1914 (O_1914,N_18210,N_18651);
or UO_1915 (O_1915,N_18954,N_18001);
or UO_1916 (O_1916,N_19015,N_19120);
nand UO_1917 (O_1917,N_18947,N_19271);
nor UO_1918 (O_1918,N_19032,N_18776);
or UO_1919 (O_1919,N_19649,N_18400);
nor UO_1920 (O_1920,N_18068,N_19145);
nor UO_1921 (O_1921,N_18500,N_19621);
nand UO_1922 (O_1922,N_19867,N_18089);
xnor UO_1923 (O_1923,N_18272,N_18543);
or UO_1924 (O_1924,N_18111,N_18708);
and UO_1925 (O_1925,N_19186,N_19179);
or UO_1926 (O_1926,N_18109,N_18558);
xor UO_1927 (O_1927,N_18978,N_19153);
xnor UO_1928 (O_1928,N_18003,N_19445);
and UO_1929 (O_1929,N_18571,N_19204);
and UO_1930 (O_1930,N_19179,N_18917);
nor UO_1931 (O_1931,N_19218,N_19058);
nand UO_1932 (O_1932,N_19347,N_18754);
and UO_1933 (O_1933,N_18195,N_19827);
nand UO_1934 (O_1934,N_19465,N_19128);
or UO_1935 (O_1935,N_19174,N_19226);
or UO_1936 (O_1936,N_18074,N_18500);
nor UO_1937 (O_1937,N_19341,N_18380);
nor UO_1938 (O_1938,N_18072,N_19247);
and UO_1939 (O_1939,N_18753,N_18763);
nand UO_1940 (O_1940,N_19908,N_18724);
and UO_1941 (O_1941,N_18580,N_19868);
and UO_1942 (O_1942,N_18866,N_19398);
nor UO_1943 (O_1943,N_18555,N_18435);
or UO_1944 (O_1944,N_19538,N_19262);
nor UO_1945 (O_1945,N_19026,N_18543);
nor UO_1946 (O_1946,N_18469,N_19354);
and UO_1947 (O_1947,N_18926,N_19876);
xor UO_1948 (O_1948,N_18449,N_18376);
and UO_1949 (O_1949,N_19641,N_18888);
or UO_1950 (O_1950,N_18398,N_19132);
nor UO_1951 (O_1951,N_19722,N_18032);
nand UO_1952 (O_1952,N_19743,N_18592);
and UO_1953 (O_1953,N_18175,N_18049);
xor UO_1954 (O_1954,N_18019,N_19356);
nor UO_1955 (O_1955,N_18833,N_18587);
and UO_1956 (O_1956,N_19694,N_18251);
or UO_1957 (O_1957,N_19132,N_19633);
xor UO_1958 (O_1958,N_18784,N_19308);
nand UO_1959 (O_1959,N_19396,N_19491);
xnor UO_1960 (O_1960,N_19744,N_18148);
and UO_1961 (O_1961,N_19341,N_19269);
and UO_1962 (O_1962,N_19566,N_18378);
nand UO_1963 (O_1963,N_18312,N_19094);
nand UO_1964 (O_1964,N_18419,N_18484);
and UO_1965 (O_1965,N_18608,N_18889);
or UO_1966 (O_1966,N_19185,N_18633);
and UO_1967 (O_1967,N_18856,N_18231);
or UO_1968 (O_1968,N_19763,N_19786);
or UO_1969 (O_1969,N_19531,N_18435);
nor UO_1970 (O_1970,N_18304,N_18100);
nand UO_1971 (O_1971,N_18696,N_18007);
and UO_1972 (O_1972,N_19112,N_19196);
and UO_1973 (O_1973,N_19822,N_18193);
and UO_1974 (O_1974,N_19789,N_18914);
nand UO_1975 (O_1975,N_19929,N_19007);
xnor UO_1976 (O_1976,N_18772,N_19613);
nor UO_1977 (O_1977,N_18704,N_18977);
and UO_1978 (O_1978,N_18865,N_18426);
nand UO_1979 (O_1979,N_18827,N_18221);
or UO_1980 (O_1980,N_18658,N_19530);
or UO_1981 (O_1981,N_18747,N_18666);
and UO_1982 (O_1982,N_19260,N_19888);
nand UO_1983 (O_1983,N_19140,N_18984);
nand UO_1984 (O_1984,N_18050,N_18636);
nor UO_1985 (O_1985,N_18019,N_19869);
or UO_1986 (O_1986,N_18859,N_18891);
nor UO_1987 (O_1987,N_19109,N_18479);
nor UO_1988 (O_1988,N_19856,N_19983);
or UO_1989 (O_1989,N_18992,N_18563);
and UO_1990 (O_1990,N_19052,N_19945);
nand UO_1991 (O_1991,N_19511,N_19119);
nor UO_1992 (O_1992,N_18698,N_19332);
and UO_1993 (O_1993,N_19167,N_18338);
nor UO_1994 (O_1994,N_19181,N_18708);
and UO_1995 (O_1995,N_18048,N_19166);
nand UO_1996 (O_1996,N_19496,N_18532);
nor UO_1997 (O_1997,N_18708,N_19814);
and UO_1998 (O_1998,N_19919,N_18989);
nand UO_1999 (O_1999,N_19810,N_18544);
xnor UO_2000 (O_2000,N_19393,N_19542);
nor UO_2001 (O_2001,N_18371,N_19126);
nor UO_2002 (O_2002,N_19856,N_19287);
xor UO_2003 (O_2003,N_18128,N_18381);
nor UO_2004 (O_2004,N_18273,N_18812);
nand UO_2005 (O_2005,N_18565,N_19565);
nand UO_2006 (O_2006,N_18715,N_19242);
nor UO_2007 (O_2007,N_18792,N_18455);
and UO_2008 (O_2008,N_18566,N_19590);
nor UO_2009 (O_2009,N_18003,N_19919);
and UO_2010 (O_2010,N_19514,N_18051);
nand UO_2011 (O_2011,N_18106,N_19594);
nor UO_2012 (O_2012,N_19016,N_18402);
or UO_2013 (O_2013,N_18391,N_19414);
nand UO_2014 (O_2014,N_19683,N_18994);
or UO_2015 (O_2015,N_18724,N_18864);
xor UO_2016 (O_2016,N_19071,N_19953);
nand UO_2017 (O_2017,N_18860,N_19154);
nand UO_2018 (O_2018,N_19164,N_18227);
and UO_2019 (O_2019,N_19190,N_19744);
nand UO_2020 (O_2020,N_18827,N_18047);
nor UO_2021 (O_2021,N_19023,N_19630);
xor UO_2022 (O_2022,N_18721,N_19870);
nor UO_2023 (O_2023,N_19922,N_18768);
and UO_2024 (O_2024,N_19162,N_19903);
nor UO_2025 (O_2025,N_19419,N_19404);
and UO_2026 (O_2026,N_19891,N_19736);
nand UO_2027 (O_2027,N_18903,N_19828);
nor UO_2028 (O_2028,N_18047,N_18449);
nor UO_2029 (O_2029,N_18932,N_18609);
or UO_2030 (O_2030,N_19271,N_18414);
nor UO_2031 (O_2031,N_19702,N_19473);
or UO_2032 (O_2032,N_18444,N_18198);
nand UO_2033 (O_2033,N_19390,N_18089);
nor UO_2034 (O_2034,N_19231,N_18857);
and UO_2035 (O_2035,N_18235,N_19363);
nand UO_2036 (O_2036,N_19217,N_18641);
or UO_2037 (O_2037,N_18082,N_19859);
nor UO_2038 (O_2038,N_18343,N_19130);
or UO_2039 (O_2039,N_19385,N_18130);
nor UO_2040 (O_2040,N_19914,N_19806);
nand UO_2041 (O_2041,N_18521,N_19876);
and UO_2042 (O_2042,N_19182,N_19122);
or UO_2043 (O_2043,N_19088,N_19265);
or UO_2044 (O_2044,N_18368,N_18892);
nand UO_2045 (O_2045,N_19268,N_19183);
or UO_2046 (O_2046,N_19523,N_19554);
nand UO_2047 (O_2047,N_18696,N_19797);
or UO_2048 (O_2048,N_18877,N_19886);
xor UO_2049 (O_2049,N_18260,N_18718);
xnor UO_2050 (O_2050,N_19315,N_19286);
nand UO_2051 (O_2051,N_18771,N_18147);
nor UO_2052 (O_2052,N_19625,N_18399);
nand UO_2053 (O_2053,N_18358,N_18863);
nand UO_2054 (O_2054,N_19814,N_18037);
and UO_2055 (O_2055,N_18392,N_19843);
and UO_2056 (O_2056,N_18560,N_18654);
or UO_2057 (O_2057,N_19965,N_18937);
or UO_2058 (O_2058,N_19185,N_19746);
and UO_2059 (O_2059,N_18729,N_18014);
and UO_2060 (O_2060,N_18229,N_19849);
nor UO_2061 (O_2061,N_18060,N_18555);
nor UO_2062 (O_2062,N_19654,N_18878);
nand UO_2063 (O_2063,N_18026,N_19392);
and UO_2064 (O_2064,N_19681,N_18603);
and UO_2065 (O_2065,N_18365,N_18445);
nand UO_2066 (O_2066,N_19681,N_18962);
or UO_2067 (O_2067,N_18923,N_19607);
xnor UO_2068 (O_2068,N_19712,N_18537);
nor UO_2069 (O_2069,N_18631,N_18489);
or UO_2070 (O_2070,N_19854,N_18551);
nand UO_2071 (O_2071,N_18625,N_18160);
and UO_2072 (O_2072,N_19161,N_18171);
and UO_2073 (O_2073,N_18806,N_18935);
nand UO_2074 (O_2074,N_18745,N_19180);
nand UO_2075 (O_2075,N_19199,N_18866);
nand UO_2076 (O_2076,N_19589,N_18911);
xor UO_2077 (O_2077,N_19826,N_19169);
or UO_2078 (O_2078,N_18863,N_19778);
nand UO_2079 (O_2079,N_19021,N_19004);
nor UO_2080 (O_2080,N_19737,N_19954);
nor UO_2081 (O_2081,N_19250,N_19991);
nor UO_2082 (O_2082,N_19714,N_18796);
nor UO_2083 (O_2083,N_18814,N_18119);
and UO_2084 (O_2084,N_19080,N_18913);
nor UO_2085 (O_2085,N_18427,N_19448);
or UO_2086 (O_2086,N_19920,N_19205);
nor UO_2087 (O_2087,N_18524,N_19248);
and UO_2088 (O_2088,N_18163,N_18836);
nand UO_2089 (O_2089,N_19970,N_19080);
or UO_2090 (O_2090,N_18019,N_18283);
xor UO_2091 (O_2091,N_18369,N_19391);
or UO_2092 (O_2092,N_18905,N_19217);
nor UO_2093 (O_2093,N_18296,N_19554);
nand UO_2094 (O_2094,N_19154,N_19209);
nand UO_2095 (O_2095,N_18900,N_19576);
nand UO_2096 (O_2096,N_18440,N_19165);
xor UO_2097 (O_2097,N_19871,N_19433);
or UO_2098 (O_2098,N_19214,N_18111);
nand UO_2099 (O_2099,N_19272,N_19644);
nand UO_2100 (O_2100,N_18872,N_19711);
and UO_2101 (O_2101,N_19417,N_19111);
nand UO_2102 (O_2102,N_18128,N_19456);
nor UO_2103 (O_2103,N_18503,N_18260);
nand UO_2104 (O_2104,N_18253,N_19287);
and UO_2105 (O_2105,N_19069,N_19202);
nor UO_2106 (O_2106,N_19986,N_18063);
and UO_2107 (O_2107,N_19249,N_19326);
nor UO_2108 (O_2108,N_19476,N_19047);
or UO_2109 (O_2109,N_18165,N_18747);
nor UO_2110 (O_2110,N_19044,N_19022);
xnor UO_2111 (O_2111,N_18012,N_18997);
or UO_2112 (O_2112,N_18071,N_18121);
nand UO_2113 (O_2113,N_18999,N_19961);
nor UO_2114 (O_2114,N_19549,N_18673);
or UO_2115 (O_2115,N_19096,N_18273);
and UO_2116 (O_2116,N_19410,N_18967);
nor UO_2117 (O_2117,N_19406,N_19387);
xor UO_2118 (O_2118,N_19486,N_19386);
nor UO_2119 (O_2119,N_18028,N_19997);
nand UO_2120 (O_2120,N_19669,N_18331);
nor UO_2121 (O_2121,N_19292,N_18637);
and UO_2122 (O_2122,N_18348,N_18505);
nor UO_2123 (O_2123,N_19186,N_19849);
nor UO_2124 (O_2124,N_19511,N_19933);
or UO_2125 (O_2125,N_19259,N_18733);
nand UO_2126 (O_2126,N_19196,N_19586);
and UO_2127 (O_2127,N_19763,N_19526);
and UO_2128 (O_2128,N_19573,N_19271);
nor UO_2129 (O_2129,N_18223,N_18027);
and UO_2130 (O_2130,N_19613,N_19875);
nand UO_2131 (O_2131,N_18272,N_19129);
nor UO_2132 (O_2132,N_18369,N_18933);
nor UO_2133 (O_2133,N_19605,N_18132);
and UO_2134 (O_2134,N_19866,N_19242);
nor UO_2135 (O_2135,N_18815,N_18616);
nand UO_2136 (O_2136,N_18319,N_18125);
nand UO_2137 (O_2137,N_19143,N_19930);
or UO_2138 (O_2138,N_18249,N_19834);
nand UO_2139 (O_2139,N_18293,N_18164);
or UO_2140 (O_2140,N_18504,N_18155);
and UO_2141 (O_2141,N_18987,N_18683);
nand UO_2142 (O_2142,N_18326,N_18592);
nand UO_2143 (O_2143,N_18703,N_19211);
nand UO_2144 (O_2144,N_19923,N_18353);
xor UO_2145 (O_2145,N_19584,N_18958);
or UO_2146 (O_2146,N_18195,N_19476);
and UO_2147 (O_2147,N_19241,N_18737);
and UO_2148 (O_2148,N_18620,N_18300);
or UO_2149 (O_2149,N_18842,N_19590);
nor UO_2150 (O_2150,N_19814,N_19594);
xnor UO_2151 (O_2151,N_19607,N_18067);
nor UO_2152 (O_2152,N_18262,N_19967);
nand UO_2153 (O_2153,N_18462,N_19360);
nor UO_2154 (O_2154,N_18393,N_19917);
and UO_2155 (O_2155,N_18889,N_18657);
or UO_2156 (O_2156,N_19320,N_18068);
nand UO_2157 (O_2157,N_19818,N_18168);
or UO_2158 (O_2158,N_19000,N_18265);
and UO_2159 (O_2159,N_19154,N_19134);
and UO_2160 (O_2160,N_18856,N_19699);
nor UO_2161 (O_2161,N_19649,N_18685);
and UO_2162 (O_2162,N_19168,N_18149);
or UO_2163 (O_2163,N_19971,N_18743);
nand UO_2164 (O_2164,N_18134,N_19861);
nor UO_2165 (O_2165,N_18117,N_19251);
nand UO_2166 (O_2166,N_19731,N_18856);
or UO_2167 (O_2167,N_19855,N_18140);
xnor UO_2168 (O_2168,N_18251,N_18280);
nand UO_2169 (O_2169,N_18023,N_18869);
nand UO_2170 (O_2170,N_18212,N_18978);
nand UO_2171 (O_2171,N_18368,N_19121);
nor UO_2172 (O_2172,N_18038,N_18943);
or UO_2173 (O_2173,N_18678,N_18622);
nand UO_2174 (O_2174,N_19716,N_19874);
nor UO_2175 (O_2175,N_19131,N_18081);
nor UO_2176 (O_2176,N_18265,N_18877);
or UO_2177 (O_2177,N_18812,N_18552);
xnor UO_2178 (O_2178,N_19553,N_19187);
or UO_2179 (O_2179,N_18501,N_18215);
nand UO_2180 (O_2180,N_19096,N_18093);
nand UO_2181 (O_2181,N_19728,N_19887);
nand UO_2182 (O_2182,N_19044,N_19131);
nor UO_2183 (O_2183,N_19063,N_19792);
nand UO_2184 (O_2184,N_19174,N_19130);
or UO_2185 (O_2185,N_19815,N_18693);
and UO_2186 (O_2186,N_19733,N_18823);
nand UO_2187 (O_2187,N_18582,N_19544);
nand UO_2188 (O_2188,N_19781,N_18266);
nand UO_2189 (O_2189,N_18580,N_19324);
and UO_2190 (O_2190,N_19527,N_18387);
nor UO_2191 (O_2191,N_19400,N_19234);
and UO_2192 (O_2192,N_18995,N_19090);
nand UO_2193 (O_2193,N_19787,N_19949);
nand UO_2194 (O_2194,N_19715,N_18302);
nand UO_2195 (O_2195,N_18879,N_18607);
nor UO_2196 (O_2196,N_18585,N_19666);
and UO_2197 (O_2197,N_19020,N_18641);
or UO_2198 (O_2198,N_19428,N_19866);
nor UO_2199 (O_2199,N_19294,N_19603);
and UO_2200 (O_2200,N_18128,N_19789);
and UO_2201 (O_2201,N_18574,N_19420);
xnor UO_2202 (O_2202,N_18070,N_18658);
nand UO_2203 (O_2203,N_19006,N_19858);
nor UO_2204 (O_2204,N_19770,N_19842);
xor UO_2205 (O_2205,N_19167,N_18729);
nand UO_2206 (O_2206,N_18637,N_18823);
xnor UO_2207 (O_2207,N_18141,N_18829);
and UO_2208 (O_2208,N_19268,N_19852);
nand UO_2209 (O_2209,N_18708,N_19765);
or UO_2210 (O_2210,N_19731,N_19077);
and UO_2211 (O_2211,N_19867,N_19828);
nand UO_2212 (O_2212,N_18999,N_18901);
and UO_2213 (O_2213,N_19711,N_19902);
nand UO_2214 (O_2214,N_19005,N_18350);
nor UO_2215 (O_2215,N_18488,N_19679);
or UO_2216 (O_2216,N_18292,N_19877);
or UO_2217 (O_2217,N_18166,N_19855);
and UO_2218 (O_2218,N_19319,N_19390);
nor UO_2219 (O_2219,N_18659,N_19717);
or UO_2220 (O_2220,N_18924,N_19979);
nand UO_2221 (O_2221,N_18314,N_18747);
nor UO_2222 (O_2222,N_18181,N_19858);
nand UO_2223 (O_2223,N_19107,N_18818);
nand UO_2224 (O_2224,N_19822,N_18042);
or UO_2225 (O_2225,N_19918,N_19964);
or UO_2226 (O_2226,N_19523,N_18777);
nand UO_2227 (O_2227,N_19112,N_18525);
nand UO_2228 (O_2228,N_19202,N_18370);
nand UO_2229 (O_2229,N_18012,N_19821);
and UO_2230 (O_2230,N_18012,N_18525);
nand UO_2231 (O_2231,N_18756,N_18093);
nor UO_2232 (O_2232,N_19666,N_18531);
nand UO_2233 (O_2233,N_19977,N_19283);
xor UO_2234 (O_2234,N_18974,N_19327);
xnor UO_2235 (O_2235,N_18228,N_18366);
and UO_2236 (O_2236,N_18402,N_18667);
and UO_2237 (O_2237,N_19997,N_19576);
nor UO_2238 (O_2238,N_18515,N_18186);
nand UO_2239 (O_2239,N_18012,N_19640);
and UO_2240 (O_2240,N_18802,N_18667);
nand UO_2241 (O_2241,N_18098,N_18469);
nand UO_2242 (O_2242,N_19353,N_18086);
nor UO_2243 (O_2243,N_19182,N_19100);
nor UO_2244 (O_2244,N_19393,N_18314);
and UO_2245 (O_2245,N_18429,N_19069);
nor UO_2246 (O_2246,N_19802,N_18123);
nand UO_2247 (O_2247,N_18439,N_19563);
nor UO_2248 (O_2248,N_19521,N_19260);
or UO_2249 (O_2249,N_18315,N_18355);
or UO_2250 (O_2250,N_19092,N_18625);
nand UO_2251 (O_2251,N_18666,N_19112);
nor UO_2252 (O_2252,N_19525,N_18418);
xor UO_2253 (O_2253,N_19197,N_18334);
nand UO_2254 (O_2254,N_19875,N_19874);
and UO_2255 (O_2255,N_18133,N_19227);
nand UO_2256 (O_2256,N_19315,N_19481);
nand UO_2257 (O_2257,N_19128,N_19029);
and UO_2258 (O_2258,N_19621,N_19353);
or UO_2259 (O_2259,N_18682,N_18880);
and UO_2260 (O_2260,N_19840,N_18928);
nor UO_2261 (O_2261,N_18910,N_18351);
nor UO_2262 (O_2262,N_19513,N_19789);
nor UO_2263 (O_2263,N_19758,N_19333);
and UO_2264 (O_2264,N_19802,N_19384);
nand UO_2265 (O_2265,N_18107,N_19581);
xnor UO_2266 (O_2266,N_18466,N_18111);
and UO_2267 (O_2267,N_19459,N_19974);
xnor UO_2268 (O_2268,N_19226,N_19611);
or UO_2269 (O_2269,N_19230,N_18192);
xnor UO_2270 (O_2270,N_18126,N_19855);
nand UO_2271 (O_2271,N_18653,N_18761);
and UO_2272 (O_2272,N_19631,N_19482);
or UO_2273 (O_2273,N_18746,N_19019);
nand UO_2274 (O_2274,N_19183,N_19228);
nor UO_2275 (O_2275,N_18475,N_18049);
xor UO_2276 (O_2276,N_19958,N_19235);
nand UO_2277 (O_2277,N_19399,N_18230);
or UO_2278 (O_2278,N_19221,N_19256);
xnor UO_2279 (O_2279,N_19180,N_19176);
nand UO_2280 (O_2280,N_19547,N_19009);
nand UO_2281 (O_2281,N_19112,N_19965);
nor UO_2282 (O_2282,N_18939,N_18308);
xor UO_2283 (O_2283,N_19731,N_19575);
xor UO_2284 (O_2284,N_19126,N_19868);
nand UO_2285 (O_2285,N_19702,N_19191);
nand UO_2286 (O_2286,N_18471,N_18156);
and UO_2287 (O_2287,N_19761,N_19386);
or UO_2288 (O_2288,N_19750,N_19636);
nor UO_2289 (O_2289,N_19796,N_19651);
or UO_2290 (O_2290,N_19361,N_19191);
nand UO_2291 (O_2291,N_18555,N_18521);
nor UO_2292 (O_2292,N_19516,N_19676);
xnor UO_2293 (O_2293,N_18526,N_18410);
nand UO_2294 (O_2294,N_19752,N_18786);
and UO_2295 (O_2295,N_18025,N_18152);
nor UO_2296 (O_2296,N_19515,N_18457);
or UO_2297 (O_2297,N_18860,N_18261);
nor UO_2298 (O_2298,N_18430,N_19067);
or UO_2299 (O_2299,N_19935,N_19032);
or UO_2300 (O_2300,N_18858,N_18886);
or UO_2301 (O_2301,N_19949,N_18190);
nand UO_2302 (O_2302,N_18464,N_19324);
or UO_2303 (O_2303,N_19028,N_18546);
and UO_2304 (O_2304,N_18251,N_18291);
and UO_2305 (O_2305,N_18568,N_18364);
nor UO_2306 (O_2306,N_18522,N_18023);
nor UO_2307 (O_2307,N_18946,N_19985);
nor UO_2308 (O_2308,N_18592,N_19004);
or UO_2309 (O_2309,N_19022,N_18935);
nor UO_2310 (O_2310,N_19251,N_19142);
or UO_2311 (O_2311,N_18880,N_19592);
or UO_2312 (O_2312,N_19936,N_19643);
nor UO_2313 (O_2313,N_19892,N_19815);
xnor UO_2314 (O_2314,N_18554,N_18907);
xnor UO_2315 (O_2315,N_19538,N_18258);
nand UO_2316 (O_2316,N_19761,N_19656);
nor UO_2317 (O_2317,N_19154,N_19944);
nand UO_2318 (O_2318,N_19257,N_18591);
xnor UO_2319 (O_2319,N_19597,N_18104);
xnor UO_2320 (O_2320,N_18642,N_19142);
and UO_2321 (O_2321,N_18781,N_19188);
or UO_2322 (O_2322,N_18750,N_18883);
and UO_2323 (O_2323,N_18873,N_18591);
nor UO_2324 (O_2324,N_18738,N_18025);
or UO_2325 (O_2325,N_18924,N_18667);
nand UO_2326 (O_2326,N_19879,N_19403);
nor UO_2327 (O_2327,N_19037,N_18802);
and UO_2328 (O_2328,N_19053,N_19214);
xnor UO_2329 (O_2329,N_19782,N_19862);
and UO_2330 (O_2330,N_18996,N_18162);
and UO_2331 (O_2331,N_18384,N_19389);
or UO_2332 (O_2332,N_18292,N_18178);
nand UO_2333 (O_2333,N_19981,N_18315);
or UO_2334 (O_2334,N_18400,N_18416);
xnor UO_2335 (O_2335,N_19429,N_18730);
nor UO_2336 (O_2336,N_19828,N_19673);
and UO_2337 (O_2337,N_19053,N_19357);
and UO_2338 (O_2338,N_19551,N_18054);
or UO_2339 (O_2339,N_19649,N_18566);
xnor UO_2340 (O_2340,N_19170,N_18138);
and UO_2341 (O_2341,N_19803,N_18263);
nor UO_2342 (O_2342,N_19191,N_18407);
nor UO_2343 (O_2343,N_18663,N_19808);
nor UO_2344 (O_2344,N_19224,N_18710);
or UO_2345 (O_2345,N_18635,N_19930);
nand UO_2346 (O_2346,N_18839,N_18611);
nor UO_2347 (O_2347,N_18208,N_19767);
and UO_2348 (O_2348,N_19843,N_19306);
or UO_2349 (O_2349,N_18665,N_18871);
or UO_2350 (O_2350,N_18436,N_19284);
or UO_2351 (O_2351,N_18440,N_18897);
and UO_2352 (O_2352,N_19824,N_19254);
nand UO_2353 (O_2353,N_18814,N_19390);
and UO_2354 (O_2354,N_19583,N_19044);
nor UO_2355 (O_2355,N_19615,N_18646);
nor UO_2356 (O_2356,N_18390,N_19025);
nand UO_2357 (O_2357,N_19021,N_18477);
nand UO_2358 (O_2358,N_18885,N_18073);
xnor UO_2359 (O_2359,N_18320,N_19613);
or UO_2360 (O_2360,N_19223,N_19262);
and UO_2361 (O_2361,N_19071,N_19243);
and UO_2362 (O_2362,N_18848,N_19800);
nand UO_2363 (O_2363,N_19598,N_18058);
nand UO_2364 (O_2364,N_18262,N_18197);
and UO_2365 (O_2365,N_18306,N_19678);
or UO_2366 (O_2366,N_19651,N_19427);
or UO_2367 (O_2367,N_18024,N_18962);
nand UO_2368 (O_2368,N_18242,N_18849);
or UO_2369 (O_2369,N_18947,N_18034);
nand UO_2370 (O_2370,N_19800,N_19773);
nor UO_2371 (O_2371,N_19322,N_18692);
xor UO_2372 (O_2372,N_18502,N_18954);
nand UO_2373 (O_2373,N_18636,N_19663);
or UO_2374 (O_2374,N_18085,N_18322);
nor UO_2375 (O_2375,N_19238,N_19261);
nor UO_2376 (O_2376,N_18790,N_18978);
nor UO_2377 (O_2377,N_19343,N_18692);
nand UO_2378 (O_2378,N_19685,N_18256);
and UO_2379 (O_2379,N_19650,N_18469);
or UO_2380 (O_2380,N_18254,N_18489);
nand UO_2381 (O_2381,N_18777,N_19558);
xnor UO_2382 (O_2382,N_19276,N_18949);
nor UO_2383 (O_2383,N_18205,N_18241);
or UO_2384 (O_2384,N_19060,N_19056);
nor UO_2385 (O_2385,N_18215,N_18711);
and UO_2386 (O_2386,N_19770,N_19456);
nand UO_2387 (O_2387,N_18573,N_18271);
and UO_2388 (O_2388,N_18676,N_19661);
or UO_2389 (O_2389,N_18642,N_18844);
and UO_2390 (O_2390,N_18225,N_18560);
xor UO_2391 (O_2391,N_19277,N_19840);
nand UO_2392 (O_2392,N_19102,N_18527);
nor UO_2393 (O_2393,N_19941,N_18298);
nand UO_2394 (O_2394,N_19280,N_18900);
nor UO_2395 (O_2395,N_19283,N_19397);
nand UO_2396 (O_2396,N_19714,N_19069);
nand UO_2397 (O_2397,N_19398,N_18948);
xnor UO_2398 (O_2398,N_19745,N_18344);
nand UO_2399 (O_2399,N_18894,N_19098);
nor UO_2400 (O_2400,N_18233,N_19051);
and UO_2401 (O_2401,N_18256,N_19705);
nand UO_2402 (O_2402,N_18398,N_18772);
and UO_2403 (O_2403,N_19935,N_19555);
nand UO_2404 (O_2404,N_18343,N_19703);
or UO_2405 (O_2405,N_19047,N_18177);
or UO_2406 (O_2406,N_18811,N_18365);
and UO_2407 (O_2407,N_18892,N_19876);
nand UO_2408 (O_2408,N_18090,N_18943);
nor UO_2409 (O_2409,N_19255,N_18961);
or UO_2410 (O_2410,N_19345,N_18049);
or UO_2411 (O_2411,N_18460,N_18201);
xnor UO_2412 (O_2412,N_19146,N_18952);
or UO_2413 (O_2413,N_18777,N_19208);
xnor UO_2414 (O_2414,N_19100,N_19532);
xnor UO_2415 (O_2415,N_18043,N_18102);
and UO_2416 (O_2416,N_18993,N_19060);
and UO_2417 (O_2417,N_19897,N_19687);
nor UO_2418 (O_2418,N_19036,N_19201);
and UO_2419 (O_2419,N_19638,N_18910);
or UO_2420 (O_2420,N_19233,N_19637);
nor UO_2421 (O_2421,N_19721,N_19179);
nand UO_2422 (O_2422,N_18723,N_19874);
xor UO_2423 (O_2423,N_19133,N_19990);
nand UO_2424 (O_2424,N_18003,N_18278);
or UO_2425 (O_2425,N_18381,N_19037);
or UO_2426 (O_2426,N_19368,N_19907);
and UO_2427 (O_2427,N_18346,N_18441);
or UO_2428 (O_2428,N_19498,N_18313);
or UO_2429 (O_2429,N_19700,N_18944);
nand UO_2430 (O_2430,N_18991,N_18542);
nand UO_2431 (O_2431,N_19409,N_19421);
or UO_2432 (O_2432,N_19445,N_18916);
nand UO_2433 (O_2433,N_18908,N_19031);
nor UO_2434 (O_2434,N_19359,N_19332);
and UO_2435 (O_2435,N_19813,N_19803);
and UO_2436 (O_2436,N_18071,N_19847);
or UO_2437 (O_2437,N_18026,N_18667);
nand UO_2438 (O_2438,N_18366,N_19649);
nand UO_2439 (O_2439,N_18379,N_18198);
and UO_2440 (O_2440,N_18812,N_19527);
and UO_2441 (O_2441,N_19312,N_19548);
nor UO_2442 (O_2442,N_19006,N_18939);
and UO_2443 (O_2443,N_18381,N_19774);
and UO_2444 (O_2444,N_18094,N_19644);
or UO_2445 (O_2445,N_18265,N_19348);
xor UO_2446 (O_2446,N_18971,N_19397);
and UO_2447 (O_2447,N_19753,N_19350);
nor UO_2448 (O_2448,N_18534,N_18294);
nor UO_2449 (O_2449,N_18594,N_18144);
nand UO_2450 (O_2450,N_19511,N_18756);
or UO_2451 (O_2451,N_18766,N_18391);
nor UO_2452 (O_2452,N_19868,N_18142);
and UO_2453 (O_2453,N_19345,N_19311);
nand UO_2454 (O_2454,N_18095,N_19201);
and UO_2455 (O_2455,N_18958,N_18331);
and UO_2456 (O_2456,N_19360,N_18235);
and UO_2457 (O_2457,N_19910,N_18996);
or UO_2458 (O_2458,N_19266,N_19109);
and UO_2459 (O_2459,N_18584,N_19248);
nand UO_2460 (O_2460,N_19365,N_19346);
and UO_2461 (O_2461,N_19319,N_18978);
or UO_2462 (O_2462,N_19023,N_18602);
nand UO_2463 (O_2463,N_19898,N_19911);
nor UO_2464 (O_2464,N_18848,N_19592);
or UO_2465 (O_2465,N_19101,N_18501);
and UO_2466 (O_2466,N_19385,N_18240);
or UO_2467 (O_2467,N_19882,N_18786);
nor UO_2468 (O_2468,N_19877,N_18241);
xnor UO_2469 (O_2469,N_19209,N_18510);
and UO_2470 (O_2470,N_18186,N_19280);
or UO_2471 (O_2471,N_19847,N_19137);
nor UO_2472 (O_2472,N_19004,N_19587);
or UO_2473 (O_2473,N_18801,N_18617);
and UO_2474 (O_2474,N_19652,N_19707);
xnor UO_2475 (O_2475,N_18165,N_19659);
or UO_2476 (O_2476,N_19850,N_19584);
or UO_2477 (O_2477,N_18136,N_19522);
nor UO_2478 (O_2478,N_19987,N_19698);
xor UO_2479 (O_2479,N_18254,N_19267);
and UO_2480 (O_2480,N_18874,N_19419);
nor UO_2481 (O_2481,N_19653,N_19159);
and UO_2482 (O_2482,N_19857,N_18883);
or UO_2483 (O_2483,N_18834,N_19332);
or UO_2484 (O_2484,N_18975,N_18295);
and UO_2485 (O_2485,N_18580,N_19216);
nand UO_2486 (O_2486,N_19689,N_18152);
nor UO_2487 (O_2487,N_19997,N_18244);
or UO_2488 (O_2488,N_19309,N_19638);
nor UO_2489 (O_2489,N_19259,N_19040);
nor UO_2490 (O_2490,N_18892,N_18250);
and UO_2491 (O_2491,N_18824,N_18914);
and UO_2492 (O_2492,N_19352,N_19416);
nand UO_2493 (O_2493,N_19098,N_19039);
xor UO_2494 (O_2494,N_18139,N_18141);
nor UO_2495 (O_2495,N_18295,N_18944);
nand UO_2496 (O_2496,N_18429,N_19731);
nand UO_2497 (O_2497,N_18556,N_18688);
or UO_2498 (O_2498,N_19021,N_19269);
and UO_2499 (O_2499,N_19811,N_19852);
endmodule