module basic_750_5000_1000_2_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2505,N_2507,N_2509,N_2510,N_2511,N_2512,N_2514,N_2515,N_2518,N_2519,N_2520,N_2521,N_2522,N_2524,N_2526,N_2529,N_2531,N_2532,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2550,N_2551,N_2552,N_2553,N_2554,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2573,N_2574,N_2577,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2635,N_2636,N_2639,N_2640,N_2641,N_2642,N_2644,N_2645,N_2646,N_2647,N_2648,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2678,N_2680,N_2681,N_2682,N_2683,N_2684,N_2686,N_2687,N_2688,N_2689,N_2691,N_2692,N_2693,N_2694,N_2695,N_2698,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2714,N_2715,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2741,N_2742,N_2743,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2767,N_2769,N_2770,N_2771,N_2772,N_2774,N_2776,N_2777,N_2778,N_2779,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2789,N_2790,N_2791,N_2792,N_2795,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2827,N_2829,N_2830,N_2833,N_2835,N_2836,N_2837,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2850,N_2851,N_2852,N_2853,N_2854,N_2856,N_2858,N_2859,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2881,N_2883,N_2884,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2897,N_2898,N_2899,N_2902,N_2903,N_2904,N_2905,N_2908,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2926,N_2927,N_2929,N_2931,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2963,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2972,N_2973,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2984,N_2985,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2997,N_2998,N_3000,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3013,N_3014,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3058,N_3060,N_3061,N_3062,N_3063,N_3064,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3075,N_3077,N_3078,N_3079,N_3081,N_3082,N_3083,N_3085,N_3087,N_3088,N_3089,N_3090,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3101,N_3102,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3112,N_3113,N_3114,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3140,N_3142,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3168,N_3170,N_3171,N_3174,N_3175,N_3176,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3209,N_3210,N_3211,N_3213,N_3214,N_3215,N_3216,N_3217,N_3220,N_3221,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3230,N_3233,N_3234,N_3236,N_3237,N_3238,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3250,N_3251,N_3254,N_3256,N_3258,N_3259,N_3260,N_3262,N_3263,N_3264,N_3265,N_3266,N_3268,N_3269,N_3270,N_3272,N_3273,N_3274,N_3275,N_3276,N_3278,N_3279,N_3280,N_3282,N_3283,N_3284,N_3285,N_3287,N_3288,N_3289,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3302,N_3304,N_3305,N_3306,N_3307,N_3308,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3327,N_3328,N_3329,N_3332,N_3333,N_3334,N_3335,N_3337,N_3338,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3356,N_3357,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3370,N_3372,N_3374,N_3375,N_3377,N_3378,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3407,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3438,N_3439,N_3441,N_3442,N_3443,N_3444,N_3445,N_3447,N_3448,N_3450,N_3451,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3462,N_3463,N_3464,N_3466,N_3467,N_3468,N_3469,N_3470,N_3472,N_3473,N_3474,N_3476,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3492,N_3495,N_3496,N_3497,N_3498,N_3500,N_3501,N_3502,N_3503,N_3505,N_3506,N_3508,N_3511,N_3512,N_3513,N_3515,N_3516,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3526,N_3527,N_3528,N_3529,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3538,N_3540,N_3541,N_3542,N_3543,N_3545,N_3546,N_3547,N_3548,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3561,N_3562,N_3565,N_3566,N_3567,N_3568,N_3569,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3581,N_3583,N_3584,N_3585,N_3586,N_3588,N_3590,N_3591,N_3592,N_3593,N_3594,N_3596,N_3597,N_3598,N_3600,N_3601,N_3602,N_3603,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3615,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3650,N_3654,N_3655,N_3656,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3682,N_3684,N_3687,N_3688,N_3689,N_3690,N_3692,N_3693,N_3694,N_3695,N_3696,N_3698,N_3699,N_3700,N_3701,N_3703,N_3705,N_3706,N_3707,N_3708,N_3709,N_3711,N_3712,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3723,N_3724,N_3725,N_3726,N_3727,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3755,N_3757,N_3758,N_3759,N_3761,N_3762,N_3763,N_3765,N_3768,N_3769,N_3770,N_3771,N_3772,N_3774,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3801,N_3802,N_3804,N_3805,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3836,N_3837,N_3838,N_3839,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3854,N_3855,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3867,N_3869,N_3871,N_3872,N_3873,N_3874,N_3876,N_3878,N_3879,N_3880,N_3882,N_3884,N_3885,N_3886,N_3889,N_3890,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3912,N_3913,N_3914,N_3915,N_3916,N_3920,N_3923,N_3924,N_3925,N_3926,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3941,N_3942,N_3943,N_3944,N_3945,N_3947,N_3948,N_3950,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3966,N_3967,N_3968,N_3970,N_3971,N_3972,N_3974,N_3975,N_3977,N_3978,N_3979,N_3980,N_3981,N_3984,N_3985,N_3987,N_3988,N_3991,N_3992,N_3993,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4004,N_4005,N_4008,N_4010,N_4013,N_4016,N_4017,N_4018,N_4020,N_4022,N_4023,N_4025,N_4026,N_4027,N_4029,N_4031,N_4033,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4042,N_4043,N_4044,N_4045,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4072,N_4073,N_4074,N_4075,N_4077,N_4078,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4120,N_4122,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4134,N_4135,N_4136,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4148,N_4149,N_4152,N_4153,N_4154,N_4155,N_4156,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4172,N_4173,N_4174,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4242,N_4243,N_4245,N_4246,N_4247,N_4249,N_4250,N_4253,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4281,N_4282,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4321,N_4322,N_4326,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4356,N_4357,N_4358,N_4359,N_4360,N_4364,N_4365,N_4366,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4377,N_4379,N_4381,N_4382,N_4383,N_4384,N_4386,N_4387,N_4388,N_4390,N_4391,N_4392,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4407,N_4408,N_4409,N_4413,N_4414,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4437,N_4438,N_4440,N_4442,N_4443,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4473,N_4474,N_4475,N_4476,N_4477,N_4479,N_4480,N_4482,N_4483,N_4485,N_4486,N_4487,N_4488,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4503,N_4504,N_4505,N_4506,N_4507,N_4509,N_4510,N_4511,N_4512,N_4513,N_4515,N_4516,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4533,N_4534,N_4535,N_4537,N_4538,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4551,N_4553,N_4554,N_4555,N_4557,N_4559,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4572,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4581,N_4582,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4623,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4645,N_4646,N_4648,N_4649,N_4650,N_4651,N_4653,N_4654,N_4655,N_4656,N_4657,N_4659,N_4660,N_4661,N_4662,N_4663,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4673,N_4674,N_4675,N_4676,N_4678,N_4680,N_4682,N_4683,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4704,N_4705,N_4706,N_4707,N_4708,N_4710,N_4711,N_4712,N_4713,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4723,N_4724,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4742,N_4744,N_4746,N_4747,N_4748,N_4751,N_4754,N_4755,N_4757,N_4758,N_4759,N_4760,N_4761,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4776,N_4778,N_4779,N_4780,N_4781,N_4783,N_4784,N_4786,N_4787,N_4788,N_4789,N_4791,N_4792,N_4794,N_4796,N_4797,N_4798,N_4799,N_4800,N_4802,N_4803,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4817,N_4819,N_4820,N_4821,N_4822,N_4823,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4837,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4853,N_4856,N_4857,N_4858,N_4859,N_4861,N_4862,N_4863,N_4864,N_4866,N_4867,N_4868,N_4869,N_4870,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4881,N_4884,N_4885,N_4886,N_4888,N_4889,N_4890,N_4891,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4906,N_4907,N_4908,N_4910,N_4912,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4931,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4945,N_4946,N_4947,N_4948,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4959,N_4960,N_4961,N_4964,N_4965,N_4966,N_4967,N_4968,N_4970,N_4971,N_4973,N_4974,N_4975,N_4976,N_4978,N_4979,N_4981,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_168,In_31);
nand U1 (N_1,In_398,In_18);
nor U2 (N_2,In_227,In_557);
or U3 (N_3,In_135,In_80);
xor U4 (N_4,In_24,In_698);
or U5 (N_5,In_79,In_43);
and U6 (N_6,In_309,In_125);
nor U7 (N_7,In_702,In_409);
and U8 (N_8,In_368,In_721);
nand U9 (N_9,In_123,In_52);
nor U10 (N_10,In_728,In_559);
xnor U11 (N_11,In_144,In_345);
and U12 (N_12,In_203,In_208);
nor U13 (N_13,In_406,In_133);
xor U14 (N_14,In_15,In_513);
nand U15 (N_15,In_556,In_419);
and U16 (N_16,In_654,In_648);
and U17 (N_17,In_548,In_141);
nor U18 (N_18,In_718,In_372);
nand U19 (N_19,In_277,In_365);
and U20 (N_20,In_418,In_480);
nand U21 (N_21,In_333,In_482);
and U22 (N_22,In_13,In_99);
nor U23 (N_23,In_514,In_349);
nor U24 (N_24,In_330,In_485);
and U25 (N_25,In_85,In_565);
nor U26 (N_26,In_222,In_447);
xor U27 (N_27,In_719,In_749);
and U28 (N_28,In_646,In_540);
nor U29 (N_29,In_645,In_744);
and U30 (N_30,In_252,In_132);
nand U31 (N_31,In_267,In_103);
nand U32 (N_32,In_561,In_490);
and U33 (N_33,In_710,In_301);
xnor U34 (N_34,In_61,In_148);
and U35 (N_35,In_190,In_36);
nand U36 (N_36,In_261,In_131);
nor U37 (N_37,In_631,In_332);
nor U38 (N_38,In_272,In_620);
xnor U39 (N_39,In_671,In_235);
nor U40 (N_40,In_126,In_165);
and U41 (N_41,In_680,In_436);
nand U42 (N_42,In_689,In_242);
or U43 (N_43,In_517,In_594);
and U44 (N_44,In_188,In_158);
nor U45 (N_45,In_285,In_88);
and U46 (N_46,In_662,In_536);
and U47 (N_47,In_236,In_380);
nand U48 (N_48,In_644,In_101);
and U49 (N_49,In_164,In_474);
nand U50 (N_50,In_588,In_128);
nor U51 (N_51,In_48,In_110);
nand U52 (N_52,In_558,In_497);
xor U53 (N_53,In_170,In_628);
nand U54 (N_54,In_218,In_467);
nand U55 (N_55,In_280,In_395);
and U56 (N_56,In_313,In_106);
xor U57 (N_57,In_414,In_475);
nand U58 (N_58,In_707,In_295);
and U59 (N_59,In_528,In_342);
and U60 (N_60,In_499,In_733);
nand U61 (N_61,In_373,In_120);
xnor U62 (N_62,In_383,In_531);
nor U63 (N_63,In_351,In_56);
nor U64 (N_64,In_745,In_529);
nand U65 (N_65,In_576,In_326);
and U66 (N_66,In_569,In_434);
nor U67 (N_67,In_509,In_274);
and U68 (N_68,In_535,In_407);
nor U69 (N_69,In_45,In_362);
nand U70 (N_70,In_5,In_316);
nor U71 (N_71,In_667,In_130);
or U72 (N_72,In_462,In_382);
or U73 (N_73,In_675,In_206);
nand U74 (N_74,In_183,In_738);
nand U75 (N_75,In_108,In_697);
and U76 (N_76,In_303,In_38);
or U77 (N_77,In_174,In_624);
or U78 (N_78,In_466,In_178);
or U79 (N_79,In_520,In_371);
and U80 (N_80,In_248,In_69);
nand U81 (N_81,In_181,In_265);
or U82 (N_82,In_622,In_118);
xor U83 (N_83,In_401,In_172);
nor U84 (N_84,In_715,In_153);
nand U85 (N_85,In_220,In_547);
or U86 (N_86,In_605,In_578);
nor U87 (N_87,In_604,In_618);
nor U88 (N_88,In_672,In_228);
nor U89 (N_89,In_636,In_384);
nor U90 (N_90,In_162,In_417);
and U91 (N_91,In_611,In_609);
and U92 (N_92,In_608,In_601);
and U93 (N_93,In_399,In_606);
or U94 (N_94,In_364,In_64);
nand U95 (N_95,In_655,In_276);
nand U96 (N_96,In_484,In_457);
nor U97 (N_97,In_93,In_35);
or U98 (N_98,In_592,In_584);
and U99 (N_99,In_129,In_59);
or U100 (N_100,In_483,In_319);
nand U101 (N_101,In_98,In_723);
nand U102 (N_102,In_633,In_302);
and U103 (N_103,In_177,In_327);
nor U104 (N_104,In_214,In_338);
nand U105 (N_105,In_508,In_20);
nor U106 (N_106,In_217,In_269);
xnor U107 (N_107,In_408,In_202);
nor U108 (N_108,In_374,In_344);
nand U109 (N_109,In_403,In_109);
nor U110 (N_110,In_534,In_353);
nor U111 (N_111,In_432,In_647);
nor U112 (N_112,In_427,In_659);
or U113 (N_113,In_17,In_113);
nand U114 (N_114,In_3,In_154);
or U115 (N_115,In_107,In_637);
or U116 (N_116,In_155,In_694);
and U117 (N_117,In_670,In_89);
nand U118 (N_118,In_652,In_375);
or U119 (N_119,In_489,In_270);
or U120 (N_120,In_640,In_521);
and U121 (N_121,In_727,In_713);
and U122 (N_122,In_264,In_431);
nor U123 (N_123,In_415,In_639);
nor U124 (N_124,In_321,In_307);
nor U125 (N_125,In_530,In_26);
or U126 (N_126,In_502,In_10);
nor U127 (N_127,In_204,In_6);
nand U128 (N_128,In_86,In_273);
xnor U129 (N_129,In_437,In_136);
or U130 (N_130,In_479,In_424);
and U131 (N_131,In_630,In_137);
nand U132 (N_132,In_200,In_615);
and U133 (N_133,In_526,In_405);
nor U134 (N_134,In_71,In_567);
or U135 (N_135,In_463,In_450);
or U136 (N_136,In_385,In_741);
xor U137 (N_137,In_39,In_552);
or U138 (N_138,In_305,In_82);
and U139 (N_139,In_614,In_68);
nand U140 (N_140,In_369,In_421);
or U141 (N_141,In_116,In_674);
xor U142 (N_142,In_735,In_230);
and U143 (N_143,In_501,In_104);
and U144 (N_144,In_145,In_564);
nand U145 (N_145,In_241,In_105);
nand U146 (N_146,In_726,In_481);
xor U147 (N_147,In_102,In_322);
and U148 (N_148,In_542,In_83);
or U149 (N_149,In_677,In_159);
nor U150 (N_150,In_711,In_658);
or U151 (N_151,In_729,In_14);
nor U152 (N_152,In_100,In_152);
xor U153 (N_153,In_247,In_323);
nand U154 (N_154,In_494,In_673);
nor U155 (N_155,In_324,In_524);
and U156 (N_156,In_669,In_394);
and U157 (N_157,In_76,In_579);
or U158 (N_158,In_90,In_549);
nand U159 (N_159,In_392,In_435);
xor U160 (N_160,In_705,In_21);
and U161 (N_161,In_532,In_32);
nand U162 (N_162,In_492,In_404);
or U163 (N_163,In_67,In_459);
and U164 (N_164,In_232,In_495);
nand U165 (N_165,In_590,In_629);
nand U166 (N_166,In_297,In_266);
nor U167 (N_167,In_681,In_439);
or U168 (N_168,In_461,In_597);
nor U169 (N_169,In_127,In_732);
nand U170 (N_170,In_456,In_198);
nor U171 (N_171,In_358,In_207);
or U172 (N_172,In_650,In_176);
or U173 (N_173,In_411,In_453);
and U174 (N_174,In_151,In_498);
or U175 (N_175,In_625,In_448);
nor U176 (N_176,In_238,In_396);
or U177 (N_177,In_237,In_317);
and U178 (N_178,In_171,In_550);
xnor U179 (N_179,In_600,In_7);
nand U180 (N_180,In_527,In_537);
or U181 (N_181,In_335,In_161);
nand U182 (N_182,In_25,In_336);
or U183 (N_183,In_746,In_286);
nor U184 (N_184,In_660,In_568);
nor U185 (N_185,In_449,In_476);
and U186 (N_186,In_229,In_97);
and U187 (N_187,In_668,In_219);
xor U188 (N_188,In_65,In_92);
or U189 (N_189,In_742,In_740);
nand U190 (N_190,In_693,In_402);
or U191 (N_191,In_271,In_470);
and U192 (N_192,In_94,In_377);
or U193 (N_193,In_337,In_391);
nor U194 (N_194,In_268,In_255);
nand U195 (N_195,In_251,In_44);
or U196 (N_196,In_512,In_641);
and U197 (N_197,In_525,In_743);
nor U198 (N_198,In_119,In_416);
or U199 (N_199,In_124,In_621);
nand U200 (N_200,In_186,In_16);
or U201 (N_201,In_653,In_246);
and U202 (N_202,In_196,In_701);
nor U203 (N_203,In_682,In_306);
and U204 (N_204,In_666,In_199);
or U205 (N_205,In_41,In_390);
nand U206 (N_206,In_685,In_638);
nand U207 (N_207,In_185,In_656);
nand U208 (N_208,In_748,In_50);
and U209 (N_209,In_341,In_360);
or U210 (N_210,In_423,In_47);
and U211 (N_211,In_379,In_503);
nand U212 (N_212,In_343,In_114);
nor U213 (N_213,In_122,In_320);
xor U214 (N_214,In_739,In_376);
xor U215 (N_215,In_197,In_4);
and U216 (N_216,In_704,In_298);
nand U217 (N_217,In_78,In_291);
nor U218 (N_218,In_573,In_292);
nand U219 (N_219,In_23,In_477);
nand U220 (N_220,In_506,In_722);
or U221 (N_221,In_239,In_279);
nand U222 (N_222,In_560,In_209);
nor U223 (N_223,In_166,In_487);
nor U224 (N_224,In_262,In_410);
or U225 (N_225,In_426,In_626);
nand U226 (N_226,In_553,In_142);
nand U227 (N_227,In_692,In_37);
or U228 (N_228,In_231,In_635);
or U229 (N_229,In_473,In_551);
xnor U230 (N_230,In_356,In_585);
nand U231 (N_231,In_486,In_62);
and U232 (N_232,In_212,In_533);
or U233 (N_233,In_554,In_308);
or U234 (N_234,In_632,In_40);
nand U235 (N_235,In_593,In_312);
nor U236 (N_236,In_596,In_706);
xor U237 (N_237,In_213,In_175);
nor U238 (N_238,In_49,In_679);
and U239 (N_239,In_731,In_224);
and U240 (N_240,In_451,In_9);
and U241 (N_241,In_205,In_77);
nand U242 (N_242,In_370,In_651);
or U243 (N_243,In_329,In_354);
nor U244 (N_244,In_357,In_304);
nand U245 (N_245,In_96,In_589);
nand U246 (N_246,In_300,In_577);
xor U247 (N_247,In_250,In_63);
and U248 (N_248,In_504,In_42);
nand U249 (N_249,In_444,In_455);
nand U250 (N_250,In_195,In_240);
or U251 (N_251,In_378,In_642);
and U252 (N_252,In_683,In_57);
or U253 (N_253,In_348,In_328);
xor U254 (N_254,In_257,In_464);
or U255 (N_255,In_623,In_574);
and U256 (N_256,In_747,In_734);
or U257 (N_257,In_215,In_602);
and U258 (N_258,In_310,In_296);
and U259 (N_259,In_189,In_446);
nand U260 (N_260,In_27,In_367);
nand U261 (N_261,In_544,In_339);
and U262 (N_262,In_516,In_422);
and U263 (N_263,In_442,In_496);
nand U264 (N_264,In_657,In_34);
and U265 (N_265,In_294,In_259);
and U266 (N_266,In_58,In_500);
nand U267 (N_267,In_182,In_393);
nand U268 (N_268,In_580,In_420);
or U269 (N_269,In_613,In_138);
xnor U270 (N_270,In_260,In_610);
xnor U271 (N_271,In_737,In_381);
and U272 (N_272,In_187,In_433);
xor U273 (N_273,In_712,In_19);
or U274 (N_274,In_290,In_676);
or U275 (N_275,In_562,In_582);
and U276 (N_276,In_688,In_717);
nand U277 (N_277,In_245,In_387);
nand U278 (N_278,In_256,In_361);
nand U279 (N_279,In_157,In_8);
nor U280 (N_280,In_334,In_73);
and U281 (N_281,In_661,In_193);
and U282 (N_282,In_507,In_95);
nor U283 (N_283,In_325,In_695);
nor U284 (N_284,In_598,In_599);
nand U285 (N_285,In_173,In_143);
nand U286 (N_286,In_425,In_440);
nand U287 (N_287,In_583,In_488);
nand U288 (N_288,In_684,In_244);
nor U289 (N_289,In_134,In_318);
and U290 (N_290,In_346,In_619);
and U291 (N_291,In_720,In_117);
xnor U292 (N_292,In_60,In_180);
nor U293 (N_293,In_716,In_288);
and U294 (N_294,In_192,In_179);
nand U295 (N_295,In_546,In_150);
or U296 (N_296,In_359,In_572);
and U297 (N_297,In_538,In_53);
and U298 (N_298,In_591,In_289);
nor U299 (N_299,In_340,In_350);
nand U300 (N_300,In_283,In_627);
nor U301 (N_301,In_581,In_115);
and U302 (N_302,In_703,In_539);
or U303 (N_303,In_445,In_81);
and U304 (N_304,In_649,In_263);
nand U305 (N_305,In_545,In_690);
and U306 (N_306,In_234,In_438);
nor U307 (N_307,In_33,In_221);
and U308 (N_308,In_147,In_612);
or U309 (N_309,In_428,In_510);
xor U310 (N_310,In_347,In_566);
and U311 (N_311,In_29,In_571);
nor U312 (N_312,In_575,In_472);
or U313 (N_313,In_730,In_412);
xor U314 (N_314,In_315,In_468);
and U315 (N_315,In_299,In_515);
and U316 (N_316,In_523,In_555);
nor U317 (N_317,In_687,In_314);
or U318 (N_318,In_441,In_11);
or U319 (N_319,In_66,In_191);
nand U320 (N_320,In_429,In_160);
nor U321 (N_321,In_281,In_2);
or U322 (N_322,In_458,In_452);
nand U323 (N_323,In_216,In_55);
nand U324 (N_324,In_478,In_696);
nand U325 (N_325,In_570,In_617);
or U326 (N_326,In_587,In_519);
xnor U327 (N_327,In_725,In_543);
or U328 (N_328,In_91,In_714);
nand U329 (N_329,In_210,In_643);
or U330 (N_330,In_184,In_22);
nor U331 (N_331,In_454,In_471);
nor U332 (N_332,In_54,In_709);
nor U333 (N_333,In_469,In_388);
nand U334 (N_334,In_194,In_686);
xor U335 (N_335,In_700,In_233);
xor U336 (N_336,In_30,In_699);
and U337 (N_337,In_603,In_140);
nor U338 (N_338,In_253,In_28);
nor U339 (N_339,In_163,In_413);
or U340 (N_340,In_287,In_465);
and U341 (N_341,In_664,In_400);
xor U342 (N_342,In_284,In_331);
nand U343 (N_343,In_121,In_258);
nand U344 (N_344,In_111,In_149);
nand U345 (N_345,In_511,In_616);
and U346 (N_346,In_595,In_74);
nand U347 (N_347,In_460,In_678);
nand U348 (N_348,In_201,In_169);
or U349 (N_349,In_505,In_541);
nor U350 (N_350,In_139,In_708);
or U351 (N_351,In_634,In_46);
nand U352 (N_352,In_0,In_563);
nand U353 (N_353,In_223,In_311);
and U354 (N_354,In_691,In_278);
nand U355 (N_355,In_491,In_665);
or U356 (N_356,In_443,In_518);
and U357 (N_357,In_243,In_249);
and U358 (N_358,In_87,In_366);
nand U359 (N_359,In_363,In_736);
or U360 (N_360,In_282,In_156);
nor U361 (N_361,In_355,In_493);
or U362 (N_362,In_386,In_397);
nand U363 (N_363,In_663,In_167);
or U364 (N_364,In_522,In_75);
nor U365 (N_365,In_586,In_1);
nor U366 (N_366,In_293,In_226);
or U367 (N_367,In_607,In_254);
or U368 (N_368,In_146,In_225);
and U369 (N_369,In_211,In_84);
nand U370 (N_370,In_51,In_352);
or U371 (N_371,In_430,In_724);
nand U372 (N_372,In_275,In_72);
or U373 (N_373,In_12,In_389);
nand U374 (N_374,In_112,In_70);
nor U375 (N_375,In_745,In_86);
nand U376 (N_376,In_342,In_263);
and U377 (N_377,In_287,In_97);
nand U378 (N_378,In_466,In_334);
and U379 (N_379,In_478,In_599);
or U380 (N_380,In_532,In_142);
and U381 (N_381,In_244,In_662);
nand U382 (N_382,In_635,In_318);
nand U383 (N_383,In_634,In_636);
nor U384 (N_384,In_589,In_182);
or U385 (N_385,In_399,In_475);
nor U386 (N_386,In_92,In_498);
nor U387 (N_387,In_591,In_256);
nor U388 (N_388,In_60,In_71);
nand U389 (N_389,In_709,In_530);
nand U390 (N_390,In_329,In_680);
or U391 (N_391,In_589,In_135);
or U392 (N_392,In_500,In_188);
or U393 (N_393,In_433,In_163);
nor U394 (N_394,In_310,In_446);
nor U395 (N_395,In_264,In_549);
nand U396 (N_396,In_642,In_13);
xor U397 (N_397,In_224,In_532);
nand U398 (N_398,In_185,In_457);
nor U399 (N_399,In_579,In_665);
nor U400 (N_400,In_448,In_728);
and U401 (N_401,In_504,In_455);
and U402 (N_402,In_152,In_214);
or U403 (N_403,In_597,In_571);
or U404 (N_404,In_15,In_542);
nand U405 (N_405,In_304,In_450);
and U406 (N_406,In_159,In_464);
nand U407 (N_407,In_653,In_532);
and U408 (N_408,In_600,In_248);
and U409 (N_409,In_339,In_555);
nand U410 (N_410,In_612,In_89);
and U411 (N_411,In_63,In_507);
nand U412 (N_412,In_562,In_155);
nand U413 (N_413,In_394,In_600);
or U414 (N_414,In_481,In_275);
or U415 (N_415,In_89,In_614);
nand U416 (N_416,In_602,In_738);
xor U417 (N_417,In_151,In_124);
and U418 (N_418,In_694,In_567);
and U419 (N_419,In_7,In_529);
or U420 (N_420,In_189,In_595);
nor U421 (N_421,In_700,In_340);
or U422 (N_422,In_607,In_744);
nor U423 (N_423,In_606,In_44);
and U424 (N_424,In_275,In_214);
and U425 (N_425,In_53,In_304);
nor U426 (N_426,In_304,In_316);
xnor U427 (N_427,In_241,In_229);
or U428 (N_428,In_347,In_444);
and U429 (N_429,In_223,In_550);
nand U430 (N_430,In_314,In_288);
xor U431 (N_431,In_497,In_200);
or U432 (N_432,In_117,In_254);
nor U433 (N_433,In_380,In_494);
nand U434 (N_434,In_476,In_42);
and U435 (N_435,In_525,In_381);
and U436 (N_436,In_284,In_235);
or U437 (N_437,In_475,In_599);
nor U438 (N_438,In_154,In_498);
xor U439 (N_439,In_492,In_732);
nand U440 (N_440,In_663,In_487);
and U441 (N_441,In_375,In_682);
and U442 (N_442,In_143,In_721);
or U443 (N_443,In_141,In_191);
nand U444 (N_444,In_644,In_331);
xor U445 (N_445,In_156,In_25);
or U446 (N_446,In_213,In_565);
or U447 (N_447,In_634,In_706);
or U448 (N_448,In_12,In_52);
and U449 (N_449,In_342,In_126);
and U450 (N_450,In_692,In_107);
xor U451 (N_451,In_380,In_678);
nor U452 (N_452,In_352,In_46);
or U453 (N_453,In_618,In_203);
nor U454 (N_454,In_628,In_389);
nand U455 (N_455,In_495,In_446);
or U456 (N_456,In_432,In_393);
and U457 (N_457,In_661,In_503);
or U458 (N_458,In_50,In_460);
nor U459 (N_459,In_275,In_615);
or U460 (N_460,In_303,In_203);
nand U461 (N_461,In_30,In_193);
and U462 (N_462,In_61,In_728);
nor U463 (N_463,In_551,In_471);
nand U464 (N_464,In_710,In_592);
nand U465 (N_465,In_297,In_263);
and U466 (N_466,In_722,In_622);
or U467 (N_467,In_62,In_135);
nand U468 (N_468,In_691,In_348);
nand U469 (N_469,In_699,In_80);
or U470 (N_470,In_45,In_273);
and U471 (N_471,In_622,In_506);
and U472 (N_472,In_97,In_44);
or U473 (N_473,In_340,In_699);
or U474 (N_474,In_230,In_524);
or U475 (N_475,In_242,In_46);
nand U476 (N_476,In_358,In_558);
nand U477 (N_477,In_80,In_597);
nor U478 (N_478,In_446,In_705);
nand U479 (N_479,In_636,In_733);
and U480 (N_480,In_529,In_548);
or U481 (N_481,In_18,In_688);
nand U482 (N_482,In_473,In_708);
and U483 (N_483,In_331,In_308);
nand U484 (N_484,In_459,In_531);
or U485 (N_485,In_330,In_56);
nor U486 (N_486,In_715,In_239);
nand U487 (N_487,In_573,In_718);
and U488 (N_488,In_615,In_302);
nand U489 (N_489,In_660,In_486);
or U490 (N_490,In_155,In_482);
and U491 (N_491,In_541,In_227);
nand U492 (N_492,In_110,In_96);
and U493 (N_493,In_272,In_407);
or U494 (N_494,In_516,In_78);
nand U495 (N_495,In_588,In_151);
and U496 (N_496,In_279,In_155);
nand U497 (N_497,In_101,In_389);
and U498 (N_498,In_277,In_172);
nand U499 (N_499,In_230,In_421);
and U500 (N_500,In_506,In_523);
xor U501 (N_501,In_624,In_457);
nor U502 (N_502,In_246,In_396);
nand U503 (N_503,In_486,In_270);
nor U504 (N_504,In_206,In_22);
nand U505 (N_505,In_728,In_349);
nor U506 (N_506,In_456,In_243);
nor U507 (N_507,In_726,In_392);
nand U508 (N_508,In_138,In_134);
and U509 (N_509,In_22,In_443);
and U510 (N_510,In_419,In_198);
nor U511 (N_511,In_272,In_630);
nor U512 (N_512,In_599,In_701);
or U513 (N_513,In_732,In_475);
nor U514 (N_514,In_502,In_0);
nor U515 (N_515,In_484,In_648);
or U516 (N_516,In_389,In_504);
and U517 (N_517,In_593,In_336);
and U518 (N_518,In_656,In_658);
nor U519 (N_519,In_721,In_192);
or U520 (N_520,In_237,In_9);
and U521 (N_521,In_232,In_420);
or U522 (N_522,In_405,In_91);
nor U523 (N_523,In_202,In_58);
xnor U524 (N_524,In_311,In_708);
and U525 (N_525,In_350,In_382);
nand U526 (N_526,In_274,In_67);
nor U527 (N_527,In_526,In_281);
or U528 (N_528,In_618,In_377);
nand U529 (N_529,In_172,In_235);
nand U530 (N_530,In_561,In_691);
and U531 (N_531,In_459,In_230);
and U532 (N_532,In_244,In_603);
nand U533 (N_533,In_269,In_96);
or U534 (N_534,In_38,In_515);
nand U535 (N_535,In_357,In_74);
nor U536 (N_536,In_630,In_207);
and U537 (N_537,In_741,In_177);
and U538 (N_538,In_59,In_81);
or U539 (N_539,In_376,In_406);
nor U540 (N_540,In_654,In_497);
xnor U541 (N_541,In_31,In_667);
xor U542 (N_542,In_287,In_453);
xor U543 (N_543,In_224,In_402);
nand U544 (N_544,In_687,In_151);
and U545 (N_545,In_312,In_85);
nand U546 (N_546,In_731,In_461);
nor U547 (N_547,In_331,In_587);
nand U548 (N_548,In_544,In_604);
and U549 (N_549,In_618,In_638);
nor U550 (N_550,In_548,In_102);
nor U551 (N_551,In_12,In_207);
nor U552 (N_552,In_197,In_591);
nand U553 (N_553,In_709,In_612);
nand U554 (N_554,In_204,In_97);
nand U555 (N_555,In_95,In_342);
and U556 (N_556,In_458,In_90);
and U557 (N_557,In_473,In_118);
or U558 (N_558,In_723,In_614);
or U559 (N_559,In_494,In_235);
nor U560 (N_560,In_186,In_534);
nand U561 (N_561,In_538,In_672);
xor U562 (N_562,In_310,In_204);
nand U563 (N_563,In_501,In_509);
nor U564 (N_564,In_75,In_64);
xor U565 (N_565,In_404,In_352);
and U566 (N_566,In_198,In_547);
or U567 (N_567,In_583,In_173);
nand U568 (N_568,In_37,In_716);
nand U569 (N_569,In_358,In_221);
or U570 (N_570,In_533,In_75);
nand U571 (N_571,In_74,In_390);
or U572 (N_572,In_270,In_352);
and U573 (N_573,In_445,In_520);
nand U574 (N_574,In_505,In_684);
xnor U575 (N_575,In_226,In_201);
nor U576 (N_576,In_454,In_607);
or U577 (N_577,In_179,In_186);
nand U578 (N_578,In_0,In_73);
and U579 (N_579,In_463,In_135);
nand U580 (N_580,In_209,In_232);
nand U581 (N_581,In_74,In_351);
nor U582 (N_582,In_11,In_531);
nor U583 (N_583,In_118,In_71);
and U584 (N_584,In_412,In_192);
or U585 (N_585,In_718,In_118);
and U586 (N_586,In_144,In_563);
and U587 (N_587,In_297,In_434);
xor U588 (N_588,In_97,In_620);
or U589 (N_589,In_609,In_532);
nand U590 (N_590,In_15,In_668);
nand U591 (N_591,In_376,In_584);
nand U592 (N_592,In_619,In_267);
nor U593 (N_593,In_499,In_328);
nand U594 (N_594,In_748,In_638);
or U595 (N_595,In_614,In_409);
nand U596 (N_596,In_472,In_224);
and U597 (N_597,In_394,In_522);
or U598 (N_598,In_233,In_530);
xnor U599 (N_599,In_651,In_463);
nor U600 (N_600,In_744,In_190);
xnor U601 (N_601,In_101,In_71);
nand U602 (N_602,In_339,In_211);
nand U603 (N_603,In_467,In_377);
nor U604 (N_604,In_135,In_378);
nand U605 (N_605,In_428,In_40);
xor U606 (N_606,In_404,In_219);
nand U607 (N_607,In_428,In_577);
nor U608 (N_608,In_126,In_144);
nor U609 (N_609,In_276,In_696);
nor U610 (N_610,In_744,In_19);
or U611 (N_611,In_718,In_393);
and U612 (N_612,In_530,In_592);
nor U613 (N_613,In_260,In_210);
nor U614 (N_614,In_54,In_513);
nand U615 (N_615,In_81,In_609);
nor U616 (N_616,In_575,In_612);
xnor U617 (N_617,In_472,In_137);
nand U618 (N_618,In_359,In_210);
nor U619 (N_619,In_452,In_9);
or U620 (N_620,In_544,In_599);
xnor U621 (N_621,In_588,In_86);
nand U622 (N_622,In_269,In_337);
nor U623 (N_623,In_239,In_648);
nand U624 (N_624,In_526,In_717);
or U625 (N_625,In_414,In_708);
or U626 (N_626,In_235,In_734);
nor U627 (N_627,In_581,In_194);
nor U628 (N_628,In_694,In_250);
nor U629 (N_629,In_310,In_707);
or U630 (N_630,In_256,In_580);
nand U631 (N_631,In_346,In_562);
nand U632 (N_632,In_244,In_18);
nand U633 (N_633,In_437,In_324);
xor U634 (N_634,In_639,In_693);
xnor U635 (N_635,In_690,In_596);
xnor U636 (N_636,In_116,In_398);
and U637 (N_637,In_335,In_162);
or U638 (N_638,In_660,In_329);
or U639 (N_639,In_323,In_431);
nor U640 (N_640,In_724,In_189);
or U641 (N_641,In_626,In_579);
nand U642 (N_642,In_424,In_417);
and U643 (N_643,In_746,In_374);
nor U644 (N_644,In_116,In_678);
and U645 (N_645,In_190,In_397);
nand U646 (N_646,In_731,In_111);
xor U647 (N_647,In_113,In_114);
or U648 (N_648,In_635,In_330);
nor U649 (N_649,In_81,In_671);
nor U650 (N_650,In_608,In_287);
nor U651 (N_651,In_661,In_592);
and U652 (N_652,In_657,In_157);
and U653 (N_653,In_454,In_507);
nand U654 (N_654,In_123,In_621);
and U655 (N_655,In_486,In_639);
nand U656 (N_656,In_409,In_15);
nand U657 (N_657,In_732,In_83);
and U658 (N_658,In_717,In_86);
and U659 (N_659,In_224,In_587);
xnor U660 (N_660,In_60,In_693);
or U661 (N_661,In_368,In_197);
nand U662 (N_662,In_350,In_56);
nor U663 (N_663,In_474,In_124);
nor U664 (N_664,In_292,In_369);
and U665 (N_665,In_113,In_482);
nand U666 (N_666,In_262,In_163);
xnor U667 (N_667,In_192,In_324);
xnor U668 (N_668,In_469,In_127);
and U669 (N_669,In_706,In_554);
nand U670 (N_670,In_617,In_665);
and U671 (N_671,In_34,In_361);
and U672 (N_672,In_448,In_198);
or U673 (N_673,In_30,In_110);
nor U674 (N_674,In_226,In_702);
and U675 (N_675,In_474,In_410);
or U676 (N_676,In_157,In_612);
nand U677 (N_677,In_378,In_445);
xor U678 (N_678,In_505,In_510);
and U679 (N_679,In_486,In_730);
nor U680 (N_680,In_212,In_285);
and U681 (N_681,In_217,In_583);
xor U682 (N_682,In_371,In_205);
nor U683 (N_683,In_476,In_408);
or U684 (N_684,In_596,In_91);
and U685 (N_685,In_617,In_304);
xor U686 (N_686,In_487,In_210);
or U687 (N_687,In_667,In_604);
and U688 (N_688,In_510,In_560);
nor U689 (N_689,In_519,In_297);
and U690 (N_690,In_57,In_175);
xnor U691 (N_691,In_360,In_167);
or U692 (N_692,In_50,In_326);
or U693 (N_693,In_55,In_687);
and U694 (N_694,In_11,In_617);
and U695 (N_695,In_195,In_237);
nand U696 (N_696,In_149,In_748);
nor U697 (N_697,In_427,In_160);
nand U698 (N_698,In_693,In_666);
nor U699 (N_699,In_610,In_432);
xnor U700 (N_700,In_657,In_138);
nor U701 (N_701,In_252,In_353);
or U702 (N_702,In_279,In_448);
nor U703 (N_703,In_311,In_569);
nand U704 (N_704,In_210,In_606);
or U705 (N_705,In_492,In_514);
nor U706 (N_706,In_255,In_281);
nor U707 (N_707,In_306,In_426);
nand U708 (N_708,In_118,In_443);
nand U709 (N_709,In_664,In_366);
and U710 (N_710,In_344,In_283);
nand U711 (N_711,In_288,In_31);
nand U712 (N_712,In_94,In_496);
or U713 (N_713,In_161,In_594);
or U714 (N_714,In_148,In_664);
and U715 (N_715,In_178,In_432);
nor U716 (N_716,In_649,In_694);
and U717 (N_717,In_601,In_723);
nand U718 (N_718,In_134,In_629);
and U719 (N_719,In_227,In_89);
nor U720 (N_720,In_367,In_154);
nor U721 (N_721,In_343,In_50);
and U722 (N_722,In_614,In_239);
nand U723 (N_723,In_470,In_113);
and U724 (N_724,In_504,In_326);
or U725 (N_725,In_501,In_220);
and U726 (N_726,In_381,In_135);
or U727 (N_727,In_110,In_327);
or U728 (N_728,In_171,In_313);
nand U729 (N_729,In_245,In_452);
and U730 (N_730,In_309,In_217);
nor U731 (N_731,In_737,In_322);
xnor U732 (N_732,In_364,In_332);
or U733 (N_733,In_648,In_510);
and U734 (N_734,In_401,In_353);
nor U735 (N_735,In_726,In_32);
xor U736 (N_736,In_127,In_502);
nor U737 (N_737,In_97,In_674);
and U738 (N_738,In_171,In_195);
nand U739 (N_739,In_269,In_739);
nand U740 (N_740,In_327,In_231);
or U741 (N_741,In_523,In_359);
nand U742 (N_742,In_481,In_86);
nor U743 (N_743,In_327,In_186);
nand U744 (N_744,In_156,In_40);
or U745 (N_745,In_613,In_86);
or U746 (N_746,In_686,In_163);
nor U747 (N_747,In_508,In_461);
or U748 (N_748,In_612,In_512);
and U749 (N_749,In_254,In_674);
or U750 (N_750,In_497,In_108);
nor U751 (N_751,In_623,In_190);
xnor U752 (N_752,In_696,In_86);
nand U753 (N_753,In_34,In_425);
and U754 (N_754,In_109,In_277);
and U755 (N_755,In_401,In_474);
or U756 (N_756,In_706,In_516);
xnor U757 (N_757,In_29,In_438);
nor U758 (N_758,In_119,In_697);
or U759 (N_759,In_180,In_715);
nor U760 (N_760,In_483,In_732);
xnor U761 (N_761,In_490,In_376);
or U762 (N_762,In_569,In_339);
nor U763 (N_763,In_246,In_13);
nor U764 (N_764,In_590,In_76);
and U765 (N_765,In_22,In_621);
nand U766 (N_766,In_205,In_721);
and U767 (N_767,In_257,In_121);
xor U768 (N_768,In_38,In_112);
and U769 (N_769,In_675,In_664);
nor U770 (N_770,In_334,In_570);
nand U771 (N_771,In_539,In_206);
and U772 (N_772,In_436,In_269);
xnor U773 (N_773,In_354,In_182);
nand U774 (N_774,In_547,In_126);
nand U775 (N_775,In_731,In_691);
or U776 (N_776,In_585,In_393);
or U777 (N_777,In_256,In_741);
or U778 (N_778,In_695,In_17);
nor U779 (N_779,In_521,In_391);
and U780 (N_780,In_320,In_569);
or U781 (N_781,In_248,In_256);
or U782 (N_782,In_225,In_541);
or U783 (N_783,In_371,In_168);
nor U784 (N_784,In_74,In_447);
nand U785 (N_785,In_642,In_113);
or U786 (N_786,In_122,In_474);
and U787 (N_787,In_557,In_609);
or U788 (N_788,In_672,In_365);
nor U789 (N_789,In_355,In_434);
nand U790 (N_790,In_730,In_69);
nor U791 (N_791,In_557,In_90);
xnor U792 (N_792,In_403,In_616);
nor U793 (N_793,In_1,In_584);
or U794 (N_794,In_659,In_278);
nor U795 (N_795,In_93,In_354);
or U796 (N_796,In_140,In_132);
and U797 (N_797,In_93,In_406);
and U798 (N_798,In_81,In_696);
xor U799 (N_799,In_419,In_486);
and U800 (N_800,In_589,In_278);
nor U801 (N_801,In_604,In_689);
and U802 (N_802,In_373,In_180);
nand U803 (N_803,In_545,In_10);
nand U804 (N_804,In_304,In_503);
nor U805 (N_805,In_45,In_334);
or U806 (N_806,In_10,In_532);
or U807 (N_807,In_87,In_299);
nor U808 (N_808,In_221,In_699);
nand U809 (N_809,In_747,In_651);
or U810 (N_810,In_550,In_151);
nand U811 (N_811,In_38,In_26);
nand U812 (N_812,In_254,In_482);
nand U813 (N_813,In_633,In_8);
nand U814 (N_814,In_248,In_467);
or U815 (N_815,In_324,In_459);
or U816 (N_816,In_250,In_433);
and U817 (N_817,In_152,In_489);
nor U818 (N_818,In_496,In_48);
nor U819 (N_819,In_591,In_284);
xor U820 (N_820,In_576,In_301);
and U821 (N_821,In_716,In_246);
nor U822 (N_822,In_46,In_362);
and U823 (N_823,In_729,In_212);
nor U824 (N_824,In_726,In_4);
or U825 (N_825,In_605,In_345);
and U826 (N_826,In_395,In_281);
and U827 (N_827,In_730,In_38);
and U828 (N_828,In_506,In_307);
or U829 (N_829,In_214,In_520);
and U830 (N_830,In_492,In_256);
or U831 (N_831,In_473,In_600);
or U832 (N_832,In_282,In_90);
nor U833 (N_833,In_88,In_381);
and U834 (N_834,In_469,In_401);
nor U835 (N_835,In_324,In_487);
and U836 (N_836,In_329,In_704);
and U837 (N_837,In_733,In_253);
or U838 (N_838,In_156,In_698);
nand U839 (N_839,In_65,In_226);
or U840 (N_840,In_212,In_112);
nand U841 (N_841,In_135,In_704);
or U842 (N_842,In_511,In_716);
nor U843 (N_843,In_361,In_54);
nand U844 (N_844,In_672,In_27);
nor U845 (N_845,In_314,In_163);
nand U846 (N_846,In_513,In_99);
nand U847 (N_847,In_109,In_450);
xor U848 (N_848,In_732,In_452);
or U849 (N_849,In_594,In_457);
nor U850 (N_850,In_683,In_533);
and U851 (N_851,In_686,In_649);
or U852 (N_852,In_26,In_682);
and U853 (N_853,In_502,In_475);
and U854 (N_854,In_602,In_406);
and U855 (N_855,In_145,In_13);
nand U856 (N_856,In_371,In_273);
and U857 (N_857,In_726,In_278);
xnor U858 (N_858,In_216,In_360);
nor U859 (N_859,In_650,In_594);
nor U860 (N_860,In_28,In_647);
or U861 (N_861,In_679,In_407);
nor U862 (N_862,In_562,In_741);
and U863 (N_863,In_737,In_25);
and U864 (N_864,In_524,In_292);
nor U865 (N_865,In_180,In_590);
nand U866 (N_866,In_96,In_615);
nor U867 (N_867,In_678,In_204);
xor U868 (N_868,In_584,In_541);
or U869 (N_869,In_510,In_725);
or U870 (N_870,In_377,In_561);
or U871 (N_871,In_319,In_341);
or U872 (N_872,In_526,In_158);
or U873 (N_873,In_472,In_292);
nor U874 (N_874,In_341,In_128);
and U875 (N_875,In_42,In_398);
and U876 (N_876,In_576,In_711);
nand U877 (N_877,In_39,In_338);
nand U878 (N_878,In_669,In_612);
and U879 (N_879,In_372,In_254);
or U880 (N_880,In_9,In_351);
nor U881 (N_881,In_622,In_391);
nor U882 (N_882,In_236,In_667);
or U883 (N_883,In_566,In_301);
and U884 (N_884,In_535,In_258);
nor U885 (N_885,In_495,In_19);
nor U886 (N_886,In_677,In_169);
or U887 (N_887,In_428,In_544);
xnor U888 (N_888,In_527,In_328);
and U889 (N_889,In_448,In_40);
and U890 (N_890,In_588,In_302);
or U891 (N_891,In_222,In_450);
nor U892 (N_892,In_536,In_291);
or U893 (N_893,In_405,In_234);
nor U894 (N_894,In_480,In_360);
xor U895 (N_895,In_275,In_698);
nand U896 (N_896,In_84,In_377);
nand U897 (N_897,In_307,In_72);
xor U898 (N_898,In_328,In_155);
or U899 (N_899,In_138,In_172);
xor U900 (N_900,In_705,In_153);
nand U901 (N_901,In_351,In_50);
nor U902 (N_902,In_48,In_153);
or U903 (N_903,In_703,In_154);
or U904 (N_904,In_199,In_593);
xnor U905 (N_905,In_318,In_268);
nor U906 (N_906,In_236,In_118);
nand U907 (N_907,In_591,In_566);
xor U908 (N_908,In_442,In_433);
or U909 (N_909,In_495,In_675);
or U910 (N_910,In_130,In_691);
or U911 (N_911,In_274,In_100);
and U912 (N_912,In_614,In_701);
xnor U913 (N_913,In_608,In_266);
and U914 (N_914,In_627,In_483);
or U915 (N_915,In_165,In_695);
or U916 (N_916,In_50,In_331);
and U917 (N_917,In_573,In_264);
nand U918 (N_918,In_494,In_133);
xnor U919 (N_919,In_521,In_99);
nor U920 (N_920,In_179,In_113);
nor U921 (N_921,In_337,In_154);
and U922 (N_922,In_607,In_52);
and U923 (N_923,In_711,In_69);
xor U924 (N_924,In_535,In_176);
or U925 (N_925,In_111,In_364);
or U926 (N_926,In_257,In_116);
or U927 (N_927,In_710,In_168);
and U928 (N_928,In_132,In_554);
nand U929 (N_929,In_466,In_203);
or U930 (N_930,In_357,In_104);
and U931 (N_931,In_286,In_622);
and U932 (N_932,In_511,In_588);
and U933 (N_933,In_528,In_524);
or U934 (N_934,In_615,In_223);
xor U935 (N_935,In_57,In_544);
nand U936 (N_936,In_7,In_671);
nand U937 (N_937,In_632,In_243);
nand U938 (N_938,In_346,In_627);
nor U939 (N_939,In_121,In_663);
nor U940 (N_940,In_365,In_504);
nor U941 (N_941,In_732,In_652);
nand U942 (N_942,In_441,In_5);
and U943 (N_943,In_740,In_233);
nor U944 (N_944,In_266,In_663);
nor U945 (N_945,In_298,In_521);
nor U946 (N_946,In_445,In_44);
or U947 (N_947,In_360,In_12);
nand U948 (N_948,In_2,In_708);
nor U949 (N_949,In_739,In_199);
nand U950 (N_950,In_286,In_441);
xnor U951 (N_951,In_297,In_344);
nor U952 (N_952,In_477,In_386);
or U953 (N_953,In_321,In_61);
xor U954 (N_954,In_633,In_162);
nand U955 (N_955,In_303,In_575);
nor U956 (N_956,In_478,In_366);
xnor U957 (N_957,In_371,In_646);
and U958 (N_958,In_38,In_83);
nor U959 (N_959,In_174,In_398);
nor U960 (N_960,In_340,In_431);
and U961 (N_961,In_61,In_365);
or U962 (N_962,In_415,In_372);
xnor U963 (N_963,In_58,In_421);
xnor U964 (N_964,In_188,In_249);
xnor U965 (N_965,In_16,In_455);
and U966 (N_966,In_341,In_686);
and U967 (N_967,In_418,In_471);
and U968 (N_968,In_686,In_563);
and U969 (N_969,In_715,In_1);
and U970 (N_970,In_564,In_666);
and U971 (N_971,In_477,In_744);
xnor U972 (N_972,In_720,In_381);
and U973 (N_973,In_218,In_677);
nor U974 (N_974,In_541,In_241);
nand U975 (N_975,In_417,In_123);
or U976 (N_976,In_187,In_742);
or U977 (N_977,In_292,In_707);
and U978 (N_978,In_317,In_285);
or U979 (N_979,In_544,In_708);
and U980 (N_980,In_434,In_486);
and U981 (N_981,In_77,In_159);
or U982 (N_982,In_651,In_371);
nand U983 (N_983,In_643,In_75);
or U984 (N_984,In_699,In_517);
or U985 (N_985,In_355,In_739);
nor U986 (N_986,In_355,In_240);
xor U987 (N_987,In_170,In_503);
nor U988 (N_988,In_402,In_340);
or U989 (N_989,In_331,In_617);
nand U990 (N_990,In_440,In_326);
xor U991 (N_991,In_580,In_601);
or U992 (N_992,In_121,In_100);
and U993 (N_993,In_352,In_302);
xnor U994 (N_994,In_159,In_120);
nand U995 (N_995,In_204,In_593);
nor U996 (N_996,In_87,In_327);
nor U997 (N_997,In_263,In_372);
and U998 (N_998,In_50,In_722);
nor U999 (N_999,In_460,In_561);
and U1000 (N_1000,In_543,In_172);
nand U1001 (N_1001,In_643,In_346);
nand U1002 (N_1002,In_736,In_742);
xor U1003 (N_1003,In_552,In_555);
nor U1004 (N_1004,In_307,In_195);
xor U1005 (N_1005,In_504,In_711);
xnor U1006 (N_1006,In_296,In_679);
nor U1007 (N_1007,In_393,In_131);
or U1008 (N_1008,In_573,In_666);
and U1009 (N_1009,In_652,In_373);
or U1010 (N_1010,In_33,In_333);
and U1011 (N_1011,In_562,In_65);
xnor U1012 (N_1012,In_232,In_211);
nor U1013 (N_1013,In_472,In_603);
or U1014 (N_1014,In_447,In_535);
or U1015 (N_1015,In_619,In_238);
nor U1016 (N_1016,In_356,In_567);
xnor U1017 (N_1017,In_356,In_294);
nor U1018 (N_1018,In_672,In_684);
or U1019 (N_1019,In_354,In_500);
nor U1020 (N_1020,In_166,In_291);
nor U1021 (N_1021,In_267,In_193);
nand U1022 (N_1022,In_714,In_594);
nor U1023 (N_1023,In_404,In_678);
nor U1024 (N_1024,In_296,In_509);
nor U1025 (N_1025,In_168,In_338);
and U1026 (N_1026,In_583,In_651);
and U1027 (N_1027,In_302,In_339);
nand U1028 (N_1028,In_700,In_568);
nand U1029 (N_1029,In_669,In_661);
and U1030 (N_1030,In_746,In_487);
or U1031 (N_1031,In_320,In_130);
or U1032 (N_1032,In_563,In_645);
nand U1033 (N_1033,In_570,In_417);
or U1034 (N_1034,In_283,In_696);
nor U1035 (N_1035,In_297,In_71);
nor U1036 (N_1036,In_733,In_676);
nor U1037 (N_1037,In_125,In_200);
or U1038 (N_1038,In_35,In_254);
nor U1039 (N_1039,In_634,In_48);
nand U1040 (N_1040,In_34,In_74);
or U1041 (N_1041,In_612,In_37);
or U1042 (N_1042,In_566,In_408);
nand U1043 (N_1043,In_565,In_305);
nand U1044 (N_1044,In_258,In_223);
or U1045 (N_1045,In_416,In_620);
and U1046 (N_1046,In_422,In_448);
nor U1047 (N_1047,In_145,In_452);
nand U1048 (N_1048,In_252,In_468);
or U1049 (N_1049,In_359,In_209);
nand U1050 (N_1050,In_341,In_581);
nor U1051 (N_1051,In_616,In_727);
nor U1052 (N_1052,In_240,In_663);
nand U1053 (N_1053,In_362,In_346);
nand U1054 (N_1054,In_454,In_658);
and U1055 (N_1055,In_642,In_497);
nand U1056 (N_1056,In_80,In_564);
and U1057 (N_1057,In_693,In_144);
xnor U1058 (N_1058,In_580,In_662);
xor U1059 (N_1059,In_512,In_148);
nor U1060 (N_1060,In_402,In_309);
and U1061 (N_1061,In_413,In_463);
nand U1062 (N_1062,In_427,In_511);
nand U1063 (N_1063,In_207,In_50);
xnor U1064 (N_1064,In_99,In_183);
xor U1065 (N_1065,In_729,In_436);
nand U1066 (N_1066,In_611,In_416);
nor U1067 (N_1067,In_39,In_685);
or U1068 (N_1068,In_202,In_529);
xor U1069 (N_1069,In_721,In_697);
or U1070 (N_1070,In_106,In_688);
nand U1071 (N_1071,In_203,In_553);
nor U1072 (N_1072,In_484,In_276);
or U1073 (N_1073,In_454,In_279);
nand U1074 (N_1074,In_34,In_204);
or U1075 (N_1075,In_746,In_422);
nor U1076 (N_1076,In_6,In_664);
nor U1077 (N_1077,In_404,In_358);
nor U1078 (N_1078,In_115,In_47);
and U1079 (N_1079,In_76,In_137);
nor U1080 (N_1080,In_550,In_501);
nand U1081 (N_1081,In_275,In_441);
or U1082 (N_1082,In_696,In_573);
or U1083 (N_1083,In_449,In_659);
or U1084 (N_1084,In_616,In_94);
nor U1085 (N_1085,In_608,In_294);
nor U1086 (N_1086,In_673,In_77);
xor U1087 (N_1087,In_187,In_719);
or U1088 (N_1088,In_433,In_497);
nand U1089 (N_1089,In_635,In_710);
and U1090 (N_1090,In_234,In_748);
nand U1091 (N_1091,In_245,In_122);
nor U1092 (N_1092,In_671,In_594);
and U1093 (N_1093,In_645,In_203);
xor U1094 (N_1094,In_349,In_270);
or U1095 (N_1095,In_191,In_239);
and U1096 (N_1096,In_239,In_665);
nor U1097 (N_1097,In_105,In_378);
nor U1098 (N_1098,In_120,In_487);
nor U1099 (N_1099,In_375,In_543);
nor U1100 (N_1100,In_160,In_565);
xnor U1101 (N_1101,In_93,In_398);
nor U1102 (N_1102,In_198,In_562);
and U1103 (N_1103,In_173,In_198);
nor U1104 (N_1104,In_448,In_278);
nand U1105 (N_1105,In_378,In_361);
and U1106 (N_1106,In_239,In_506);
nand U1107 (N_1107,In_298,In_738);
nand U1108 (N_1108,In_88,In_87);
nand U1109 (N_1109,In_634,In_607);
nor U1110 (N_1110,In_388,In_412);
nand U1111 (N_1111,In_208,In_237);
or U1112 (N_1112,In_522,In_413);
xor U1113 (N_1113,In_83,In_656);
xnor U1114 (N_1114,In_633,In_581);
nand U1115 (N_1115,In_245,In_707);
or U1116 (N_1116,In_622,In_364);
nand U1117 (N_1117,In_83,In_563);
nand U1118 (N_1118,In_481,In_717);
or U1119 (N_1119,In_715,In_491);
xor U1120 (N_1120,In_495,In_218);
xnor U1121 (N_1121,In_696,In_519);
nor U1122 (N_1122,In_203,In_141);
nand U1123 (N_1123,In_326,In_745);
xnor U1124 (N_1124,In_705,In_223);
and U1125 (N_1125,In_355,In_314);
xor U1126 (N_1126,In_414,In_177);
or U1127 (N_1127,In_318,In_139);
nand U1128 (N_1128,In_125,In_639);
nand U1129 (N_1129,In_454,In_719);
nand U1130 (N_1130,In_423,In_5);
nor U1131 (N_1131,In_342,In_684);
and U1132 (N_1132,In_535,In_85);
or U1133 (N_1133,In_556,In_497);
and U1134 (N_1134,In_470,In_214);
or U1135 (N_1135,In_200,In_256);
and U1136 (N_1136,In_547,In_506);
or U1137 (N_1137,In_217,In_428);
nand U1138 (N_1138,In_264,In_101);
and U1139 (N_1139,In_699,In_573);
nand U1140 (N_1140,In_496,In_369);
nor U1141 (N_1141,In_664,In_133);
nor U1142 (N_1142,In_342,In_42);
nor U1143 (N_1143,In_451,In_739);
and U1144 (N_1144,In_78,In_559);
or U1145 (N_1145,In_461,In_421);
nor U1146 (N_1146,In_454,In_199);
and U1147 (N_1147,In_111,In_224);
and U1148 (N_1148,In_695,In_534);
and U1149 (N_1149,In_293,In_178);
or U1150 (N_1150,In_81,In_505);
and U1151 (N_1151,In_394,In_138);
nand U1152 (N_1152,In_679,In_259);
nor U1153 (N_1153,In_272,In_633);
xnor U1154 (N_1154,In_491,In_25);
xnor U1155 (N_1155,In_568,In_492);
and U1156 (N_1156,In_242,In_555);
or U1157 (N_1157,In_475,In_419);
nand U1158 (N_1158,In_248,In_67);
xnor U1159 (N_1159,In_498,In_632);
nand U1160 (N_1160,In_609,In_273);
xor U1161 (N_1161,In_131,In_364);
or U1162 (N_1162,In_101,In_273);
xor U1163 (N_1163,In_333,In_104);
or U1164 (N_1164,In_278,In_69);
or U1165 (N_1165,In_537,In_385);
or U1166 (N_1166,In_590,In_347);
and U1167 (N_1167,In_86,In_402);
nand U1168 (N_1168,In_699,In_300);
nand U1169 (N_1169,In_319,In_348);
nor U1170 (N_1170,In_514,In_489);
nor U1171 (N_1171,In_640,In_446);
and U1172 (N_1172,In_172,In_334);
nor U1173 (N_1173,In_669,In_181);
or U1174 (N_1174,In_245,In_119);
nand U1175 (N_1175,In_500,In_491);
nand U1176 (N_1176,In_634,In_407);
or U1177 (N_1177,In_460,In_114);
and U1178 (N_1178,In_326,In_231);
or U1179 (N_1179,In_747,In_412);
or U1180 (N_1180,In_89,In_189);
nand U1181 (N_1181,In_25,In_289);
nor U1182 (N_1182,In_299,In_633);
or U1183 (N_1183,In_61,In_665);
or U1184 (N_1184,In_136,In_452);
nor U1185 (N_1185,In_298,In_73);
or U1186 (N_1186,In_191,In_9);
and U1187 (N_1187,In_214,In_51);
nor U1188 (N_1188,In_240,In_377);
or U1189 (N_1189,In_657,In_428);
or U1190 (N_1190,In_252,In_552);
xnor U1191 (N_1191,In_37,In_564);
nand U1192 (N_1192,In_625,In_544);
or U1193 (N_1193,In_647,In_266);
nor U1194 (N_1194,In_484,In_724);
and U1195 (N_1195,In_26,In_280);
nor U1196 (N_1196,In_624,In_102);
nand U1197 (N_1197,In_392,In_82);
and U1198 (N_1198,In_304,In_228);
nand U1199 (N_1199,In_587,In_49);
or U1200 (N_1200,In_406,In_537);
nor U1201 (N_1201,In_677,In_326);
xnor U1202 (N_1202,In_637,In_258);
nor U1203 (N_1203,In_720,In_222);
nor U1204 (N_1204,In_123,In_573);
or U1205 (N_1205,In_720,In_10);
xor U1206 (N_1206,In_519,In_569);
xor U1207 (N_1207,In_263,In_314);
and U1208 (N_1208,In_601,In_25);
nor U1209 (N_1209,In_352,In_209);
nor U1210 (N_1210,In_429,In_690);
and U1211 (N_1211,In_103,In_301);
and U1212 (N_1212,In_535,In_582);
or U1213 (N_1213,In_119,In_181);
nor U1214 (N_1214,In_41,In_451);
and U1215 (N_1215,In_77,In_55);
and U1216 (N_1216,In_352,In_518);
nor U1217 (N_1217,In_330,In_745);
nor U1218 (N_1218,In_655,In_54);
nand U1219 (N_1219,In_270,In_577);
or U1220 (N_1220,In_390,In_53);
xor U1221 (N_1221,In_628,In_234);
nor U1222 (N_1222,In_533,In_77);
nor U1223 (N_1223,In_611,In_733);
and U1224 (N_1224,In_518,In_331);
nor U1225 (N_1225,In_23,In_300);
nand U1226 (N_1226,In_646,In_470);
or U1227 (N_1227,In_443,In_400);
nor U1228 (N_1228,In_557,In_323);
nor U1229 (N_1229,In_479,In_747);
nor U1230 (N_1230,In_470,In_412);
or U1231 (N_1231,In_466,In_268);
nor U1232 (N_1232,In_227,In_569);
nand U1233 (N_1233,In_132,In_599);
or U1234 (N_1234,In_59,In_190);
nor U1235 (N_1235,In_227,In_697);
nor U1236 (N_1236,In_229,In_531);
and U1237 (N_1237,In_132,In_592);
and U1238 (N_1238,In_261,In_737);
or U1239 (N_1239,In_84,In_591);
nor U1240 (N_1240,In_505,In_348);
and U1241 (N_1241,In_302,In_581);
nand U1242 (N_1242,In_190,In_647);
nor U1243 (N_1243,In_419,In_705);
or U1244 (N_1244,In_532,In_678);
nand U1245 (N_1245,In_333,In_410);
nand U1246 (N_1246,In_41,In_701);
nand U1247 (N_1247,In_706,In_682);
and U1248 (N_1248,In_703,In_363);
xnor U1249 (N_1249,In_156,In_182);
and U1250 (N_1250,In_290,In_535);
or U1251 (N_1251,In_287,In_144);
and U1252 (N_1252,In_503,In_654);
nand U1253 (N_1253,In_414,In_85);
nand U1254 (N_1254,In_26,In_152);
nor U1255 (N_1255,In_17,In_167);
and U1256 (N_1256,In_657,In_565);
nand U1257 (N_1257,In_207,In_641);
nor U1258 (N_1258,In_3,In_258);
or U1259 (N_1259,In_450,In_624);
nand U1260 (N_1260,In_637,In_109);
nor U1261 (N_1261,In_687,In_748);
or U1262 (N_1262,In_169,In_697);
xnor U1263 (N_1263,In_250,In_728);
nor U1264 (N_1264,In_554,In_63);
nand U1265 (N_1265,In_337,In_357);
and U1266 (N_1266,In_389,In_23);
or U1267 (N_1267,In_537,In_456);
nand U1268 (N_1268,In_513,In_276);
nand U1269 (N_1269,In_322,In_555);
nand U1270 (N_1270,In_62,In_453);
and U1271 (N_1271,In_249,In_186);
nand U1272 (N_1272,In_366,In_139);
and U1273 (N_1273,In_728,In_26);
xnor U1274 (N_1274,In_361,In_393);
nor U1275 (N_1275,In_391,In_372);
and U1276 (N_1276,In_594,In_461);
nor U1277 (N_1277,In_442,In_109);
nand U1278 (N_1278,In_338,In_110);
nor U1279 (N_1279,In_494,In_205);
and U1280 (N_1280,In_606,In_276);
and U1281 (N_1281,In_701,In_106);
nor U1282 (N_1282,In_36,In_695);
xnor U1283 (N_1283,In_361,In_575);
and U1284 (N_1284,In_82,In_350);
and U1285 (N_1285,In_179,In_718);
nor U1286 (N_1286,In_743,In_37);
or U1287 (N_1287,In_498,In_612);
and U1288 (N_1288,In_257,In_49);
or U1289 (N_1289,In_521,In_281);
and U1290 (N_1290,In_707,In_497);
nand U1291 (N_1291,In_707,In_606);
nor U1292 (N_1292,In_725,In_508);
nor U1293 (N_1293,In_134,In_611);
nand U1294 (N_1294,In_412,In_440);
nor U1295 (N_1295,In_674,In_303);
nor U1296 (N_1296,In_401,In_383);
and U1297 (N_1297,In_311,In_418);
nand U1298 (N_1298,In_467,In_422);
nor U1299 (N_1299,In_12,In_125);
and U1300 (N_1300,In_177,In_604);
or U1301 (N_1301,In_632,In_589);
and U1302 (N_1302,In_680,In_204);
nor U1303 (N_1303,In_125,In_505);
and U1304 (N_1304,In_268,In_300);
and U1305 (N_1305,In_109,In_365);
or U1306 (N_1306,In_270,In_470);
or U1307 (N_1307,In_262,In_651);
and U1308 (N_1308,In_198,In_657);
or U1309 (N_1309,In_665,In_230);
nor U1310 (N_1310,In_495,In_713);
xnor U1311 (N_1311,In_149,In_292);
and U1312 (N_1312,In_643,In_84);
or U1313 (N_1313,In_670,In_114);
or U1314 (N_1314,In_274,In_539);
xor U1315 (N_1315,In_327,In_449);
and U1316 (N_1316,In_555,In_696);
nor U1317 (N_1317,In_187,In_307);
nand U1318 (N_1318,In_154,In_400);
nor U1319 (N_1319,In_284,In_635);
nor U1320 (N_1320,In_505,In_372);
and U1321 (N_1321,In_548,In_294);
nor U1322 (N_1322,In_511,In_666);
nor U1323 (N_1323,In_518,In_639);
nor U1324 (N_1324,In_710,In_19);
and U1325 (N_1325,In_492,In_664);
nand U1326 (N_1326,In_386,In_535);
and U1327 (N_1327,In_270,In_110);
xnor U1328 (N_1328,In_443,In_531);
nor U1329 (N_1329,In_150,In_443);
nor U1330 (N_1330,In_593,In_694);
or U1331 (N_1331,In_260,In_232);
and U1332 (N_1332,In_279,In_619);
nand U1333 (N_1333,In_224,In_628);
or U1334 (N_1334,In_639,In_80);
or U1335 (N_1335,In_392,In_132);
or U1336 (N_1336,In_693,In_514);
or U1337 (N_1337,In_683,In_679);
or U1338 (N_1338,In_734,In_102);
xnor U1339 (N_1339,In_22,In_175);
xor U1340 (N_1340,In_568,In_36);
nor U1341 (N_1341,In_251,In_586);
nor U1342 (N_1342,In_83,In_651);
and U1343 (N_1343,In_455,In_120);
or U1344 (N_1344,In_103,In_251);
or U1345 (N_1345,In_633,In_374);
nor U1346 (N_1346,In_131,In_534);
and U1347 (N_1347,In_19,In_279);
xor U1348 (N_1348,In_321,In_686);
nand U1349 (N_1349,In_709,In_221);
nor U1350 (N_1350,In_92,In_207);
or U1351 (N_1351,In_497,In_438);
and U1352 (N_1352,In_25,In_705);
nor U1353 (N_1353,In_580,In_150);
nor U1354 (N_1354,In_315,In_291);
or U1355 (N_1355,In_567,In_744);
and U1356 (N_1356,In_268,In_562);
or U1357 (N_1357,In_508,In_260);
nor U1358 (N_1358,In_497,In_181);
nor U1359 (N_1359,In_39,In_726);
nand U1360 (N_1360,In_263,In_411);
and U1361 (N_1361,In_344,In_441);
nor U1362 (N_1362,In_384,In_729);
or U1363 (N_1363,In_607,In_465);
or U1364 (N_1364,In_469,In_369);
nor U1365 (N_1365,In_624,In_65);
nor U1366 (N_1366,In_741,In_111);
nor U1367 (N_1367,In_425,In_502);
and U1368 (N_1368,In_87,In_680);
nor U1369 (N_1369,In_521,In_161);
nor U1370 (N_1370,In_258,In_188);
and U1371 (N_1371,In_167,In_37);
or U1372 (N_1372,In_484,In_726);
xor U1373 (N_1373,In_473,In_352);
or U1374 (N_1374,In_369,In_132);
nor U1375 (N_1375,In_659,In_729);
nand U1376 (N_1376,In_649,In_372);
and U1377 (N_1377,In_101,In_366);
or U1378 (N_1378,In_427,In_277);
or U1379 (N_1379,In_177,In_691);
nand U1380 (N_1380,In_9,In_406);
nand U1381 (N_1381,In_206,In_425);
and U1382 (N_1382,In_457,In_652);
nand U1383 (N_1383,In_475,In_155);
nor U1384 (N_1384,In_154,In_341);
nor U1385 (N_1385,In_642,In_10);
or U1386 (N_1386,In_541,In_747);
or U1387 (N_1387,In_424,In_130);
or U1388 (N_1388,In_24,In_254);
nand U1389 (N_1389,In_250,In_417);
nand U1390 (N_1390,In_537,In_0);
or U1391 (N_1391,In_377,In_608);
and U1392 (N_1392,In_611,In_126);
xnor U1393 (N_1393,In_192,In_661);
nor U1394 (N_1394,In_104,In_60);
or U1395 (N_1395,In_449,In_0);
and U1396 (N_1396,In_479,In_377);
and U1397 (N_1397,In_345,In_51);
and U1398 (N_1398,In_369,In_375);
nor U1399 (N_1399,In_355,In_120);
nand U1400 (N_1400,In_136,In_393);
and U1401 (N_1401,In_497,In_289);
and U1402 (N_1402,In_658,In_471);
nand U1403 (N_1403,In_701,In_303);
or U1404 (N_1404,In_660,In_747);
or U1405 (N_1405,In_600,In_80);
nand U1406 (N_1406,In_682,In_54);
xor U1407 (N_1407,In_430,In_641);
and U1408 (N_1408,In_727,In_66);
nand U1409 (N_1409,In_378,In_428);
nor U1410 (N_1410,In_204,In_685);
nand U1411 (N_1411,In_78,In_493);
and U1412 (N_1412,In_78,In_370);
nand U1413 (N_1413,In_149,In_233);
nand U1414 (N_1414,In_739,In_603);
and U1415 (N_1415,In_461,In_579);
nand U1416 (N_1416,In_230,In_454);
nand U1417 (N_1417,In_157,In_545);
xnor U1418 (N_1418,In_345,In_555);
nor U1419 (N_1419,In_284,In_424);
nor U1420 (N_1420,In_37,In_446);
and U1421 (N_1421,In_474,In_357);
nand U1422 (N_1422,In_361,In_490);
and U1423 (N_1423,In_85,In_658);
xnor U1424 (N_1424,In_161,In_151);
nor U1425 (N_1425,In_458,In_465);
nand U1426 (N_1426,In_88,In_675);
nand U1427 (N_1427,In_451,In_441);
nand U1428 (N_1428,In_584,In_510);
or U1429 (N_1429,In_127,In_569);
nand U1430 (N_1430,In_708,In_1);
nand U1431 (N_1431,In_200,In_584);
or U1432 (N_1432,In_230,In_68);
or U1433 (N_1433,In_191,In_67);
or U1434 (N_1434,In_340,In_584);
and U1435 (N_1435,In_166,In_739);
nand U1436 (N_1436,In_68,In_96);
nor U1437 (N_1437,In_131,In_22);
nor U1438 (N_1438,In_671,In_89);
nand U1439 (N_1439,In_504,In_665);
and U1440 (N_1440,In_673,In_323);
xnor U1441 (N_1441,In_154,In_171);
nor U1442 (N_1442,In_502,In_159);
and U1443 (N_1443,In_670,In_301);
and U1444 (N_1444,In_211,In_404);
or U1445 (N_1445,In_233,In_122);
or U1446 (N_1446,In_466,In_645);
and U1447 (N_1447,In_605,In_531);
and U1448 (N_1448,In_283,In_616);
and U1449 (N_1449,In_338,In_550);
nor U1450 (N_1450,In_540,In_626);
or U1451 (N_1451,In_2,In_206);
and U1452 (N_1452,In_550,In_407);
or U1453 (N_1453,In_456,In_215);
nor U1454 (N_1454,In_615,In_222);
nor U1455 (N_1455,In_100,In_160);
nand U1456 (N_1456,In_547,In_695);
or U1457 (N_1457,In_185,In_430);
nor U1458 (N_1458,In_264,In_355);
and U1459 (N_1459,In_650,In_579);
nor U1460 (N_1460,In_60,In_335);
and U1461 (N_1461,In_312,In_106);
nand U1462 (N_1462,In_547,In_535);
nor U1463 (N_1463,In_627,In_568);
and U1464 (N_1464,In_88,In_100);
xor U1465 (N_1465,In_521,In_383);
nor U1466 (N_1466,In_329,In_706);
and U1467 (N_1467,In_501,In_96);
and U1468 (N_1468,In_662,In_313);
and U1469 (N_1469,In_620,In_717);
nand U1470 (N_1470,In_526,In_375);
and U1471 (N_1471,In_52,In_158);
nand U1472 (N_1472,In_381,In_18);
xor U1473 (N_1473,In_712,In_341);
xor U1474 (N_1474,In_723,In_238);
and U1475 (N_1475,In_591,In_74);
or U1476 (N_1476,In_457,In_717);
nand U1477 (N_1477,In_496,In_121);
nor U1478 (N_1478,In_286,In_156);
or U1479 (N_1479,In_523,In_339);
and U1480 (N_1480,In_324,In_424);
and U1481 (N_1481,In_73,In_679);
xor U1482 (N_1482,In_640,In_140);
nor U1483 (N_1483,In_118,In_206);
and U1484 (N_1484,In_165,In_315);
or U1485 (N_1485,In_439,In_318);
nor U1486 (N_1486,In_559,In_238);
or U1487 (N_1487,In_503,In_443);
and U1488 (N_1488,In_12,In_483);
nor U1489 (N_1489,In_331,In_285);
nor U1490 (N_1490,In_314,In_215);
or U1491 (N_1491,In_682,In_258);
and U1492 (N_1492,In_270,In_219);
or U1493 (N_1493,In_581,In_33);
nand U1494 (N_1494,In_241,In_390);
nor U1495 (N_1495,In_82,In_267);
nand U1496 (N_1496,In_691,In_140);
nor U1497 (N_1497,In_723,In_545);
or U1498 (N_1498,In_333,In_356);
nor U1499 (N_1499,In_510,In_283);
nand U1500 (N_1500,In_543,In_713);
nand U1501 (N_1501,In_258,In_209);
xor U1502 (N_1502,In_175,In_609);
nand U1503 (N_1503,In_120,In_739);
and U1504 (N_1504,In_372,In_200);
xnor U1505 (N_1505,In_157,In_154);
xnor U1506 (N_1506,In_256,In_249);
nand U1507 (N_1507,In_473,In_336);
xor U1508 (N_1508,In_329,In_14);
and U1509 (N_1509,In_478,In_479);
nor U1510 (N_1510,In_575,In_153);
nor U1511 (N_1511,In_451,In_720);
xnor U1512 (N_1512,In_721,In_631);
nand U1513 (N_1513,In_710,In_234);
or U1514 (N_1514,In_710,In_86);
or U1515 (N_1515,In_131,In_745);
nor U1516 (N_1516,In_245,In_312);
or U1517 (N_1517,In_294,In_725);
nand U1518 (N_1518,In_75,In_333);
xor U1519 (N_1519,In_0,In_198);
or U1520 (N_1520,In_593,In_25);
nor U1521 (N_1521,In_386,In_62);
nand U1522 (N_1522,In_628,In_124);
nor U1523 (N_1523,In_73,In_402);
or U1524 (N_1524,In_378,In_107);
nand U1525 (N_1525,In_723,In_302);
nor U1526 (N_1526,In_459,In_44);
xnor U1527 (N_1527,In_347,In_7);
nor U1528 (N_1528,In_38,In_465);
nand U1529 (N_1529,In_581,In_624);
or U1530 (N_1530,In_666,In_143);
or U1531 (N_1531,In_698,In_341);
xor U1532 (N_1532,In_11,In_306);
nand U1533 (N_1533,In_242,In_738);
or U1534 (N_1534,In_116,In_371);
nand U1535 (N_1535,In_180,In_460);
nor U1536 (N_1536,In_77,In_214);
nor U1537 (N_1537,In_343,In_428);
xnor U1538 (N_1538,In_714,In_119);
nor U1539 (N_1539,In_611,In_227);
or U1540 (N_1540,In_699,In_260);
or U1541 (N_1541,In_45,In_26);
or U1542 (N_1542,In_527,In_495);
or U1543 (N_1543,In_11,In_399);
or U1544 (N_1544,In_105,In_399);
nor U1545 (N_1545,In_115,In_177);
and U1546 (N_1546,In_63,In_576);
or U1547 (N_1547,In_341,In_565);
xor U1548 (N_1548,In_648,In_586);
nor U1549 (N_1549,In_10,In_82);
xor U1550 (N_1550,In_50,In_490);
nor U1551 (N_1551,In_222,In_66);
xnor U1552 (N_1552,In_218,In_137);
nand U1553 (N_1553,In_570,In_335);
nor U1554 (N_1554,In_499,In_476);
nand U1555 (N_1555,In_188,In_453);
nand U1556 (N_1556,In_361,In_136);
and U1557 (N_1557,In_343,In_403);
and U1558 (N_1558,In_210,In_383);
nand U1559 (N_1559,In_54,In_37);
and U1560 (N_1560,In_224,In_689);
nor U1561 (N_1561,In_426,In_327);
nor U1562 (N_1562,In_383,In_506);
and U1563 (N_1563,In_30,In_117);
and U1564 (N_1564,In_315,In_138);
xor U1565 (N_1565,In_77,In_395);
nand U1566 (N_1566,In_320,In_55);
and U1567 (N_1567,In_507,In_313);
nor U1568 (N_1568,In_645,In_15);
and U1569 (N_1569,In_481,In_623);
or U1570 (N_1570,In_38,In_43);
nor U1571 (N_1571,In_186,In_564);
or U1572 (N_1572,In_20,In_537);
xnor U1573 (N_1573,In_136,In_424);
nor U1574 (N_1574,In_312,In_272);
nand U1575 (N_1575,In_10,In_701);
or U1576 (N_1576,In_687,In_49);
nor U1577 (N_1577,In_70,In_18);
nand U1578 (N_1578,In_164,In_440);
xor U1579 (N_1579,In_103,In_215);
nor U1580 (N_1580,In_5,In_230);
nand U1581 (N_1581,In_156,In_361);
and U1582 (N_1582,In_412,In_720);
nand U1583 (N_1583,In_41,In_264);
or U1584 (N_1584,In_242,In_37);
or U1585 (N_1585,In_198,In_161);
nand U1586 (N_1586,In_170,In_232);
and U1587 (N_1587,In_692,In_399);
nand U1588 (N_1588,In_560,In_535);
nand U1589 (N_1589,In_736,In_704);
nand U1590 (N_1590,In_538,In_457);
and U1591 (N_1591,In_743,In_2);
or U1592 (N_1592,In_241,In_712);
nor U1593 (N_1593,In_169,In_603);
nand U1594 (N_1594,In_309,In_626);
nand U1595 (N_1595,In_274,In_330);
nand U1596 (N_1596,In_523,In_684);
nand U1597 (N_1597,In_468,In_385);
nor U1598 (N_1598,In_699,In_188);
nand U1599 (N_1599,In_473,In_581);
nand U1600 (N_1600,In_133,In_367);
and U1601 (N_1601,In_737,In_582);
or U1602 (N_1602,In_315,In_26);
and U1603 (N_1603,In_489,In_194);
nor U1604 (N_1604,In_312,In_270);
nor U1605 (N_1605,In_293,In_747);
and U1606 (N_1606,In_308,In_336);
and U1607 (N_1607,In_174,In_311);
nor U1608 (N_1608,In_348,In_740);
or U1609 (N_1609,In_418,In_394);
nand U1610 (N_1610,In_619,In_110);
nor U1611 (N_1611,In_722,In_377);
or U1612 (N_1612,In_575,In_120);
and U1613 (N_1613,In_548,In_429);
nand U1614 (N_1614,In_693,In_302);
or U1615 (N_1615,In_665,In_212);
and U1616 (N_1616,In_281,In_31);
nand U1617 (N_1617,In_286,In_300);
or U1618 (N_1618,In_697,In_516);
or U1619 (N_1619,In_166,In_445);
or U1620 (N_1620,In_270,In_23);
nand U1621 (N_1621,In_79,In_550);
nor U1622 (N_1622,In_593,In_376);
nand U1623 (N_1623,In_377,In_638);
or U1624 (N_1624,In_405,In_286);
and U1625 (N_1625,In_617,In_248);
or U1626 (N_1626,In_133,In_583);
and U1627 (N_1627,In_540,In_247);
nor U1628 (N_1628,In_136,In_627);
nand U1629 (N_1629,In_743,In_77);
and U1630 (N_1630,In_683,In_20);
or U1631 (N_1631,In_479,In_740);
nor U1632 (N_1632,In_596,In_331);
nor U1633 (N_1633,In_288,In_282);
nor U1634 (N_1634,In_737,In_419);
and U1635 (N_1635,In_278,In_48);
nor U1636 (N_1636,In_54,In_358);
or U1637 (N_1637,In_141,In_453);
and U1638 (N_1638,In_622,In_669);
or U1639 (N_1639,In_43,In_152);
nor U1640 (N_1640,In_189,In_123);
nand U1641 (N_1641,In_278,In_553);
or U1642 (N_1642,In_246,In_453);
xnor U1643 (N_1643,In_248,In_491);
or U1644 (N_1644,In_347,In_171);
nor U1645 (N_1645,In_162,In_26);
xnor U1646 (N_1646,In_725,In_256);
or U1647 (N_1647,In_716,In_286);
and U1648 (N_1648,In_674,In_565);
or U1649 (N_1649,In_697,In_389);
or U1650 (N_1650,In_687,In_394);
xor U1651 (N_1651,In_126,In_387);
or U1652 (N_1652,In_277,In_194);
or U1653 (N_1653,In_440,In_434);
or U1654 (N_1654,In_399,In_158);
or U1655 (N_1655,In_178,In_207);
xnor U1656 (N_1656,In_442,In_210);
and U1657 (N_1657,In_235,In_723);
nand U1658 (N_1658,In_621,In_183);
and U1659 (N_1659,In_31,In_344);
or U1660 (N_1660,In_740,In_136);
or U1661 (N_1661,In_600,In_2);
and U1662 (N_1662,In_108,In_460);
and U1663 (N_1663,In_597,In_120);
nor U1664 (N_1664,In_347,In_238);
and U1665 (N_1665,In_604,In_690);
or U1666 (N_1666,In_646,In_542);
nand U1667 (N_1667,In_666,In_434);
nor U1668 (N_1668,In_322,In_136);
and U1669 (N_1669,In_415,In_49);
and U1670 (N_1670,In_94,In_109);
and U1671 (N_1671,In_63,In_573);
nor U1672 (N_1672,In_212,In_563);
nand U1673 (N_1673,In_158,In_745);
xnor U1674 (N_1674,In_127,In_420);
nor U1675 (N_1675,In_309,In_614);
and U1676 (N_1676,In_526,In_463);
and U1677 (N_1677,In_89,In_249);
nor U1678 (N_1678,In_490,In_28);
and U1679 (N_1679,In_211,In_466);
or U1680 (N_1680,In_57,In_29);
and U1681 (N_1681,In_97,In_192);
and U1682 (N_1682,In_504,In_105);
and U1683 (N_1683,In_39,In_180);
and U1684 (N_1684,In_569,In_128);
and U1685 (N_1685,In_195,In_182);
or U1686 (N_1686,In_189,In_618);
or U1687 (N_1687,In_400,In_641);
and U1688 (N_1688,In_16,In_183);
and U1689 (N_1689,In_357,In_0);
nand U1690 (N_1690,In_519,In_499);
xnor U1691 (N_1691,In_519,In_303);
and U1692 (N_1692,In_682,In_416);
and U1693 (N_1693,In_503,In_125);
or U1694 (N_1694,In_408,In_429);
nand U1695 (N_1695,In_649,In_316);
and U1696 (N_1696,In_38,In_569);
or U1697 (N_1697,In_388,In_480);
nor U1698 (N_1698,In_20,In_362);
or U1699 (N_1699,In_20,In_714);
or U1700 (N_1700,In_59,In_590);
or U1701 (N_1701,In_506,In_185);
and U1702 (N_1702,In_191,In_363);
nand U1703 (N_1703,In_466,In_258);
or U1704 (N_1704,In_344,In_549);
and U1705 (N_1705,In_176,In_700);
and U1706 (N_1706,In_1,In_187);
nor U1707 (N_1707,In_688,In_555);
xor U1708 (N_1708,In_567,In_368);
nand U1709 (N_1709,In_94,In_216);
or U1710 (N_1710,In_391,In_52);
xor U1711 (N_1711,In_731,In_59);
nor U1712 (N_1712,In_483,In_194);
and U1713 (N_1713,In_650,In_293);
and U1714 (N_1714,In_604,In_663);
nor U1715 (N_1715,In_687,In_611);
and U1716 (N_1716,In_279,In_371);
nor U1717 (N_1717,In_478,In_146);
or U1718 (N_1718,In_100,In_489);
nand U1719 (N_1719,In_214,In_369);
and U1720 (N_1720,In_544,In_713);
nor U1721 (N_1721,In_557,In_618);
nor U1722 (N_1722,In_102,In_440);
and U1723 (N_1723,In_64,In_696);
xor U1724 (N_1724,In_167,In_338);
or U1725 (N_1725,In_146,In_530);
nand U1726 (N_1726,In_518,In_71);
nor U1727 (N_1727,In_472,In_307);
nand U1728 (N_1728,In_10,In_293);
nand U1729 (N_1729,In_5,In_512);
nand U1730 (N_1730,In_245,In_328);
xor U1731 (N_1731,In_700,In_495);
or U1732 (N_1732,In_553,In_199);
nor U1733 (N_1733,In_184,In_583);
and U1734 (N_1734,In_659,In_357);
nor U1735 (N_1735,In_343,In_522);
nand U1736 (N_1736,In_230,In_181);
nand U1737 (N_1737,In_12,In_249);
nand U1738 (N_1738,In_702,In_498);
xnor U1739 (N_1739,In_21,In_175);
and U1740 (N_1740,In_384,In_587);
nand U1741 (N_1741,In_229,In_200);
or U1742 (N_1742,In_41,In_75);
and U1743 (N_1743,In_163,In_571);
nand U1744 (N_1744,In_328,In_659);
and U1745 (N_1745,In_32,In_254);
nand U1746 (N_1746,In_297,In_134);
or U1747 (N_1747,In_143,In_148);
nand U1748 (N_1748,In_615,In_241);
and U1749 (N_1749,In_172,In_215);
and U1750 (N_1750,In_546,In_216);
nand U1751 (N_1751,In_90,In_265);
nor U1752 (N_1752,In_453,In_442);
and U1753 (N_1753,In_496,In_259);
nor U1754 (N_1754,In_435,In_10);
or U1755 (N_1755,In_508,In_270);
nand U1756 (N_1756,In_664,In_629);
and U1757 (N_1757,In_456,In_715);
or U1758 (N_1758,In_669,In_288);
nor U1759 (N_1759,In_126,In_669);
xor U1760 (N_1760,In_522,In_33);
or U1761 (N_1761,In_531,In_695);
nand U1762 (N_1762,In_207,In_102);
nor U1763 (N_1763,In_246,In_564);
and U1764 (N_1764,In_138,In_408);
nand U1765 (N_1765,In_29,In_675);
nand U1766 (N_1766,In_543,In_513);
xor U1767 (N_1767,In_372,In_627);
nand U1768 (N_1768,In_302,In_445);
nor U1769 (N_1769,In_744,In_544);
nor U1770 (N_1770,In_225,In_665);
and U1771 (N_1771,In_687,In_96);
or U1772 (N_1772,In_234,In_129);
or U1773 (N_1773,In_173,In_515);
or U1774 (N_1774,In_556,In_77);
xnor U1775 (N_1775,In_397,In_370);
and U1776 (N_1776,In_181,In_300);
nand U1777 (N_1777,In_132,In_613);
nor U1778 (N_1778,In_700,In_630);
nand U1779 (N_1779,In_570,In_114);
nand U1780 (N_1780,In_334,In_438);
and U1781 (N_1781,In_211,In_342);
nor U1782 (N_1782,In_188,In_728);
and U1783 (N_1783,In_395,In_534);
nor U1784 (N_1784,In_650,In_364);
nand U1785 (N_1785,In_11,In_319);
nand U1786 (N_1786,In_63,In_126);
and U1787 (N_1787,In_591,In_701);
nand U1788 (N_1788,In_116,In_693);
or U1789 (N_1789,In_637,In_269);
and U1790 (N_1790,In_120,In_303);
nand U1791 (N_1791,In_113,In_155);
or U1792 (N_1792,In_489,In_678);
nand U1793 (N_1793,In_238,In_453);
or U1794 (N_1794,In_602,In_379);
and U1795 (N_1795,In_118,In_240);
and U1796 (N_1796,In_557,In_451);
or U1797 (N_1797,In_441,In_555);
or U1798 (N_1798,In_600,In_603);
nor U1799 (N_1799,In_189,In_544);
and U1800 (N_1800,In_63,In_632);
and U1801 (N_1801,In_278,In_535);
or U1802 (N_1802,In_71,In_174);
or U1803 (N_1803,In_117,In_26);
nand U1804 (N_1804,In_252,In_314);
nand U1805 (N_1805,In_217,In_243);
and U1806 (N_1806,In_20,In_293);
nor U1807 (N_1807,In_230,In_468);
nand U1808 (N_1808,In_389,In_188);
nor U1809 (N_1809,In_502,In_446);
nand U1810 (N_1810,In_36,In_648);
nor U1811 (N_1811,In_409,In_40);
and U1812 (N_1812,In_108,In_164);
or U1813 (N_1813,In_672,In_644);
nand U1814 (N_1814,In_238,In_469);
or U1815 (N_1815,In_548,In_336);
nand U1816 (N_1816,In_100,In_76);
nand U1817 (N_1817,In_673,In_356);
or U1818 (N_1818,In_588,In_310);
or U1819 (N_1819,In_287,In_293);
and U1820 (N_1820,In_187,In_732);
nand U1821 (N_1821,In_449,In_672);
and U1822 (N_1822,In_343,In_253);
or U1823 (N_1823,In_108,In_270);
or U1824 (N_1824,In_537,In_336);
or U1825 (N_1825,In_108,In_176);
nand U1826 (N_1826,In_225,In_101);
or U1827 (N_1827,In_230,In_253);
xor U1828 (N_1828,In_393,In_740);
and U1829 (N_1829,In_52,In_166);
nand U1830 (N_1830,In_322,In_612);
and U1831 (N_1831,In_230,In_334);
or U1832 (N_1832,In_419,In_232);
nor U1833 (N_1833,In_355,In_435);
and U1834 (N_1834,In_107,In_500);
nor U1835 (N_1835,In_57,In_55);
nand U1836 (N_1836,In_208,In_605);
xor U1837 (N_1837,In_129,In_140);
nor U1838 (N_1838,In_71,In_572);
xor U1839 (N_1839,In_89,In_478);
or U1840 (N_1840,In_517,In_229);
nand U1841 (N_1841,In_483,In_704);
nor U1842 (N_1842,In_41,In_483);
or U1843 (N_1843,In_559,In_18);
nor U1844 (N_1844,In_481,In_137);
nor U1845 (N_1845,In_416,In_513);
or U1846 (N_1846,In_132,In_612);
or U1847 (N_1847,In_84,In_398);
nand U1848 (N_1848,In_174,In_374);
and U1849 (N_1849,In_341,In_523);
and U1850 (N_1850,In_64,In_539);
nor U1851 (N_1851,In_363,In_525);
xnor U1852 (N_1852,In_295,In_152);
nor U1853 (N_1853,In_290,In_466);
or U1854 (N_1854,In_625,In_603);
nor U1855 (N_1855,In_413,In_340);
and U1856 (N_1856,In_331,In_139);
and U1857 (N_1857,In_339,In_402);
xnor U1858 (N_1858,In_153,In_749);
xnor U1859 (N_1859,In_196,In_4);
and U1860 (N_1860,In_250,In_245);
and U1861 (N_1861,In_600,In_267);
and U1862 (N_1862,In_40,In_653);
or U1863 (N_1863,In_180,In_712);
nand U1864 (N_1864,In_546,In_466);
nor U1865 (N_1865,In_307,In_446);
or U1866 (N_1866,In_551,In_217);
nand U1867 (N_1867,In_82,In_206);
xnor U1868 (N_1868,In_441,In_410);
xor U1869 (N_1869,In_435,In_737);
or U1870 (N_1870,In_183,In_41);
and U1871 (N_1871,In_411,In_293);
nand U1872 (N_1872,In_482,In_559);
and U1873 (N_1873,In_276,In_206);
nor U1874 (N_1874,In_305,In_317);
or U1875 (N_1875,In_520,In_489);
or U1876 (N_1876,In_679,In_232);
and U1877 (N_1877,In_412,In_709);
or U1878 (N_1878,In_310,In_264);
nand U1879 (N_1879,In_459,In_584);
nand U1880 (N_1880,In_512,In_243);
nor U1881 (N_1881,In_441,In_200);
or U1882 (N_1882,In_227,In_471);
and U1883 (N_1883,In_598,In_593);
nand U1884 (N_1884,In_360,In_140);
and U1885 (N_1885,In_527,In_184);
nand U1886 (N_1886,In_493,In_172);
nor U1887 (N_1887,In_407,In_471);
and U1888 (N_1888,In_572,In_461);
and U1889 (N_1889,In_619,In_180);
and U1890 (N_1890,In_738,In_663);
or U1891 (N_1891,In_635,In_459);
and U1892 (N_1892,In_569,In_16);
nand U1893 (N_1893,In_608,In_153);
nand U1894 (N_1894,In_5,In_255);
nand U1895 (N_1895,In_559,In_552);
or U1896 (N_1896,In_447,In_70);
and U1897 (N_1897,In_197,In_109);
or U1898 (N_1898,In_556,In_718);
nor U1899 (N_1899,In_384,In_709);
and U1900 (N_1900,In_569,In_210);
or U1901 (N_1901,In_260,In_433);
nand U1902 (N_1902,In_689,In_550);
and U1903 (N_1903,In_260,In_497);
and U1904 (N_1904,In_326,In_113);
nor U1905 (N_1905,In_438,In_100);
and U1906 (N_1906,In_24,In_289);
or U1907 (N_1907,In_502,In_654);
nor U1908 (N_1908,In_86,In_252);
nor U1909 (N_1909,In_522,In_327);
and U1910 (N_1910,In_199,In_188);
or U1911 (N_1911,In_4,In_466);
nand U1912 (N_1912,In_322,In_497);
nor U1913 (N_1913,In_692,In_259);
nor U1914 (N_1914,In_668,In_198);
nor U1915 (N_1915,In_178,In_220);
and U1916 (N_1916,In_28,In_734);
and U1917 (N_1917,In_189,In_362);
xnor U1918 (N_1918,In_578,In_65);
and U1919 (N_1919,In_309,In_247);
nor U1920 (N_1920,In_136,In_564);
nand U1921 (N_1921,In_252,In_632);
nor U1922 (N_1922,In_394,In_285);
nor U1923 (N_1923,In_618,In_445);
and U1924 (N_1924,In_399,In_242);
and U1925 (N_1925,In_202,In_645);
or U1926 (N_1926,In_2,In_519);
or U1927 (N_1927,In_35,In_309);
nor U1928 (N_1928,In_248,In_234);
or U1929 (N_1929,In_567,In_75);
and U1930 (N_1930,In_680,In_134);
nor U1931 (N_1931,In_641,In_676);
nand U1932 (N_1932,In_560,In_231);
and U1933 (N_1933,In_200,In_501);
and U1934 (N_1934,In_674,In_688);
nor U1935 (N_1935,In_456,In_220);
nand U1936 (N_1936,In_90,In_412);
nor U1937 (N_1937,In_550,In_264);
nand U1938 (N_1938,In_204,In_247);
or U1939 (N_1939,In_91,In_38);
nor U1940 (N_1940,In_380,In_165);
nand U1941 (N_1941,In_134,In_48);
xor U1942 (N_1942,In_94,In_466);
nand U1943 (N_1943,In_711,In_425);
and U1944 (N_1944,In_195,In_553);
nor U1945 (N_1945,In_652,In_256);
and U1946 (N_1946,In_64,In_560);
nor U1947 (N_1947,In_727,In_248);
and U1948 (N_1948,In_745,In_535);
nor U1949 (N_1949,In_225,In_344);
nand U1950 (N_1950,In_583,In_589);
xor U1951 (N_1951,In_687,In_224);
nand U1952 (N_1952,In_145,In_640);
nand U1953 (N_1953,In_560,In_138);
nor U1954 (N_1954,In_541,In_211);
nand U1955 (N_1955,In_50,In_354);
nor U1956 (N_1956,In_114,In_517);
and U1957 (N_1957,In_310,In_482);
or U1958 (N_1958,In_128,In_593);
xor U1959 (N_1959,In_494,In_654);
and U1960 (N_1960,In_297,In_459);
nor U1961 (N_1961,In_118,In_351);
or U1962 (N_1962,In_239,In_243);
nand U1963 (N_1963,In_208,In_449);
or U1964 (N_1964,In_525,In_555);
xnor U1965 (N_1965,In_631,In_564);
nor U1966 (N_1966,In_87,In_406);
or U1967 (N_1967,In_706,In_73);
nand U1968 (N_1968,In_491,In_357);
xnor U1969 (N_1969,In_407,In_224);
nand U1970 (N_1970,In_153,In_555);
nor U1971 (N_1971,In_480,In_458);
nor U1972 (N_1972,In_138,In_25);
nand U1973 (N_1973,In_18,In_128);
and U1974 (N_1974,In_616,In_430);
nor U1975 (N_1975,In_452,In_361);
nand U1976 (N_1976,In_271,In_661);
nand U1977 (N_1977,In_424,In_707);
nand U1978 (N_1978,In_645,In_99);
nand U1979 (N_1979,In_348,In_534);
nand U1980 (N_1980,In_701,In_169);
and U1981 (N_1981,In_518,In_154);
and U1982 (N_1982,In_601,In_696);
nand U1983 (N_1983,In_162,In_308);
or U1984 (N_1984,In_426,In_495);
and U1985 (N_1985,In_569,In_623);
and U1986 (N_1986,In_59,In_94);
nand U1987 (N_1987,In_60,In_447);
and U1988 (N_1988,In_443,In_0);
or U1989 (N_1989,In_703,In_377);
or U1990 (N_1990,In_160,In_348);
or U1991 (N_1991,In_309,In_290);
xor U1992 (N_1992,In_116,In_160);
nor U1993 (N_1993,In_352,In_175);
and U1994 (N_1994,In_203,In_68);
nor U1995 (N_1995,In_218,In_666);
or U1996 (N_1996,In_29,In_295);
and U1997 (N_1997,In_258,In_157);
nand U1998 (N_1998,In_168,In_522);
or U1999 (N_1999,In_375,In_393);
nor U2000 (N_2000,In_241,In_609);
xnor U2001 (N_2001,In_545,In_252);
nor U2002 (N_2002,In_118,In_685);
nand U2003 (N_2003,In_455,In_450);
nor U2004 (N_2004,In_54,In_101);
nor U2005 (N_2005,In_45,In_468);
or U2006 (N_2006,In_150,In_649);
nand U2007 (N_2007,In_185,In_159);
xnor U2008 (N_2008,In_210,In_292);
nor U2009 (N_2009,In_6,In_53);
or U2010 (N_2010,In_14,In_659);
or U2011 (N_2011,In_235,In_37);
nor U2012 (N_2012,In_73,In_300);
nor U2013 (N_2013,In_499,In_6);
xnor U2014 (N_2014,In_458,In_608);
nor U2015 (N_2015,In_86,In_666);
and U2016 (N_2016,In_622,In_459);
nand U2017 (N_2017,In_678,In_437);
and U2018 (N_2018,In_438,In_142);
nor U2019 (N_2019,In_154,In_150);
nor U2020 (N_2020,In_364,In_105);
or U2021 (N_2021,In_402,In_562);
or U2022 (N_2022,In_316,In_317);
nand U2023 (N_2023,In_59,In_51);
or U2024 (N_2024,In_407,In_394);
or U2025 (N_2025,In_308,In_498);
nor U2026 (N_2026,In_669,In_745);
nand U2027 (N_2027,In_502,In_285);
and U2028 (N_2028,In_383,In_545);
nor U2029 (N_2029,In_388,In_468);
nand U2030 (N_2030,In_566,In_480);
nand U2031 (N_2031,In_417,In_476);
or U2032 (N_2032,In_176,In_157);
and U2033 (N_2033,In_406,In_220);
and U2034 (N_2034,In_366,In_567);
xnor U2035 (N_2035,In_33,In_424);
or U2036 (N_2036,In_690,In_631);
or U2037 (N_2037,In_629,In_179);
xor U2038 (N_2038,In_670,In_568);
or U2039 (N_2039,In_53,In_516);
nor U2040 (N_2040,In_76,In_577);
nand U2041 (N_2041,In_36,In_165);
nor U2042 (N_2042,In_158,In_224);
or U2043 (N_2043,In_329,In_324);
nand U2044 (N_2044,In_64,In_512);
or U2045 (N_2045,In_39,In_496);
and U2046 (N_2046,In_130,In_110);
or U2047 (N_2047,In_692,In_80);
nor U2048 (N_2048,In_57,In_174);
or U2049 (N_2049,In_470,In_555);
nor U2050 (N_2050,In_670,In_297);
or U2051 (N_2051,In_738,In_477);
or U2052 (N_2052,In_33,In_547);
nand U2053 (N_2053,In_43,In_587);
nor U2054 (N_2054,In_521,In_105);
xnor U2055 (N_2055,In_168,In_145);
nand U2056 (N_2056,In_380,In_686);
nand U2057 (N_2057,In_158,In_459);
xnor U2058 (N_2058,In_528,In_446);
xor U2059 (N_2059,In_255,In_464);
nor U2060 (N_2060,In_712,In_460);
nor U2061 (N_2061,In_302,In_49);
nand U2062 (N_2062,In_639,In_373);
xnor U2063 (N_2063,In_732,In_575);
and U2064 (N_2064,In_67,In_480);
and U2065 (N_2065,In_3,In_128);
nor U2066 (N_2066,In_404,In_33);
and U2067 (N_2067,In_10,In_415);
nor U2068 (N_2068,In_524,In_151);
xnor U2069 (N_2069,In_569,In_408);
xor U2070 (N_2070,In_563,In_677);
nor U2071 (N_2071,In_672,In_396);
or U2072 (N_2072,In_152,In_212);
nand U2073 (N_2073,In_709,In_316);
nand U2074 (N_2074,In_445,In_510);
nand U2075 (N_2075,In_398,In_489);
nand U2076 (N_2076,In_167,In_372);
and U2077 (N_2077,In_210,In_694);
nor U2078 (N_2078,In_475,In_698);
or U2079 (N_2079,In_285,In_253);
or U2080 (N_2080,In_639,In_399);
and U2081 (N_2081,In_581,In_152);
and U2082 (N_2082,In_570,In_498);
nor U2083 (N_2083,In_349,In_135);
nand U2084 (N_2084,In_407,In_183);
and U2085 (N_2085,In_152,In_84);
nor U2086 (N_2086,In_512,In_253);
xor U2087 (N_2087,In_428,In_269);
or U2088 (N_2088,In_251,In_18);
xor U2089 (N_2089,In_57,In_384);
xnor U2090 (N_2090,In_612,In_127);
xor U2091 (N_2091,In_483,In_318);
nand U2092 (N_2092,In_47,In_330);
and U2093 (N_2093,In_258,In_460);
nand U2094 (N_2094,In_558,In_240);
nor U2095 (N_2095,In_743,In_147);
and U2096 (N_2096,In_6,In_638);
nor U2097 (N_2097,In_332,In_317);
or U2098 (N_2098,In_137,In_86);
or U2099 (N_2099,In_563,In_238);
nor U2100 (N_2100,In_620,In_543);
nor U2101 (N_2101,In_106,In_172);
nand U2102 (N_2102,In_398,In_92);
or U2103 (N_2103,In_382,In_651);
xnor U2104 (N_2104,In_717,In_387);
nand U2105 (N_2105,In_44,In_418);
nor U2106 (N_2106,In_294,In_739);
xnor U2107 (N_2107,In_496,In_387);
and U2108 (N_2108,In_133,In_741);
nor U2109 (N_2109,In_57,In_737);
nand U2110 (N_2110,In_406,In_192);
and U2111 (N_2111,In_54,In_246);
or U2112 (N_2112,In_335,In_552);
nand U2113 (N_2113,In_374,In_214);
or U2114 (N_2114,In_206,In_727);
and U2115 (N_2115,In_163,In_601);
and U2116 (N_2116,In_395,In_53);
nor U2117 (N_2117,In_146,In_173);
nor U2118 (N_2118,In_88,In_529);
nor U2119 (N_2119,In_158,In_43);
nor U2120 (N_2120,In_272,In_287);
and U2121 (N_2121,In_300,In_450);
xor U2122 (N_2122,In_741,In_443);
and U2123 (N_2123,In_207,In_451);
and U2124 (N_2124,In_162,In_658);
nand U2125 (N_2125,In_740,In_738);
nor U2126 (N_2126,In_527,In_185);
nand U2127 (N_2127,In_281,In_235);
nand U2128 (N_2128,In_140,In_165);
or U2129 (N_2129,In_353,In_78);
nand U2130 (N_2130,In_106,In_516);
nor U2131 (N_2131,In_162,In_391);
nor U2132 (N_2132,In_448,In_86);
and U2133 (N_2133,In_363,In_2);
or U2134 (N_2134,In_403,In_250);
or U2135 (N_2135,In_519,In_509);
xor U2136 (N_2136,In_351,In_682);
nand U2137 (N_2137,In_746,In_588);
nand U2138 (N_2138,In_446,In_551);
and U2139 (N_2139,In_746,In_452);
nand U2140 (N_2140,In_418,In_528);
or U2141 (N_2141,In_312,In_197);
or U2142 (N_2142,In_277,In_655);
xnor U2143 (N_2143,In_543,In_722);
nand U2144 (N_2144,In_533,In_147);
nor U2145 (N_2145,In_215,In_513);
nand U2146 (N_2146,In_94,In_744);
nand U2147 (N_2147,In_183,In_234);
xnor U2148 (N_2148,In_552,In_54);
and U2149 (N_2149,In_517,In_133);
nor U2150 (N_2150,In_507,In_506);
nand U2151 (N_2151,In_134,In_172);
nor U2152 (N_2152,In_339,In_389);
or U2153 (N_2153,In_436,In_132);
nand U2154 (N_2154,In_56,In_7);
or U2155 (N_2155,In_600,In_690);
nand U2156 (N_2156,In_283,In_317);
and U2157 (N_2157,In_588,In_462);
or U2158 (N_2158,In_566,In_386);
or U2159 (N_2159,In_436,In_33);
or U2160 (N_2160,In_278,In_703);
and U2161 (N_2161,In_50,In_119);
or U2162 (N_2162,In_162,In_295);
nor U2163 (N_2163,In_318,In_523);
nand U2164 (N_2164,In_174,In_2);
nand U2165 (N_2165,In_2,In_41);
and U2166 (N_2166,In_677,In_241);
and U2167 (N_2167,In_110,In_290);
and U2168 (N_2168,In_381,In_116);
or U2169 (N_2169,In_420,In_475);
nor U2170 (N_2170,In_525,In_611);
and U2171 (N_2171,In_426,In_565);
and U2172 (N_2172,In_143,In_380);
nor U2173 (N_2173,In_138,In_114);
and U2174 (N_2174,In_664,In_39);
and U2175 (N_2175,In_404,In_648);
nand U2176 (N_2176,In_37,In_157);
nand U2177 (N_2177,In_346,In_542);
and U2178 (N_2178,In_439,In_362);
or U2179 (N_2179,In_377,In_469);
and U2180 (N_2180,In_411,In_608);
nand U2181 (N_2181,In_217,In_415);
nor U2182 (N_2182,In_346,In_379);
nand U2183 (N_2183,In_440,In_738);
or U2184 (N_2184,In_261,In_318);
nand U2185 (N_2185,In_450,In_695);
or U2186 (N_2186,In_274,In_600);
xnor U2187 (N_2187,In_94,In_222);
nor U2188 (N_2188,In_504,In_644);
nor U2189 (N_2189,In_330,In_98);
or U2190 (N_2190,In_697,In_43);
and U2191 (N_2191,In_131,In_541);
nor U2192 (N_2192,In_378,In_70);
nor U2193 (N_2193,In_46,In_181);
xnor U2194 (N_2194,In_51,In_429);
or U2195 (N_2195,In_570,In_379);
or U2196 (N_2196,In_320,In_170);
nor U2197 (N_2197,In_129,In_611);
or U2198 (N_2198,In_9,In_72);
and U2199 (N_2199,In_314,In_82);
or U2200 (N_2200,In_632,In_449);
nor U2201 (N_2201,In_529,In_369);
and U2202 (N_2202,In_246,In_405);
nor U2203 (N_2203,In_170,In_324);
nand U2204 (N_2204,In_488,In_656);
or U2205 (N_2205,In_474,In_472);
nor U2206 (N_2206,In_73,In_179);
or U2207 (N_2207,In_736,In_129);
nand U2208 (N_2208,In_190,In_517);
and U2209 (N_2209,In_119,In_298);
and U2210 (N_2210,In_330,In_22);
nor U2211 (N_2211,In_296,In_101);
nor U2212 (N_2212,In_643,In_124);
or U2213 (N_2213,In_605,In_572);
or U2214 (N_2214,In_293,In_447);
and U2215 (N_2215,In_236,In_512);
nand U2216 (N_2216,In_220,In_310);
or U2217 (N_2217,In_1,In_369);
or U2218 (N_2218,In_655,In_693);
xnor U2219 (N_2219,In_445,In_580);
or U2220 (N_2220,In_406,In_71);
xor U2221 (N_2221,In_358,In_271);
nand U2222 (N_2222,In_228,In_439);
nand U2223 (N_2223,In_5,In_80);
nor U2224 (N_2224,In_320,In_197);
and U2225 (N_2225,In_441,In_93);
nor U2226 (N_2226,In_459,In_35);
nor U2227 (N_2227,In_156,In_498);
or U2228 (N_2228,In_408,In_54);
nor U2229 (N_2229,In_646,In_654);
xnor U2230 (N_2230,In_496,In_278);
nand U2231 (N_2231,In_653,In_446);
or U2232 (N_2232,In_700,In_683);
nand U2233 (N_2233,In_194,In_38);
nor U2234 (N_2234,In_465,In_168);
or U2235 (N_2235,In_187,In_467);
or U2236 (N_2236,In_700,In_34);
or U2237 (N_2237,In_151,In_305);
xor U2238 (N_2238,In_329,In_234);
or U2239 (N_2239,In_89,In_315);
nor U2240 (N_2240,In_529,In_594);
nor U2241 (N_2241,In_680,In_643);
nand U2242 (N_2242,In_570,In_326);
or U2243 (N_2243,In_33,In_743);
and U2244 (N_2244,In_214,In_624);
or U2245 (N_2245,In_629,In_449);
xor U2246 (N_2246,In_207,In_465);
and U2247 (N_2247,In_497,In_745);
nor U2248 (N_2248,In_24,In_665);
and U2249 (N_2249,In_222,In_674);
nor U2250 (N_2250,In_189,In_75);
or U2251 (N_2251,In_571,In_134);
or U2252 (N_2252,In_371,In_446);
or U2253 (N_2253,In_220,In_185);
nor U2254 (N_2254,In_699,In_542);
or U2255 (N_2255,In_292,In_203);
nand U2256 (N_2256,In_245,In_581);
nand U2257 (N_2257,In_634,In_134);
and U2258 (N_2258,In_396,In_9);
xnor U2259 (N_2259,In_83,In_434);
or U2260 (N_2260,In_309,In_552);
or U2261 (N_2261,In_745,In_401);
nand U2262 (N_2262,In_696,In_375);
and U2263 (N_2263,In_516,In_439);
or U2264 (N_2264,In_746,In_269);
nor U2265 (N_2265,In_179,In_1);
and U2266 (N_2266,In_105,In_299);
nor U2267 (N_2267,In_585,In_312);
and U2268 (N_2268,In_715,In_375);
or U2269 (N_2269,In_737,In_268);
nand U2270 (N_2270,In_634,In_743);
and U2271 (N_2271,In_401,In_655);
nor U2272 (N_2272,In_210,In_445);
nand U2273 (N_2273,In_586,In_96);
and U2274 (N_2274,In_178,In_714);
nand U2275 (N_2275,In_305,In_41);
nor U2276 (N_2276,In_69,In_680);
or U2277 (N_2277,In_391,In_736);
nand U2278 (N_2278,In_230,In_210);
and U2279 (N_2279,In_127,In_584);
xor U2280 (N_2280,In_205,In_191);
nor U2281 (N_2281,In_456,In_357);
nand U2282 (N_2282,In_697,In_601);
nor U2283 (N_2283,In_627,In_620);
nand U2284 (N_2284,In_349,In_483);
and U2285 (N_2285,In_611,In_747);
nor U2286 (N_2286,In_15,In_442);
and U2287 (N_2287,In_28,In_111);
nor U2288 (N_2288,In_707,In_210);
nand U2289 (N_2289,In_607,In_294);
nand U2290 (N_2290,In_608,In_484);
or U2291 (N_2291,In_238,In_362);
or U2292 (N_2292,In_20,In_620);
or U2293 (N_2293,In_591,In_363);
nor U2294 (N_2294,In_47,In_600);
xor U2295 (N_2295,In_724,In_689);
nand U2296 (N_2296,In_374,In_663);
nand U2297 (N_2297,In_685,In_144);
xnor U2298 (N_2298,In_356,In_213);
nor U2299 (N_2299,In_309,In_477);
nor U2300 (N_2300,In_562,In_699);
nand U2301 (N_2301,In_699,In_230);
nand U2302 (N_2302,In_440,In_172);
nand U2303 (N_2303,In_405,In_437);
and U2304 (N_2304,In_80,In_643);
nand U2305 (N_2305,In_677,In_111);
or U2306 (N_2306,In_614,In_357);
nor U2307 (N_2307,In_98,In_26);
nand U2308 (N_2308,In_272,In_419);
nor U2309 (N_2309,In_234,In_244);
nor U2310 (N_2310,In_352,In_61);
or U2311 (N_2311,In_378,In_202);
and U2312 (N_2312,In_203,In_253);
xnor U2313 (N_2313,In_548,In_170);
nor U2314 (N_2314,In_75,In_564);
and U2315 (N_2315,In_105,In_456);
or U2316 (N_2316,In_237,In_479);
nor U2317 (N_2317,In_398,In_378);
and U2318 (N_2318,In_670,In_118);
nand U2319 (N_2319,In_203,In_487);
and U2320 (N_2320,In_234,In_152);
and U2321 (N_2321,In_337,In_6);
or U2322 (N_2322,In_343,In_17);
nor U2323 (N_2323,In_646,In_531);
and U2324 (N_2324,In_615,In_46);
and U2325 (N_2325,In_559,In_671);
nor U2326 (N_2326,In_120,In_245);
nor U2327 (N_2327,In_411,In_197);
nor U2328 (N_2328,In_638,In_492);
nor U2329 (N_2329,In_333,In_118);
or U2330 (N_2330,In_658,In_15);
nand U2331 (N_2331,In_437,In_250);
nor U2332 (N_2332,In_188,In_144);
or U2333 (N_2333,In_746,In_503);
nand U2334 (N_2334,In_721,In_180);
nor U2335 (N_2335,In_69,In_234);
nor U2336 (N_2336,In_10,In_3);
nand U2337 (N_2337,In_205,In_388);
or U2338 (N_2338,In_360,In_118);
xor U2339 (N_2339,In_336,In_294);
nand U2340 (N_2340,In_81,In_362);
nand U2341 (N_2341,In_670,In_574);
nand U2342 (N_2342,In_279,In_506);
nand U2343 (N_2343,In_274,In_738);
or U2344 (N_2344,In_352,In_340);
or U2345 (N_2345,In_506,In_147);
and U2346 (N_2346,In_479,In_378);
and U2347 (N_2347,In_725,In_314);
nand U2348 (N_2348,In_447,In_118);
and U2349 (N_2349,In_46,In_341);
and U2350 (N_2350,In_513,In_594);
nand U2351 (N_2351,In_132,In_353);
or U2352 (N_2352,In_686,In_385);
or U2353 (N_2353,In_497,In_545);
xor U2354 (N_2354,In_53,In_374);
xor U2355 (N_2355,In_342,In_442);
nand U2356 (N_2356,In_143,In_459);
and U2357 (N_2357,In_556,In_337);
nand U2358 (N_2358,In_348,In_636);
nand U2359 (N_2359,In_352,In_555);
or U2360 (N_2360,In_661,In_133);
nor U2361 (N_2361,In_90,In_570);
or U2362 (N_2362,In_95,In_321);
or U2363 (N_2363,In_391,In_664);
or U2364 (N_2364,In_571,In_201);
nand U2365 (N_2365,In_415,In_201);
or U2366 (N_2366,In_133,In_304);
nand U2367 (N_2367,In_668,In_718);
xnor U2368 (N_2368,In_138,In_328);
and U2369 (N_2369,In_49,In_275);
and U2370 (N_2370,In_154,In_377);
or U2371 (N_2371,In_661,In_276);
nand U2372 (N_2372,In_302,In_650);
nor U2373 (N_2373,In_698,In_601);
or U2374 (N_2374,In_205,In_203);
nor U2375 (N_2375,In_539,In_586);
nand U2376 (N_2376,In_662,In_208);
or U2377 (N_2377,In_16,In_79);
xnor U2378 (N_2378,In_615,In_377);
nand U2379 (N_2379,In_98,In_175);
xnor U2380 (N_2380,In_449,In_184);
nand U2381 (N_2381,In_540,In_743);
nand U2382 (N_2382,In_78,In_145);
nand U2383 (N_2383,In_294,In_601);
nor U2384 (N_2384,In_573,In_125);
or U2385 (N_2385,In_746,In_397);
xnor U2386 (N_2386,In_126,In_214);
or U2387 (N_2387,In_660,In_55);
or U2388 (N_2388,In_721,In_373);
nor U2389 (N_2389,In_583,In_207);
xnor U2390 (N_2390,In_86,In_274);
or U2391 (N_2391,In_542,In_524);
or U2392 (N_2392,In_29,In_122);
or U2393 (N_2393,In_180,In_119);
nand U2394 (N_2394,In_620,In_274);
nor U2395 (N_2395,In_184,In_550);
or U2396 (N_2396,In_591,In_40);
xnor U2397 (N_2397,In_69,In_79);
nand U2398 (N_2398,In_605,In_420);
nor U2399 (N_2399,In_253,In_749);
nor U2400 (N_2400,In_588,In_510);
and U2401 (N_2401,In_507,In_52);
nand U2402 (N_2402,In_283,In_555);
nor U2403 (N_2403,In_538,In_631);
nor U2404 (N_2404,In_299,In_481);
nand U2405 (N_2405,In_27,In_230);
and U2406 (N_2406,In_507,In_185);
or U2407 (N_2407,In_252,In_705);
or U2408 (N_2408,In_517,In_207);
xnor U2409 (N_2409,In_688,In_316);
nor U2410 (N_2410,In_243,In_458);
and U2411 (N_2411,In_460,In_739);
or U2412 (N_2412,In_697,In_602);
xor U2413 (N_2413,In_725,In_56);
or U2414 (N_2414,In_464,In_168);
or U2415 (N_2415,In_399,In_549);
or U2416 (N_2416,In_540,In_660);
nand U2417 (N_2417,In_209,In_370);
and U2418 (N_2418,In_583,In_316);
and U2419 (N_2419,In_133,In_628);
or U2420 (N_2420,In_196,In_715);
nand U2421 (N_2421,In_116,In_660);
or U2422 (N_2422,In_372,In_314);
xor U2423 (N_2423,In_622,In_67);
or U2424 (N_2424,In_403,In_687);
and U2425 (N_2425,In_158,In_486);
nand U2426 (N_2426,In_369,In_423);
nand U2427 (N_2427,In_423,In_593);
xnor U2428 (N_2428,In_516,In_141);
and U2429 (N_2429,In_720,In_577);
nand U2430 (N_2430,In_35,In_370);
nand U2431 (N_2431,In_502,In_42);
nand U2432 (N_2432,In_606,In_462);
and U2433 (N_2433,In_614,In_11);
nor U2434 (N_2434,In_722,In_361);
or U2435 (N_2435,In_590,In_190);
nor U2436 (N_2436,In_695,In_200);
nor U2437 (N_2437,In_9,In_450);
xor U2438 (N_2438,In_323,In_497);
nor U2439 (N_2439,In_278,In_662);
nand U2440 (N_2440,In_685,In_554);
nand U2441 (N_2441,In_339,In_732);
nand U2442 (N_2442,In_358,In_637);
or U2443 (N_2443,In_451,In_606);
nor U2444 (N_2444,In_497,In_262);
and U2445 (N_2445,In_673,In_579);
and U2446 (N_2446,In_97,In_588);
or U2447 (N_2447,In_243,In_517);
and U2448 (N_2448,In_563,In_228);
or U2449 (N_2449,In_596,In_274);
nand U2450 (N_2450,In_128,In_153);
and U2451 (N_2451,In_681,In_346);
nor U2452 (N_2452,In_15,In_139);
or U2453 (N_2453,In_225,In_121);
nand U2454 (N_2454,In_275,In_69);
xnor U2455 (N_2455,In_57,In_471);
or U2456 (N_2456,In_434,In_727);
nor U2457 (N_2457,In_640,In_468);
nor U2458 (N_2458,In_463,In_748);
or U2459 (N_2459,In_273,In_274);
nor U2460 (N_2460,In_489,In_710);
xor U2461 (N_2461,In_300,In_111);
and U2462 (N_2462,In_464,In_432);
nand U2463 (N_2463,In_435,In_537);
and U2464 (N_2464,In_617,In_625);
xor U2465 (N_2465,In_646,In_189);
nor U2466 (N_2466,In_533,In_551);
and U2467 (N_2467,In_502,In_696);
nor U2468 (N_2468,In_582,In_71);
nor U2469 (N_2469,In_493,In_273);
and U2470 (N_2470,In_55,In_38);
and U2471 (N_2471,In_406,In_495);
or U2472 (N_2472,In_166,In_214);
or U2473 (N_2473,In_384,In_238);
or U2474 (N_2474,In_663,In_543);
and U2475 (N_2475,In_257,In_741);
nor U2476 (N_2476,In_441,In_184);
xnor U2477 (N_2477,In_632,In_350);
or U2478 (N_2478,In_504,In_122);
nor U2479 (N_2479,In_714,In_156);
or U2480 (N_2480,In_332,In_350);
xnor U2481 (N_2481,In_134,In_620);
or U2482 (N_2482,In_355,In_460);
nor U2483 (N_2483,In_196,In_600);
nor U2484 (N_2484,In_171,In_381);
nand U2485 (N_2485,In_416,In_445);
nand U2486 (N_2486,In_680,In_708);
or U2487 (N_2487,In_324,In_581);
xnor U2488 (N_2488,In_98,In_401);
nor U2489 (N_2489,In_150,In_217);
and U2490 (N_2490,In_178,In_125);
and U2491 (N_2491,In_661,In_6);
or U2492 (N_2492,In_509,In_470);
and U2493 (N_2493,In_18,In_736);
xnor U2494 (N_2494,In_485,In_663);
and U2495 (N_2495,In_398,In_67);
and U2496 (N_2496,In_553,In_248);
nand U2497 (N_2497,In_120,In_89);
and U2498 (N_2498,In_513,In_166);
or U2499 (N_2499,In_457,In_501);
and U2500 (N_2500,N_65,N_276);
or U2501 (N_2501,N_1876,N_363);
nor U2502 (N_2502,N_2176,N_1020);
or U2503 (N_2503,N_1626,N_1557);
and U2504 (N_2504,N_1358,N_959);
or U2505 (N_2505,N_2425,N_2138);
and U2506 (N_2506,N_1912,N_1476);
and U2507 (N_2507,N_1695,N_988);
nor U2508 (N_2508,N_1605,N_639);
or U2509 (N_2509,N_371,N_1811);
nand U2510 (N_2510,N_1861,N_617);
nand U2511 (N_2511,N_1266,N_1933);
nand U2512 (N_2512,N_2487,N_1437);
or U2513 (N_2513,N_2091,N_991);
and U2514 (N_2514,N_1706,N_1508);
and U2515 (N_2515,N_1113,N_1349);
or U2516 (N_2516,N_2270,N_960);
xnor U2517 (N_2517,N_243,N_378);
nor U2518 (N_2518,N_500,N_1640);
nor U2519 (N_2519,N_2128,N_1218);
xnor U2520 (N_2520,N_2348,N_2253);
nand U2521 (N_2521,N_1857,N_161);
or U2522 (N_2522,N_2498,N_246);
nor U2523 (N_2523,N_2324,N_633);
xnor U2524 (N_2524,N_21,N_2135);
and U2525 (N_2525,N_2130,N_2032);
xnor U2526 (N_2526,N_1973,N_1918);
or U2527 (N_2527,N_682,N_1169);
or U2528 (N_2528,N_2318,N_2342);
or U2529 (N_2529,N_1592,N_1726);
xnor U2530 (N_2530,N_514,N_261);
or U2531 (N_2531,N_2462,N_2394);
nand U2532 (N_2532,N_1504,N_2048);
nor U2533 (N_2533,N_293,N_518);
nand U2534 (N_2534,N_1791,N_2315);
nand U2535 (N_2535,N_977,N_740);
and U2536 (N_2536,N_1549,N_551);
xnor U2537 (N_2537,N_928,N_874);
and U2538 (N_2538,N_461,N_655);
and U2539 (N_2539,N_521,N_140);
or U2540 (N_2540,N_1075,N_1324);
or U2541 (N_2541,N_1907,N_1537);
xor U2542 (N_2542,N_1170,N_1021);
and U2543 (N_2543,N_1301,N_813);
and U2544 (N_2544,N_1931,N_41);
and U2545 (N_2545,N_632,N_1087);
and U2546 (N_2546,N_1765,N_359);
or U2547 (N_2547,N_116,N_305);
or U2548 (N_2548,N_793,N_772);
or U2549 (N_2549,N_70,N_1018);
nand U2550 (N_2550,N_473,N_75);
xnor U2551 (N_2551,N_221,N_525);
nor U2552 (N_2552,N_2037,N_1274);
nand U2553 (N_2553,N_1243,N_1828);
nor U2554 (N_2554,N_522,N_468);
xor U2555 (N_2555,N_47,N_2145);
or U2556 (N_2556,N_260,N_1397);
nand U2557 (N_2557,N_1875,N_1685);
nor U2558 (N_2558,N_332,N_12);
nor U2559 (N_2559,N_155,N_318);
xnor U2560 (N_2560,N_1402,N_636);
and U2561 (N_2561,N_382,N_1011);
nor U2562 (N_2562,N_104,N_274);
nand U2563 (N_2563,N_1763,N_257);
nor U2564 (N_2564,N_2167,N_1375);
or U2565 (N_2565,N_1153,N_1328);
and U2566 (N_2566,N_1280,N_786);
nor U2567 (N_2567,N_2075,N_109);
or U2568 (N_2568,N_567,N_1500);
nor U2569 (N_2569,N_267,N_590);
nand U2570 (N_2570,N_1787,N_73);
and U2571 (N_2571,N_903,N_1817);
nor U2572 (N_2572,N_1968,N_1072);
nor U2573 (N_2573,N_2300,N_2197);
and U2574 (N_2574,N_2426,N_1942);
nor U2575 (N_2575,N_1834,N_728);
nor U2576 (N_2576,N_346,N_1486);
or U2577 (N_2577,N_212,N_1454);
nand U2578 (N_2578,N_238,N_1228);
nand U2579 (N_2579,N_1330,N_1693);
or U2580 (N_2580,N_1841,N_701);
nand U2581 (N_2581,N_1434,N_1022);
xnor U2582 (N_2582,N_1989,N_1095);
nor U2583 (N_2583,N_1300,N_571);
and U2584 (N_2584,N_58,N_125);
nor U2585 (N_2585,N_54,N_2148);
and U2586 (N_2586,N_232,N_1479);
nand U2587 (N_2587,N_2183,N_19);
or U2588 (N_2588,N_123,N_1269);
and U2589 (N_2589,N_1611,N_26);
and U2590 (N_2590,N_846,N_1908);
and U2591 (N_2591,N_887,N_979);
nand U2592 (N_2592,N_1248,N_2217);
nor U2593 (N_2593,N_338,N_896);
and U2594 (N_2594,N_533,N_1591);
nor U2595 (N_2595,N_1576,N_1452);
or U2596 (N_2596,N_1085,N_2186);
or U2597 (N_2597,N_1847,N_618);
and U2598 (N_2598,N_2356,N_1029);
or U2599 (N_2599,N_62,N_357);
nor U2600 (N_2600,N_2435,N_491);
and U2601 (N_2601,N_1713,N_537);
nand U2602 (N_2602,N_1383,N_2257);
nand U2603 (N_2603,N_615,N_727);
or U2604 (N_2604,N_2361,N_366);
and U2605 (N_2605,N_910,N_474);
nand U2606 (N_2606,N_900,N_1762);
xnor U2607 (N_2607,N_483,N_1715);
and U2608 (N_2608,N_817,N_2499);
or U2609 (N_2609,N_5,N_1356);
or U2610 (N_2610,N_1172,N_2073);
nor U2611 (N_2611,N_983,N_1894);
nand U2612 (N_2612,N_1319,N_2364);
nand U2613 (N_2613,N_2280,N_1002);
nor U2614 (N_2614,N_1914,N_3);
and U2615 (N_2615,N_2164,N_2005);
nor U2616 (N_2616,N_2424,N_2255);
and U2617 (N_2617,N_139,N_87);
nor U2618 (N_2618,N_170,N_2235);
or U2619 (N_2619,N_1167,N_1975);
or U2620 (N_2620,N_2294,N_1325);
nor U2621 (N_2621,N_511,N_1831);
and U2622 (N_2622,N_766,N_1642);
xnor U2623 (N_2623,N_148,N_469);
nand U2624 (N_2624,N_2093,N_370);
nand U2625 (N_2625,N_224,N_179);
nand U2626 (N_2626,N_465,N_1039);
nand U2627 (N_2627,N_2132,N_547);
and U2628 (N_2628,N_2427,N_194);
nor U2629 (N_2629,N_1806,N_2021);
or U2630 (N_2630,N_2221,N_1065);
or U2631 (N_2631,N_1,N_872);
or U2632 (N_2632,N_953,N_1886);
or U2633 (N_2633,N_1601,N_1524);
nor U2634 (N_2634,N_250,N_1044);
nand U2635 (N_2635,N_132,N_29);
or U2636 (N_2636,N_1921,N_1850);
or U2637 (N_2637,N_2036,N_1543);
nand U2638 (N_2638,N_773,N_815);
and U2639 (N_2639,N_287,N_957);
xnor U2640 (N_2640,N_171,N_2468);
xor U2641 (N_2641,N_1106,N_669);
or U2642 (N_2642,N_133,N_334);
nand U2643 (N_2643,N_2219,N_1988);
or U2644 (N_2644,N_311,N_858);
xnor U2645 (N_2645,N_2063,N_1037);
nand U2646 (N_2646,N_1822,N_2284);
nand U2647 (N_2647,N_820,N_427);
nor U2648 (N_2648,N_1070,N_2391);
or U2649 (N_2649,N_320,N_2290);
nand U2650 (N_2650,N_195,N_1023);
and U2651 (N_2651,N_1845,N_1751);
and U2652 (N_2652,N_690,N_2430);
and U2653 (N_2653,N_2188,N_253);
or U2654 (N_2654,N_1802,N_2311);
or U2655 (N_2655,N_1635,N_1938);
or U2656 (N_2656,N_2367,N_621);
or U2657 (N_2657,N_1949,N_2377);
nand U2658 (N_2658,N_993,N_1374);
nand U2659 (N_2659,N_2136,N_752);
and U2660 (N_2660,N_559,N_1798);
nand U2661 (N_2661,N_169,N_2309);
xor U2662 (N_2662,N_1177,N_442);
nand U2663 (N_2663,N_1441,N_1317);
or U2664 (N_2664,N_723,N_1760);
and U2665 (N_2665,N_118,N_738);
xor U2666 (N_2666,N_386,N_905);
and U2667 (N_2667,N_583,N_2368);
nand U2668 (N_2668,N_1745,N_1796);
nand U2669 (N_2669,N_542,N_698);
and U2670 (N_2670,N_8,N_2258);
or U2671 (N_2671,N_2068,N_672);
xor U2672 (N_2672,N_2343,N_2001);
nor U2673 (N_2673,N_201,N_143);
nor U2674 (N_2674,N_845,N_1493);
nand U2675 (N_2675,N_278,N_1048);
and U2676 (N_2676,N_784,N_2259);
nor U2677 (N_2677,N_1547,N_647);
nand U2678 (N_2678,N_59,N_891);
or U2679 (N_2679,N_251,N_1308);
xnor U2680 (N_2680,N_1080,N_455);
nand U2681 (N_2681,N_966,N_436);
xnor U2682 (N_2682,N_906,N_1323);
nand U2683 (N_2683,N_38,N_1136);
nand U2684 (N_2684,N_981,N_1928);
nand U2685 (N_2685,N_2023,N_875);
nor U2686 (N_2686,N_2440,N_1285);
nor U2687 (N_2687,N_1016,N_1904);
xnor U2688 (N_2688,N_1945,N_1940);
nor U2689 (N_2689,N_708,N_785);
nand U2690 (N_2690,N_1423,N_605);
and U2691 (N_2691,N_31,N_1736);
xor U2692 (N_2692,N_753,N_1499);
nand U2693 (N_2693,N_331,N_829);
and U2694 (N_2694,N_2011,N_265);
and U2695 (N_2695,N_877,N_2305);
xnor U2696 (N_2696,N_641,N_2140);
nand U2697 (N_2697,N_271,N_1162);
xor U2698 (N_2698,N_2481,N_1719);
or U2699 (N_2699,N_2269,N_831);
nor U2700 (N_2700,N_1922,N_105);
nor U2701 (N_2701,N_1226,N_980);
nor U2702 (N_2702,N_627,N_1830);
nor U2703 (N_2703,N_184,N_2155);
xnor U2704 (N_2704,N_1270,N_1478);
nor U2705 (N_2705,N_2121,N_2473);
or U2706 (N_2706,N_1316,N_1755);
nand U2707 (N_2707,N_1345,N_965);
nand U2708 (N_2708,N_866,N_2325);
nor U2709 (N_2709,N_941,N_1497);
nand U2710 (N_2710,N_403,N_1871);
nand U2711 (N_2711,N_1502,N_1146);
nand U2712 (N_2712,N_803,N_396);
nand U2713 (N_2713,N_2019,N_1916);
xnor U2714 (N_2714,N_218,N_2218);
xnor U2715 (N_2715,N_1887,N_827);
nor U2716 (N_2716,N_272,N_1665);
nand U2717 (N_2717,N_1128,N_266);
nand U2718 (N_2718,N_1978,N_931);
nand U2719 (N_2719,N_1003,N_2224);
or U2720 (N_2720,N_187,N_2228);
nand U2721 (N_2721,N_2483,N_1141);
or U2722 (N_2722,N_2264,N_660);
or U2723 (N_2723,N_1560,N_1032);
and U2724 (N_2724,N_225,N_95);
nor U2725 (N_2725,N_1326,N_946);
and U2726 (N_2726,N_2388,N_2112);
or U2727 (N_2727,N_611,N_799);
nor U2728 (N_2728,N_1006,N_1027);
nand U2729 (N_2729,N_864,N_1976);
and U2730 (N_2730,N_592,N_870);
nand U2731 (N_2731,N_1779,N_2243);
nand U2732 (N_2732,N_750,N_317);
nor U2733 (N_2733,N_1766,N_2213);
and U2734 (N_2734,N_1009,N_2098);
nand U2735 (N_2735,N_1111,N_2191);
nand U2736 (N_2736,N_2071,N_1463);
nor U2737 (N_2737,N_2107,N_854);
and U2738 (N_2738,N_178,N_1951);
xnor U2739 (N_2739,N_1073,N_1086);
nor U2740 (N_2740,N_1137,N_2190);
nor U2741 (N_2741,N_1564,N_2436);
or U2742 (N_2742,N_2281,N_247);
xor U2743 (N_2743,N_973,N_323);
nor U2744 (N_2744,N_984,N_630);
or U2745 (N_2745,N_254,N_1151);
or U2746 (N_2746,N_2118,N_2072);
and U2747 (N_2747,N_2474,N_154);
nor U2748 (N_2748,N_1298,N_2469);
and U2749 (N_2749,N_1281,N_702);
nand U2750 (N_2750,N_1740,N_1898);
nand U2751 (N_2751,N_2094,N_421);
and U2752 (N_2752,N_1821,N_2015);
nand U2753 (N_2753,N_1874,N_411);
and U2754 (N_2754,N_2334,N_1220);
or U2755 (N_2755,N_1679,N_353);
nand U2756 (N_2756,N_2248,N_86);
and U2757 (N_2757,N_1173,N_1772);
or U2758 (N_2758,N_230,N_1789);
or U2759 (N_2759,N_602,N_2331);
nand U2760 (N_2760,N_2082,N_2042);
nor U2761 (N_2761,N_1292,N_942);
and U2762 (N_2762,N_2491,N_1692);
nor U2763 (N_2763,N_433,N_2156);
nand U2764 (N_2764,N_1004,N_1716);
nor U2765 (N_2765,N_2030,N_2446);
or U2766 (N_2766,N_1707,N_1117);
or U2767 (N_2767,N_1133,N_2344);
nand U2768 (N_2768,N_352,N_613);
nor U2769 (N_2769,N_2204,N_622);
nor U2770 (N_2770,N_1149,N_2053);
or U2771 (N_2771,N_1013,N_1401);
or U2772 (N_2772,N_398,N_1371);
nand U2773 (N_2773,N_1484,N_2234);
or U2774 (N_2774,N_640,N_493);
and U2775 (N_2775,N_2395,N_1333);
xor U2776 (N_2776,N_1334,N_2151);
or U2777 (N_2777,N_1844,N_956);
nor U2778 (N_2778,N_1064,N_1473);
nand U2779 (N_2779,N_2389,N_594);
xor U2780 (N_2780,N_1846,N_7);
nand U2781 (N_2781,N_1235,N_2060);
or U2782 (N_2782,N_2495,N_130);
nand U2783 (N_2783,N_1671,N_1498);
and U2784 (N_2784,N_724,N_1739);
or U2785 (N_2785,N_1122,N_479);
nor U2786 (N_2786,N_2406,N_309);
and U2787 (N_2787,N_901,N_2051);
nand U2788 (N_2788,N_924,N_573);
xor U2789 (N_2789,N_1666,N_2116);
or U2790 (N_2790,N_591,N_907);
or U2791 (N_2791,N_177,N_1572);
xor U2792 (N_2792,N_328,N_1824);
nor U2793 (N_2793,N_2025,N_685);
xnor U2794 (N_2794,N_743,N_2285);
or U2795 (N_2795,N_1534,N_1078);
nand U2796 (N_2796,N_1691,N_1678);
nand U2797 (N_2797,N_2332,N_108);
and U2798 (N_2798,N_2404,N_2421);
xnor U2799 (N_2799,N_1418,N_1287);
nor U2800 (N_2800,N_1362,N_1110);
or U2801 (N_2801,N_85,N_2307);
nand U2802 (N_2802,N_1066,N_2077);
nor U2803 (N_2803,N_1741,N_2102);
nor U2804 (N_2804,N_149,N_68);
nand U2805 (N_2805,N_2454,N_197);
xnor U2806 (N_2806,N_1361,N_1494);
nor U2807 (N_2807,N_1115,N_836);
xor U2808 (N_2808,N_1756,N_175);
nand U2809 (N_2809,N_1247,N_1757);
nor U2810 (N_2810,N_1651,N_2049);
and U2811 (N_2811,N_308,N_152);
nor U2812 (N_2812,N_2439,N_2316);
nor U2813 (N_2813,N_1419,N_1276);
nor U2814 (N_2814,N_998,N_2292);
xnor U2815 (N_2815,N_563,N_781);
and U2816 (N_2816,N_516,N_1878);
nor U2817 (N_2817,N_1142,N_1105);
xor U2818 (N_2818,N_1033,N_1184);
nor U2819 (N_2819,N_2423,N_1744);
xnor U2820 (N_2820,N_968,N_709);
and U2821 (N_2821,N_2268,N_1879);
xnor U2822 (N_2822,N_294,N_2397);
nor U2823 (N_2823,N_2414,N_284);
nor U2824 (N_2824,N_607,N_519);
nand U2825 (N_2825,N_37,N_2407);
or U2826 (N_2826,N_992,N_2383);
or U2827 (N_2827,N_662,N_1536);
nor U2828 (N_2828,N_1015,N_1134);
nor U2829 (N_2829,N_385,N_34);
nand U2830 (N_2830,N_2146,N_1414);
nor U2831 (N_2831,N_415,N_1465);
or U2832 (N_2832,N_2222,N_1725);
and U2833 (N_2833,N_499,N_1781);
nand U2834 (N_2834,N_2058,N_847);
and U2835 (N_2835,N_470,N_1246);
and U2836 (N_2836,N_1118,N_1208);
or U2837 (N_2837,N_400,N_964);
nor U2838 (N_2838,N_1785,N_1188);
or U2839 (N_2839,N_277,N_2003);
nand U2840 (N_2840,N_2143,N_2413);
nor U2841 (N_2841,N_1863,N_1299);
and U2842 (N_2842,N_2119,N_1081);
nor U2843 (N_2843,N_2067,N_768);
or U2844 (N_2844,N_1820,N_2434);
nor U2845 (N_2845,N_2247,N_1152);
xnor U2846 (N_2846,N_1377,N_1223);
and U2847 (N_2847,N_1225,N_72);
nand U2848 (N_2848,N_731,N_1838);
nor U2849 (N_2849,N_2341,N_498);
and U2850 (N_2850,N_623,N_2412);
nand U2851 (N_2851,N_733,N_477);
or U2852 (N_2852,N_10,N_1379);
nand U2853 (N_2853,N_2452,N_1747);
xor U2854 (N_2854,N_1311,N_585);
xnor U2855 (N_2855,N_2338,N_1239);
nand U2856 (N_2856,N_577,N_2340);
xnor U2857 (N_2857,N_1742,N_2131);
and U2858 (N_2858,N_1631,N_1539);
and U2859 (N_2859,N_2443,N_297);
nand U2860 (N_2860,N_190,N_1034);
nand U2861 (N_2861,N_1800,N_2056);
and U2862 (N_2862,N_2239,N_716);
nor U2863 (N_2863,N_2327,N_612);
xor U2864 (N_2864,N_1643,N_1659);
nand U2865 (N_2865,N_674,N_2245);
nand U2866 (N_2866,N_1185,N_1495);
or U2867 (N_2867,N_288,N_2225);
nor U2868 (N_2868,N_673,N_2124);
and U2869 (N_2869,N_1718,N_216);
nand U2870 (N_2870,N_1815,N_546);
or U2871 (N_2871,N_2366,N_2192);
and U2872 (N_2872,N_1909,N_2357);
and U2873 (N_2873,N_1438,N_1077);
or U2874 (N_2874,N_1565,N_2162);
nor U2875 (N_2875,N_44,N_98);
nand U2876 (N_2876,N_2139,N_406);
or U2877 (N_2877,N_186,N_1813);
or U2878 (N_2878,N_729,N_1937);
or U2879 (N_2879,N_715,N_295);
or U2880 (N_2880,N_1060,N_310);
nand U2881 (N_2881,N_1343,N_330);
nand U2882 (N_2882,N_1114,N_1112);
nor U2883 (N_2883,N_2321,N_264);
or U2884 (N_2884,N_688,N_241);
nor U2885 (N_2885,N_1131,N_1069);
nor U2886 (N_2886,N_1602,N_1517);
and U2887 (N_2887,N_1271,N_1786);
xnor U2888 (N_2888,N_1624,N_1108);
nand U2889 (N_2889,N_157,N_168);
nand U2890 (N_2890,N_1203,N_687);
or U2891 (N_2891,N_1250,N_579);
and U2892 (N_2892,N_115,N_30);
xnor U2893 (N_2893,N_191,N_1544);
nor U2894 (N_2894,N_1145,N_1888);
and U2895 (N_2895,N_2158,N_678);
or U2896 (N_2896,N_1840,N_492);
nor U2897 (N_2897,N_325,N_1296);
or U2898 (N_2898,N_1620,N_783);
and U2899 (N_2899,N_2198,N_1157);
xor U2900 (N_2900,N_2057,N_217);
xnor U2901 (N_2901,N_2043,N_391);
and U2902 (N_2902,N_600,N_163);
and U2903 (N_2903,N_200,N_855);
xor U2904 (N_2904,N_2010,N_1373);
xor U2905 (N_2905,N_1934,N_696);
nand U2906 (N_2906,N_555,N_1451);
nor U2907 (N_2907,N_439,N_1364);
nand U2908 (N_2908,N_2438,N_684);
and U2909 (N_2909,N_444,N_2265);
nand U2910 (N_2910,N_1853,N_1297);
or U2911 (N_2911,N_2034,N_2374);
or U2912 (N_2912,N_1783,N_298);
or U2913 (N_2913,N_1868,N_1974);
and U2914 (N_2914,N_1955,N_1552);
xnor U2915 (N_2915,N_162,N_2018);
and U2916 (N_2916,N_188,N_1284);
and U2917 (N_2917,N_628,N_1551);
nor U2918 (N_2918,N_951,N_596);
and U2919 (N_2919,N_919,N_262);
and U2920 (N_2920,N_850,N_1190);
and U2921 (N_2921,N_1354,N_2287);
or U2922 (N_2922,N_1369,N_759);
nor U2923 (N_2923,N_2352,N_1618);
nand U2924 (N_2924,N_1542,N_176);
nand U2925 (N_2925,N_2154,N_868);
and U2926 (N_2926,N_544,N_46);
nand U2927 (N_2927,N_1697,N_2471);
and U2928 (N_2928,N_653,N_510);
and U2929 (N_2929,N_2310,N_2196);
and U2930 (N_2930,N_686,N_535);
xnor U2931 (N_2931,N_1014,N_1279);
nand U2932 (N_2932,N_1610,N_2086);
nor U2933 (N_2933,N_1729,N_2184);
nor U2934 (N_2934,N_1683,N_1573);
nand U2935 (N_2935,N_426,N_80);
xnor U2936 (N_2936,N_1689,N_1468);
and U2937 (N_2937,N_1776,N_1843);
or U2938 (N_2938,N_2223,N_570);
nand U2939 (N_2939,N_438,N_1723);
nand U2940 (N_2940,N_713,N_970);
xor U2941 (N_2941,N_997,N_2460);
nor U2942 (N_2942,N_2323,N_1049);
and U2943 (N_2943,N_2293,N_1035);
nor U2944 (N_2944,N_456,N_381);
nor U2945 (N_2945,N_955,N_865);
and U2946 (N_2946,N_540,N_1667);
nand U2947 (N_2947,N_839,N_823);
nor U2948 (N_2948,N_597,N_27);
nand U2949 (N_2949,N_2161,N_1807);
and U2950 (N_2950,N_1481,N_1529);
or U2951 (N_2951,N_1489,N_2220);
nand U2952 (N_2952,N_101,N_646);
nand U2953 (N_2953,N_464,N_2013);
or U2954 (N_2954,N_1612,N_828);
or U2955 (N_2955,N_392,N_167);
nor U2956 (N_2956,N_897,N_915);
and U2957 (N_2957,N_1771,N_1905);
and U2958 (N_2958,N_1480,N_884);
nand U2959 (N_2959,N_146,N_1261);
nand U2960 (N_2960,N_1943,N_2142);
nor U2961 (N_2961,N_1047,N_578);
and U2962 (N_2962,N_707,N_206);
and U2963 (N_2963,N_1230,N_520);
nor U2964 (N_2964,N_529,N_365);
nor U2965 (N_2965,N_895,N_1946);
nand U2966 (N_2966,N_890,N_79);
nor U2967 (N_2967,N_1063,N_1986);
nand U2968 (N_2968,N_393,N_2444);
nand U2969 (N_2969,N_2458,N_747);
and U2970 (N_2970,N_336,N_982);
or U2971 (N_2971,N_292,N_2026);
nor U2972 (N_2972,N_1192,N_654);
and U2973 (N_2973,N_180,N_402);
or U2974 (N_2974,N_1553,N_985);
nand U2975 (N_2975,N_671,N_113);
nand U2976 (N_2976,N_2000,N_1242);
and U2977 (N_2977,N_205,N_704);
xnor U2978 (N_2978,N_650,N_742);
or U2979 (N_2979,N_844,N_818);
xnor U2980 (N_2980,N_1351,N_39);
and U2981 (N_2981,N_1926,N_122);
nand U2982 (N_2982,N_2267,N_15);
nor U2983 (N_2983,N_703,N_1604);
and U2984 (N_2984,N_598,N_871);
or U2985 (N_2985,N_390,N_2153);
or U2986 (N_2986,N_952,N_2047);
and U2987 (N_2987,N_364,N_2169);
or U2988 (N_2988,N_1211,N_307);
nand U2989 (N_2989,N_349,N_372);
or U2990 (N_2990,N_2163,N_252);
or U2991 (N_2991,N_620,N_719);
nor U2992 (N_2992,N_1808,N_2402);
nand U2993 (N_2993,N_1554,N_1139);
nand U2994 (N_2994,N_860,N_629);
and U2995 (N_2995,N_1872,N_1059);
nor U2996 (N_2996,N_971,N_2100);
or U2997 (N_2997,N_48,N_2240);
nand U2998 (N_2998,N_405,N_2306);
and U2999 (N_2999,N_2195,N_1200);
or U3000 (N_3000,N_2451,N_1124);
nand U3001 (N_3001,N_351,N_2350);
xor U3002 (N_3002,N_2,N_1525);
nand U3003 (N_3003,N_222,N_1599);
nand U3004 (N_3004,N_1915,N_1099);
and U3005 (N_3005,N_213,N_681);
and U3006 (N_3006,N_2006,N_1550);
nor U3007 (N_3007,N_1570,N_458);
nor U3008 (N_3008,N_1140,N_1555);
or U3009 (N_3009,N_748,N_1094);
xor U3010 (N_3010,N_2493,N_527);
nor U3011 (N_3011,N_2479,N_172);
or U3012 (N_3012,N_638,N_1273);
or U3013 (N_3013,N_2429,N_1953);
and U3014 (N_3014,N_1265,N_501);
nand U3015 (N_3015,N_380,N_593);
or U3016 (N_3016,N_568,N_78);
nand U3017 (N_3017,N_2486,N_100);
nor U3018 (N_3018,N_487,N_1455);
and U3019 (N_3019,N_668,N_220);
nand U3020 (N_3020,N_142,N_1393);
or U3021 (N_3021,N_649,N_582);
and U3022 (N_3022,N_144,N_562);
and U3023 (N_3023,N_746,N_45);
or U3024 (N_3024,N_1470,N_1982);
nor U3025 (N_3025,N_327,N_81);
nor U3026 (N_3026,N_1743,N_1731);
nor U3027 (N_3027,N_1215,N_948);
and U3028 (N_3028,N_451,N_303);
or U3029 (N_3029,N_333,N_2482);
nor U3030 (N_3030,N_699,N_2096);
or U3031 (N_3031,N_2382,N_635);
nand U3032 (N_3032,N_677,N_420);
nor U3033 (N_3033,N_1198,N_2279);
nor U3034 (N_3034,N_1045,N_2016);
nor U3035 (N_3035,N_1538,N_401);
nor U3036 (N_3036,N_202,N_782);
nor U3037 (N_3037,N_2392,N_2205);
nor U3038 (N_3038,N_1224,N_2433);
nand U3039 (N_3039,N_1335,N_730);
and U3040 (N_3040,N_838,N_2097);
and U3041 (N_3041,N_1346,N_2230);
and U3042 (N_3042,N_1129,N_697);
or U3043 (N_3043,N_1302,N_1439);
or U3044 (N_3044,N_1390,N_2372);
nand U3045 (N_3045,N_181,N_2303);
nor U3046 (N_3046,N_859,N_56);
or U3047 (N_3047,N_1597,N_812);
nor U3048 (N_3048,N_2211,N_24);
nand U3049 (N_3049,N_1019,N_737);
nor U3050 (N_3050,N_1368,N_676);
nor U3051 (N_3051,N_2398,N_1232);
and U3052 (N_3052,N_1036,N_534);
nand U3053 (N_3053,N_1410,N_778);
or U3054 (N_3054,N_1866,N_2083);
nand U3055 (N_3055,N_2050,N_976);
nor U3056 (N_3056,N_1594,N_1431);
xor U3057 (N_3057,N_1089,N_495);
nor U3058 (N_3058,N_862,N_2066);
nand U3059 (N_3059,N_1407,N_1130);
or U3060 (N_3060,N_430,N_1983);
nor U3061 (N_3061,N_379,N_1206);
and U3062 (N_3062,N_1176,N_610);
nor U3063 (N_3063,N_1630,N_228);
or U3064 (N_3064,N_777,N_76);
and U3065 (N_3065,N_1711,N_1286);
or U3066 (N_3066,N_1753,N_2173);
nand U3067 (N_3067,N_1897,N_929);
nand U3068 (N_3068,N_625,N_2062);
nor U3069 (N_3069,N_1471,N_819);
nand U3070 (N_3070,N_478,N_826);
or U3071 (N_3071,N_926,N_588);
nor U3072 (N_3072,N_1491,N_1429);
nand U3073 (N_3073,N_60,N_925);
nor U3074 (N_3074,N_804,N_648);
nor U3075 (N_3075,N_2496,N_2202);
nor U3076 (N_3076,N_2059,N_2246);
and U3077 (N_3077,N_1645,N_2411);
nor U3078 (N_3078,N_324,N_880);
nand U3079 (N_3079,N_505,N_1984);
and U3080 (N_3080,N_1522,N_429);
or U3081 (N_3081,N_2009,N_2232);
and U3082 (N_3082,N_506,N_64);
or U3083 (N_3083,N_1312,N_314);
and U3084 (N_3084,N_1282,N_1458);
and U3085 (N_3085,N_1865,N_1617);
nand U3086 (N_3086,N_1428,N_347);
or U3087 (N_3087,N_878,N_1588);
nand U3088 (N_3088,N_962,N_1629);
or U3089 (N_3089,N_526,N_1994);
nand U3090 (N_3090,N_1327,N_2319);
and U3091 (N_3091,N_714,N_987);
or U3092 (N_3092,N_198,N_136);
and U3093 (N_3093,N_1165,N_383);
and U3094 (N_3094,N_659,N_1202);
nand U3095 (N_3095,N_1295,N_2302);
nor U3096 (N_3096,N_1780,N_1990);
and U3097 (N_3097,N_1854,N_399);
nand U3098 (N_3098,N_1180,N_1969);
nor U3099 (N_3099,N_899,N_2045);
and U3100 (N_3100,N_2046,N_0);
nand U3101 (N_3101,N_2378,N_2365);
and U3102 (N_3102,N_1858,N_2249);
and U3103 (N_3103,N_938,N_2110);
nor U3104 (N_3104,N_1043,N_1126);
xor U3105 (N_3105,N_1639,N_1699);
nor U3106 (N_3106,N_475,N_825);
nand U3107 (N_3107,N_2490,N_606);
or U3108 (N_3108,N_404,N_33);
xnor U3109 (N_3109,N_1566,N_2420);
and U3110 (N_3110,N_1205,N_358);
nor U3111 (N_3111,N_1950,N_2113);
or U3112 (N_3112,N_2384,N_1892);
nor U3113 (N_3113,N_645,N_967);
nor U3114 (N_3114,N_1240,N_1443);
nand U3115 (N_3115,N_1911,N_507);
or U3116 (N_3116,N_285,N_211);
xor U3117 (N_3117,N_1616,N_249);
xor U3118 (N_3118,N_1456,N_1159);
and U3119 (N_3119,N_97,N_1026);
and U3120 (N_3120,N_340,N_1448);
or U3121 (N_3121,N_2126,N_601);
nand U3122 (N_3122,N_1816,N_1530);
and U3123 (N_3123,N_1728,N_1656);
or U3124 (N_3124,N_1450,N_1930);
or U3125 (N_3125,N_2238,N_150);
or U3126 (N_3126,N_1359,N_1520);
and U3127 (N_3127,N_239,N_735);
nor U3128 (N_3128,N_9,N_1754);
xnor U3129 (N_3129,N_453,N_193);
or U3130 (N_3130,N_1187,N_440);
or U3131 (N_3131,N_102,N_1233);
nor U3132 (N_3132,N_1805,N_739);
and U3133 (N_3133,N_675,N_1580);
or U3134 (N_3134,N_343,N_797);
xor U3135 (N_3135,N_435,N_2330);
and U3136 (N_3136,N_204,N_1427);
xor U3137 (N_3137,N_756,N_637);
nand U3138 (N_3138,N_1322,N_2061);
nand U3139 (N_3139,N_2298,N_1347);
nand U3140 (N_3140,N_1143,N_1890);
nand U3141 (N_3141,N_972,N_425);
nor U3142 (N_3142,N_2274,N_1827);
or U3143 (N_3143,N_1156,N_1913);
nand U3144 (N_3144,N_700,N_103);
and U3145 (N_3145,N_2177,N_236);
or U3146 (N_3146,N_1608,N_545);
nor U3147 (N_3147,N_1088,N_861);
or U3148 (N_3148,N_2129,N_1353);
nor U3149 (N_3149,N_2203,N_1182);
xnor U3150 (N_3150,N_1814,N_1884);
xnor U3151 (N_3151,N_89,N_1793);
nor U3152 (N_3152,N_1721,N_1531);
nand U3153 (N_3153,N_1648,N_1724);
and U3154 (N_3154,N_892,N_1163);
xnor U3155 (N_3155,N_414,N_1216);
nor U3156 (N_3156,N_1394,N_564);
nand U3157 (N_3157,N_1199,N_2109);
nor U3158 (N_3158,N_651,N_2179);
nor U3159 (N_3159,N_1510,N_1584);
nand U3160 (N_3160,N_745,N_248);
nand U3161 (N_3161,N_842,N_2456);
or U3162 (N_3162,N_1160,N_1966);
or U3163 (N_3163,N_1829,N_1971);
nor U3164 (N_3164,N_166,N_1462);
xnor U3165 (N_3165,N_1264,N_2379);
nor U3166 (N_3166,N_2080,N_1768);
nor U3167 (N_3167,N_376,N_1511);
or U3168 (N_3168,N_418,N_2422);
xnor U3169 (N_3169,N_1251,N_1249);
nor U3170 (N_3170,N_2076,N_1384);
nand U3171 (N_3171,N_1363,N_57);
nand U3172 (N_3172,N_99,N_1686);
or U3173 (N_3173,N_807,N_20);
nand U3174 (N_3174,N_1365,N_1939);
nand U3175 (N_3175,N_2104,N_51);
nand U3176 (N_3176,N_2296,N_1416);
or U3177 (N_3177,N_1031,N_2078);
or U3178 (N_3178,N_1132,N_853);
or U3179 (N_3179,N_2428,N_502);
nand U3180 (N_3180,N_569,N_2295);
nand U3181 (N_3181,N_360,N_35);
nand U3182 (N_3182,N_43,N_587);
and U3183 (N_3183,N_1116,N_1799);
and U3184 (N_3184,N_2201,N_1360);
and U3185 (N_3185,N_387,N_790);
nand U3186 (N_3186,N_1698,N_883);
nand U3187 (N_3187,N_1746,N_1501);
nand U3188 (N_3188,N_299,N_912);
xor U3189 (N_3189,N_1650,N_575);
and U3190 (N_3190,N_2494,N_156);
and U3191 (N_3191,N_1392,N_1010);
nand U3192 (N_3192,N_512,N_1352);
nor U3193 (N_3193,N_355,N_270);
nand U3194 (N_3194,N_2276,N_1997);
nand U3195 (N_3195,N_74,N_2170);
nor U3196 (N_3196,N_1174,N_765);
or U3197 (N_3197,N_2346,N_886);
nand U3198 (N_3198,N_2108,N_1670);
xnor U3199 (N_3199,N_1154,N_1899);
nand U3200 (N_3200,N_192,N_1881);
nor U3201 (N_3201,N_755,N_164);
nand U3202 (N_3202,N_2418,N_2380);
nand U3203 (N_3203,N_1411,N_189);
nand U3204 (N_3204,N_2193,N_2004);
nand U3205 (N_3205,N_1674,N_841);
and U3206 (N_3206,N_1869,N_1647);
xor U3207 (N_3207,N_554,N_963);
xnor U3208 (N_3208,N_300,N_223);
or U3209 (N_3209,N_2092,N_940);
or U3210 (N_3210,N_1348,N_1730);
nand U3211 (N_3211,N_490,N_1076);
and U3212 (N_3212,N_1103,N_1405);
nor U3213 (N_3213,N_2029,N_1492);
and U3214 (N_3214,N_694,N_329);
nand U3215 (N_3215,N_2165,N_1842);
or U3216 (N_3216,N_2027,N_2081);
xnor U3217 (N_3217,N_1254,N_94);
and U3218 (N_3218,N_408,N_2308);
or U3219 (N_3219,N_788,N_2114);
nand U3220 (N_3220,N_2210,N_536);
nor U3221 (N_3221,N_1613,N_1687);
xor U3222 (N_3222,N_851,N_2074);
or U3223 (N_3223,N_1677,N_996);
or U3224 (N_3224,N_2012,N_922);
nand U3225 (N_3225,N_2301,N_1622);
and U3226 (N_3226,N_943,N_1229);
or U3227 (N_3227,N_1102,N_1475);
or U3228 (N_3228,N_913,N_2465);
nor U3229 (N_3229,N_809,N_1158);
and U3230 (N_3230,N_1548,N_927);
nand U3231 (N_3231,N_93,N_1100);
or U3232 (N_3232,N_1959,N_2272);
or U3233 (N_3233,N_234,N_898);
and U3234 (N_3234,N_1797,N_447);
nand U3235 (N_3235,N_302,N_1773);
nand U3236 (N_3236,N_634,N_2401);
xor U3237 (N_3237,N_1446,N_1469);
or U3238 (N_3238,N_1258,N_259);
nand U3239 (N_3239,N_760,N_2152);
nor U3240 (N_3240,N_508,N_2054);
nor U3241 (N_3241,N_1150,N_2263);
or U3242 (N_3242,N_280,N_767);
nor U3243 (N_3243,N_1889,N_2064);
or U3244 (N_3244,N_726,N_2111);
nand U3245 (N_3245,N_2065,N_705);
nor U3246 (N_3246,N_397,N_1579);
nor U3247 (N_3247,N_1556,N_2489);
and U3248 (N_3248,N_1341,N_196);
xnor U3249 (N_3249,N_1409,N_1000);
nand U3250 (N_3250,N_377,N_2122);
or U3251 (N_3251,N_933,N_950);
or U3252 (N_3252,N_876,N_1749);
and U3253 (N_3253,N_2447,N_1929);
and U3254 (N_3254,N_2326,N_1819);
and U3255 (N_3255,N_1412,N_774);
nand U3256 (N_3256,N_1398,N_832);
or U3257 (N_3257,N_661,N_1306);
nand U3258 (N_3258,N_1709,N_1148);
nand U3259 (N_3259,N_28,N_2336);
and U3260 (N_3260,N_2475,N_1703);
xnor U3261 (N_3261,N_1241,N_1571);
or U3262 (N_3262,N_2031,N_1155);
and U3263 (N_3263,N_463,N_1025);
nor U3264 (N_3264,N_1424,N_1710);
or U3265 (N_3265,N_1944,N_2415);
or U3266 (N_3266,N_1386,N_462);
and U3267 (N_3267,N_509,N_834);
nor U3268 (N_3268,N_2206,N_1204);
nand U3269 (N_3269,N_1998,N_974);
or U3270 (N_3270,N_2087,N_1696);
nand U3271 (N_3271,N_2369,N_466);
and U3272 (N_3272,N_1222,N_16);
or U3273 (N_3273,N_2322,N_1058);
nor U3274 (N_3274,N_821,N_296);
nand U3275 (N_3275,N_419,N_428);
or U3276 (N_3276,N_1574,N_437);
nor U3277 (N_3277,N_1873,N_1053);
or U3278 (N_3278,N_1268,N_242);
xnor U3279 (N_3279,N_2393,N_2445);
nand U3280 (N_3280,N_550,N_619);
and U3281 (N_3281,N_256,N_2212);
and U3282 (N_3282,N_608,N_1523);
nor U3283 (N_3283,N_1586,N_2345);
nand U3284 (N_3284,N_904,N_1483);
nor U3285 (N_3285,N_787,N_315);
and U3286 (N_3286,N_1259,N_664);
nor U3287 (N_3287,N_2419,N_339);
nor U3288 (N_3288,N_1782,N_1965);
xor U3289 (N_3289,N_2329,N_1851);
or U3290 (N_3290,N_2416,N_1091);
nand U3291 (N_3291,N_431,N_1050);
or U3292 (N_3292,N_1967,N_485);
or U3293 (N_3293,N_2052,N_106);
nor U3294 (N_3294,N_2022,N_367);
or U3295 (N_3295,N_1444,N_131);
or U3296 (N_3296,N_90,N_595);
nand U3297 (N_3297,N_1684,N_644);
and U3298 (N_3298,N_1987,N_2085);
nor U3299 (N_3299,N_665,N_2070);
nor U3300 (N_3300,N_693,N_1862);
nor U3301 (N_3301,N_165,N_744);
nand U3302 (N_3302,N_894,N_580);
nand U3303 (N_3303,N_810,N_233);
nand U3304 (N_3304,N_921,N_1669);
or U3305 (N_3305,N_843,N_1957);
and U3306 (N_3306,N_1396,N_524);
or U3307 (N_3307,N_322,N_145);
nand U3308 (N_3308,N_1700,N_806);
or U3309 (N_3309,N_1561,N_63);
or U3310 (N_3310,N_471,N_1307);
nand U3311 (N_3311,N_712,N_1474);
or U3312 (N_3312,N_1303,N_801);
nand U3313 (N_3313,N_824,N_237);
nor U3314 (N_3314,N_936,N_137);
or U3315 (N_3315,N_2095,N_1774);
nand U3316 (N_3316,N_1109,N_1466);
nor U3317 (N_3317,N_52,N_1752);
and U3318 (N_3318,N_800,N_1127);
nor U3319 (N_3319,N_1910,N_1748);
nand U3320 (N_3320,N_1040,N_1310);
xnor U3321 (N_3321,N_120,N_2466);
nor U3322 (N_3322,N_2459,N_2127);
xor U3323 (N_3323,N_497,N_2185);
nor U3324 (N_3324,N_2390,N_1896);
and U3325 (N_3325,N_2288,N_2463);
nor U3326 (N_3326,N_1186,N_944);
and U3327 (N_3327,N_657,N_486);
nand U3328 (N_3328,N_643,N_114);
nor U3329 (N_3329,N_69,N_2476);
nand U3330 (N_3330,N_1680,N_448);
and U3331 (N_3331,N_2457,N_1496);
nor U3332 (N_3332,N_1238,N_978);
or U3333 (N_3333,N_530,N_1598);
nor U3334 (N_3334,N_1404,N_1593);
nor U3335 (N_3335,N_1614,N_736);
and U3336 (N_3336,N_450,N_2484);
or U3337 (N_3337,N_666,N_771);
nor U3338 (N_3338,N_454,N_1644);
nor U3339 (N_3339,N_117,N_683);
xor U3340 (N_3340,N_457,N_1342);
nand U3341 (N_3341,N_1464,N_1417);
xor U3342 (N_3342,N_718,N_77);
nor U3343 (N_3343,N_1606,N_717);
nand U3344 (N_3344,N_1304,N_1291);
or U3345 (N_3345,N_2339,N_112);
and U3346 (N_3346,N_2157,N_1672);
nor U3347 (N_3347,N_480,N_2044);
nand U3348 (N_3348,N_174,N_1430);
and U3349 (N_3349,N_749,N_4);
and U3350 (N_3350,N_1372,N_245);
nor U3351 (N_3351,N_1924,N_467);
and U3352 (N_3352,N_2236,N_1262);
and U3353 (N_3353,N_1054,N_504);
nor U3354 (N_3354,N_1795,N_732);
xor U3355 (N_3355,N_2448,N_1197);
or U3356 (N_3356,N_2199,N_893);
and U3357 (N_3357,N_2149,N_14);
or U3358 (N_3358,N_920,N_1288);
and U3359 (N_3359,N_1925,N_1378);
xnor U3360 (N_3360,N_881,N_1422);
nor U3361 (N_3361,N_159,N_2178);
and U3362 (N_3362,N_599,N_1055);
and U3363 (N_3363,N_1357,N_1207);
nand U3364 (N_3364,N_1625,N_2137);
and U3365 (N_3365,N_1559,N_830);
or U3366 (N_3366,N_111,N_361);
nor U3367 (N_3367,N_496,N_2105);
nor U3368 (N_3368,N_2277,N_494);
nor U3369 (N_3369,N_1337,N_2488);
nor U3370 (N_3370,N_413,N_2478);
or U3371 (N_3371,N_2405,N_61);
nand U3372 (N_3372,N_1903,N_1848);
nand U3373 (N_3373,N_1859,N_1900);
nand U3374 (N_3374,N_1275,N_1350);
nand U3375 (N_3375,N_1812,N_517);
xor U3376 (N_3376,N_255,N_1977);
nor U3377 (N_3377,N_1367,N_822);
and U3378 (N_3378,N_2442,N_1440);
nand U3379 (N_3379,N_1619,N_1999);
and U3380 (N_3380,N_263,N_975);
or U3381 (N_3381,N_1195,N_84);
nand U3382 (N_3382,N_1329,N_1964);
or U3383 (N_3383,N_1540,N_2090);
and U3384 (N_3384,N_1447,N_1963);
nand U3385 (N_3385,N_219,N_1201);
and U3386 (N_3386,N_2038,N_2266);
and U3387 (N_3387,N_2069,N_1558);
nor U3388 (N_3388,N_2189,N_2275);
and U3389 (N_3389,N_326,N_761);
nor U3390 (N_3390,N_2375,N_1005);
nand U3391 (N_3391,N_2417,N_667);
and U3392 (N_3392,N_867,N_1546);
or U3393 (N_3393,N_869,N_1628);
or U3394 (N_3394,N_319,N_1826);
nor U3395 (N_3395,N_1252,N_663);
or U3396 (N_3396,N_209,N_2250);
and U3397 (N_3397,N_1532,N_11);
nor U3398 (N_3398,N_2262,N_1992);
nand U3399 (N_3399,N_1575,N_1518);
nor U3400 (N_3400,N_1567,N_1609);
nor U3401 (N_3401,N_814,N_301);
or U3402 (N_3402,N_1717,N_321);
and U3403 (N_3403,N_670,N_362);
xnor U3404 (N_3404,N_911,N_2227);
or U3405 (N_3405,N_775,N_1688);
and U3406 (N_3406,N_55,N_40);
and U3407 (N_3407,N_581,N_135);
nor U3408 (N_3408,N_460,N_1956);
xor U3409 (N_3409,N_2134,N_1801);
or U3410 (N_3410,N_2472,N_1449);
nor U3411 (N_3411,N_2174,N_720);
nand U3412 (N_3412,N_1568,N_354);
nor U3413 (N_3413,N_1958,N_441);
and U3414 (N_3414,N_2297,N_1257);
xor U3415 (N_3415,N_1727,N_999);
and U3416 (N_3416,N_2033,N_1321);
or U3417 (N_3417,N_2349,N_127);
and U3418 (N_3418,N_445,N_1093);
nand U3419 (N_3419,N_1294,N_1395);
and U3420 (N_3420,N_1512,N_312);
or U3421 (N_3421,N_2286,N_1860);
nor U3422 (N_3422,N_954,N_1212);
and U3423 (N_3423,N_2385,N_1733);
or U3424 (N_3424,N_1832,N_1885);
nor U3425 (N_3425,N_389,N_231);
or U3426 (N_3426,N_235,N_1104);
nor U3427 (N_3427,N_1017,N_2399);
or U3428 (N_3428,N_423,N_1272);
nand U3429 (N_3429,N_2437,N_279);
nor U3430 (N_3430,N_107,N_1880);
and U3431 (N_3431,N_680,N_1877);
nor U3432 (N_3432,N_13,N_1804);
or U3433 (N_3433,N_1339,N_1587);
nor U3434 (N_3434,N_434,N_1569);
nor U3435 (N_3435,N_2207,N_1682);
nor U3436 (N_3436,N_2144,N_1366);
or U3437 (N_3437,N_1784,N_2215);
or U3438 (N_3438,N_1883,N_945);
and U3439 (N_3439,N_1221,N_290);
or U3440 (N_3440,N_42,N_1485);
xor U3441 (N_3441,N_1526,N_1320);
nor U3442 (N_3442,N_1660,N_1961);
and U3443 (N_3443,N_882,N_412);
or U3444 (N_3444,N_1803,N_794);
and U3445 (N_3445,N_110,N_306);
nor U3446 (N_3446,N_1734,N_1627);
or U3447 (N_3447,N_1704,N_96);
or U3448 (N_3448,N_2084,N_1581);
nor U3449 (N_3449,N_158,N_1759);
nor U3450 (N_3450,N_1818,N_2289);
xnor U3451 (N_3451,N_215,N_914);
and U3452 (N_3452,N_407,N_1636);
nor U3453 (N_3453,N_203,N_1260);
and U3454 (N_3454,N_754,N_689);
nor U3455 (N_3455,N_1722,N_2371);
xnor U3456 (N_3456,N_388,N_1936);
nand U3457 (N_3457,N_1867,N_416);
and U3458 (N_3458,N_1436,N_1948);
nor U3459 (N_3459,N_2180,N_1332);
and U3460 (N_3460,N_6,N_557);
and U3461 (N_3461,N_50,N_1336);
and U3462 (N_3462,N_1051,N_2017);
xor U3463 (N_3463,N_2314,N_1490);
nor U3464 (N_3464,N_1227,N_566);
nor U3465 (N_3465,N_1653,N_1024);
xnor U3466 (N_3466,N_989,N_1096);
and U3467 (N_3467,N_2450,N_837);
nand U3468 (N_3468,N_2353,N_1435);
and U3469 (N_3469,N_835,N_1046);
and U3470 (N_3470,N_1600,N_523);
xor U3471 (N_3471,N_147,N_2244);
nor U3472 (N_3472,N_802,N_1960);
nand U3473 (N_3473,N_2441,N_66);
or U3474 (N_3474,N_53,N_1891);
nor U3475 (N_3475,N_711,N_1209);
nand U3476 (N_3476,N_1917,N_2041);
and U3477 (N_3477,N_1513,N_1790);
and U3478 (N_3478,N_2123,N_2103);
nor U3479 (N_3479,N_335,N_1331);
and U3480 (N_3480,N_1183,N_1413);
or U3481 (N_3481,N_1562,N_1690);
nor U3482 (N_3482,N_1632,N_1382);
nand U3483 (N_3483,N_432,N_384);
and U3484 (N_3484,N_67,N_574);
xor U3485 (N_3485,N_1758,N_1985);
and U3486 (N_3486,N_1244,N_226);
nand U3487 (N_3487,N_1792,N_1123);
or U3488 (N_3488,N_808,N_1507);
nand U3489 (N_3489,N_1420,N_2175);
or U3490 (N_3490,N_1767,N_2147);
or U3491 (N_3491,N_1460,N_879);
and U3492 (N_3492,N_1293,N_1705);
nand U3493 (N_3493,N_1980,N_2358);
nand U3494 (N_3494,N_532,N_2337);
nor U3495 (N_3495,N_572,N_2320);
xor U3496 (N_3496,N_848,N_128);
or U3497 (N_3497,N_1038,N_1714);
nand U3498 (N_3498,N_356,N_576);
nand U3499 (N_3499,N_2014,N_374);
nand U3500 (N_3500,N_1179,N_1519);
nor U3501 (N_3501,N_990,N_863);
nand U3502 (N_3502,N_337,N_2171);
and U3503 (N_3503,N_1514,N_2317);
nand U3504 (N_3504,N_1338,N_1972);
xor U3505 (N_3505,N_2480,N_1901);
nor U3506 (N_3506,N_949,N_269);
xnor U3507 (N_3507,N_1895,N_1735);
or U3508 (N_3508,N_969,N_840);
nand U3509 (N_3509,N_2020,N_1623);
nand U3510 (N_3510,N_2200,N_1487);
and U3511 (N_3511,N_281,N_1445);
nor U3512 (N_3512,N_2226,N_1101);
or U3513 (N_3513,N_917,N_995);
nand U3514 (N_3514,N_1649,N_1472);
or U3515 (N_3515,N_1582,N_1855);
xor U3516 (N_3516,N_1107,N_958);
nand U3517 (N_3517,N_986,N_443);
xnor U3518 (N_3518,N_2233,N_489);
and U3519 (N_3519,N_1245,N_1119);
or U3520 (N_3520,N_2088,N_1425);
or U3521 (N_3521,N_2141,N_23);
nand U3522 (N_3522,N_1506,N_1253);
and U3523 (N_3523,N_1421,N_1057);
or U3524 (N_3524,N_1837,N_1309);
nor U3525 (N_3525,N_1661,N_1638);
and U3526 (N_3526,N_1720,N_934);
or U3527 (N_3527,N_780,N_1527);
and U3528 (N_3528,N_344,N_565);
or U3529 (N_3529,N_1509,N_1399);
or U3530 (N_3530,N_769,N_214);
nor U3531 (N_3531,N_616,N_240);
xor U3532 (N_3532,N_126,N_153);
xnor U3533 (N_3533,N_1432,N_1919);
nor U3534 (N_3534,N_1442,N_2256);
or U3535 (N_3535,N_2172,N_1426);
or U3536 (N_3536,N_1255,N_2497);
nand U3537 (N_3537,N_2485,N_1902);
nand U3538 (N_3538,N_2261,N_561);
and U3539 (N_3539,N_1090,N_1488);
or U3540 (N_3540,N_2312,N_539);
nor U3541 (N_3541,N_2260,N_119);
and U3542 (N_3542,N_2335,N_1981);
and U3543 (N_3543,N_1219,N_1189);
and U3544 (N_3544,N_2278,N_227);
xnor U3545 (N_3545,N_652,N_2363);
and U3546 (N_3546,N_1008,N_1708);
xnor U3547 (N_3547,N_1750,N_1196);
nand U3548 (N_3548,N_2492,N_1563);
or U3549 (N_3549,N_1387,N_395);
or U3550 (N_3550,N_543,N_1457);
and U3551 (N_3551,N_1164,N_2099);
xor U3552 (N_3552,N_2431,N_2242);
and U3553 (N_3553,N_2408,N_751);
nor U3554 (N_3554,N_1596,N_2028);
nand U3555 (N_3555,N_373,N_32);
nor U3556 (N_3556,N_558,N_341);
nand U3557 (N_3557,N_2007,N_2362);
or U3558 (N_3558,N_1168,N_1315);
xnor U3559 (N_3559,N_923,N_1681);
nor U3560 (N_3560,N_1675,N_2370);
nand U3561 (N_3561,N_816,N_1595);
or U3562 (N_3562,N_1231,N_1603);
nor U3563 (N_3563,N_1217,N_1181);
or U3564 (N_3564,N_1652,N_394);
and U3565 (N_3565,N_2040,N_1097);
and U3566 (N_3566,N_1415,N_908);
or U3567 (N_3567,N_1135,N_947);
and U3568 (N_3568,N_1388,N_1941);
nor U3569 (N_3569,N_199,N_417);
nor U3570 (N_3570,N_409,N_1712);
or U3571 (N_3571,N_2166,N_1668);
or U3572 (N_3572,N_857,N_1676);
nor U3573 (N_3573,N_1068,N_1993);
and U3574 (N_3574,N_2125,N_1236);
and U3575 (N_3575,N_1380,N_151);
xnor U3576 (N_3576,N_1663,N_1893);
and U3577 (N_3577,N_692,N_2453);
nor U3578 (N_3578,N_1482,N_1920);
nand U3579 (N_3579,N_679,N_1646);
nor U3580 (N_3580,N_1833,N_1083);
nand U3581 (N_3581,N_1389,N_1467);
xnor U3582 (N_3582,N_513,N_1585);
nor U3583 (N_3583,N_2101,N_1761);
or U3584 (N_3584,N_183,N_1277);
nand U3585 (N_3585,N_2328,N_642);
nand U3586 (N_3586,N_1082,N_626);
nand U3587 (N_3587,N_1079,N_609);
or U3588 (N_3588,N_2373,N_1979);
or U3589 (N_3589,N_603,N_1175);
nand U3590 (N_3590,N_1864,N_1535);
or U3591 (N_3591,N_1856,N_1701);
nor U3592 (N_3592,N_1810,N_1028);
nor U3593 (N_3593,N_2079,N_885);
nand U3594 (N_3594,N_2282,N_1590);
nand U3595 (N_3595,N_1290,N_706);
or U3596 (N_3596,N_1870,N_2359);
nand U3597 (N_3597,N_1528,N_1370);
or U3598 (N_3598,N_721,N_589);
nor U3599 (N_3599,N_348,N_631);
or U3600 (N_3600,N_796,N_229);
and U3601 (N_3601,N_658,N_1210);
and U3602 (N_3602,N_410,N_763);
or U3603 (N_3603,N_1052,N_1737);
or U3604 (N_3604,N_2024,N_614);
and U3605 (N_3605,N_2313,N_1125);
or U3606 (N_3606,N_1355,N_2467);
or U3607 (N_3607,N_1927,N_88);
nor U3608 (N_3608,N_2187,N_889);
nand U3609 (N_3609,N_2237,N_2133);
and U3610 (N_3610,N_779,N_71);
xnor U3611 (N_3611,N_291,N_1400);
nand U3612 (N_3612,N_1970,N_1521);
and U3613 (N_3613,N_1770,N_734);
or U3614 (N_3614,N_1403,N_375);
or U3615 (N_3615,N_2449,N_541);
nor U3616 (N_3616,N_2410,N_1084);
nand U3617 (N_3617,N_273,N_134);
and U3618 (N_3618,N_560,N_275);
and U3619 (N_3619,N_1583,N_2194);
nor U3620 (N_3620,N_795,N_244);
xnor U3621 (N_3621,N_472,N_515);
nand U3622 (N_3622,N_1477,N_2477);
or U3623 (N_3623,N_1962,N_268);
or U3624 (N_3624,N_833,N_2461);
or U3625 (N_3625,N_2333,N_1171);
nand U3626 (N_3626,N_1732,N_994);
or U3627 (N_3627,N_939,N_811);
nand U3628 (N_3628,N_2182,N_1061);
nand U3629 (N_3629,N_345,N_1637);
and U3630 (N_3630,N_2039,N_1615);
nor U3631 (N_3631,N_961,N_138);
or U3632 (N_3632,N_2181,N_762);
nor U3633 (N_3633,N_725,N_452);
and U3634 (N_3634,N_1461,N_121);
and U3635 (N_3635,N_36,N_2387);
nor U3636 (N_3636,N_1995,N_1041);
or U3637 (N_3637,N_1515,N_2432);
or U3638 (N_3638,N_2089,N_446);
or U3639 (N_3639,N_1144,N_1825);
and U3640 (N_3640,N_1283,N_1453);
xnor U3641 (N_3641,N_789,N_282);
nor U3642 (N_3642,N_2251,N_2291);
nor U3643 (N_3643,N_932,N_1067);
and U3644 (N_3644,N_2002,N_369);
or U3645 (N_3645,N_2283,N_1657);
nor U3646 (N_3646,N_1777,N_92);
nand U3647 (N_3647,N_1318,N_1932);
nand U3648 (N_3648,N_2376,N_18);
nor U3649 (N_3649,N_82,N_2106);
or U3650 (N_3650,N_1256,N_22);
or U3651 (N_3651,N_1589,N_283);
or U3652 (N_3652,N_1263,N_1385);
nor U3653 (N_3653,N_604,N_792);
xnor U3654 (N_3654,N_1344,N_2115);
or U3655 (N_3655,N_1237,N_798);
nor U3656 (N_3656,N_476,N_1121);
nor U3657 (N_3657,N_2386,N_449);
nand U3658 (N_3658,N_1545,N_805);
nor U3659 (N_3659,N_1769,N_1340);
and U3660 (N_3660,N_1836,N_909);
xnor U3661 (N_3661,N_1194,N_1662);
nor U3662 (N_3662,N_2229,N_1120);
and U3663 (N_3663,N_481,N_129);
or U3664 (N_3664,N_764,N_1213);
nor U3665 (N_3665,N_1381,N_141);
nor U3666 (N_3666,N_1042,N_1835);
nor U3667 (N_3667,N_1738,N_2347);
nand U3668 (N_3668,N_791,N_553);
nand U3669 (N_3669,N_538,N_1658);
nand U3670 (N_3670,N_1664,N_2252);
nor U3671 (N_3671,N_1794,N_1655);
or U3672 (N_3672,N_528,N_691);
and U3673 (N_3673,N_548,N_1991);
nand U3674 (N_3674,N_1607,N_1074);
and U3675 (N_3675,N_2455,N_1882);
nor U3676 (N_3676,N_549,N_459);
nor U3677 (N_3677,N_556,N_1007);
nor U3678 (N_3678,N_1702,N_422);
nand U3679 (N_3679,N_1161,N_1459);
xor U3680 (N_3680,N_1505,N_1641);
nand U3681 (N_3681,N_552,N_17);
nand U3682 (N_3682,N_2117,N_1056);
and U3683 (N_3683,N_586,N_888);
or U3684 (N_3684,N_1071,N_856);
nand U3685 (N_3685,N_2351,N_937);
nand U3686 (N_3686,N_1178,N_849);
and U3687 (N_3687,N_2254,N_2355);
and U3688 (N_3688,N_2231,N_1012);
or U3689 (N_3689,N_2360,N_424);
xor U3690 (N_3690,N_1314,N_1533);
and U3691 (N_3691,N_1621,N_208);
nand U3692 (N_3692,N_1234,N_531);
nor U3693 (N_3693,N_1823,N_2035);
nand U3694 (N_3694,N_2354,N_25);
nor U3695 (N_3695,N_1166,N_2381);
nand U3696 (N_3696,N_1849,N_1694);
and U3697 (N_3697,N_1138,N_1996);
nand U3698 (N_3698,N_918,N_770);
and U3699 (N_3699,N_2120,N_1788);
nor U3700 (N_3700,N_2271,N_258);
and U3701 (N_3701,N_1267,N_2208);
and U3702 (N_3702,N_182,N_758);
or U3703 (N_3703,N_656,N_710);
or U3704 (N_3704,N_624,N_2160);
or U3705 (N_3705,N_1098,N_1634);
or U3706 (N_3706,N_1935,N_286);
nor U3707 (N_3707,N_1191,N_1313);
and U3708 (N_3708,N_207,N_1764);
or U3709 (N_3709,N_1516,N_930);
nor U3710 (N_3710,N_1578,N_2241);
nand U3711 (N_3711,N_2273,N_1092);
nor U3712 (N_3712,N_757,N_1954);
nand U3713 (N_3713,N_91,N_83);
and U3714 (N_3714,N_160,N_1503);
nand U3715 (N_3715,N_1305,N_1193);
or U3716 (N_3716,N_1673,N_2403);
and U3717 (N_3717,N_776,N_488);
nor U3718 (N_3718,N_368,N_2400);
and U3719 (N_3719,N_1947,N_2396);
and U3720 (N_3720,N_2470,N_1433);
and U3721 (N_3721,N_503,N_2209);
xor U3722 (N_3722,N_2008,N_49);
or U3723 (N_3723,N_1775,N_2216);
or U3724 (N_3724,N_484,N_2304);
and U3725 (N_3725,N_1289,N_289);
nand U3726 (N_3726,N_173,N_2159);
xor U3727 (N_3727,N_1952,N_2214);
nor U3728 (N_3728,N_722,N_2299);
nor U3729 (N_3729,N_873,N_1809);
nor U3730 (N_3730,N_316,N_2464);
or U3731 (N_3731,N_1001,N_2168);
and U3732 (N_3732,N_916,N_482);
nand U3733 (N_3733,N_1778,N_124);
xnor U3734 (N_3734,N_1406,N_2409);
xnor U3735 (N_3735,N_1839,N_185);
or U3736 (N_3736,N_1541,N_313);
nand U3737 (N_3737,N_1214,N_2055);
nand U3738 (N_3738,N_1654,N_1408);
or U3739 (N_3739,N_1391,N_350);
nand U3740 (N_3740,N_1577,N_1030);
nor U3741 (N_3741,N_210,N_1852);
and U3742 (N_3742,N_342,N_1147);
and U3743 (N_3743,N_852,N_584);
nand U3744 (N_3744,N_741,N_1923);
nor U3745 (N_3745,N_1376,N_1906);
nor U3746 (N_3746,N_304,N_1633);
xnor U3747 (N_3747,N_1062,N_695);
and U3748 (N_3748,N_2150,N_1278);
or U3749 (N_3749,N_935,N_902);
or U3750 (N_3750,N_1316,N_1884);
or U3751 (N_3751,N_1173,N_455);
and U3752 (N_3752,N_458,N_193);
nand U3753 (N_3753,N_2157,N_1691);
nand U3754 (N_3754,N_1407,N_5);
or U3755 (N_3755,N_796,N_2033);
nand U3756 (N_3756,N_1436,N_2069);
nor U3757 (N_3757,N_2212,N_1339);
nand U3758 (N_3758,N_633,N_1199);
and U3759 (N_3759,N_589,N_1304);
nor U3760 (N_3760,N_1810,N_305);
nor U3761 (N_3761,N_509,N_2332);
and U3762 (N_3762,N_1317,N_1613);
nand U3763 (N_3763,N_1182,N_635);
nor U3764 (N_3764,N_2036,N_906);
xnor U3765 (N_3765,N_325,N_50);
nand U3766 (N_3766,N_2150,N_906);
nand U3767 (N_3767,N_2132,N_1739);
or U3768 (N_3768,N_1296,N_1345);
xor U3769 (N_3769,N_192,N_2085);
xnor U3770 (N_3770,N_773,N_2111);
nand U3771 (N_3771,N_2329,N_722);
nor U3772 (N_3772,N_222,N_10);
or U3773 (N_3773,N_189,N_1788);
xor U3774 (N_3774,N_432,N_1027);
nand U3775 (N_3775,N_334,N_302);
or U3776 (N_3776,N_1942,N_1404);
nand U3777 (N_3777,N_1602,N_1121);
nand U3778 (N_3778,N_2441,N_806);
or U3779 (N_3779,N_1194,N_1158);
nor U3780 (N_3780,N_1124,N_384);
nand U3781 (N_3781,N_1755,N_356);
xor U3782 (N_3782,N_1986,N_819);
and U3783 (N_3783,N_2015,N_1591);
or U3784 (N_3784,N_831,N_539);
or U3785 (N_3785,N_2151,N_1991);
nor U3786 (N_3786,N_1823,N_1555);
and U3787 (N_3787,N_2396,N_1332);
nand U3788 (N_3788,N_867,N_1493);
nand U3789 (N_3789,N_2186,N_1592);
nor U3790 (N_3790,N_2105,N_432);
or U3791 (N_3791,N_1528,N_1029);
and U3792 (N_3792,N_565,N_131);
nor U3793 (N_3793,N_2201,N_1654);
and U3794 (N_3794,N_2,N_1207);
nand U3795 (N_3795,N_1060,N_601);
or U3796 (N_3796,N_1755,N_403);
or U3797 (N_3797,N_1996,N_105);
nor U3798 (N_3798,N_799,N_2209);
and U3799 (N_3799,N_770,N_1114);
nor U3800 (N_3800,N_221,N_374);
nand U3801 (N_3801,N_570,N_2197);
nor U3802 (N_3802,N_2409,N_2207);
and U3803 (N_3803,N_992,N_1320);
nor U3804 (N_3804,N_1364,N_224);
nor U3805 (N_3805,N_65,N_1910);
or U3806 (N_3806,N_1452,N_1287);
and U3807 (N_3807,N_1319,N_961);
or U3808 (N_3808,N_1944,N_1253);
xor U3809 (N_3809,N_2476,N_372);
nand U3810 (N_3810,N_995,N_2304);
nand U3811 (N_3811,N_1297,N_917);
or U3812 (N_3812,N_958,N_1681);
nor U3813 (N_3813,N_565,N_1652);
nand U3814 (N_3814,N_1099,N_2467);
xor U3815 (N_3815,N_1901,N_1540);
and U3816 (N_3816,N_969,N_1649);
nor U3817 (N_3817,N_1976,N_2186);
and U3818 (N_3818,N_1455,N_1083);
or U3819 (N_3819,N_185,N_114);
and U3820 (N_3820,N_1413,N_2118);
nand U3821 (N_3821,N_2422,N_2341);
or U3822 (N_3822,N_2116,N_1542);
nand U3823 (N_3823,N_451,N_1317);
xnor U3824 (N_3824,N_1089,N_2478);
or U3825 (N_3825,N_1787,N_2082);
or U3826 (N_3826,N_414,N_1848);
xor U3827 (N_3827,N_541,N_2471);
nand U3828 (N_3828,N_1815,N_1179);
xnor U3829 (N_3829,N_1977,N_1941);
or U3830 (N_3830,N_1995,N_2163);
nand U3831 (N_3831,N_2029,N_727);
or U3832 (N_3832,N_1636,N_49);
xor U3833 (N_3833,N_1939,N_2071);
or U3834 (N_3834,N_2493,N_1077);
nand U3835 (N_3835,N_1271,N_1825);
and U3836 (N_3836,N_1880,N_2098);
nand U3837 (N_3837,N_2037,N_2401);
nor U3838 (N_3838,N_920,N_2232);
and U3839 (N_3839,N_954,N_640);
nor U3840 (N_3840,N_170,N_1128);
and U3841 (N_3841,N_1285,N_35);
and U3842 (N_3842,N_707,N_569);
or U3843 (N_3843,N_2374,N_1193);
nor U3844 (N_3844,N_316,N_1913);
nor U3845 (N_3845,N_1202,N_1130);
and U3846 (N_3846,N_1835,N_1631);
nor U3847 (N_3847,N_1977,N_1049);
or U3848 (N_3848,N_2128,N_1629);
and U3849 (N_3849,N_1435,N_26);
or U3850 (N_3850,N_613,N_2429);
nor U3851 (N_3851,N_231,N_529);
or U3852 (N_3852,N_1921,N_1808);
or U3853 (N_3853,N_1677,N_713);
or U3854 (N_3854,N_988,N_53);
and U3855 (N_3855,N_129,N_398);
nand U3856 (N_3856,N_273,N_1486);
or U3857 (N_3857,N_1146,N_812);
and U3858 (N_3858,N_404,N_2226);
or U3859 (N_3859,N_784,N_1140);
and U3860 (N_3860,N_384,N_126);
or U3861 (N_3861,N_564,N_685);
nand U3862 (N_3862,N_2389,N_1040);
or U3863 (N_3863,N_933,N_1141);
xor U3864 (N_3864,N_2031,N_2499);
nand U3865 (N_3865,N_1559,N_207);
and U3866 (N_3866,N_2492,N_641);
nand U3867 (N_3867,N_1371,N_716);
and U3868 (N_3868,N_270,N_2169);
or U3869 (N_3869,N_2165,N_1496);
nor U3870 (N_3870,N_303,N_2387);
or U3871 (N_3871,N_2479,N_478);
or U3872 (N_3872,N_2287,N_1937);
or U3873 (N_3873,N_2253,N_1060);
nor U3874 (N_3874,N_58,N_2358);
and U3875 (N_3875,N_353,N_2200);
or U3876 (N_3876,N_1092,N_752);
nor U3877 (N_3877,N_98,N_880);
nor U3878 (N_3878,N_550,N_1213);
nor U3879 (N_3879,N_2467,N_1657);
xor U3880 (N_3880,N_962,N_845);
nor U3881 (N_3881,N_1826,N_139);
and U3882 (N_3882,N_2134,N_461);
nand U3883 (N_3883,N_2463,N_137);
nor U3884 (N_3884,N_1385,N_1812);
nand U3885 (N_3885,N_798,N_686);
nor U3886 (N_3886,N_1820,N_1979);
or U3887 (N_3887,N_1112,N_1058);
or U3888 (N_3888,N_2223,N_2283);
or U3889 (N_3889,N_1694,N_1424);
nor U3890 (N_3890,N_486,N_1897);
xor U3891 (N_3891,N_2099,N_1167);
and U3892 (N_3892,N_2439,N_575);
and U3893 (N_3893,N_1109,N_2487);
xnor U3894 (N_3894,N_394,N_1193);
or U3895 (N_3895,N_2312,N_2417);
or U3896 (N_3896,N_321,N_1636);
nor U3897 (N_3897,N_1607,N_1446);
xor U3898 (N_3898,N_1370,N_696);
and U3899 (N_3899,N_1936,N_150);
or U3900 (N_3900,N_598,N_2485);
nand U3901 (N_3901,N_292,N_580);
nor U3902 (N_3902,N_882,N_1588);
or U3903 (N_3903,N_1655,N_756);
or U3904 (N_3904,N_468,N_574);
nand U3905 (N_3905,N_719,N_2454);
or U3906 (N_3906,N_2379,N_1564);
and U3907 (N_3907,N_880,N_1301);
nand U3908 (N_3908,N_1067,N_1059);
or U3909 (N_3909,N_2280,N_1170);
or U3910 (N_3910,N_290,N_1921);
nor U3911 (N_3911,N_1595,N_2434);
xor U3912 (N_3912,N_1221,N_1148);
nor U3913 (N_3913,N_221,N_1447);
or U3914 (N_3914,N_172,N_1722);
nand U3915 (N_3915,N_509,N_581);
xor U3916 (N_3916,N_181,N_1100);
or U3917 (N_3917,N_590,N_945);
xor U3918 (N_3918,N_158,N_443);
nor U3919 (N_3919,N_2450,N_2050);
xnor U3920 (N_3920,N_2251,N_816);
nor U3921 (N_3921,N_1481,N_2328);
or U3922 (N_3922,N_811,N_2372);
or U3923 (N_3923,N_1976,N_1639);
nand U3924 (N_3924,N_1488,N_1697);
or U3925 (N_3925,N_1792,N_1587);
nor U3926 (N_3926,N_2355,N_1623);
nor U3927 (N_3927,N_300,N_2254);
nor U3928 (N_3928,N_2029,N_477);
nor U3929 (N_3929,N_1018,N_473);
nand U3930 (N_3930,N_820,N_1565);
nor U3931 (N_3931,N_633,N_768);
nor U3932 (N_3932,N_1248,N_2211);
nor U3933 (N_3933,N_1730,N_908);
nand U3934 (N_3934,N_1318,N_1902);
and U3935 (N_3935,N_135,N_388);
or U3936 (N_3936,N_5,N_485);
or U3937 (N_3937,N_1298,N_2130);
or U3938 (N_3938,N_693,N_283);
or U3939 (N_3939,N_1209,N_2234);
and U3940 (N_3940,N_2495,N_274);
or U3941 (N_3941,N_1163,N_574);
and U3942 (N_3942,N_1757,N_500);
or U3943 (N_3943,N_72,N_2296);
and U3944 (N_3944,N_714,N_1363);
and U3945 (N_3945,N_2092,N_415);
nand U3946 (N_3946,N_136,N_1462);
nand U3947 (N_3947,N_324,N_1007);
xor U3948 (N_3948,N_147,N_23);
and U3949 (N_3949,N_980,N_847);
nand U3950 (N_3950,N_1291,N_1870);
or U3951 (N_3951,N_1838,N_1199);
and U3952 (N_3952,N_547,N_2410);
nor U3953 (N_3953,N_644,N_847);
nand U3954 (N_3954,N_2097,N_898);
nand U3955 (N_3955,N_1446,N_1977);
and U3956 (N_3956,N_753,N_1429);
or U3957 (N_3957,N_2302,N_158);
or U3958 (N_3958,N_1254,N_856);
nor U3959 (N_3959,N_848,N_1014);
nor U3960 (N_3960,N_2078,N_1702);
nor U3961 (N_3961,N_2489,N_1603);
and U3962 (N_3962,N_1348,N_394);
nand U3963 (N_3963,N_529,N_552);
nand U3964 (N_3964,N_561,N_1032);
or U3965 (N_3965,N_208,N_1107);
nor U3966 (N_3966,N_538,N_675);
nand U3967 (N_3967,N_1606,N_72);
nor U3968 (N_3968,N_1746,N_144);
nand U3969 (N_3969,N_938,N_1254);
nand U3970 (N_3970,N_44,N_2133);
nand U3971 (N_3971,N_1928,N_1884);
and U3972 (N_3972,N_13,N_2059);
xor U3973 (N_3973,N_554,N_1318);
nor U3974 (N_3974,N_1639,N_1814);
or U3975 (N_3975,N_1660,N_1747);
xnor U3976 (N_3976,N_162,N_1274);
xnor U3977 (N_3977,N_2383,N_25);
nand U3978 (N_3978,N_1644,N_1853);
nor U3979 (N_3979,N_2252,N_80);
nor U3980 (N_3980,N_804,N_2030);
xor U3981 (N_3981,N_1399,N_1013);
and U3982 (N_3982,N_2341,N_628);
xnor U3983 (N_3983,N_456,N_10);
nand U3984 (N_3984,N_173,N_1913);
or U3985 (N_3985,N_1316,N_2389);
nand U3986 (N_3986,N_72,N_2136);
or U3987 (N_3987,N_2259,N_2044);
nor U3988 (N_3988,N_1693,N_2225);
or U3989 (N_3989,N_2204,N_900);
or U3990 (N_3990,N_1651,N_1516);
or U3991 (N_3991,N_696,N_1293);
or U3992 (N_3992,N_49,N_208);
and U3993 (N_3993,N_1672,N_1976);
nand U3994 (N_3994,N_1970,N_1374);
or U3995 (N_3995,N_2112,N_2193);
nand U3996 (N_3996,N_335,N_942);
and U3997 (N_3997,N_1318,N_481);
and U3998 (N_3998,N_36,N_453);
nor U3999 (N_3999,N_1333,N_1378);
nand U4000 (N_4000,N_1982,N_1089);
nor U4001 (N_4001,N_1390,N_1835);
or U4002 (N_4002,N_64,N_1283);
xnor U4003 (N_4003,N_720,N_2490);
xor U4004 (N_4004,N_480,N_128);
xnor U4005 (N_4005,N_1074,N_1441);
nor U4006 (N_4006,N_471,N_51);
nor U4007 (N_4007,N_2432,N_1943);
or U4008 (N_4008,N_96,N_63);
nor U4009 (N_4009,N_1691,N_1696);
or U4010 (N_4010,N_2252,N_1422);
and U4011 (N_4011,N_276,N_144);
or U4012 (N_4012,N_758,N_1883);
nor U4013 (N_4013,N_985,N_960);
xnor U4014 (N_4014,N_2245,N_1925);
and U4015 (N_4015,N_419,N_1837);
nor U4016 (N_4016,N_2381,N_885);
and U4017 (N_4017,N_347,N_2409);
nand U4018 (N_4018,N_2148,N_768);
or U4019 (N_4019,N_828,N_1547);
and U4020 (N_4020,N_2292,N_729);
nand U4021 (N_4021,N_1544,N_1002);
xor U4022 (N_4022,N_2211,N_949);
and U4023 (N_4023,N_1997,N_1888);
nand U4024 (N_4024,N_2134,N_151);
nor U4025 (N_4025,N_588,N_239);
or U4026 (N_4026,N_1358,N_2001);
or U4027 (N_4027,N_2171,N_1);
and U4028 (N_4028,N_1000,N_1869);
nand U4029 (N_4029,N_303,N_636);
nor U4030 (N_4030,N_433,N_1559);
or U4031 (N_4031,N_2162,N_954);
and U4032 (N_4032,N_1766,N_2456);
nor U4033 (N_4033,N_2455,N_444);
nand U4034 (N_4034,N_1672,N_1153);
and U4035 (N_4035,N_1518,N_831);
and U4036 (N_4036,N_539,N_369);
or U4037 (N_4037,N_1568,N_1658);
nor U4038 (N_4038,N_650,N_206);
or U4039 (N_4039,N_527,N_116);
xor U4040 (N_4040,N_2259,N_2267);
nor U4041 (N_4041,N_628,N_2251);
or U4042 (N_4042,N_584,N_573);
or U4043 (N_4043,N_1859,N_21);
nand U4044 (N_4044,N_1159,N_178);
and U4045 (N_4045,N_1074,N_2007);
nor U4046 (N_4046,N_2366,N_663);
nor U4047 (N_4047,N_2184,N_1645);
nand U4048 (N_4048,N_2451,N_1515);
nand U4049 (N_4049,N_1851,N_2173);
or U4050 (N_4050,N_508,N_1294);
and U4051 (N_4051,N_2059,N_2047);
and U4052 (N_4052,N_1896,N_2467);
and U4053 (N_4053,N_652,N_937);
nand U4054 (N_4054,N_1057,N_1996);
and U4055 (N_4055,N_1595,N_447);
nor U4056 (N_4056,N_50,N_2401);
or U4057 (N_4057,N_1910,N_1141);
or U4058 (N_4058,N_8,N_1923);
and U4059 (N_4059,N_2105,N_1534);
or U4060 (N_4060,N_619,N_1142);
nor U4061 (N_4061,N_771,N_511);
or U4062 (N_4062,N_1963,N_867);
nor U4063 (N_4063,N_698,N_2328);
xnor U4064 (N_4064,N_352,N_415);
nor U4065 (N_4065,N_2370,N_2385);
xnor U4066 (N_4066,N_1280,N_2113);
and U4067 (N_4067,N_239,N_1526);
and U4068 (N_4068,N_2222,N_683);
or U4069 (N_4069,N_132,N_2346);
and U4070 (N_4070,N_1737,N_1772);
nor U4071 (N_4071,N_2043,N_361);
and U4072 (N_4072,N_1081,N_95);
nor U4073 (N_4073,N_327,N_2186);
or U4074 (N_4074,N_2251,N_1470);
nand U4075 (N_4075,N_1654,N_2198);
nor U4076 (N_4076,N_1757,N_617);
and U4077 (N_4077,N_1065,N_1090);
nand U4078 (N_4078,N_786,N_602);
nor U4079 (N_4079,N_1479,N_2028);
nor U4080 (N_4080,N_983,N_1679);
nor U4081 (N_4081,N_386,N_762);
nand U4082 (N_4082,N_1762,N_141);
and U4083 (N_4083,N_392,N_1363);
nor U4084 (N_4084,N_137,N_2016);
and U4085 (N_4085,N_2151,N_2141);
nand U4086 (N_4086,N_1121,N_2093);
or U4087 (N_4087,N_1484,N_286);
nor U4088 (N_4088,N_2116,N_1727);
or U4089 (N_4089,N_1549,N_871);
xor U4090 (N_4090,N_2027,N_978);
or U4091 (N_4091,N_2363,N_650);
nand U4092 (N_4092,N_1277,N_413);
nand U4093 (N_4093,N_1564,N_156);
or U4094 (N_4094,N_442,N_2312);
and U4095 (N_4095,N_87,N_1696);
nor U4096 (N_4096,N_2472,N_1845);
or U4097 (N_4097,N_793,N_2419);
nor U4098 (N_4098,N_871,N_1982);
nor U4099 (N_4099,N_1823,N_46);
or U4100 (N_4100,N_1777,N_1613);
and U4101 (N_4101,N_1827,N_1948);
and U4102 (N_4102,N_1064,N_1058);
xor U4103 (N_4103,N_2363,N_2238);
or U4104 (N_4104,N_323,N_2356);
nor U4105 (N_4105,N_2229,N_1555);
nand U4106 (N_4106,N_1474,N_1310);
nor U4107 (N_4107,N_1657,N_745);
and U4108 (N_4108,N_907,N_603);
or U4109 (N_4109,N_879,N_692);
or U4110 (N_4110,N_1990,N_1405);
nand U4111 (N_4111,N_1023,N_2297);
nand U4112 (N_4112,N_2467,N_187);
nand U4113 (N_4113,N_2081,N_1400);
or U4114 (N_4114,N_380,N_1441);
nor U4115 (N_4115,N_825,N_2041);
nand U4116 (N_4116,N_1004,N_2110);
or U4117 (N_4117,N_1114,N_1865);
xor U4118 (N_4118,N_1045,N_2298);
and U4119 (N_4119,N_794,N_1117);
or U4120 (N_4120,N_223,N_1909);
nor U4121 (N_4121,N_116,N_669);
and U4122 (N_4122,N_1281,N_700);
and U4123 (N_4123,N_1722,N_1860);
nor U4124 (N_4124,N_203,N_425);
nand U4125 (N_4125,N_2194,N_573);
and U4126 (N_4126,N_1282,N_67);
nor U4127 (N_4127,N_1638,N_1681);
nand U4128 (N_4128,N_607,N_2195);
nor U4129 (N_4129,N_2063,N_1690);
or U4130 (N_4130,N_1778,N_628);
and U4131 (N_4131,N_893,N_1623);
nand U4132 (N_4132,N_383,N_1920);
xor U4133 (N_4133,N_1198,N_2351);
and U4134 (N_4134,N_651,N_33);
nor U4135 (N_4135,N_671,N_2037);
nor U4136 (N_4136,N_2201,N_348);
and U4137 (N_4137,N_673,N_1838);
and U4138 (N_4138,N_2146,N_1282);
and U4139 (N_4139,N_976,N_1845);
nand U4140 (N_4140,N_1456,N_773);
xnor U4141 (N_4141,N_697,N_262);
and U4142 (N_4142,N_247,N_1213);
xnor U4143 (N_4143,N_1944,N_1446);
and U4144 (N_4144,N_364,N_12);
or U4145 (N_4145,N_1828,N_2292);
xnor U4146 (N_4146,N_872,N_2090);
nand U4147 (N_4147,N_479,N_2380);
and U4148 (N_4148,N_1148,N_330);
xor U4149 (N_4149,N_576,N_304);
nand U4150 (N_4150,N_2130,N_2063);
nor U4151 (N_4151,N_1166,N_1520);
nor U4152 (N_4152,N_2287,N_138);
xor U4153 (N_4153,N_1885,N_1578);
nand U4154 (N_4154,N_2385,N_652);
nor U4155 (N_4155,N_238,N_1091);
nand U4156 (N_4156,N_2476,N_1801);
or U4157 (N_4157,N_1433,N_359);
nand U4158 (N_4158,N_772,N_1506);
or U4159 (N_4159,N_2026,N_1304);
nand U4160 (N_4160,N_389,N_1896);
nand U4161 (N_4161,N_638,N_2020);
or U4162 (N_4162,N_1806,N_1372);
or U4163 (N_4163,N_71,N_186);
nor U4164 (N_4164,N_2494,N_2251);
and U4165 (N_4165,N_440,N_713);
nor U4166 (N_4166,N_2347,N_1829);
nor U4167 (N_4167,N_902,N_919);
xnor U4168 (N_4168,N_1737,N_2387);
and U4169 (N_4169,N_113,N_1728);
nor U4170 (N_4170,N_1260,N_841);
and U4171 (N_4171,N_1381,N_1097);
nand U4172 (N_4172,N_1331,N_2039);
nor U4173 (N_4173,N_2243,N_322);
nor U4174 (N_4174,N_709,N_638);
or U4175 (N_4175,N_1477,N_1077);
nand U4176 (N_4176,N_2285,N_1423);
nor U4177 (N_4177,N_669,N_2293);
nor U4178 (N_4178,N_784,N_2060);
nand U4179 (N_4179,N_1596,N_1825);
or U4180 (N_4180,N_218,N_902);
or U4181 (N_4181,N_1157,N_1464);
nand U4182 (N_4182,N_1242,N_2167);
or U4183 (N_4183,N_2257,N_1479);
nand U4184 (N_4184,N_1446,N_1423);
nand U4185 (N_4185,N_2324,N_923);
and U4186 (N_4186,N_849,N_2115);
nor U4187 (N_4187,N_1811,N_931);
xor U4188 (N_4188,N_32,N_1352);
or U4189 (N_4189,N_1961,N_1848);
and U4190 (N_4190,N_2008,N_635);
nand U4191 (N_4191,N_91,N_2191);
or U4192 (N_4192,N_2070,N_1914);
nor U4193 (N_4193,N_1385,N_2328);
or U4194 (N_4194,N_629,N_851);
nand U4195 (N_4195,N_358,N_2156);
or U4196 (N_4196,N_521,N_2346);
nand U4197 (N_4197,N_911,N_2362);
and U4198 (N_4198,N_2323,N_1132);
nand U4199 (N_4199,N_2037,N_1204);
nand U4200 (N_4200,N_2328,N_1195);
nor U4201 (N_4201,N_1956,N_1480);
or U4202 (N_4202,N_350,N_1367);
nand U4203 (N_4203,N_1529,N_520);
or U4204 (N_4204,N_507,N_1058);
nor U4205 (N_4205,N_2319,N_1307);
nor U4206 (N_4206,N_1672,N_2326);
nand U4207 (N_4207,N_2354,N_675);
nor U4208 (N_4208,N_226,N_1216);
nand U4209 (N_4209,N_1922,N_746);
nor U4210 (N_4210,N_251,N_2082);
nor U4211 (N_4211,N_248,N_447);
nand U4212 (N_4212,N_72,N_1193);
or U4213 (N_4213,N_2479,N_2231);
nand U4214 (N_4214,N_572,N_2487);
nand U4215 (N_4215,N_114,N_1321);
and U4216 (N_4216,N_2298,N_1034);
or U4217 (N_4217,N_502,N_763);
xor U4218 (N_4218,N_225,N_1605);
or U4219 (N_4219,N_1876,N_828);
nor U4220 (N_4220,N_239,N_1627);
xnor U4221 (N_4221,N_1071,N_1657);
and U4222 (N_4222,N_1349,N_1456);
nor U4223 (N_4223,N_835,N_526);
nand U4224 (N_4224,N_983,N_2075);
nand U4225 (N_4225,N_186,N_1633);
and U4226 (N_4226,N_2295,N_1489);
nor U4227 (N_4227,N_1099,N_290);
or U4228 (N_4228,N_1175,N_470);
or U4229 (N_4229,N_1834,N_992);
or U4230 (N_4230,N_1254,N_2380);
and U4231 (N_4231,N_674,N_2047);
nand U4232 (N_4232,N_1095,N_1755);
and U4233 (N_4233,N_124,N_847);
nand U4234 (N_4234,N_2227,N_1113);
nand U4235 (N_4235,N_1757,N_489);
and U4236 (N_4236,N_154,N_2443);
or U4237 (N_4237,N_1166,N_1796);
or U4238 (N_4238,N_118,N_67);
nand U4239 (N_4239,N_180,N_2157);
xnor U4240 (N_4240,N_2392,N_1672);
nand U4241 (N_4241,N_415,N_323);
or U4242 (N_4242,N_869,N_2062);
and U4243 (N_4243,N_1213,N_2293);
nand U4244 (N_4244,N_2182,N_167);
nor U4245 (N_4245,N_1278,N_1312);
nor U4246 (N_4246,N_1427,N_916);
and U4247 (N_4247,N_1335,N_280);
and U4248 (N_4248,N_686,N_1117);
and U4249 (N_4249,N_1714,N_304);
and U4250 (N_4250,N_1651,N_1900);
or U4251 (N_4251,N_331,N_830);
nor U4252 (N_4252,N_1597,N_816);
xnor U4253 (N_4253,N_2003,N_1924);
or U4254 (N_4254,N_1725,N_1704);
and U4255 (N_4255,N_1738,N_665);
or U4256 (N_4256,N_1174,N_2066);
or U4257 (N_4257,N_879,N_87);
nor U4258 (N_4258,N_330,N_1080);
and U4259 (N_4259,N_653,N_957);
xor U4260 (N_4260,N_389,N_2209);
or U4261 (N_4261,N_928,N_839);
xor U4262 (N_4262,N_1006,N_610);
nand U4263 (N_4263,N_1633,N_1463);
nor U4264 (N_4264,N_782,N_917);
and U4265 (N_4265,N_2449,N_1362);
xnor U4266 (N_4266,N_2383,N_2119);
and U4267 (N_4267,N_396,N_1998);
nand U4268 (N_4268,N_1725,N_1364);
nor U4269 (N_4269,N_1251,N_1397);
xor U4270 (N_4270,N_871,N_1191);
nand U4271 (N_4271,N_232,N_2457);
nor U4272 (N_4272,N_1308,N_618);
xor U4273 (N_4273,N_773,N_1653);
or U4274 (N_4274,N_701,N_386);
or U4275 (N_4275,N_2303,N_626);
nand U4276 (N_4276,N_1910,N_2467);
or U4277 (N_4277,N_931,N_2108);
or U4278 (N_4278,N_2272,N_2266);
or U4279 (N_4279,N_310,N_569);
nor U4280 (N_4280,N_2006,N_1308);
nand U4281 (N_4281,N_1070,N_1595);
and U4282 (N_4282,N_2461,N_2286);
nor U4283 (N_4283,N_417,N_1867);
nor U4284 (N_4284,N_1266,N_1920);
xor U4285 (N_4285,N_1915,N_103);
or U4286 (N_4286,N_923,N_460);
or U4287 (N_4287,N_405,N_721);
nor U4288 (N_4288,N_1628,N_631);
or U4289 (N_4289,N_1946,N_2018);
or U4290 (N_4290,N_2235,N_995);
nor U4291 (N_4291,N_1729,N_1597);
nor U4292 (N_4292,N_491,N_435);
nand U4293 (N_4293,N_1754,N_2008);
nor U4294 (N_4294,N_1477,N_846);
or U4295 (N_4295,N_1813,N_1677);
and U4296 (N_4296,N_2121,N_191);
and U4297 (N_4297,N_1913,N_2189);
nand U4298 (N_4298,N_2475,N_2009);
xor U4299 (N_4299,N_553,N_625);
nand U4300 (N_4300,N_252,N_1299);
or U4301 (N_4301,N_2264,N_1978);
nor U4302 (N_4302,N_2118,N_2311);
or U4303 (N_4303,N_1054,N_1986);
nor U4304 (N_4304,N_143,N_542);
and U4305 (N_4305,N_2159,N_726);
and U4306 (N_4306,N_2083,N_1086);
nand U4307 (N_4307,N_1465,N_806);
xor U4308 (N_4308,N_2242,N_1516);
and U4309 (N_4309,N_2181,N_1455);
nand U4310 (N_4310,N_22,N_78);
nor U4311 (N_4311,N_1832,N_584);
nand U4312 (N_4312,N_653,N_1735);
xor U4313 (N_4313,N_2100,N_1223);
nor U4314 (N_4314,N_814,N_1734);
or U4315 (N_4315,N_1556,N_191);
xnor U4316 (N_4316,N_1794,N_2202);
xnor U4317 (N_4317,N_904,N_2469);
nand U4318 (N_4318,N_1511,N_2058);
nand U4319 (N_4319,N_1346,N_1705);
or U4320 (N_4320,N_1312,N_217);
nand U4321 (N_4321,N_1451,N_1384);
xnor U4322 (N_4322,N_16,N_120);
or U4323 (N_4323,N_1829,N_1769);
nor U4324 (N_4324,N_1040,N_1482);
xnor U4325 (N_4325,N_1668,N_2233);
nand U4326 (N_4326,N_985,N_1706);
nand U4327 (N_4327,N_475,N_1117);
nand U4328 (N_4328,N_942,N_1602);
and U4329 (N_4329,N_726,N_2103);
xnor U4330 (N_4330,N_463,N_2023);
and U4331 (N_4331,N_2194,N_2332);
or U4332 (N_4332,N_556,N_920);
xnor U4333 (N_4333,N_2265,N_455);
xnor U4334 (N_4334,N_2289,N_1703);
and U4335 (N_4335,N_2171,N_557);
nor U4336 (N_4336,N_692,N_1453);
nand U4337 (N_4337,N_1015,N_2419);
and U4338 (N_4338,N_2048,N_1242);
and U4339 (N_4339,N_7,N_333);
nand U4340 (N_4340,N_1553,N_2398);
nand U4341 (N_4341,N_883,N_2407);
or U4342 (N_4342,N_1010,N_2473);
nor U4343 (N_4343,N_2274,N_2032);
and U4344 (N_4344,N_2092,N_1820);
or U4345 (N_4345,N_2206,N_905);
nand U4346 (N_4346,N_1763,N_980);
nor U4347 (N_4347,N_1461,N_782);
or U4348 (N_4348,N_1945,N_1570);
nand U4349 (N_4349,N_991,N_1001);
nor U4350 (N_4350,N_762,N_1986);
nand U4351 (N_4351,N_766,N_2095);
nor U4352 (N_4352,N_2026,N_1129);
or U4353 (N_4353,N_1674,N_1921);
nand U4354 (N_4354,N_137,N_739);
nor U4355 (N_4355,N_2061,N_43);
nand U4356 (N_4356,N_834,N_2387);
xor U4357 (N_4357,N_2193,N_1841);
nor U4358 (N_4358,N_873,N_50);
nor U4359 (N_4359,N_2461,N_669);
and U4360 (N_4360,N_1859,N_215);
and U4361 (N_4361,N_1148,N_525);
nand U4362 (N_4362,N_178,N_245);
nand U4363 (N_4363,N_2114,N_425);
nand U4364 (N_4364,N_1163,N_1769);
or U4365 (N_4365,N_781,N_157);
and U4366 (N_4366,N_996,N_1436);
nand U4367 (N_4367,N_449,N_466);
or U4368 (N_4368,N_600,N_132);
or U4369 (N_4369,N_629,N_1365);
nor U4370 (N_4370,N_344,N_36);
or U4371 (N_4371,N_2235,N_795);
nand U4372 (N_4372,N_1406,N_2182);
and U4373 (N_4373,N_2339,N_210);
and U4374 (N_4374,N_1936,N_1635);
nand U4375 (N_4375,N_2200,N_614);
and U4376 (N_4376,N_1492,N_1767);
nor U4377 (N_4377,N_1760,N_1445);
or U4378 (N_4378,N_2434,N_1026);
and U4379 (N_4379,N_388,N_1239);
or U4380 (N_4380,N_680,N_442);
or U4381 (N_4381,N_1454,N_1621);
nor U4382 (N_4382,N_1666,N_1612);
and U4383 (N_4383,N_1237,N_2062);
nand U4384 (N_4384,N_2456,N_1547);
and U4385 (N_4385,N_1056,N_1244);
nor U4386 (N_4386,N_623,N_35);
and U4387 (N_4387,N_399,N_223);
or U4388 (N_4388,N_339,N_1427);
or U4389 (N_4389,N_2353,N_88);
xor U4390 (N_4390,N_263,N_2359);
nand U4391 (N_4391,N_1307,N_1977);
and U4392 (N_4392,N_1309,N_464);
and U4393 (N_4393,N_107,N_243);
or U4394 (N_4394,N_2244,N_2052);
nor U4395 (N_4395,N_1449,N_467);
and U4396 (N_4396,N_2125,N_2415);
nor U4397 (N_4397,N_1462,N_1624);
or U4398 (N_4398,N_1674,N_1975);
and U4399 (N_4399,N_422,N_821);
nand U4400 (N_4400,N_2305,N_54);
and U4401 (N_4401,N_1210,N_2499);
nor U4402 (N_4402,N_1246,N_1971);
and U4403 (N_4403,N_2144,N_1484);
and U4404 (N_4404,N_2414,N_529);
nor U4405 (N_4405,N_2136,N_629);
or U4406 (N_4406,N_350,N_631);
or U4407 (N_4407,N_1779,N_2202);
nand U4408 (N_4408,N_114,N_1378);
nor U4409 (N_4409,N_2451,N_667);
nor U4410 (N_4410,N_82,N_734);
nor U4411 (N_4411,N_1276,N_868);
nor U4412 (N_4412,N_1911,N_1412);
nor U4413 (N_4413,N_2447,N_556);
or U4414 (N_4414,N_1067,N_329);
nor U4415 (N_4415,N_370,N_1638);
and U4416 (N_4416,N_1937,N_240);
nor U4417 (N_4417,N_40,N_1503);
nand U4418 (N_4418,N_1268,N_2351);
nor U4419 (N_4419,N_572,N_212);
nand U4420 (N_4420,N_483,N_1325);
or U4421 (N_4421,N_1164,N_954);
and U4422 (N_4422,N_1283,N_615);
xor U4423 (N_4423,N_844,N_59);
nand U4424 (N_4424,N_1522,N_300);
or U4425 (N_4425,N_158,N_2247);
nor U4426 (N_4426,N_2359,N_1943);
nor U4427 (N_4427,N_33,N_1643);
nand U4428 (N_4428,N_1339,N_2188);
nand U4429 (N_4429,N_786,N_950);
and U4430 (N_4430,N_1431,N_946);
or U4431 (N_4431,N_2104,N_1288);
nor U4432 (N_4432,N_1274,N_1867);
nor U4433 (N_4433,N_961,N_1739);
and U4434 (N_4434,N_2470,N_2116);
and U4435 (N_4435,N_1550,N_442);
nand U4436 (N_4436,N_2298,N_833);
nand U4437 (N_4437,N_490,N_784);
nor U4438 (N_4438,N_1696,N_1098);
xnor U4439 (N_4439,N_414,N_1034);
or U4440 (N_4440,N_782,N_2280);
or U4441 (N_4441,N_802,N_642);
and U4442 (N_4442,N_1822,N_1374);
or U4443 (N_4443,N_62,N_883);
nor U4444 (N_4444,N_2220,N_216);
nand U4445 (N_4445,N_2335,N_296);
nand U4446 (N_4446,N_2463,N_652);
nor U4447 (N_4447,N_741,N_368);
nor U4448 (N_4448,N_1576,N_2275);
and U4449 (N_4449,N_2190,N_1760);
and U4450 (N_4450,N_724,N_776);
xnor U4451 (N_4451,N_805,N_1953);
xor U4452 (N_4452,N_790,N_77);
nand U4453 (N_4453,N_2483,N_2012);
nand U4454 (N_4454,N_1040,N_425);
nand U4455 (N_4455,N_1309,N_1975);
nand U4456 (N_4456,N_1720,N_1599);
and U4457 (N_4457,N_1050,N_516);
and U4458 (N_4458,N_1395,N_1426);
nor U4459 (N_4459,N_90,N_1331);
and U4460 (N_4460,N_346,N_348);
nand U4461 (N_4461,N_2475,N_1967);
or U4462 (N_4462,N_81,N_1483);
nor U4463 (N_4463,N_714,N_1545);
or U4464 (N_4464,N_2426,N_2376);
and U4465 (N_4465,N_2029,N_1957);
and U4466 (N_4466,N_1620,N_833);
nand U4467 (N_4467,N_652,N_617);
and U4468 (N_4468,N_2210,N_1965);
or U4469 (N_4469,N_1040,N_2089);
and U4470 (N_4470,N_2274,N_596);
and U4471 (N_4471,N_1602,N_808);
or U4472 (N_4472,N_1139,N_2034);
nand U4473 (N_4473,N_2273,N_62);
nor U4474 (N_4474,N_1546,N_1578);
nand U4475 (N_4475,N_2023,N_961);
nand U4476 (N_4476,N_623,N_709);
nand U4477 (N_4477,N_2269,N_2140);
nand U4478 (N_4478,N_1740,N_1505);
nor U4479 (N_4479,N_176,N_1215);
and U4480 (N_4480,N_380,N_995);
or U4481 (N_4481,N_1575,N_866);
and U4482 (N_4482,N_442,N_1915);
nor U4483 (N_4483,N_1497,N_958);
and U4484 (N_4484,N_2175,N_2310);
nor U4485 (N_4485,N_2365,N_1952);
nand U4486 (N_4486,N_1926,N_251);
and U4487 (N_4487,N_2281,N_369);
and U4488 (N_4488,N_139,N_1193);
nand U4489 (N_4489,N_4,N_69);
nor U4490 (N_4490,N_389,N_316);
xor U4491 (N_4491,N_2416,N_1168);
xnor U4492 (N_4492,N_2327,N_1959);
nand U4493 (N_4493,N_675,N_964);
or U4494 (N_4494,N_2472,N_776);
and U4495 (N_4495,N_1777,N_2494);
nor U4496 (N_4496,N_1916,N_1285);
and U4497 (N_4497,N_888,N_682);
and U4498 (N_4498,N_2008,N_1781);
or U4499 (N_4499,N_667,N_1133);
nand U4500 (N_4500,N_1884,N_1232);
or U4501 (N_4501,N_1027,N_1717);
nor U4502 (N_4502,N_1234,N_3);
nor U4503 (N_4503,N_1332,N_214);
and U4504 (N_4504,N_1912,N_2064);
nand U4505 (N_4505,N_1613,N_2399);
and U4506 (N_4506,N_2122,N_1597);
nor U4507 (N_4507,N_1502,N_2100);
nor U4508 (N_4508,N_1376,N_2136);
and U4509 (N_4509,N_2359,N_1960);
nand U4510 (N_4510,N_1754,N_57);
nor U4511 (N_4511,N_2411,N_309);
nand U4512 (N_4512,N_646,N_1652);
nand U4513 (N_4513,N_664,N_1938);
or U4514 (N_4514,N_143,N_2055);
and U4515 (N_4515,N_902,N_1942);
nand U4516 (N_4516,N_1810,N_1293);
nor U4517 (N_4517,N_2183,N_1953);
nand U4518 (N_4518,N_1961,N_1629);
or U4519 (N_4519,N_683,N_2331);
and U4520 (N_4520,N_1710,N_398);
nand U4521 (N_4521,N_442,N_917);
nor U4522 (N_4522,N_1266,N_1218);
and U4523 (N_4523,N_271,N_1140);
nor U4524 (N_4524,N_2425,N_1851);
and U4525 (N_4525,N_103,N_1464);
nor U4526 (N_4526,N_2301,N_347);
or U4527 (N_4527,N_120,N_304);
or U4528 (N_4528,N_805,N_1325);
nand U4529 (N_4529,N_1331,N_1148);
and U4530 (N_4530,N_518,N_105);
or U4531 (N_4531,N_416,N_519);
or U4532 (N_4532,N_1751,N_1974);
nand U4533 (N_4533,N_1420,N_939);
and U4534 (N_4534,N_1350,N_2451);
nand U4535 (N_4535,N_2473,N_1340);
and U4536 (N_4536,N_1823,N_1198);
nand U4537 (N_4537,N_990,N_868);
or U4538 (N_4538,N_1418,N_1911);
or U4539 (N_4539,N_795,N_434);
nor U4540 (N_4540,N_144,N_1702);
or U4541 (N_4541,N_949,N_1435);
xor U4542 (N_4542,N_325,N_2321);
nor U4543 (N_4543,N_1734,N_85);
or U4544 (N_4544,N_2414,N_1);
nor U4545 (N_4545,N_689,N_1373);
nor U4546 (N_4546,N_1701,N_1590);
and U4547 (N_4547,N_1185,N_2406);
nand U4548 (N_4548,N_54,N_300);
nor U4549 (N_4549,N_2454,N_1667);
or U4550 (N_4550,N_613,N_2143);
nand U4551 (N_4551,N_1025,N_27);
nand U4552 (N_4552,N_1157,N_767);
and U4553 (N_4553,N_1225,N_1498);
xnor U4554 (N_4554,N_2087,N_1513);
xnor U4555 (N_4555,N_742,N_1919);
nand U4556 (N_4556,N_1418,N_2473);
or U4557 (N_4557,N_1614,N_1172);
or U4558 (N_4558,N_830,N_494);
xor U4559 (N_4559,N_1409,N_1834);
and U4560 (N_4560,N_628,N_1274);
and U4561 (N_4561,N_272,N_1846);
or U4562 (N_4562,N_435,N_340);
nand U4563 (N_4563,N_2386,N_589);
and U4564 (N_4564,N_2311,N_1497);
nor U4565 (N_4565,N_1514,N_1734);
and U4566 (N_4566,N_1178,N_1716);
and U4567 (N_4567,N_79,N_2206);
or U4568 (N_4568,N_454,N_1214);
nand U4569 (N_4569,N_2029,N_1125);
nand U4570 (N_4570,N_523,N_1083);
or U4571 (N_4571,N_813,N_2314);
nand U4572 (N_4572,N_633,N_2465);
nand U4573 (N_4573,N_986,N_1490);
and U4574 (N_4574,N_1711,N_2422);
nor U4575 (N_4575,N_1361,N_2179);
or U4576 (N_4576,N_741,N_2194);
or U4577 (N_4577,N_672,N_671);
and U4578 (N_4578,N_1961,N_2432);
or U4579 (N_4579,N_1607,N_2226);
and U4580 (N_4580,N_633,N_1135);
and U4581 (N_4581,N_17,N_1930);
nand U4582 (N_4582,N_299,N_113);
or U4583 (N_4583,N_1571,N_2031);
nor U4584 (N_4584,N_1493,N_1271);
and U4585 (N_4585,N_2246,N_2111);
or U4586 (N_4586,N_487,N_2410);
nor U4587 (N_4587,N_2041,N_120);
nor U4588 (N_4588,N_1518,N_1042);
and U4589 (N_4589,N_229,N_2464);
xor U4590 (N_4590,N_2209,N_1873);
nor U4591 (N_4591,N_2219,N_1138);
and U4592 (N_4592,N_34,N_442);
nor U4593 (N_4593,N_2014,N_8);
xnor U4594 (N_4594,N_12,N_1832);
nand U4595 (N_4595,N_192,N_896);
nand U4596 (N_4596,N_1029,N_1121);
xnor U4597 (N_4597,N_2383,N_946);
xnor U4598 (N_4598,N_397,N_873);
nor U4599 (N_4599,N_787,N_542);
nand U4600 (N_4600,N_1577,N_1687);
nor U4601 (N_4601,N_916,N_355);
or U4602 (N_4602,N_159,N_1398);
nor U4603 (N_4603,N_756,N_985);
or U4604 (N_4604,N_1664,N_1730);
or U4605 (N_4605,N_2447,N_902);
nand U4606 (N_4606,N_1468,N_99);
xnor U4607 (N_4607,N_1331,N_997);
and U4608 (N_4608,N_770,N_1044);
nor U4609 (N_4609,N_1096,N_1554);
nand U4610 (N_4610,N_18,N_65);
xor U4611 (N_4611,N_1236,N_681);
or U4612 (N_4612,N_1343,N_1755);
nand U4613 (N_4613,N_1732,N_2412);
nor U4614 (N_4614,N_1053,N_1096);
nand U4615 (N_4615,N_427,N_1339);
xor U4616 (N_4616,N_1705,N_1164);
nand U4617 (N_4617,N_2098,N_2180);
nand U4618 (N_4618,N_1,N_1246);
or U4619 (N_4619,N_1289,N_115);
nand U4620 (N_4620,N_1981,N_2020);
xnor U4621 (N_4621,N_389,N_1228);
or U4622 (N_4622,N_2259,N_600);
and U4623 (N_4623,N_1620,N_1431);
nor U4624 (N_4624,N_1628,N_498);
nand U4625 (N_4625,N_197,N_105);
nor U4626 (N_4626,N_854,N_1414);
or U4627 (N_4627,N_317,N_24);
nor U4628 (N_4628,N_1502,N_1553);
xnor U4629 (N_4629,N_1674,N_2139);
nor U4630 (N_4630,N_2474,N_511);
nor U4631 (N_4631,N_1439,N_2392);
nor U4632 (N_4632,N_55,N_1080);
nand U4633 (N_4633,N_1060,N_1473);
nor U4634 (N_4634,N_1847,N_1151);
nand U4635 (N_4635,N_2246,N_1077);
nor U4636 (N_4636,N_2487,N_1919);
and U4637 (N_4637,N_1419,N_1294);
nand U4638 (N_4638,N_91,N_2027);
and U4639 (N_4639,N_2340,N_2387);
nor U4640 (N_4640,N_852,N_672);
nand U4641 (N_4641,N_769,N_382);
nand U4642 (N_4642,N_1429,N_1512);
or U4643 (N_4643,N_1165,N_1054);
and U4644 (N_4644,N_2065,N_2346);
nor U4645 (N_4645,N_2246,N_648);
xor U4646 (N_4646,N_2471,N_134);
nand U4647 (N_4647,N_2322,N_435);
nor U4648 (N_4648,N_2288,N_1648);
or U4649 (N_4649,N_102,N_622);
and U4650 (N_4650,N_180,N_1337);
and U4651 (N_4651,N_2265,N_2340);
or U4652 (N_4652,N_622,N_2394);
nand U4653 (N_4653,N_71,N_695);
nand U4654 (N_4654,N_1705,N_74);
or U4655 (N_4655,N_1785,N_692);
xnor U4656 (N_4656,N_618,N_2388);
nor U4657 (N_4657,N_1754,N_333);
nand U4658 (N_4658,N_1522,N_759);
or U4659 (N_4659,N_218,N_2388);
or U4660 (N_4660,N_1216,N_947);
and U4661 (N_4661,N_1166,N_447);
nand U4662 (N_4662,N_479,N_1537);
or U4663 (N_4663,N_2299,N_251);
or U4664 (N_4664,N_1536,N_78);
or U4665 (N_4665,N_1275,N_68);
nand U4666 (N_4666,N_676,N_2161);
nor U4667 (N_4667,N_1564,N_1989);
nand U4668 (N_4668,N_93,N_1991);
xnor U4669 (N_4669,N_913,N_50);
nand U4670 (N_4670,N_777,N_1751);
nand U4671 (N_4671,N_984,N_1415);
nand U4672 (N_4672,N_1130,N_295);
or U4673 (N_4673,N_1423,N_2466);
and U4674 (N_4674,N_694,N_1535);
nand U4675 (N_4675,N_41,N_1656);
nand U4676 (N_4676,N_889,N_2145);
nand U4677 (N_4677,N_1772,N_2280);
xnor U4678 (N_4678,N_504,N_1990);
xnor U4679 (N_4679,N_2130,N_1048);
or U4680 (N_4680,N_2214,N_1205);
xnor U4681 (N_4681,N_2212,N_2005);
xnor U4682 (N_4682,N_1267,N_1018);
nand U4683 (N_4683,N_1202,N_1078);
nand U4684 (N_4684,N_1570,N_367);
nor U4685 (N_4685,N_1199,N_586);
nand U4686 (N_4686,N_1585,N_1135);
or U4687 (N_4687,N_1874,N_384);
and U4688 (N_4688,N_537,N_836);
nor U4689 (N_4689,N_1211,N_593);
nor U4690 (N_4690,N_1638,N_748);
nand U4691 (N_4691,N_1404,N_515);
or U4692 (N_4692,N_1769,N_1355);
or U4693 (N_4693,N_1900,N_395);
and U4694 (N_4694,N_469,N_1607);
and U4695 (N_4695,N_834,N_2029);
and U4696 (N_4696,N_1875,N_1517);
and U4697 (N_4697,N_887,N_365);
or U4698 (N_4698,N_749,N_990);
nor U4699 (N_4699,N_706,N_2128);
or U4700 (N_4700,N_2300,N_13);
nor U4701 (N_4701,N_904,N_85);
nand U4702 (N_4702,N_2168,N_1063);
and U4703 (N_4703,N_1299,N_722);
and U4704 (N_4704,N_830,N_807);
nor U4705 (N_4705,N_613,N_466);
xor U4706 (N_4706,N_85,N_1470);
nand U4707 (N_4707,N_1906,N_157);
and U4708 (N_4708,N_495,N_1588);
or U4709 (N_4709,N_978,N_805);
or U4710 (N_4710,N_1982,N_767);
and U4711 (N_4711,N_1764,N_1090);
nor U4712 (N_4712,N_636,N_1510);
nand U4713 (N_4713,N_1438,N_140);
nor U4714 (N_4714,N_1936,N_574);
or U4715 (N_4715,N_1176,N_1627);
nand U4716 (N_4716,N_1867,N_1119);
and U4717 (N_4717,N_1888,N_899);
and U4718 (N_4718,N_1715,N_674);
or U4719 (N_4719,N_747,N_778);
nor U4720 (N_4720,N_1232,N_1581);
xnor U4721 (N_4721,N_477,N_741);
nor U4722 (N_4722,N_125,N_1074);
nor U4723 (N_4723,N_541,N_2130);
and U4724 (N_4724,N_158,N_2400);
xor U4725 (N_4725,N_921,N_981);
and U4726 (N_4726,N_432,N_1727);
and U4727 (N_4727,N_1253,N_773);
and U4728 (N_4728,N_1842,N_744);
xnor U4729 (N_4729,N_2299,N_1196);
nor U4730 (N_4730,N_1853,N_1425);
nand U4731 (N_4731,N_997,N_2355);
nand U4732 (N_4732,N_465,N_715);
or U4733 (N_4733,N_2077,N_1365);
or U4734 (N_4734,N_197,N_2062);
xnor U4735 (N_4735,N_2384,N_2403);
xor U4736 (N_4736,N_2271,N_742);
nand U4737 (N_4737,N_2233,N_144);
and U4738 (N_4738,N_477,N_1907);
nor U4739 (N_4739,N_920,N_657);
and U4740 (N_4740,N_175,N_1820);
nor U4741 (N_4741,N_204,N_2103);
xnor U4742 (N_4742,N_1875,N_1772);
nor U4743 (N_4743,N_1066,N_1742);
and U4744 (N_4744,N_2116,N_994);
nor U4745 (N_4745,N_351,N_949);
nor U4746 (N_4746,N_2452,N_1391);
nor U4747 (N_4747,N_1744,N_2371);
and U4748 (N_4748,N_1416,N_636);
and U4749 (N_4749,N_1611,N_1874);
nor U4750 (N_4750,N_2177,N_708);
nand U4751 (N_4751,N_243,N_1396);
and U4752 (N_4752,N_1346,N_2411);
xnor U4753 (N_4753,N_792,N_2143);
nand U4754 (N_4754,N_328,N_1384);
and U4755 (N_4755,N_41,N_2019);
nor U4756 (N_4756,N_409,N_1924);
xor U4757 (N_4757,N_2405,N_898);
or U4758 (N_4758,N_554,N_1760);
or U4759 (N_4759,N_219,N_1242);
or U4760 (N_4760,N_830,N_235);
and U4761 (N_4761,N_1186,N_2484);
and U4762 (N_4762,N_2268,N_834);
nand U4763 (N_4763,N_373,N_1640);
and U4764 (N_4764,N_131,N_297);
nand U4765 (N_4765,N_479,N_205);
or U4766 (N_4766,N_906,N_875);
or U4767 (N_4767,N_97,N_1526);
nor U4768 (N_4768,N_467,N_1600);
nor U4769 (N_4769,N_1322,N_374);
and U4770 (N_4770,N_1185,N_2403);
and U4771 (N_4771,N_2463,N_802);
and U4772 (N_4772,N_772,N_2482);
nand U4773 (N_4773,N_1785,N_1809);
xor U4774 (N_4774,N_59,N_422);
or U4775 (N_4775,N_2371,N_550);
and U4776 (N_4776,N_32,N_1045);
or U4777 (N_4777,N_1918,N_327);
and U4778 (N_4778,N_557,N_648);
xnor U4779 (N_4779,N_2382,N_1679);
or U4780 (N_4780,N_1564,N_1450);
xor U4781 (N_4781,N_2103,N_323);
and U4782 (N_4782,N_2247,N_261);
nand U4783 (N_4783,N_640,N_1206);
and U4784 (N_4784,N_2469,N_2449);
and U4785 (N_4785,N_1958,N_1551);
xnor U4786 (N_4786,N_122,N_2464);
and U4787 (N_4787,N_1175,N_1304);
nand U4788 (N_4788,N_900,N_1072);
nand U4789 (N_4789,N_1005,N_2463);
or U4790 (N_4790,N_871,N_1899);
or U4791 (N_4791,N_885,N_2142);
nand U4792 (N_4792,N_317,N_1181);
nor U4793 (N_4793,N_1443,N_419);
nor U4794 (N_4794,N_1519,N_968);
or U4795 (N_4795,N_1944,N_722);
and U4796 (N_4796,N_1814,N_671);
nand U4797 (N_4797,N_96,N_1559);
nand U4798 (N_4798,N_2120,N_1602);
or U4799 (N_4799,N_2386,N_1891);
or U4800 (N_4800,N_2387,N_147);
or U4801 (N_4801,N_1601,N_1442);
and U4802 (N_4802,N_2253,N_1510);
or U4803 (N_4803,N_737,N_2375);
xnor U4804 (N_4804,N_776,N_2212);
and U4805 (N_4805,N_602,N_285);
or U4806 (N_4806,N_2154,N_782);
and U4807 (N_4807,N_1698,N_2284);
nor U4808 (N_4808,N_593,N_1333);
or U4809 (N_4809,N_1027,N_2092);
and U4810 (N_4810,N_2364,N_379);
and U4811 (N_4811,N_410,N_1558);
xor U4812 (N_4812,N_1199,N_846);
nand U4813 (N_4813,N_1134,N_905);
nor U4814 (N_4814,N_88,N_1565);
or U4815 (N_4815,N_1665,N_1149);
nand U4816 (N_4816,N_253,N_391);
nand U4817 (N_4817,N_1490,N_1401);
nand U4818 (N_4818,N_171,N_1417);
nor U4819 (N_4819,N_2444,N_1540);
nor U4820 (N_4820,N_1403,N_2141);
or U4821 (N_4821,N_3,N_330);
nand U4822 (N_4822,N_2147,N_2464);
or U4823 (N_4823,N_1113,N_302);
and U4824 (N_4824,N_138,N_501);
or U4825 (N_4825,N_667,N_822);
or U4826 (N_4826,N_1489,N_3);
or U4827 (N_4827,N_270,N_2477);
or U4828 (N_4828,N_2464,N_612);
and U4829 (N_4829,N_2311,N_705);
and U4830 (N_4830,N_35,N_823);
nand U4831 (N_4831,N_2383,N_1563);
or U4832 (N_4832,N_637,N_721);
xnor U4833 (N_4833,N_1639,N_640);
or U4834 (N_4834,N_948,N_552);
xor U4835 (N_4835,N_1322,N_1901);
or U4836 (N_4836,N_778,N_441);
nor U4837 (N_4837,N_785,N_1772);
nor U4838 (N_4838,N_1104,N_1468);
or U4839 (N_4839,N_1351,N_1008);
or U4840 (N_4840,N_319,N_1427);
xor U4841 (N_4841,N_1345,N_574);
and U4842 (N_4842,N_1989,N_759);
nor U4843 (N_4843,N_297,N_10);
nor U4844 (N_4844,N_1868,N_1089);
or U4845 (N_4845,N_2309,N_788);
and U4846 (N_4846,N_560,N_2047);
and U4847 (N_4847,N_2468,N_1256);
or U4848 (N_4848,N_995,N_438);
xor U4849 (N_4849,N_1913,N_223);
nor U4850 (N_4850,N_886,N_649);
or U4851 (N_4851,N_1522,N_1403);
nor U4852 (N_4852,N_400,N_1849);
nor U4853 (N_4853,N_2015,N_2185);
or U4854 (N_4854,N_352,N_1867);
and U4855 (N_4855,N_1626,N_2350);
xnor U4856 (N_4856,N_982,N_2272);
or U4857 (N_4857,N_1030,N_1208);
and U4858 (N_4858,N_2375,N_1236);
xnor U4859 (N_4859,N_83,N_1401);
or U4860 (N_4860,N_2398,N_844);
nor U4861 (N_4861,N_1928,N_1601);
xor U4862 (N_4862,N_1358,N_1879);
or U4863 (N_4863,N_1069,N_944);
nand U4864 (N_4864,N_1804,N_2067);
nor U4865 (N_4865,N_1755,N_769);
or U4866 (N_4866,N_1245,N_2121);
or U4867 (N_4867,N_2178,N_2410);
or U4868 (N_4868,N_2472,N_426);
nor U4869 (N_4869,N_1811,N_2390);
nand U4870 (N_4870,N_2389,N_472);
nor U4871 (N_4871,N_166,N_2149);
nand U4872 (N_4872,N_1125,N_1556);
nor U4873 (N_4873,N_1061,N_1181);
and U4874 (N_4874,N_1556,N_1943);
or U4875 (N_4875,N_2422,N_696);
or U4876 (N_4876,N_2069,N_356);
nand U4877 (N_4877,N_1010,N_1767);
nand U4878 (N_4878,N_2241,N_1170);
nand U4879 (N_4879,N_1269,N_1393);
and U4880 (N_4880,N_2016,N_1779);
and U4881 (N_4881,N_1218,N_2018);
nor U4882 (N_4882,N_2312,N_1811);
nand U4883 (N_4883,N_2294,N_672);
xor U4884 (N_4884,N_1175,N_2269);
xnor U4885 (N_4885,N_1552,N_685);
nand U4886 (N_4886,N_1199,N_2014);
or U4887 (N_4887,N_1170,N_357);
nor U4888 (N_4888,N_287,N_1849);
or U4889 (N_4889,N_1237,N_697);
and U4890 (N_4890,N_920,N_984);
nor U4891 (N_4891,N_691,N_935);
nor U4892 (N_4892,N_708,N_628);
nor U4893 (N_4893,N_1667,N_2155);
or U4894 (N_4894,N_522,N_1907);
nor U4895 (N_4895,N_1526,N_101);
nor U4896 (N_4896,N_972,N_2273);
nand U4897 (N_4897,N_1744,N_203);
xor U4898 (N_4898,N_81,N_3);
nand U4899 (N_4899,N_1918,N_2010);
and U4900 (N_4900,N_2389,N_346);
xor U4901 (N_4901,N_405,N_566);
or U4902 (N_4902,N_1521,N_1794);
nand U4903 (N_4903,N_1415,N_2013);
xnor U4904 (N_4904,N_76,N_992);
and U4905 (N_4905,N_136,N_380);
nand U4906 (N_4906,N_831,N_294);
nor U4907 (N_4907,N_480,N_774);
nor U4908 (N_4908,N_675,N_1226);
nand U4909 (N_4909,N_209,N_553);
and U4910 (N_4910,N_233,N_541);
xor U4911 (N_4911,N_874,N_2234);
nor U4912 (N_4912,N_180,N_1963);
nor U4913 (N_4913,N_1947,N_698);
or U4914 (N_4914,N_622,N_11);
or U4915 (N_4915,N_2491,N_415);
nor U4916 (N_4916,N_1614,N_1659);
and U4917 (N_4917,N_249,N_413);
or U4918 (N_4918,N_1864,N_166);
and U4919 (N_4919,N_490,N_1867);
nand U4920 (N_4920,N_123,N_1518);
nand U4921 (N_4921,N_248,N_1036);
or U4922 (N_4922,N_2424,N_2293);
nand U4923 (N_4923,N_1538,N_547);
nand U4924 (N_4924,N_1572,N_320);
xnor U4925 (N_4925,N_2199,N_1893);
and U4926 (N_4926,N_2481,N_1058);
or U4927 (N_4927,N_2109,N_1287);
or U4928 (N_4928,N_1957,N_1396);
nand U4929 (N_4929,N_1906,N_170);
nand U4930 (N_4930,N_2482,N_153);
and U4931 (N_4931,N_694,N_1289);
nor U4932 (N_4932,N_1715,N_891);
or U4933 (N_4933,N_2220,N_1164);
nand U4934 (N_4934,N_2497,N_2330);
nor U4935 (N_4935,N_887,N_2028);
and U4936 (N_4936,N_2078,N_918);
xor U4937 (N_4937,N_1800,N_120);
and U4938 (N_4938,N_2442,N_1470);
and U4939 (N_4939,N_2377,N_576);
or U4940 (N_4940,N_43,N_934);
nor U4941 (N_4941,N_185,N_808);
nand U4942 (N_4942,N_803,N_523);
xor U4943 (N_4943,N_1138,N_1108);
or U4944 (N_4944,N_2480,N_1826);
or U4945 (N_4945,N_706,N_2340);
nand U4946 (N_4946,N_1567,N_597);
nand U4947 (N_4947,N_1477,N_1921);
nand U4948 (N_4948,N_1891,N_1004);
or U4949 (N_4949,N_1619,N_2054);
xnor U4950 (N_4950,N_2413,N_2151);
or U4951 (N_4951,N_2406,N_35);
nand U4952 (N_4952,N_1939,N_1405);
nand U4953 (N_4953,N_342,N_686);
nand U4954 (N_4954,N_869,N_327);
and U4955 (N_4955,N_2447,N_590);
and U4956 (N_4956,N_106,N_245);
xnor U4957 (N_4957,N_926,N_907);
nand U4958 (N_4958,N_1692,N_1782);
nor U4959 (N_4959,N_466,N_2052);
or U4960 (N_4960,N_2331,N_1932);
or U4961 (N_4961,N_1919,N_2177);
nand U4962 (N_4962,N_1264,N_2464);
xor U4963 (N_4963,N_518,N_902);
or U4964 (N_4964,N_2346,N_675);
and U4965 (N_4965,N_2270,N_26);
nor U4966 (N_4966,N_2248,N_1242);
nand U4967 (N_4967,N_394,N_2481);
nand U4968 (N_4968,N_919,N_2264);
or U4969 (N_4969,N_725,N_300);
or U4970 (N_4970,N_1691,N_1759);
nor U4971 (N_4971,N_425,N_1999);
nand U4972 (N_4972,N_524,N_201);
and U4973 (N_4973,N_726,N_1771);
nor U4974 (N_4974,N_569,N_1356);
nor U4975 (N_4975,N_1559,N_1192);
nor U4976 (N_4976,N_108,N_1298);
and U4977 (N_4977,N_691,N_2208);
nor U4978 (N_4978,N_1547,N_1668);
nand U4979 (N_4979,N_1152,N_2442);
nor U4980 (N_4980,N_377,N_703);
nor U4981 (N_4981,N_1739,N_2094);
or U4982 (N_4982,N_2479,N_1932);
and U4983 (N_4983,N_1206,N_190);
nor U4984 (N_4984,N_1344,N_755);
or U4985 (N_4985,N_1289,N_600);
nand U4986 (N_4986,N_1754,N_991);
or U4987 (N_4987,N_2275,N_6);
and U4988 (N_4988,N_1650,N_1815);
and U4989 (N_4989,N_1848,N_629);
nor U4990 (N_4990,N_1126,N_1133);
nand U4991 (N_4991,N_2359,N_174);
and U4992 (N_4992,N_666,N_1788);
or U4993 (N_4993,N_490,N_1787);
nand U4994 (N_4994,N_1764,N_153);
or U4995 (N_4995,N_504,N_2028);
or U4996 (N_4996,N_2108,N_1212);
nor U4997 (N_4997,N_2253,N_1206);
nand U4998 (N_4998,N_1678,N_1515);
nor U4999 (N_4999,N_616,N_2254);
and UO_0 (O_0,N_2603,N_4513);
nand UO_1 (O_1,N_2863,N_3605);
xor UO_2 (O_2,N_3518,N_4853);
or UO_3 (O_3,N_3294,N_2548);
nor UO_4 (O_4,N_4670,N_2815);
and UO_5 (O_5,N_4245,N_3992);
xor UO_6 (O_6,N_3185,N_4113);
or UO_7 (O_7,N_4130,N_4974);
and UO_8 (O_8,N_4504,N_3158);
and UO_9 (O_9,N_4420,N_3321);
nand UO_10 (O_10,N_3863,N_4945);
nor UO_11 (O_11,N_4961,N_4414);
xnor UO_12 (O_12,N_3541,N_2850);
or UO_13 (O_13,N_3630,N_3230);
nand UO_14 (O_14,N_3523,N_2504);
or UO_15 (O_15,N_4939,N_3224);
nor UO_16 (O_16,N_4674,N_2777);
or UO_17 (O_17,N_2941,N_4168);
nand UO_18 (O_18,N_4356,N_3679);
nor UO_19 (O_19,N_3724,N_2730);
nor UO_20 (O_20,N_3316,N_3195);
and UO_21 (O_21,N_2606,N_3553);
or UO_22 (O_22,N_4946,N_4810);
nand UO_23 (O_23,N_2536,N_4900);
nor UO_24 (O_24,N_2554,N_3771);
xor UO_25 (O_25,N_3315,N_4984);
and UO_26 (O_26,N_2802,N_3357);
nor UO_27 (O_27,N_3869,N_3841);
and UO_28 (O_28,N_4027,N_4935);
nand UO_29 (O_29,N_3283,N_4043);
xor UO_30 (O_30,N_4213,N_3188);
or UO_31 (O_31,N_4392,N_4620);
and UO_32 (O_32,N_2680,N_3532);
and UO_33 (O_33,N_3817,N_3362);
and UO_34 (O_34,N_4802,N_2952);
nor UO_35 (O_35,N_4845,N_3522);
and UO_36 (O_36,N_3439,N_3628);
nor UO_37 (O_37,N_3804,N_3133);
nand UO_38 (O_38,N_4720,N_2552);
or UO_39 (O_39,N_4728,N_4022);
xnor UO_40 (O_40,N_3967,N_2591);
or UO_41 (O_41,N_2894,N_3545);
xor UO_42 (O_42,N_3128,N_2976);
nand UO_43 (O_43,N_2597,N_2753);
or UO_44 (O_44,N_3737,N_2613);
nor UO_45 (O_45,N_2568,N_4187);
nor UO_46 (O_46,N_4960,N_2584);
or UO_47 (O_47,N_2703,N_4302);
nand UO_48 (O_48,N_2632,N_3310);
or UO_49 (O_49,N_3820,N_4091);
and UO_50 (O_50,N_2969,N_3245);
nand UO_51 (O_51,N_4396,N_4633);
nor UO_52 (O_52,N_2899,N_4582);
or UO_53 (O_53,N_4273,N_2563);
and UO_54 (O_54,N_3738,N_2521);
and UO_55 (O_55,N_4074,N_4625);
nand UO_56 (O_56,N_3401,N_4370);
and UO_57 (O_57,N_3624,N_4454);
nand UO_58 (O_58,N_2734,N_2866);
nand UO_59 (O_59,N_3341,N_4614);
or UO_60 (O_60,N_3247,N_3396);
nand UO_61 (O_61,N_4986,N_2938);
nand UO_62 (O_62,N_3772,N_4357);
nor UO_63 (O_63,N_3468,N_3814);
nor UO_64 (O_64,N_3166,N_4886);
nor UO_65 (O_65,N_3160,N_4084);
or UO_66 (O_66,N_3345,N_4428);
nand UO_67 (O_67,N_3473,N_3010);
nor UO_68 (O_68,N_3113,N_4085);
nor UO_69 (O_69,N_3931,N_4268);
nand UO_70 (O_70,N_3398,N_3744);
nor UO_71 (O_71,N_3819,N_4149);
and UO_72 (O_72,N_2902,N_3700);
and UO_73 (O_73,N_3526,N_3592);
nand UO_74 (O_74,N_3210,N_4145);
nor UO_75 (O_75,N_3574,N_4056);
or UO_76 (O_76,N_2825,N_3181);
or UO_77 (O_77,N_3520,N_3045);
nor UO_78 (O_78,N_3385,N_4899);
nor UO_79 (O_79,N_3977,N_4894);
nand UO_80 (O_80,N_2547,N_4331);
or UO_81 (O_81,N_3782,N_4088);
or UO_82 (O_82,N_3250,N_4281);
nand UO_83 (O_83,N_4475,N_4713);
or UO_84 (O_84,N_3622,N_2854);
nor UO_85 (O_85,N_3913,N_4100);
or UO_86 (O_86,N_4226,N_4827);
or UO_87 (O_87,N_3603,N_4553);
nor UO_88 (O_88,N_3675,N_2935);
nor UO_89 (O_89,N_4417,N_3300);
and UO_90 (O_90,N_3213,N_3939);
or UO_91 (O_91,N_4884,N_3384);
or UO_92 (O_92,N_4242,N_3950);
and UO_93 (O_93,N_4381,N_2522);
and UO_94 (O_94,N_4293,N_3741);
or UO_95 (O_95,N_2764,N_4624);
nor UO_96 (O_96,N_4282,N_4530);
and UO_97 (O_97,N_3944,N_3855);
and UO_98 (O_98,N_2770,N_4186);
and UO_99 (O_99,N_3747,N_2827);
or UO_100 (O_100,N_4727,N_3458);
and UO_101 (O_101,N_4761,N_3088);
and UO_102 (O_102,N_4192,N_4630);
xnor UO_103 (O_103,N_4044,N_4010);
nand UO_104 (O_104,N_4321,N_2960);
nand UO_105 (O_105,N_4759,N_3156);
xnor UO_106 (O_106,N_3008,N_3621);
nor UO_107 (O_107,N_4366,N_2982);
nand UO_108 (O_108,N_4249,N_2994);
or UO_109 (O_109,N_3656,N_3081);
or UO_110 (O_110,N_3061,N_2887);
and UO_111 (O_111,N_2908,N_3162);
or UO_112 (O_112,N_4017,N_2569);
xor UO_113 (O_113,N_3907,N_4416);
and UO_114 (O_114,N_4103,N_4055);
or UO_115 (O_115,N_3102,N_3389);
nand UO_116 (O_116,N_3478,N_3118);
nand UO_117 (O_117,N_3180,N_4528);
and UO_118 (O_118,N_2845,N_4052);
or UO_119 (O_119,N_3256,N_2822);
and UO_120 (O_120,N_2737,N_2884);
nand UO_121 (O_121,N_4593,N_3129);
nand UO_122 (O_122,N_3463,N_4985);
nand UO_123 (O_123,N_3849,N_4646);
or UO_124 (O_124,N_4906,N_2720);
and UO_125 (O_125,N_3995,N_3936);
nand UO_126 (O_126,N_3665,N_4161);
nand UO_127 (O_127,N_2503,N_2799);
or UO_128 (O_128,N_4893,N_3588);
nand UO_129 (O_129,N_3405,N_3757);
nand UO_130 (O_130,N_4219,N_4518);
nand UO_131 (O_131,N_2787,N_4109);
nor UO_132 (O_132,N_4702,N_4295);
nand UO_133 (O_133,N_4967,N_2813);
and UO_134 (O_134,N_3220,N_4262);
xnor UO_135 (O_135,N_4285,N_2712);
and UO_136 (O_136,N_4708,N_4527);
xor UO_137 (O_137,N_4606,N_3619);
and UO_138 (O_138,N_2747,N_4350);
nor UO_139 (O_139,N_2812,N_2784);
or UO_140 (O_140,N_3769,N_4538);
nand UO_141 (O_141,N_4953,N_4451);
or UO_142 (O_142,N_2988,N_4399);
or UO_143 (O_143,N_3876,N_4666);
nand UO_144 (O_144,N_3018,N_2668);
nand UO_145 (O_145,N_2816,N_3546);
nor UO_146 (O_146,N_4269,N_4063);
or UO_147 (O_147,N_3305,N_3930);
nor UO_148 (O_148,N_3689,N_2942);
nand UO_149 (O_149,N_4143,N_2519);
nor UO_150 (O_150,N_3497,N_4768);
nand UO_151 (O_151,N_2727,N_4694);
and UO_152 (O_152,N_4609,N_4405);
and UO_153 (O_153,N_4431,N_4372);
and UO_154 (O_154,N_3703,N_4699);
nand UO_155 (O_155,N_3847,N_3112);
and UO_156 (O_156,N_4919,N_2625);
and UO_157 (O_157,N_2934,N_2655);
nor UO_158 (O_158,N_2746,N_3641);
or UO_159 (O_159,N_3898,N_3658);
xor UO_160 (O_160,N_2526,N_3272);
nor UO_161 (O_161,N_3009,N_4912);
xnor UO_162 (O_162,N_2642,N_4065);
and UO_163 (O_163,N_3368,N_3938);
and UO_164 (O_164,N_4803,N_4231);
nand UO_165 (O_165,N_4343,N_3645);
xnor UO_166 (O_166,N_3561,N_4223);
or UO_167 (O_167,N_4008,N_3635);
nor UO_168 (O_168,N_3671,N_3712);
and UO_169 (O_169,N_4989,N_3016);
nand UO_170 (O_170,N_3372,N_3496);
and UO_171 (O_171,N_4170,N_2915);
nor UO_172 (O_172,N_4276,N_2931);
xor UO_173 (O_173,N_4638,N_4077);
nand UO_174 (O_174,N_4051,N_4574);
and UO_175 (O_175,N_4526,N_4612);
nand UO_176 (O_176,N_4832,N_3238);
nor UO_177 (O_177,N_4049,N_4503);
or UO_178 (O_178,N_3388,N_3266);
nand UO_179 (O_179,N_3033,N_4937);
and UO_180 (O_180,N_3715,N_4062);
or UO_181 (O_181,N_4983,N_4379);
and UO_182 (O_182,N_3611,N_4924);
or UO_183 (O_183,N_3058,N_4408);
nand UO_184 (O_184,N_4443,N_3171);
nor UO_185 (O_185,N_3822,N_4797);
nand UO_186 (O_186,N_2583,N_2710);
xor UO_187 (O_187,N_4297,N_3324);
nor UO_188 (O_188,N_3299,N_3034);
nor UO_189 (O_189,N_4619,N_4844);
and UO_190 (O_190,N_4304,N_3956);
nand UO_191 (O_191,N_2949,N_4469);
nor UO_192 (O_192,N_4765,N_4771);
nand UO_193 (O_193,N_2514,N_3743);
and UO_194 (O_194,N_4164,N_3205);
nand UO_195 (O_195,N_3914,N_2532);
nand UO_196 (O_196,N_4811,N_4987);
nand UO_197 (O_197,N_2836,N_4964);
or UO_198 (O_198,N_2824,N_2851);
or UO_199 (O_199,N_2858,N_3157);
and UO_200 (O_200,N_3327,N_3435);
or UO_201 (O_201,N_3674,N_2619);
xor UO_202 (O_202,N_2856,N_2599);
nor UO_203 (O_203,N_4822,N_4457);
nand UO_204 (O_204,N_4442,N_3433);
or UO_205 (O_205,N_4979,N_4485);
xnor UO_206 (O_206,N_3456,N_3991);
nand UO_207 (O_207,N_2987,N_4115);
or UO_208 (O_208,N_3547,N_3566);
and UO_209 (O_209,N_4733,N_3540);
nor UO_210 (O_210,N_4075,N_2742);
or UO_211 (O_211,N_4641,N_4496);
or UO_212 (O_212,N_3445,N_3079);
nor UO_213 (O_213,N_4823,N_3270);
or UO_214 (O_214,N_4715,N_4755);
or UO_215 (O_215,N_2715,N_2963);
or UO_216 (O_216,N_3575,N_3122);
nor UO_217 (O_217,N_4601,N_4332);
nor UO_218 (O_218,N_2829,N_3259);
nand UO_219 (O_219,N_4347,N_4596);
and UO_220 (O_220,N_4018,N_3706);
and UO_221 (O_221,N_4004,N_3457);
nor UO_222 (O_222,N_4541,N_3460);
or UO_223 (O_223,N_4807,N_4559);
or UO_224 (O_224,N_3816,N_2722);
nand UO_225 (O_225,N_4106,N_4791);
and UO_226 (O_226,N_3090,N_4794);
nand UO_227 (O_227,N_3469,N_2608);
nor UO_228 (O_228,N_4851,N_2754);
nand UO_229 (O_229,N_2652,N_3484);
xnor UO_230 (O_230,N_3901,N_2587);
and UO_231 (O_231,N_4423,N_4232);
and UO_232 (O_232,N_4275,N_4458);
or UO_233 (O_233,N_4267,N_4025);
and UO_234 (O_234,N_2956,N_3732);
and UO_235 (O_235,N_2757,N_4477);
nand UO_236 (O_236,N_3607,N_4543);
and UO_237 (O_237,N_2590,N_4305);
and UO_238 (O_238,N_3291,N_3485);
nand UO_239 (O_239,N_3778,N_4453);
or UO_240 (O_240,N_3695,N_4828);
or UO_241 (O_241,N_2600,N_4692);
and UO_242 (O_242,N_3786,N_4456);
nand UO_243 (O_243,N_3909,N_2872);
nor UO_244 (O_244,N_3837,N_4258);
and UO_245 (O_245,N_4642,N_3447);
or UO_246 (O_246,N_3610,N_3844);
nor UO_247 (O_247,N_3170,N_3165);
nor UO_248 (O_248,N_3548,N_3236);
nand UO_249 (O_249,N_4510,N_3443);
nor UO_250 (O_250,N_4691,N_3438);
and UO_251 (O_251,N_2707,N_3954);
nand UO_252 (O_252,N_2911,N_3501);
xor UO_253 (O_253,N_4549,N_4166);
or UO_254 (O_254,N_3859,N_4994);
xor UO_255 (O_255,N_2843,N_3970);
nand UO_256 (O_256,N_4617,N_4169);
or UO_257 (O_257,N_4798,N_4901);
and UO_258 (O_258,N_3066,N_4590);
or UO_259 (O_259,N_3503,N_2659);
xor UO_260 (O_260,N_4648,N_2678);
and UO_261 (O_261,N_4839,N_4497);
nor UO_262 (O_262,N_4923,N_4789);
or UO_263 (O_263,N_4227,N_4398);
nor UO_264 (O_264,N_3828,N_3414);
nand UO_265 (O_265,N_2890,N_2708);
nand UO_266 (O_266,N_3805,N_3296);
nand UO_267 (O_267,N_4190,N_4512);
xnor UO_268 (O_268,N_2876,N_4300);
and UO_269 (O_269,N_4039,N_3192);
or UO_270 (O_270,N_4959,N_3818);
or UO_271 (O_271,N_3246,N_4922);
or UO_272 (O_272,N_4388,N_3958);
and UO_273 (O_273,N_3676,N_4162);
nor UO_274 (O_274,N_3933,N_2859);
or UO_275 (O_275,N_3618,N_4493);
nor UO_276 (O_276,N_3851,N_2965);
nand UO_277 (O_277,N_4033,N_2743);
nor UO_278 (O_278,N_4146,N_3135);
nand UO_279 (O_279,N_3101,N_2847);
nor UO_280 (O_280,N_3638,N_4483);
and UO_281 (O_281,N_2700,N_4659);
nor UO_282 (O_282,N_4344,N_4799);
or UO_283 (O_283,N_3972,N_4778);
and UO_284 (O_284,N_3854,N_2620);
nand UO_285 (O_285,N_4000,N_2631);
or UO_286 (O_286,N_3536,N_4656);
nor UO_287 (O_287,N_2940,N_3390);
or UO_288 (O_288,N_4718,N_3726);
nand UO_289 (O_289,N_4037,N_3882);
or UO_290 (O_290,N_4448,N_3402);
and UO_291 (O_291,N_4846,N_2912);
and UO_292 (O_292,N_4490,N_4345);
nor UO_293 (O_293,N_4661,N_3030);
or UO_294 (O_294,N_3382,N_3350);
or UO_295 (O_295,N_4296,N_4888);
xnor UO_296 (O_296,N_4933,N_4289);
or UO_297 (O_297,N_4222,N_4592);
and UO_298 (O_298,N_3788,N_3583);
xor UO_299 (O_299,N_4565,N_3812);
and UO_300 (O_300,N_2616,N_4135);
nor UO_301 (O_301,N_3041,N_3749);
nand UO_302 (O_302,N_3556,N_3323);
or UO_303 (O_303,N_4754,N_3196);
xor UO_304 (O_304,N_4196,N_4938);
and UO_305 (O_305,N_2817,N_4736);
or UO_306 (O_306,N_3953,N_3397);
xor UO_307 (O_307,N_3506,N_3421);
or UO_308 (O_308,N_2535,N_3317);
nor UO_309 (O_309,N_2647,N_3998);
nand UO_310 (O_310,N_4198,N_4383);
nand UO_311 (O_311,N_4632,N_4307);
nor UO_312 (O_312,N_4346,N_2502);
nand UO_313 (O_313,N_2995,N_4421);
nand UO_314 (O_314,N_4724,N_3488);
and UO_315 (O_315,N_2875,N_2674);
and UO_316 (O_316,N_3739,N_4413);
xnor UO_317 (O_317,N_3426,N_3123);
xor UO_318 (O_318,N_3237,N_3842);
xnor UO_319 (O_319,N_2990,N_3669);
nand UO_320 (O_320,N_4516,N_3590);
nand UO_321 (O_321,N_3762,N_2852);
nor UO_322 (O_322,N_3225,N_4988);
nand UO_323 (O_323,N_4349,N_3687);
or UO_324 (O_324,N_3625,N_2726);
nand UO_325 (O_325,N_4318,N_3810);
or UO_326 (O_326,N_4118,N_4926);
xnor UO_327 (O_327,N_4339,N_4564);
xor UO_328 (O_328,N_4315,N_3344);
nor UO_329 (O_329,N_3746,N_3971);
nand UO_330 (O_330,N_4603,N_4608);
nor UO_331 (O_331,N_3131,N_4981);
or UO_332 (O_332,N_4707,N_3029);
nand UO_333 (O_333,N_2531,N_2913);
and UO_334 (O_334,N_4487,N_4438);
or UO_335 (O_335,N_3719,N_2640);
or UO_336 (O_336,N_4358,N_3792);
nand UO_337 (O_337,N_4758,N_3314);
xnor UO_338 (O_338,N_3428,N_2683);
or UO_339 (O_339,N_2546,N_3612);
nand UO_340 (O_340,N_3516,N_3821);
and UO_341 (O_341,N_3740,N_4178);
nor UO_342 (O_342,N_4869,N_3054);
nand UO_343 (O_343,N_4569,N_4998);
xor UO_344 (O_344,N_4382,N_3311);
xor UO_345 (O_345,N_4867,N_2791);
nor UO_346 (O_346,N_2518,N_3343);
and UO_347 (O_347,N_3774,N_3318);
nor UO_348 (O_348,N_3798,N_4563);
xor UO_349 (O_349,N_2749,N_3025);
or UO_350 (O_350,N_4667,N_4480);
or UO_351 (O_351,N_4447,N_4947);
or UO_352 (O_352,N_3801,N_2837);
and UO_353 (O_353,N_4627,N_3942);
nor UO_354 (O_354,N_4430,N_2577);
and UO_355 (O_355,N_2550,N_4341);
xnor UO_356 (O_356,N_4494,N_4461);
nand UO_357 (O_357,N_4096,N_3279);
nand UO_358 (O_358,N_3134,N_3904);
or UO_359 (O_359,N_3356,N_2779);
nand UO_360 (O_360,N_2873,N_3955);
nor UO_361 (O_361,N_2732,N_4127);
nor UO_362 (O_362,N_2898,N_2762);
nand UO_363 (O_363,N_3244,N_3062);
or UO_364 (O_364,N_4533,N_3052);
or UO_365 (O_365,N_3699,N_4792);
and UO_366 (O_366,N_2760,N_4148);
xor UO_367 (O_367,N_3896,N_3333);
or UO_368 (O_368,N_4086,N_4045);
and UO_369 (O_369,N_4813,N_3643);
and UO_370 (O_370,N_3696,N_3403);
and UO_371 (O_371,N_3945,N_3519);
xnor UO_372 (O_372,N_4271,N_4843);
and UO_373 (O_373,N_3660,N_2641);
nand UO_374 (O_374,N_4584,N_4819);
and UO_375 (O_375,N_3897,N_3273);
nor UO_376 (O_376,N_4020,N_4204);
nand UO_377 (O_377,N_3429,N_4531);
nor UO_378 (O_378,N_3718,N_4083);
or UO_379 (O_379,N_4914,N_4931);
and UO_380 (O_380,N_3092,N_3234);
and UO_381 (O_381,N_3095,N_4465);
xor UO_382 (O_382,N_4706,N_4495);
xor UO_383 (O_383,N_3666,N_3021);
xnor UO_384 (O_384,N_4460,N_4599);
or UO_385 (O_385,N_3690,N_3207);
or UO_386 (O_386,N_4311,N_2752);
or UO_387 (O_387,N_4240,N_4856);
nand UO_388 (O_388,N_2721,N_2741);
xnor UO_389 (O_389,N_4221,N_3551);
xnor UO_390 (O_390,N_4548,N_2992);
nand UO_391 (O_391,N_2650,N_4685);
nor UO_392 (O_392,N_3534,N_4435);
nor UO_393 (O_393,N_4537,N_4274);
nor UO_394 (O_394,N_4329,N_3892);
and UO_395 (O_395,N_3573,N_2756);
nor UO_396 (O_396,N_4409,N_3263);
nand UO_397 (O_397,N_2633,N_3895);
or UO_398 (O_398,N_3200,N_3500);
nor UO_399 (O_399,N_4189,N_4956);
and UO_400 (O_400,N_4831,N_2692);
nand UO_401 (O_401,N_3581,N_3078);
and UO_402 (O_402,N_4837,N_4167);
nand UO_403 (O_403,N_4976,N_4029);
or UO_404 (O_404,N_4247,N_3916);
or UO_405 (O_405,N_4298,N_3861);
nand UO_406 (O_406,N_4940,N_2883);
and UO_407 (O_407,N_4842,N_2702);
xnor UO_408 (O_408,N_3027,N_2586);
and UO_409 (O_409,N_4260,N_3932);
nor UO_410 (O_410,N_2653,N_4224);
and UO_411 (O_411,N_4566,N_4663);
and UO_412 (O_412,N_2657,N_2759);
or UO_413 (O_413,N_4814,N_4309);
nor UO_414 (O_414,N_3374,N_3032);
or UO_415 (O_415,N_4746,N_2681);
nand UO_416 (O_416,N_3417,N_3751);
nor UO_417 (O_417,N_4507,N_4763);
nor UO_418 (O_418,N_4800,N_3584);
nand UO_419 (O_419,N_4072,N_4738);
nand UO_420 (O_420,N_3640,N_4520);
nand UO_421 (O_421,N_4760,N_4114);
nor UO_422 (O_422,N_2991,N_2945);
nand UO_423 (O_423,N_4449,N_2645);
or UO_424 (O_424,N_3019,N_3492);
nor UO_425 (O_425,N_3182,N_3906);
or UO_426 (O_426,N_3217,N_4359);
nor UO_427 (O_427,N_4594,N_3620);
nor UO_428 (O_428,N_4117,N_4781);
or UO_429 (O_429,N_3194,N_3673);
nor UO_430 (O_430,N_3899,N_4129);
nor UO_431 (O_431,N_3975,N_3585);
nor UO_432 (O_432,N_3634,N_3340);
or UO_433 (O_433,N_4154,N_4821);
or UO_434 (O_434,N_3462,N_2557);
nor UO_435 (O_435,N_3383,N_2705);
and UO_436 (O_436,N_4312,N_4711);
nand UO_437 (O_437,N_3924,N_2682);
or UO_438 (O_438,N_4978,N_4655);
nand UO_439 (O_439,N_3874,N_3902);
xnor UO_440 (O_440,N_4857,N_3834);
nand UO_441 (O_441,N_2573,N_2977);
and UO_442 (O_442,N_3571,N_2654);
nand UO_443 (O_443,N_3793,N_3422);
or UO_444 (O_444,N_4206,N_2588);
and UO_445 (O_445,N_3132,N_4773);
xnor UO_446 (O_446,N_4731,N_4723);
nor UO_447 (O_447,N_3780,N_4588);
nand UO_448 (O_448,N_3727,N_2735);
nand UO_449 (O_449,N_4654,N_2505);
xor UO_450 (O_450,N_3597,N_4205);
and UO_451 (O_451,N_4214,N_3872);
nand UO_452 (O_452,N_3486,N_4185);
xor UO_453 (O_453,N_3569,N_3183);
and UO_454 (O_454,N_3831,N_3114);
xor UO_455 (O_455,N_4534,N_4155);
nor UO_456 (O_456,N_3176,N_2724);
or UO_457 (O_457,N_3394,N_3601);
xor UO_458 (O_458,N_3006,N_4488);
or UO_459 (O_459,N_4834,N_4522);
nand UO_460 (O_460,N_3020,N_3147);
or UO_461 (O_461,N_2897,N_3203);
nand UO_462 (O_462,N_4629,N_2672);
nand UO_463 (O_463,N_2520,N_4073);
nor UO_464 (O_464,N_4783,N_2801);
nor UO_465 (O_465,N_2545,N_4328);
nand UO_466 (O_466,N_3365,N_4611);
nand UO_467 (O_467,N_4669,N_3168);
nand UO_468 (O_468,N_4519,N_2543);
nand UO_469 (O_469,N_4132,N_4470);
xnor UO_470 (O_470,N_4476,N_3479);
xnor UO_471 (O_471,N_2895,N_3487);
nand UO_472 (O_472,N_3701,N_3215);
nand UO_473 (O_473,N_4890,N_3796);
nand UO_474 (O_474,N_3750,N_4885);
and UO_475 (O_475,N_2975,N_4861);
and UO_476 (O_476,N_3400,N_2629);
nor UO_477 (O_477,N_4047,N_2512);
xor UO_478 (O_478,N_3789,N_2954);
and UO_479 (O_479,N_2886,N_2840);
or UO_480 (O_480,N_4153,N_4874);
nor UO_481 (O_481,N_2795,N_3705);
nand UO_482 (O_482,N_3572,N_3427);
and UO_483 (O_483,N_3688,N_4403);
nand UO_484 (O_484,N_3606,N_3053);
or UO_485 (O_485,N_4751,N_2750);
and UO_486 (O_486,N_3243,N_2919);
xnor UO_487 (O_487,N_4764,N_4673);
and UO_488 (O_488,N_3338,N_2604);
nor UO_489 (O_489,N_3352,N_2921);
nor UO_490 (O_490,N_3632,N_4089);
and UO_491 (O_491,N_2675,N_4915);
or UO_492 (O_492,N_3885,N_4054);
and UO_493 (O_493,N_2943,N_3017);
nand UO_494 (O_494,N_4523,N_2755);
or UO_495 (O_495,N_3777,N_3337);
and UO_496 (O_496,N_3716,N_4440);
and UO_497 (O_497,N_4184,N_4545);
and UO_498 (O_498,N_4122,N_4698);
nand UO_499 (O_499,N_4286,N_3364);
or UO_500 (O_500,N_3005,N_3511);
nor UO_501 (O_501,N_3312,N_2892);
and UO_502 (O_502,N_4134,N_3758);
or UO_503 (O_503,N_3997,N_4492);
nor UO_504 (O_504,N_4253,N_4770);
and UO_505 (O_505,N_3284,N_3125);
or UO_506 (O_506,N_4936,N_2689);
nand UO_507 (O_507,N_4235,N_4917);
nor UO_508 (O_508,N_4099,N_3282);
and UO_509 (O_509,N_2804,N_3322);
nor UO_510 (O_510,N_3555,N_4144);
nand UO_511 (O_511,N_4891,N_2970);
and UO_512 (O_512,N_4929,N_2973);
nor UO_513 (O_513,N_2582,N_3867);
nor UO_514 (O_514,N_4322,N_4090);
or UO_515 (O_515,N_3698,N_3752);
or UO_516 (O_516,N_3890,N_4575);
nor UO_517 (O_517,N_4208,N_3120);
and UO_518 (O_518,N_4462,N_2544);
nand UO_519 (O_519,N_2864,N_4256);
xor UO_520 (O_520,N_3889,N_4059);
or UO_521 (O_521,N_2950,N_3529);
or UO_522 (O_522,N_3046,N_3784);
and UO_523 (O_523,N_4990,N_4554);
and UO_524 (O_524,N_3014,N_3678);
and UO_525 (O_525,N_4216,N_3037);
nand UO_526 (O_526,N_4651,N_4767);
and UO_527 (O_527,N_4610,N_4270);
and UO_528 (O_528,N_4397,N_3535);
nand UO_529 (O_529,N_4158,N_4491);
nand UO_530 (O_530,N_4278,N_4326);
or UO_531 (O_531,N_2958,N_3077);
or UO_532 (O_532,N_4352,N_3646);
or UO_533 (O_533,N_2868,N_2733);
nor UO_534 (O_534,N_4236,N_3360);
or UO_535 (O_535,N_4618,N_4371);
and UO_536 (O_536,N_4604,N_4136);
or UO_537 (O_537,N_2841,N_3662);
nor UO_538 (O_538,N_4365,N_2927);
nand UO_539 (O_539,N_3370,N_4419);
or UO_540 (O_540,N_4784,N_3920);
or UO_541 (O_541,N_4474,N_3567);
and UO_542 (O_542,N_4557,N_3110);
nand UO_543 (O_543,N_4303,N_4683);
or UO_544 (O_544,N_4112,N_4038);
nand UO_545 (O_545,N_3334,N_3948);
nor UO_546 (O_546,N_3593,N_3378);
or UO_547 (O_547,N_3083,N_4690);
and UO_548 (O_548,N_4156,N_3910);
or UO_549 (O_549,N_3961,N_3984);
xor UO_550 (O_550,N_4904,N_4968);
and UO_551 (O_551,N_2661,N_2916);
nand UO_552 (O_552,N_3404,N_4092);
nor UO_553 (O_553,N_4266,N_3146);
and UO_554 (O_554,N_3164,N_4013);
xor UO_555 (O_555,N_4586,N_3807);
and UO_556 (O_556,N_2556,N_4970);
or UO_557 (O_557,N_3328,N_4820);
xnor UO_558 (O_558,N_3431,N_2639);
nand UO_559 (O_559,N_3785,N_3227);
nand UO_560 (O_560,N_4688,N_3276);
nand UO_561 (O_561,N_2888,N_2946);
or UO_562 (O_562,N_3467,N_3680);
or UO_563 (O_563,N_3979,N_4468);
and UO_564 (O_564,N_3295,N_4766);
nand UO_565 (O_565,N_4665,N_4446);
and UO_566 (O_566,N_3251,N_2951);
nand UO_567 (O_567,N_4384,N_3297);
nor UO_568 (O_568,N_4402,N_2914);
nand UO_569 (O_569,N_4234,N_2811);
xnor UO_570 (O_570,N_3069,N_4598);
nand UO_571 (O_571,N_3064,N_3850);
and UO_572 (O_572,N_3304,N_3670);
or UO_573 (O_573,N_3152,N_3302);
nor UO_574 (O_574,N_3407,N_4696);
nand UO_575 (O_575,N_3050,N_4850);
xnor UO_576 (O_576,N_4228,N_4866);
nor UO_577 (O_577,N_2646,N_3221);
or UO_578 (O_578,N_2879,N_3049);
xnor UO_579 (O_579,N_3483,N_2839);
or UO_580 (O_580,N_4455,N_4110);
nand UO_581 (O_581,N_4643,N_3142);
nand UO_582 (O_582,N_3981,N_3615);
nor UO_583 (O_583,N_4237,N_4070);
and UO_584 (O_584,N_4250,N_4473);
nor UO_585 (O_585,N_3391,N_3905);
and UO_586 (O_586,N_3022,N_2593);
xor UO_587 (O_587,N_3963,N_3527);
and UO_588 (O_588,N_3490,N_4841);
xnor UO_589 (O_589,N_4287,N_3966);
nor UO_590 (O_590,N_3964,N_3175);
nor UO_591 (O_591,N_3934,N_2596);
or UO_592 (O_592,N_2842,N_2628);
or UO_593 (O_593,N_2961,N_3035);
nand UO_594 (O_594,N_4464,N_4433);
and UO_595 (O_595,N_4466,N_3642);
xnor UO_596 (O_596,N_3836,N_3783);
xor UO_597 (O_597,N_4591,N_4515);
or UO_598 (O_598,N_3655,N_4862);
nand UO_599 (O_599,N_3361,N_4732);
or UO_600 (O_600,N_4163,N_4215);
and UO_601 (O_601,N_4607,N_2904);
nand UO_602 (O_602,N_4097,N_4525);
nand UO_603 (O_603,N_4639,N_2846);
or UO_604 (O_604,N_2778,N_4314);
or UO_605 (O_605,N_4902,N_3048);
or UO_606 (O_606,N_3377,N_3832);
or UO_607 (O_607,N_3248,N_3104);
nand UO_608 (O_608,N_4211,N_3240);
or UO_609 (O_609,N_4057,N_3228);
nor UO_610 (O_610,N_2538,N_4966);
or UO_611 (O_611,N_4631,N_4191);
nor UO_612 (O_612,N_4772,N_4040);
and UO_613 (O_613,N_4201,N_3366);
nand UO_614 (O_614,N_3633,N_3258);
or UO_615 (O_615,N_2959,N_4060);
and UO_616 (O_616,N_2622,N_2862);
nor UO_617 (O_617,N_3515,N_4128);
or UO_618 (O_618,N_3811,N_3332);
nand UO_619 (O_619,N_3307,N_3993);
nand UO_620 (O_620,N_4081,N_3594);
nand UO_621 (O_621,N_3830,N_2955);
or UO_622 (O_622,N_4336,N_3459);
nor UO_623 (O_623,N_4082,N_3039);
nand UO_624 (O_624,N_3576,N_2997);
xnor UO_625 (O_625,N_4188,N_4600);
xnor UO_626 (O_626,N_2729,N_4567);
nor UO_627 (O_627,N_3087,N_3415);
nand UO_628 (O_628,N_2819,N_4511);
and UO_629 (O_629,N_3094,N_4220);
and UO_630 (O_630,N_4535,N_3533);
or UO_631 (O_631,N_3694,N_4653);
and UO_632 (O_632,N_4870,N_4141);
xnor UO_633 (O_633,N_2968,N_3734);
or UO_634 (O_634,N_3893,N_4719);
xnor UO_635 (O_635,N_4335,N_4479);
and UO_636 (O_636,N_2786,N_4182);
xnor UO_637 (O_637,N_4812,N_3846);
nand UO_638 (O_638,N_4437,N_2607);
or UO_639 (O_639,N_3725,N_3233);
nand UO_640 (O_640,N_3568,N_2944);
nand UO_641 (O_641,N_3524,N_3288);
or UO_642 (O_642,N_3894,N_2806);
nor UO_643 (O_643,N_4925,N_4023);
and UO_644 (O_644,N_2728,N_2644);
nand UO_645 (O_645,N_2771,N_3833);
and UO_646 (O_646,N_2922,N_4348);
or UO_647 (O_647,N_4080,N_3359);
or UO_648 (O_648,N_3795,N_2800);
xnor UO_649 (O_649,N_3843,N_4229);
and UO_650 (O_650,N_2809,N_4306);
and UO_651 (O_651,N_4210,N_4374);
nor UO_652 (O_652,N_3664,N_4671);
nand UO_653 (O_653,N_3060,N_3349);
or UO_654 (O_654,N_3002,N_3293);
or UO_655 (O_655,N_2665,N_4078);
and UO_656 (O_656,N_4815,N_4160);
and UO_657 (O_657,N_4662,N_2910);
nand UO_658 (O_658,N_3481,N_3085);
nor UO_659 (O_659,N_2648,N_4048);
nor UO_660 (O_660,N_4927,N_3935);
or UO_661 (O_661,N_3071,N_4849);
or UO_662 (O_662,N_3287,N_4628);
nand UO_663 (O_663,N_4159,N_3161);
and UO_664 (O_664,N_2774,N_4279);
xnor UO_665 (O_665,N_2989,N_4505);
or UO_666 (O_666,N_4993,N_2510);
and UO_667 (O_667,N_4176,N_2595);
nor UO_668 (O_668,N_2559,N_3412);
or UO_669 (O_669,N_3808,N_2551);
nor UO_670 (O_670,N_4225,N_2660);
nand UO_671 (O_671,N_2688,N_3242);
xnor UO_672 (O_672,N_4401,N_3860);
or UO_673 (O_673,N_4737,N_2611);
nand UO_674 (O_674,N_3026,N_3145);
or UO_675 (O_675,N_3214,N_3838);
or UO_676 (O_676,N_3968,N_3186);
nor UO_677 (O_677,N_2937,N_4195);
nand UO_678 (O_678,N_2830,N_3639);
or UO_679 (O_679,N_4877,N_4657);
and UO_680 (O_680,N_3707,N_4317);
and UO_681 (O_681,N_4742,N_4701);
xor UO_682 (O_682,N_3254,N_2694);
or UO_683 (O_683,N_4107,N_4907);
or UO_684 (O_684,N_4547,N_3420);
nor UO_685 (O_685,N_4848,N_4506);
or UO_686 (O_686,N_4427,N_3187);
or UO_687 (O_687,N_3184,N_2869);
nand UO_688 (O_688,N_4200,N_2617);
nand UO_689 (O_689,N_3093,N_3392);
and UO_690 (O_690,N_3096,N_2805);
or UO_691 (O_691,N_2814,N_4542);
nor UO_692 (O_692,N_2540,N_4868);
nand UO_693 (O_693,N_2566,N_3395);
xnor UO_694 (O_694,N_4716,N_4218);
nor UO_695 (O_695,N_2585,N_3292);
or UO_696 (O_696,N_4524,N_4053);
nand UO_697 (O_697,N_3542,N_3591);
nor UO_698 (O_698,N_3351,N_2893);
xnor UO_699 (O_699,N_3723,N_3609);
and UO_700 (O_700,N_3959,N_4509);
nor UO_701 (O_701,N_3862,N_3974);
or UO_702 (O_702,N_3608,N_3451);
nor UO_703 (O_703,N_4634,N_2594);
nand UO_704 (O_704,N_3124,N_3498);
nand UO_705 (O_705,N_3602,N_3823);
or UO_706 (O_706,N_4955,N_3912);
nand UO_707 (O_707,N_2792,N_4808);
nand UO_708 (O_708,N_2553,N_4375);
nor UO_709 (O_709,N_3692,N_3677);
and UO_710 (O_710,N_4377,N_4292);
or UO_711 (O_711,N_4272,N_3996);
or UO_712 (O_712,N_3929,N_4194);
nand UO_713 (O_713,N_4066,N_4787);
or UO_714 (O_714,N_2711,N_2979);
and UO_715 (O_715,N_2844,N_4521);
or UO_716 (O_716,N_4424,N_3631);
nand UO_717 (O_717,N_3325,N_4579);
nor UO_718 (O_718,N_4997,N_4910);
nor UO_719 (O_719,N_3150,N_4031);
nor UO_720 (O_720,N_3693,N_4660);
xor UO_721 (O_721,N_3476,N_3482);
nor UO_722 (O_722,N_2980,N_3748);
nand UO_723 (O_723,N_3063,N_3216);
nand UO_724 (O_724,N_4105,N_3274);
nand UO_725 (O_725,N_2870,N_4616);
and UO_726 (O_726,N_3845,N_3241);
or UO_727 (O_727,N_2656,N_4064);
nor UO_728 (O_728,N_2758,N_3148);
nor UO_729 (O_729,N_3260,N_4678);
nand UO_730 (O_730,N_3733,N_2581);
nand UO_731 (O_731,N_4833,N_2534);
or UO_732 (O_732,N_3763,N_3865);
xnor UO_733 (O_733,N_2891,N_3298);
nor UO_734 (O_734,N_3425,N_2601);
and UO_735 (O_735,N_3768,N_4952);
nand UO_736 (O_736,N_4636,N_3436);
and UO_737 (O_737,N_3629,N_2614);
and UO_738 (O_738,N_2798,N_3794);
and UO_739 (O_739,N_2881,N_2998);
nor UO_740 (O_740,N_3495,N_4697);
xnor UO_741 (O_741,N_3736,N_2687);
and UO_742 (O_742,N_4005,N_4354);
nor UO_743 (O_743,N_2984,N_4407);
or UO_744 (O_744,N_4830,N_4920);
or UO_745 (O_745,N_2917,N_4265);
nand UO_746 (O_746,N_3280,N_3558);
or UO_747 (O_747,N_3410,N_2782);
nand UO_748 (O_748,N_4568,N_2718);
or UO_749 (O_749,N_4288,N_3206);
nand UO_750 (O_750,N_4942,N_4921);
or UO_751 (O_751,N_2598,N_2761);
nand UO_752 (O_752,N_4881,N_2558);
and UO_753 (O_753,N_4640,N_2731);
or UO_754 (O_754,N_3505,N_2820);
and UO_755 (O_755,N_4826,N_3626);
nor UO_756 (O_756,N_3179,N_3708);
xor UO_757 (O_757,N_2853,N_4181);
or UO_758 (O_758,N_4895,N_2565);
or UO_759 (O_759,N_4602,N_3197);
and UO_760 (O_760,N_3489,N_4498);
xor UO_761 (O_761,N_2763,N_3320);
and UO_762 (O_762,N_4650,N_3163);
or UO_763 (O_763,N_3189,N_3848);
and UO_764 (O_764,N_3770,N_2524);
nand UO_765 (O_765,N_4780,N_2751);
xor UO_766 (O_766,N_3923,N_3720);
and UO_767 (O_767,N_4710,N_3880);
nand UO_768 (O_768,N_3153,N_4675);
or UO_769 (O_769,N_2947,N_4739);
nor UO_770 (O_770,N_3684,N_4965);
nand UO_771 (O_771,N_4319,N_3432);
or UO_772 (O_772,N_4847,N_4139);
nand UO_773 (O_773,N_4486,N_2736);
nor UO_774 (O_774,N_3809,N_4277);
nor UO_775 (O_775,N_2537,N_2515);
and UO_776 (O_776,N_4687,N_3202);
nor UO_777 (O_777,N_2667,N_2848);
nand UO_778 (O_778,N_2723,N_2772);
and UO_779 (O_779,N_2695,N_4050);
nand UO_780 (O_780,N_4174,N_3466);
nand UO_781 (O_781,N_4429,N_4948);
nand UO_782 (O_782,N_2542,N_4042);
and UO_783 (O_783,N_4391,N_4104);
and UO_784 (O_784,N_4835,N_4776);
nor UO_785 (O_785,N_2903,N_3411);
and UO_786 (O_786,N_2789,N_2985);
or UO_787 (O_787,N_3363,N_3802);
nand UO_788 (O_788,N_3644,N_3174);
or UO_789 (O_789,N_4310,N_4230);
and UO_790 (O_790,N_4615,N_4695);
xor UO_791 (O_791,N_4897,N_4390);
nand UO_792 (O_792,N_3089,N_3136);
nor UO_793 (O_793,N_3441,N_2926);
nand UO_794 (O_794,N_3791,N_3075);
xor UO_795 (O_795,N_4621,N_3268);
xnor UO_796 (O_796,N_4950,N_3105);
nor UO_797 (O_797,N_4111,N_4996);
and UO_798 (O_798,N_4740,N_2664);
nor UO_799 (O_799,N_4908,N_3508);
nor UO_800 (O_800,N_4142,N_2706);
nand UO_801 (O_801,N_3329,N_3423);
and UO_802 (O_802,N_3190,N_4330);
xor UO_803 (O_803,N_4757,N_3140);
or UO_804 (O_804,N_3661,N_3211);
and UO_805 (O_805,N_3827,N_2580);
and UO_806 (O_806,N_3731,N_3925);
nor UO_807 (O_807,N_3988,N_4995);
nor UO_808 (O_808,N_4338,N_4682);
or UO_809 (O_809,N_4152,N_4858);
or UO_810 (O_810,N_2635,N_3413);
or UO_811 (O_811,N_3908,N_3209);
and UO_812 (O_812,N_3442,N_3647);
and UO_813 (O_813,N_4173,N_4069);
and UO_814 (O_814,N_4395,N_3829);
and UO_815 (O_815,N_4689,N_3659);
and UO_816 (O_816,N_2571,N_4676);
or UO_817 (O_817,N_3047,N_4058);
nand UO_818 (O_818,N_3306,N_3878);
xnor UO_819 (O_819,N_4068,N_3098);
nor UO_820 (O_820,N_3036,N_2790);
nor UO_821 (O_821,N_4587,N_3031);
nor UO_822 (O_822,N_2924,N_4001);
xnor UO_823 (O_823,N_3600,N_4308);
xnor UO_824 (O_824,N_4916,N_2748);
and UO_825 (O_825,N_3787,N_3672);
and UO_826 (O_826,N_4180,N_4928);
nor UO_827 (O_827,N_2560,N_3565);
and UO_828 (O_828,N_3455,N_2605);
nor UO_829 (O_829,N_4233,N_3013);
nand UO_830 (O_830,N_3765,N_2574);
xor UO_831 (O_831,N_2874,N_4373);
and UO_832 (O_832,N_2500,N_3313);
nand UO_833 (O_833,N_3903,N_3285);
xnor UO_834 (O_834,N_3108,N_2529);
nor UO_835 (O_835,N_4769,N_2781);
and UO_836 (O_836,N_2776,N_2621);
nor UO_837 (O_837,N_4257,N_4101);
nand UO_838 (O_838,N_3051,N_4623);
nor UO_839 (O_839,N_3617,N_4898);
nand UO_840 (O_840,N_4585,N_4212);
nand UO_841 (O_841,N_4903,N_3448);
and UO_842 (O_842,N_3068,N_4434);
nor UO_843 (O_843,N_3474,N_4209);
nor UO_844 (O_844,N_3367,N_3636);
nor UO_845 (O_845,N_2821,N_4261);
or UO_846 (O_846,N_3450,N_2684);
nand UO_847 (O_847,N_4467,N_3472);
nor UO_848 (O_848,N_4061,N_4333);
nor UO_849 (O_849,N_3623,N_2693);
and UO_850 (O_850,N_2636,N_3776);
or UO_851 (O_851,N_4294,N_3067);
nand UO_852 (O_852,N_3926,N_3755);
xnor UO_853 (O_853,N_4786,N_3947);
xnor UO_854 (O_854,N_2567,N_3044);
nand UO_855 (O_855,N_2936,N_4878);
nand UO_856 (O_856,N_3987,N_3003);
and UO_857 (O_857,N_2658,N_4864);
nor UO_858 (O_858,N_4172,N_4581);
nand UO_859 (O_859,N_4704,N_3824);
nor UO_860 (O_860,N_2981,N_4259);
nor UO_861 (O_861,N_2719,N_4875);
nor UO_862 (O_862,N_4705,N_2579);
nand UO_863 (O_863,N_4873,N_2592);
or UO_864 (O_864,N_3082,N_2835);
and UO_865 (O_865,N_3444,N_2627);
and UO_866 (O_866,N_2972,N_4299);
nor UO_867 (O_867,N_3056,N_4263);
nand UO_868 (O_868,N_3663,N_2663);
and UO_869 (O_869,N_4203,N_4576);
and UO_870 (O_870,N_3109,N_4360);
nor UO_871 (O_871,N_4316,N_4193);
nor UO_872 (O_872,N_2923,N_3464);
xor UO_873 (O_873,N_4918,N_4788);
nor UO_874 (O_874,N_2564,N_3839);
or UO_875 (O_875,N_3055,N_3381);
nand UO_876 (O_876,N_3409,N_4829);
nand UO_877 (O_877,N_4098,N_4386);
and UO_878 (O_878,N_4387,N_4896);
and UO_879 (O_879,N_4035,N_3864);
nor UO_880 (O_880,N_4334,N_4595);
and UO_881 (O_881,N_4351,N_3038);
nand UO_882 (O_882,N_3957,N_4337);
nor UO_883 (O_883,N_3753,N_2810);
nor UO_884 (O_884,N_3761,N_3264);
and UO_885 (O_885,N_3375,N_3521);
or UO_886 (O_886,N_2939,N_2967);
and UO_887 (O_887,N_4501,N_3000);
nand UO_888 (O_888,N_3151,N_3226);
and UO_889 (O_889,N_4717,N_4500);
or UO_890 (O_890,N_2626,N_3513);
xor UO_891 (O_891,N_3552,N_4680);
and UO_892 (O_892,N_4353,N_4876);
and UO_893 (O_893,N_4555,N_3717);
and UO_894 (O_894,N_4120,N_4400);
or UO_895 (O_895,N_3980,N_3107);
xor UO_896 (O_896,N_4645,N_4199);
nor UO_897 (O_897,N_4482,N_4116);
nor UO_898 (O_898,N_4544,N_3586);
or UO_899 (O_899,N_2615,N_3155);
and UO_900 (O_900,N_2612,N_2767);
xnor UO_901 (O_901,N_4284,N_2867);
and UO_902 (O_902,N_3781,N_3538);
nor UO_903 (O_903,N_2691,N_3873);
nand UO_904 (O_904,N_3562,N_4726);
or UO_905 (O_905,N_3667,N_3204);
or UO_906 (O_906,N_4735,N_4036);
and UO_907 (O_907,N_2978,N_3531);
nand UO_908 (O_908,N_2671,N_3099);
nand UO_909 (O_909,N_3682,N_4730);
and UO_910 (O_910,N_3943,N_2541);
and UO_911 (O_911,N_3399,N_3223);
and UO_912 (O_912,N_2666,N_4734);
and UO_913 (O_913,N_4578,N_2920);
nor UO_914 (O_914,N_3550,N_4450);
or UO_915 (O_915,N_3879,N_3886);
nand UO_916 (O_916,N_2948,N_2725);
nand UO_917 (O_917,N_3502,N_4668);
nor UO_918 (O_918,N_3648,N_4747);
nand UO_919 (O_919,N_4165,N_3557);
xnor UO_920 (O_920,N_3985,N_3962);
nor UO_921 (O_921,N_3159,N_3007);
nand UO_922 (O_922,N_2673,N_4463);
xor UO_923 (O_923,N_4067,N_4649);
nor UO_924 (O_924,N_2957,N_3825);
xnor UO_925 (O_925,N_3040,N_3598);
nor UO_926 (O_926,N_4779,N_4140);
nor UO_927 (O_927,N_3797,N_3262);
and UO_928 (O_928,N_2701,N_2511);
or UO_929 (O_929,N_3480,N_2833);
nor UO_930 (O_930,N_3201,N_3937);
nand UO_931 (O_931,N_4577,N_3269);
or UO_932 (O_932,N_3960,N_4546);
nand UO_933 (O_933,N_3999,N_4954);
nor UO_934 (O_934,N_3416,N_4202);
nand UO_935 (O_935,N_2878,N_4108);
nand UO_936 (O_936,N_3596,N_4093);
or UO_937 (O_937,N_4562,N_4859);
or UO_938 (O_938,N_3289,N_4941);
nor UO_939 (O_939,N_4809,N_3149);
nand UO_940 (O_940,N_2539,N_3554);
nor UO_941 (O_941,N_3278,N_4729);
nand UO_942 (O_942,N_4540,N_4239);
xnor UO_943 (O_943,N_4840,N_3130);
nor UO_944 (O_944,N_3191,N_4572);
xnor UO_945 (O_945,N_4796,N_4179);
nand UO_946 (O_946,N_3915,N_2966);
or UO_947 (O_947,N_4422,N_3070);
or UO_948 (O_948,N_4016,N_4992);
nor UO_949 (O_949,N_3265,N_3354);
and UO_950 (O_950,N_4971,N_2823);
xor UO_951 (O_951,N_3470,N_2609);
nand UO_952 (O_952,N_2865,N_3308);
xnor UO_953 (O_953,N_2561,N_3884);
nor UO_954 (O_954,N_4364,N_3121);
and UO_955 (O_955,N_4499,N_3512);
nor UO_956 (O_956,N_3543,N_3742);
nor UO_957 (O_957,N_3711,N_4551);
xor UO_958 (O_958,N_2785,N_4432);
nand UO_959 (O_959,N_3709,N_2877);
or UO_960 (O_960,N_3042,N_3900);
or UO_961 (O_961,N_4369,N_2803);
and UO_962 (O_962,N_2509,N_3654);
nand UO_963 (O_963,N_4529,N_3424);
and UO_964 (O_964,N_2905,N_4934);
nand UO_965 (O_965,N_4238,N_3759);
and UO_966 (O_966,N_4975,N_2783);
nor UO_967 (O_967,N_3978,N_3813);
or UO_968 (O_968,N_3335,N_3097);
nand UO_969 (O_969,N_4177,N_4744);
xnor UO_970 (O_970,N_3434,N_4700);
nor UO_971 (O_971,N_2929,N_4637);
and UO_972 (O_972,N_4217,N_4686);
nand UO_973 (O_973,N_4243,N_4589);
and UO_974 (O_974,N_2704,N_3779);
xnor UO_975 (O_975,N_4973,N_4138);
nand UO_976 (O_976,N_2676,N_2765);
xnor UO_977 (O_977,N_2686,N_2993);
and UO_978 (O_978,N_3275,N_4418);
or UO_979 (O_979,N_4999,N_3119);
nand UO_980 (O_980,N_3028,N_2570);
nand UO_981 (O_981,N_3871,N_3004);
nor UO_982 (O_982,N_2618,N_3730);
or UO_983 (O_983,N_4951,N_2602);
or UO_984 (O_984,N_3735,N_3353);
nor UO_985 (O_985,N_3193,N_2889);
nand UO_986 (O_986,N_3342,N_2562);
or UO_987 (O_987,N_4712,N_2738);
or UO_988 (O_988,N_3650,N_3393);
nor UO_989 (O_989,N_4991,N_3852);
and UO_990 (O_990,N_4026,N_4131);
and UO_991 (O_991,N_4246,N_2709);
and UO_992 (O_992,N_2714,N_4748);
nand UO_993 (O_993,N_4817,N_2769);
or UO_994 (O_994,N_2953,N_2630);
nand UO_995 (O_995,N_2507,N_4889);
nand UO_996 (O_996,N_3386,N_4404);
nand UO_997 (O_997,N_4863,N_3528);
and UO_998 (O_998,N_2698,N_2670);
nand UO_999 (O_999,N_4342,N_3941);
endmodule