module basic_2000_20000_2500_25_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nand U0 (N_0,In_677,In_319);
or U1 (N_1,In_289,In_329);
and U2 (N_2,In_450,In_656);
or U3 (N_3,In_1095,In_160);
nand U4 (N_4,In_179,In_1336);
or U5 (N_5,In_1052,In_771);
or U6 (N_6,In_103,In_731);
nor U7 (N_7,In_609,In_899);
and U8 (N_8,In_1508,In_1833);
and U9 (N_9,In_1427,In_933);
xnor U10 (N_10,In_353,In_1730);
and U11 (N_11,In_1039,In_1432);
and U12 (N_12,In_119,In_682);
nand U13 (N_13,In_1641,In_589);
xnor U14 (N_14,In_424,In_146);
or U15 (N_15,In_565,In_243);
or U16 (N_16,In_1572,In_1585);
nand U17 (N_17,In_1248,In_1586);
nor U18 (N_18,In_703,In_18);
xnor U19 (N_19,In_960,In_1458);
nor U20 (N_20,In_1822,In_1199);
nor U21 (N_21,In_988,In_952);
nand U22 (N_22,In_1081,In_1546);
nand U23 (N_23,In_72,In_554);
nor U24 (N_24,In_1009,In_549);
nor U25 (N_25,In_1754,In_1204);
xnor U26 (N_26,In_1741,In_645);
nand U27 (N_27,In_1459,In_1973);
nand U28 (N_28,In_1981,In_1088);
and U29 (N_29,In_1571,In_903);
or U30 (N_30,In_1467,In_1104);
xnor U31 (N_31,In_1715,In_620);
or U32 (N_32,In_520,In_1147);
nand U33 (N_33,In_576,In_1817);
nor U34 (N_34,In_485,In_1538);
xnor U35 (N_35,In_762,In_1513);
nor U36 (N_36,In_754,In_1232);
or U37 (N_37,In_1835,In_1540);
xnor U38 (N_38,In_744,In_764);
xnor U39 (N_39,In_1672,In_1728);
and U40 (N_40,In_1289,In_1486);
nor U41 (N_41,In_702,In_522);
xnor U42 (N_42,In_937,In_1396);
and U43 (N_43,In_971,In_1062);
nor U44 (N_44,In_1316,In_1587);
and U45 (N_45,In_990,In_281);
nand U46 (N_46,In_743,In_157);
and U47 (N_47,In_1605,In_1071);
xor U48 (N_48,In_77,In_1383);
xor U49 (N_49,In_679,In_241);
nor U50 (N_50,In_951,In_732);
xnor U51 (N_51,In_524,In_1620);
nor U52 (N_52,In_330,In_367);
xnor U53 (N_53,In_1602,In_1043);
or U54 (N_54,In_507,In_1610);
nor U55 (N_55,In_253,In_807);
nor U56 (N_56,In_1580,In_368);
nor U57 (N_57,In_151,In_908);
or U58 (N_58,In_1409,In_1826);
nor U59 (N_59,In_815,In_1420);
nor U60 (N_60,In_130,In_1665);
xor U61 (N_61,In_1435,In_1193);
and U62 (N_62,In_700,In_847);
nor U63 (N_63,In_1830,In_844);
nor U64 (N_64,In_1206,In_787);
nor U65 (N_65,In_1123,In_356);
nand U66 (N_66,In_757,In_427);
xnor U67 (N_67,In_1405,In_285);
xor U68 (N_68,In_291,In_1058);
xor U69 (N_69,In_1891,In_715);
nand U70 (N_70,In_1170,In_1178);
nand U71 (N_71,In_148,In_1213);
nand U72 (N_72,In_850,In_347);
and U73 (N_73,In_704,In_102);
nand U74 (N_74,In_409,In_1113);
nor U75 (N_75,In_1331,In_88);
nand U76 (N_76,In_261,In_803);
or U77 (N_77,In_768,In_606);
xnor U78 (N_78,In_1977,In_931);
or U79 (N_79,In_67,In_949);
nand U80 (N_80,In_1898,In_1385);
nand U81 (N_81,In_328,In_813);
xor U82 (N_82,In_1463,In_523);
or U83 (N_83,In_9,In_1839);
nand U84 (N_84,In_1687,In_115);
and U85 (N_85,In_1475,In_1288);
or U86 (N_86,In_1964,In_76);
and U87 (N_87,In_766,In_1812);
xor U88 (N_88,In_1311,In_598);
and U89 (N_89,In_602,In_597);
and U90 (N_90,In_1386,In_379);
nor U91 (N_91,In_1746,In_265);
nand U92 (N_92,In_63,In_840);
nor U93 (N_93,In_1425,In_1258);
nor U94 (N_94,In_529,In_294);
or U95 (N_95,In_1134,In_939);
nor U96 (N_96,In_519,In_1483);
xor U97 (N_97,In_1364,In_61);
xnor U98 (N_98,In_790,In_1266);
nand U99 (N_99,In_249,In_1411);
and U100 (N_100,In_1517,In_1324);
or U101 (N_101,In_1367,In_1647);
xor U102 (N_102,In_1196,In_1584);
nor U103 (N_103,In_1806,In_438);
or U104 (N_104,In_852,In_23);
and U105 (N_105,In_1956,In_1033);
xnor U106 (N_106,In_239,In_87);
nand U107 (N_107,In_1124,In_1706);
or U108 (N_108,In_479,In_675);
nor U109 (N_109,In_1775,In_380);
or U110 (N_110,In_1923,In_1855);
nand U111 (N_111,In_1582,In_145);
or U112 (N_112,In_1748,In_1673);
xor U113 (N_113,In_987,In_1328);
nand U114 (N_114,In_517,In_767);
and U115 (N_115,In_162,In_1980);
and U116 (N_116,In_1892,In_513);
nor U117 (N_117,In_1278,In_68);
xor U118 (N_118,In_1360,In_1086);
xor U119 (N_119,In_372,In_1184);
xor U120 (N_120,In_64,In_1410);
and U121 (N_121,In_1355,In_45);
or U122 (N_122,In_1859,In_1257);
nor U123 (N_123,In_1623,In_439);
nor U124 (N_124,In_1187,In_366);
nand U125 (N_125,In_591,In_678);
xnor U126 (N_126,In_1177,In_1281);
and U127 (N_127,In_363,In_1828);
nand U128 (N_128,In_1708,In_301);
nor U129 (N_129,In_1814,In_378);
xnor U130 (N_130,In_318,In_20);
and U131 (N_131,In_575,In_1998);
and U132 (N_132,In_494,In_240);
xor U133 (N_133,In_599,In_1496);
and U134 (N_134,In_12,In_1210);
xor U135 (N_135,In_968,In_935);
nor U136 (N_136,In_1153,In_1029);
xor U137 (N_137,In_891,In_1389);
and U138 (N_138,In_1918,In_1046);
or U139 (N_139,In_1938,In_296);
nor U140 (N_140,In_770,In_642);
or U141 (N_141,In_706,In_460);
or U142 (N_142,In_1294,In_1987);
nand U143 (N_143,In_459,In_644);
xnor U144 (N_144,In_1900,In_653);
or U145 (N_145,In_1909,In_396);
nand U146 (N_146,In_1890,In_1293);
and U147 (N_147,In_1295,In_568);
and U148 (N_148,In_49,In_564);
and U149 (N_149,In_1151,In_622);
nor U150 (N_150,In_587,In_1116);
nand U151 (N_151,In_426,In_863);
and U152 (N_152,In_1704,In_1303);
and U153 (N_153,In_810,In_540);
xor U154 (N_154,In_1152,In_569);
nor U155 (N_155,In_462,In_1207);
nand U156 (N_156,In_917,In_997);
and U157 (N_157,In_545,In_1035);
or U158 (N_158,In_1406,In_583);
xor U159 (N_159,In_637,In_1698);
xnor U160 (N_160,In_1764,In_71);
or U161 (N_161,In_1504,In_884);
nand U162 (N_162,In_1310,In_672);
and U163 (N_163,In_1108,In_1651);
nand U164 (N_164,In_1543,In_1209);
nor U165 (N_165,In_1725,In_785);
nand U166 (N_166,In_1001,In_550);
and U167 (N_167,In_324,In_862);
and U168 (N_168,In_259,In_335);
and U169 (N_169,In_1276,In_1143);
xor U170 (N_170,In_106,In_267);
nand U171 (N_171,In_1264,In_1531);
and U172 (N_172,In_295,In_1352);
and U173 (N_173,In_1417,In_34);
and U174 (N_174,In_432,In_616);
xnor U175 (N_175,In_487,In_342);
or U176 (N_176,In_1073,In_410);
nor U177 (N_177,In_1963,In_1597);
or U178 (N_178,In_1723,In_475);
and U179 (N_179,In_1302,In_974);
or U180 (N_180,In_1041,In_390);
and U181 (N_181,In_167,In_729);
and U182 (N_182,In_947,In_633);
and U183 (N_183,In_761,In_1809);
and U184 (N_184,In_360,In_256);
nand U185 (N_185,In_1524,In_447);
or U186 (N_186,In_1785,In_1888);
or U187 (N_187,In_871,In_1707);
nand U188 (N_188,In_73,In_796);
and U189 (N_189,In_1811,In_463);
and U190 (N_190,In_1896,In_1864);
xor U191 (N_191,In_870,In_1881);
nand U192 (N_192,In_1493,In_1093);
nand U193 (N_193,In_758,In_1136);
nor U194 (N_194,In_1721,In_824);
and U195 (N_195,In_1755,In_999);
nand U196 (N_196,In_639,In_1569);
nand U197 (N_197,In_1150,In_1115);
nand U198 (N_198,In_1823,In_443);
or U199 (N_199,In_1091,In_1479);
nor U200 (N_200,In_1004,In_629);
or U201 (N_201,In_1323,In_492);
nand U202 (N_202,In_1300,In_506);
and U203 (N_203,In_1022,In_1766);
or U204 (N_204,In_1819,In_1270);
or U205 (N_205,In_340,In_797);
and U206 (N_206,In_1173,In_825);
nor U207 (N_207,In_407,In_1622);
or U208 (N_208,In_571,In_1915);
nand U209 (N_209,In_214,In_478);
nor U210 (N_210,In_229,In_287);
or U211 (N_211,In_1846,In_536);
nand U212 (N_212,In_1244,In_880);
nand U213 (N_213,In_901,In_1101);
xnor U214 (N_214,In_906,In_1959);
and U215 (N_215,In_538,In_1922);
xor U216 (N_216,In_521,In_1606);
or U217 (N_217,In_283,In_1590);
and U218 (N_218,In_1481,In_322);
or U219 (N_219,In_781,In_1130);
and U220 (N_220,In_1473,In_1533);
or U221 (N_221,In_1221,In_472);
nor U222 (N_222,In_890,In_775);
nor U223 (N_223,In_313,In_1263);
and U224 (N_224,In_1714,In_1110);
xor U225 (N_225,In_1502,In_331);
or U226 (N_226,In_1445,In_1327);
and U227 (N_227,In_858,In_1953);
or U228 (N_228,In_694,In_165);
nand U229 (N_229,In_236,In_1433);
nor U230 (N_230,In_1333,In_1906);
nor U231 (N_231,In_708,In_636);
nand U232 (N_232,In_1374,In_1464);
nand U233 (N_233,In_975,In_1015);
nand U234 (N_234,In_39,In_1026);
and U235 (N_235,In_47,In_1735);
and U236 (N_236,In_801,In_865);
or U237 (N_237,In_250,In_1060);
xnor U238 (N_238,In_1985,In_1008);
nor U239 (N_239,In_1949,In_941);
and U240 (N_240,In_210,In_965);
nand U241 (N_241,In_829,In_1802);
and U242 (N_242,In_627,In_65);
xnor U243 (N_243,In_446,In_1972);
or U244 (N_244,In_1391,In_1373);
nand U245 (N_245,In_1231,In_1522);
nand U246 (N_246,In_486,In_1684);
or U247 (N_247,In_31,In_375);
or U248 (N_248,In_437,In_269);
nand U249 (N_249,In_730,In_878);
nor U250 (N_250,In_1681,In_725);
and U251 (N_251,In_1075,In_1089);
or U252 (N_252,In_1003,In_126);
and U253 (N_253,In_535,In_1349);
xor U254 (N_254,In_36,In_1913);
nor U255 (N_255,In_274,In_1051);
nand U256 (N_256,In_430,In_1028);
and U257 (N_257,In_1379,In_452);
nand U258 (N_258,In_784,In_371);
nor U259 (N_259,In_1381,In_307);
and U260 (N_260,In_384,In_1233);
xor U261 (N_261,In_147,In_1719);
nor U262 (N_262,In_1343,In_352);
and U263 (N_263,In_503,In_1678);
and U264 (N_264,In_1872,In_1511);
xnor U265 (N_265,In_741,In_1924);
and U266 (N_266,In_348,In_1514);
or U267 (N_267,In_1534,In_936);
and U268 (N_268,In_734,In_1198);
nor U269 (N_269,In_212,In_433);
and U270 (N_270,In_640,In_817);
or U271 (N_271,In_1808,In_1422);
nor U272 (N_272,In_687,In_1774);
or U273 (N_273,In_1220,In_1960);
xnor U274 (N_274,In_816,In_1176);
nand U275 (N_275,In_41,In_1611);
and U276 (N_276,In_448,In_772);
xnor U277 (N_277,In_125,In_1350);
nor U278 (N_278,In_266,In_733);
nand U279 (N_279,In_1717,In_1377);
nand U280 (N_280,In_418,In_861);
and U281 (N_281,In_320,In_1224);
nand U282 (N_282,In_288,In_1341);
nand U283 (N_283,In_950,In_1693);
nand U284 (N_284,In_664,In_1287);
xnor U285 (N_285,In_337,In_263);
nand U286 (N_286,In_79,In_1055);
or U287 (N_287,In_1098,In_684);
and U288 (N_288,In_1157,In_834);
xor U289 (N_289,In_495,In_680);
nor U290 (N_290,In_1642,In_831);
xor U291 (N_291,In_1042,In_1132);
xor U292 (N_292,In_1471,In_1813);
nor U293 (N_293,In_794,In_1418);
xnor U294 (N_294,In_195,In_820);
or U295 (N_295,In_1975,In_979);
and U296 (N_296,In_303,In_1125);
or U297 (N_297,In_833,In_1056);
nand U298 (N_298,In_1696,In_873);
and U299 (N_299,In_980,In_805);
nor U300 (N_300,In_465,In_670);
nand U301 (N_301,In_127,In_1709);
or U302 (N_302,In_1625,In_930);
nand U303 (N_303,In_132,In_455);
nor U304 (N_304,In_996,In_74);
and U305 (N_305,In_305,In_1144);
nand U306 (N_306,In_1469,In_1428);
and U307 (N_307,In_46,In_1792);
or U308 (N_308,In_1013,In_783);
and U309 (N_309,In_1731,In_1592);
nor U310 (N_310,In_1279,In_1771);
nand U311 (N_311,In_894,In_1549);
nand U312 (N_312,In_1186,In_117);
xor U313 (N_313,In_1273,In_932);
and U314 (N_314,In_235,In_1114);
nor U315 (N_315,In_1423,In_1604);
nor U316 (N_316,In_808,In_1416);
or U317 (N_317,In_216,In_1810);
and U318 (N_318,In_774,In_449);
nor U319 (N_319,In_1478,In_864);
or U320 (N_320,In_251,In_481);
nand U321 (N_321,In_1,In_209);
and U322 (N_322,In_1181,In_1019);
or U323 (N_323,In_1850,In_237);
or U324 (N_324,In_89,In_1776);
nor U325 (N_325,In_421,In_621);
or U326 (N_326,In_888,In_525);
or U327 (N_327,In_1883,In_192);
xnor U328 (N_328,In_50,In_60);
nand U329 (N_329,In_1129,In_144);
or U330 (N_330,In_8,In_1105);
nand U331 (N_331,In_1241,In_218);
and U332 (N_332,In_1634,In_856);
and U333 (N_333,In_1908,In_696);
and U334 (N_334,In_1847,In_1635);
nor U335 (N_335,In_848,In_860);
nand U336 (N_336,In_184,In_1803);
xor U337 (N_337,In_1402,In_1163);
nor U338 (N_338,In_1050,In_128);
nor U339 (N_339,In_791,In_1756);
or U340 (N_340,In_1548,In_809);
nand U341 (N_341,In_13,In_362);
xor U342 (N_342,In_139,In_1120);
or U343 (N_343,In_516,In_596);
nor U344 (N_344,In_1370,In_542);
nor U345 (N_345,In_812,In_1205);
xor U346 (N_346,In_1702,In_818);
nor U347 (N_347,In_1466,In_1137);
xor U348 (N_348,In_713,In_1138);
nand U349 (N_349,In_155,In_1260);
nor U350 (N_350,In_647,In_1457);
or U351 (N_351,In_1397,In_961);
xnor U352 (N_352,In_1061,In_976);
nand U353 (N_353,In_1139,In_1485);
nand U354 (N_354,In_993,In_193);
xor U355 (N_355,In_1919,In_1660);
xor U356 (N_356,In_95,In_1939);
xnor U357 (N_357,In_84,In_1948);
or U358 (N_358,In_793,In_55);
nand U359 (N_359,In_755,In_1069);
nand U360 (N_360,In_62,In_1037);
xnor U361 (N_361,In_491,In_518);
xor U362 (N_362,In_345,In_918);
nand U363 (N_363,In_1099,In_1412);
nand U364 (N_364,In_1577,In_1542);
nand U365 (N_365,In_1000,In_1145);
xor U366 (N_366,In_257,In_1309);
and U367 (N_367,In_532,In_1886);
nand U368 (N_368,In_1259,In_1955);
or U369 (N_369,In_1269,In_412);
nor U370 (N_370,In_215,In_35);
or U371 (N_371,In_1904,In_1284);
nand U372 (N_372,In_1109,In_323);
xnor U373 (N_373,In_1195,In_1525);
nor U374 (N_374,In_879,In_1413);
nor U375 (N_375,In_207,In_293);
and U376 (N_376,In_534,In_314);
nand U377 (N_377,In_1995,In_1646);
or U378 (N_378,In_1166,In_304);
nor U379 (N_379,In_185,In_1640);
xor U380 (N_380,In_164,In_1111);
or U381 (N_381,In_1112,In_1768);
nor U382 (N_382,In_116,In_1334);
nor U383 (N_383,In_966,In_1535);
and U384 (N_384,In_255,In_1873);
xnor U385 (N_385,In_1994,In_1280);
nor U386 (N_386,In_618,In_721);
and U387 (N_387,In_502,In_1690);
xnor U388 (N_388,In_1361,In_1047);
xor U389 (N_389,In_1313,In_1645);
xnor U390 (N_390,In_1197,In_1976);
and U391 (N_391,In_1487,In_1871);
or U392 (N_392,In_377,In_559);
or U393 (N_393,In_198,In_1371);
and U394 (N_394,In_1758,In_248);
or U395 (N_395,In_150,In_1650);
and U396 (N_396,In_252,In_466);
nand U397 (N_397,In_1285,In_714);
nand U398 (N_398,In_83,In_1638);
nand U399 (N_399,In_302,In_1308);
nand U400 (N_400,In_814,In_909);
nor U401 (N_401,In_1796,In_1807);
nand U402 (N_402,In_282,In_1330);
xnor U403 (N_403,In_14,In_928);
nor U404 (N_404,In_1038,In_381);
or U405 (N_405,In_1880,In_1668);
xnor U406 (N_406,In_44,In_638);
or U407 (N_407,In_1786,In_1214);
nor U408 (N_408,In_1724,In_1040);
nor U409 (N_409,In_399,In_910);
xnor U410 (N_410,In_468,In_1100);
nor U411 (N_411,In_799,In_919);
xor U412 (N_412,In_1729,In_349);
and U413 (N_413,In_121,In_436);
xor U414 (N_414,In_228,In_1434);
nor U415 (N_415,In_557,In_417);
and U416 (N_416,In_1793,In_1789);
nand U417 (N_417,In_469,In_1921);
xor U418 (N_418,In_1993,In_32);
or U419 (N_419,In_386,In_1399);
or U420 (N_420,In_792,In_99);
nor U421 (N_421,In_582,In_1765);
or U422 (N_422,In_511,In_1320);
or U423 (N_423,In_1282,In_226);
nand U424 (N_424,In_1866,In_1378);
xor U425 (N_425,In_70,In_355);
or U426 (N_426,In_1201,In_977);
nand U427 (N_427,In_1146,In_1984);
nand U428 (N_428,In_290,In_956);
nand U429 (N_429,In_1107,In_1601);
nor U430 (N_430,In_722,In_1652);
nand U431 (N_431,In_1523,In_38);
xnor U432 (N_432,In_53,In_1854);
nand U433 (N_433,In_1421,In_1682);
nor U434 (N_434,In_1031,In_1318);
xnor U435 (N_435,In_1074,In_510);
nor U436 (N_436,In_134,In_509);
nand U437 (N_437,In_254,In_312);
and U438 (N_438,In_658,In_854);
nand U439 (N_439,In_382,In_1470);
nor U440 (N_440,In_1217,In_649);
nand U441 (N_441,In_998,In_1154);
nor U442 (N_442,In_1226,In_1692);
nand U443 (N_443,In_619,In_1261);
and U444 (N_444,In_1718,In_666);
and U445 (N_445,In_1080,In_777);
and U446 (N_446,In_660,In_1740);
nand U447 (N_447,In_78,In_1680);
and U448 (N_448,In_912,In_881);
nor U449 (N_449,In_1363,In_346);
nor U450 (N_450,In_1321,In_1551);
and U451 (N_451,In_1727,In_836);
or U452 (N_452,In_1893,In_1907);
nand U453 (N_453,In_1700,In_234);
xor U454 (N_454,In_556,In_58);
xor U455 (N_455,In_1618,In_539);
nand U456 (N_456,In_477,In_140);
nor U457 (N_457,In_720,In_1011);
xor U458 (N_458,In_563,In_152);
nor U459 (N_459,In_659,In_1797);
nand U460 (N_460,In_635,In_668);
and U461 (N_461,In_357,In_911);
nand U462 (N_462,In_625,In_258);
nand U463 (N_463,In_868,In_1431);
and U464 (N_464,In_1372,In_1856);
nor U465 (N_465,In_1347,In_1503);
or U466 (N_466,In_172,In_92);
nand U467 (N_467,In_482,In_650);
or U468 (N_468,In_1745,In_415);
xor U469 (N_469,In_686,In_1547);
nand U470 (N_470,In_779,In_1843);
or U471 (N_471,In_1490,In_268);
and U472 (N_472,In_222,In_1663);
and U473 (N_473,In_1667,In_1895);
nor U474 (N_474,In_1553,In_1818);
nor U475 (N_475,In_1390,In_1770);
nor U476 (N_476,In_1720,In_1501);
nor U477 (N_477,In_1865,In_719);
and U478 (N_478,In_364,In_838);
nand U479 (N_479,In_1928,In_505);
and U480 (N_480,In_711,In_1694);
and U481 (N_481,In_821,In_1030);
or U482 (N_482,In_661,In_105);
or U483 (N_483,In_1131,In_365);
xnor U484 (N_484,In_1229,In_1165);
nor U485 (N_485,In_351,In_336);
and U486 (N_486,In_1510,In_875);
or U487 (N_487,In_978,In_1581);
and U488 (N_488,In_1455,In_1012);
xnor U489 (N_489,In_1169,In_1978);
xor U490 (N_490,In_1526,In_1674);
nand U491 (N_491,In_1262,In_42);
and U492 (N_492,In_1317,In_1057);
nor U493 (N_493,In_1376,In_855);
or U494 (N_494,In_897,In_749);
nor U495 (N_495,In_16,In_1219);
xor U496 (N_496,In_19,In_1801);
nor U497 (N_497,In_1699,In_1512);
nand U498 (N_498,In_773,In_199);
or U499 (N_499,In_343,In_851);
nand U500 (N_500,In_1600,In_1782);
xnor U501 (N_501,In_562,In_311);
nand U502 (N_502,In_107,In_789);
nor U503 (N_503,In_1852,In_1899);
nand U504 (N_504,In_332,In_1747);
xnor U505 (N_505,In_819,In_727);
nand U506 (N_506,In_857,In_1988);
nor U507 (N_507,In_444,In_1827);
and U508 (N_508,In_769,In_1816);
xnor U509 (N_509,In_1480,In_1362);
nand U510 (N_510,In_402,In_1676);
or U511 (N_511,In_270,In_849);
and U512 (N_512,In_1240,In_484);
or U513 (N_513,In_1783,In_1049);
nor U514 (N_514,In_1382,In_1910);
and U515 (N_515,In_1256,In_1439);
nor U516 (N_516,In_138,In_497);
nand U517 (N_517,In_1744,In_1245);
or U518 (N_518,In_286,In_531);
nor U519 (N_519,In_470,In_943);
and U520 (N_520,In_1837,In_921);
or U521 (N_521,In_1286,In_1726);
or U522 (N_522,In_657,In_1944);
and U523 (N_523,In_1495,In_1140);
nand U524 (N_524,In_867,In_1338);
and U525 (N_525,In_142,In_604);
nand U526 (N_526,In_1453,In_1788);
nand U527 (N_527,In_547,In_1966);
nor U528 (N_528,In_944,In_843);
and U529 (N_529,In_953,In_1448);
and U530 (N_530,In_1778,In_723);
nand U531 (N_531,In_1326,In_1067);
or U532 (N_532,In_1474,In_166);
nand U533 (N_533,In_405,In_1820);
nor U534 (N_534,In_986,In_853);
or U535 (N_535,In_317,In_665);
nor U536 (N_536,In_922,In_1934);
xor U537 (N_537,In_1685,In_208);
nand U538 (N_538,In_788,In_300);
nand U539 (N_539,In_1016,In_1175);
nand U540 (N_540,In_1763,In_196);
nor U541 (N_541,In_605,In_994);
or U542 (N_542,In_1753,In_588);
and U543 (N_543,In_1380,In_227);
or U544 (N_544,In_242,In_1017);
nor U545 (N_545,In_308,In_630);
xor U546 (N_546,In_1952,In_846);
or U547 (N_547,In_411,In_1456);
and U548 (N_548,In_1686,In_581);
and U549 (N_549,In_493,In_190);
nor U550 (N_550,In_981,In_276);
nand U551 (N_551,In_1247,In_1243);
and U552 (N_552,In_643,In_498);
xnor U553 (N_553,In_688,In_1312);
nand U554 (N_554,In_738,In_1662);
or U555 (N_555,In_544,In_1624);
nor U556 (N_556,In_1917,In_663);
or U557 (N_557,In_1521,In_530);
nand U558 (N_558,In_1621,In_1767);
nor U559 (N_559,In_1133,In_973);
and U560 (N_560,In_1626,In_1879);
or U561 (N_561,In_1578,In_902);
xnor U562 (N_562,In_1527,In_397);
nor U563 (N_563,In_907,In_223);
and U564 (N_564,In_1999,In_955);
xnor U565 (N_565,In_1957,In_428);
xnor U566 (N_566,In_1387,In_245);
and U567 (N_567,In_1691,In_1465);
nor U568 (N_568,In_1654,In_354);
or U569 (N_569,In_1781,In_648);
and U570 (N_570,In_1616,In_113);
and U571 (N_571,In_59,In_101);
or U572 (N_572,In_392,In_1794);
and U573 (N_573,In_763,In_701);
nor U574 (N_574,In_1838,In_1002);
nand U575 (N_575,In_1078,In_1519);
nand U576 (N_576,In_1943,In_1218);
and U577 (N_577,In_995,In_1161);
or U578 (N_578,In_1780,In_400);
or U579 (N_579,In_654,In_1927);
xor U580 (N_580,In_120,In_188);
nor U581 (N_581,In_1443,In_889);
and U582 (N_582,In_1695,In_326);
nand U583 (N_583,In_24,In_413);
nand U584 (N_584,In_698,In_1940);
and U585 (N_585,In_1158,In_1554);
or U586 (N_586,In_1882,In_938);
or U587 (N_587,In_54,In_641);
nand U588 (N_588,In_262,In_1292);
and U589 (N_589,In_191,In_1969);
or U590 (N_590,In_1595,In_691);
or U591 (N_591,In_1126,In_1395);
nand U592 (N_592,In_1348,In_440);
xor U593 (N_593,In_1965,In_1254);
and U594 (N_594,In_1346,In_1862);
xnor U595 (N_595,In_610,In_233);
xor U596 (N_596,In_1760,In_1054);
or U597 (N_597,In_398,In_623);
or U598 (N_598,In_823,In_601);
xnor U599 (N_599,In_954,In_1593);
and U600 (N_600,In_284,In_33);
nand U601 (N_601,In_1649,In_201);
nor U602 (N_602,In_1267,In_1743);
or U603 (N_603,In_118,In_1345);
and U604 (N_604,In_1945,In_667);
nand U605 (N_605,In_1122,In_592);
or U606 (N_606,In_646,In_874);
xor U607 (N_607,In_454,In_1036);
nor U608 (N_608,In_1627,In_435);
xor U609 (N_609,In_272,In_391);
and U610 (N_610,In_1958,In_5);
nor U611 (N_611,In_527,In_1064);
or U612 (N_612,In_1799,In_1875);
nor U613 (N_613,In_1954,In_709);
and U614 (N_614,In_43,In_972);
nand U615 (N_615,In_1712,In_1732);
xnor U616 (N_616,In_674,In_1222);
xnor U617 (N_617,In_1555,In_887);
nor U618 (N_618,In_1162,In_501);
and U619 (N_619,In_1815,In_934);
xor U620 (N_620,In_1507,In_558);
or U621 (N_621,In_989,In_1738);
nor U622 (N_622,In_175,In_203);
xor U623 (N_623,In_1983,In_1096);
and U624 (N_624,In_181,In_561);
nand U625 (N_625,In_182,In_80);
xor U626 (N_626,In_171,In_1561);
xor U627 (N_627,In_1191,In_1669);
nor U628 (N_628,In_1941,In_798);
and U629 (N_629,In_1857,In_1291);
nand U630 (N_630,In_1946,In_1772);
or U631 (N_631,In_1171,In_1576);
nor U632 (N_632,In_946,In_992);
nor U633 (N_633,In_90,In_483);
nand U634 (N_634,In_48,In_219);
nor U635 (N_635,In_280,In_552);
xnor U636 (N_636,In_1034,In_1203);
and U637 (N_637,In_1583,In_309);
and U638 (N_638,In_776,In_123);
nor U639 (N_639,In_1683,In_1032);
nor U640 (N_640,In_244,In_1018);
nand U641 (N_641,In_1020,In_29);
and U642 (N_642,In_1566,In_149);
or U643 (N_643,In_197,In_1023);
nand U644 (N_644,In_299,In_835);
nand U645 (N_645,In_705,In_726);
xnor U646 (N_646,In_1190,In_156);
and U647 (N_647,In_94,In_1394);
xnor U648 (N_648,In_1619,In_1407);
and U649 (N_649,In_1167,In_10);
nand U650 (N_650,In_1200,In_1798);
nor U651 (N_651,In_1460,In_877);
or U652 (N_652,In_315,In_1550);
xnor U653 (N_653,In_260,In_566);
and U654 (N_654,In_278,In_1500);
or U655 (N_655,In_480,In_1188);
and U656 (N_656,In_1202,In_238);
nand U657 (N_657,In_1446,In_1436);
xnor U658 (N_658,In_983,In_1183);
xor U659 (N_659,In_1449,In_316);
or U660 (N_660,In_133,In_1148);
nand U661 (N_661,In_756,In_1440);
nor U662 (N_662,In_1306,In_1516);
and U663 (N_663,In_1916,In_350);
nor U664 (N_664,In_1869,In_628);
or U665 (N_665,In_374,In_499);
xnor U666 (N_666,In_1863,In_442);
nor U667 (N_667,In_111,In_963);
or U668 (N_668,In_325,In_40);
or U669 (N_669,In_1488,In_129);
or U670 (N_670,In_692,In_1118);
xnor U671 (N_671,In_1588,In_1025);
or U672 (N_672,In_1824,In_1530);
xor U673 (N_673,In_1250,In_514);
xor U674 (N_674,In_1461,In_298);
xnor U675 (N_675,In_608,In_1567);
or U676 (N_676,In_689,In_1845);
nor U677 (N_677,In_204,In_573);
or U678 (N_678,In_1679,In_1357);
xor U679 (N_679,In_1414,In_508);
nor U680 (N_680,In_1990,In_6);
nand U681 (N_681,In_1769,In_441);
and U682 (N_682,In_1565,In_496);
nand U683 (N_683,In_822,In_408);
nor U684 (N_684,In_388,In_590);
or U685 (N_685,In_473,In_1734);
and U686 (N_686,In_1024,In_612);
and U687 (N_687,In_1298,In_1563);
nand U688 (N_688,In_1441,In_1442);
and U689 (N_689,In_231,In_1570);
xnor U690 (N_690,In_1903,In_1403);
or U691 (N_691,In_1914,In_1598);
nor U692 (N_692,In_1805,In_488);
and U693 (N_693,In_1825,In_914);
nand U694 (N_694,In_895,In_991);
nor U695 (N_695,In_872,In_178);
or U696 (N_696,In_1437,In_1991);
nand U697 (N_697,In_1947,In_724);
nand U698 (N_698,In_177,In_1520);
and U699 (N_699,In_143,In_1630);
nand U700 (N_700,In_1613,In_1450);
nor U701 (N_701,In_1185,In_1239);
or U702 (N_702,In_112,In_1053);
nor U703 (N_703,In_1761,In_1784);
or U704 (N_704,In_1426,In_1935);
and U705 (N_705,In_420,In_1609);
xnor U706 (N_706,In_1636,In_603);
or U707 (N_707,In_1629,In_1705);
and U708 (N_708,In_1083,In_1415);
xor U709 (N_709,In_104,In_1800);
nand U710 (N_710,In_750,In_1697);
nand U711 (N_711,In_389,In_586);
xnor U712 (N_712,In_567,In_297);
nor U713 (N_713,In_1424,In_740);
nand U714 (N_714,In_1141,In_737);
and U715 (N_715,In_383,In_802);
nand U716 (N_716,In_806,In_964);
xnor U717 (N_717,In_334,In_1579);
or U718 (N_718,In_742,In_1102);
and U719 (N_719,In_69,In_1614);
nor U720 (N_720,In_1885,In_1063);
nand U721 (N_721,In_1268,In_1494);
or U722 (N_722,In_736,In_1290);
or U723 (N_723,In_141,In_1452);
and U724 (N_724,In_1354,In_1097);
nand U725 (N_725,In_86,In_4);
xor U726 (N_726,In_1006,In_611);
xnor U727 (N_727,In_699,In_1388);
nand U728 (N_728,In_327,In_180);
nor U729 (N_729,In_51,In_1305);
nand U730 (N_730,In_273,In_1762);
and U731 (N_731,In_456,In_537);
or U732 (N_732,In_1164,In_1359);
xnor U733 (N_733,In_458,In_292);
and U734 (N_734,In_339,In_1322);
nand U735 (N_735,In_1670,In_1821);
nor U736 (N_736,In_173,In_707);
nor U737 (N_737,In_414,In_896);
xnor U738 (N_738,In_1677,In_1779);
nor U739 (N_739,In_1556,In_1643);
nor U740 (N_740,In_394,In_135);
and U741 (N_741,In_595,In_1518);
nand U742 (N_742,In_1575,In_3);
and U743 (N_743,In_1860,In_114);
or U744 (N_744,In_28,In_153);
xor U745 (N_745,In_341,In_1274);
or U746 (N_746,In_7,In_1631);
or U747 (N_747,In_1489,In_1045);
and U748 (N_748,In_685,In_1119);
and U749 (N_749,In_1849,In_423);
nor U750 (N_750,In_1180,In_1216);
nor U751 (N_751,In_445,In_306);
xnor U752 (N_752,In_1401,In_338);
nand U753 (N_753,In_669,In_1255);
xnor U754 (N_754,In_1014,In_969);
xor U755 (N_755,In_925,In_1589);
nand U756 (N_756,In_461,In_1238);
nor U757 (N_757,In_213,In_1315);
xnor U758 (N_758,In_898,In_369);
xor U759 (N_759,In_577,In_916);
and U760 (N_760,In_224,In_170);
nor U761 (N_761,In_310,In_555);
and U762 (N_762,In_913,In_403);
nor U763 (N_763,In_1982,In_1319);
nor U764 (N_764,In_1876,In_1369);
nand U765 (N_765,In_1749,In_1509);
nand U766 (N_766,In_1861,In_1454);
or U767 (N_767,In_1633,In_1968);
nand U768 (N_768,In_22,In_1942);
and U769 (N_769,In_617,In_75);
nand U770 (N_770,In_800,In_1393);
nor U771 (N_771,In_457,In_1848);
nor U772 (N_772,In_1536,In_1648);
and U773 (N_773,In_474,In_1703);
nor U774 (N_774,In_886,In_885);
and U775 (N_775,In_220,In_489);
xor U776 (N_776,In_560,In_673);
or U777 (N_777,In_526,In_778);
xor U778 (N_778,In_652,In_1544);
nor U779 (N_779,In_1552,In_1832);
or U780 (N_780,In_137,In_1836);
and U781 (N_781,In_631,In_982);
nor U782 (N_782,In_1644,In_161);
or U783 (N_783,In_464,In_804);
nand U784 (N_784,In_21,In_759);
xor U785 (N_785,In_1666,In_1568);
nand U786 (N_786,In_169,In_1121);
nor U787 (N_787,In_1573,In_1079);
xnor U788 (N_788,In_1742,In_230);
xnor U789 (N_789,In_551,In_1777);
or U790 (N_790,In_1737,In_1252);
nand U791 (N_791,In_923,In_1375);
xor U792 (N_792,In_1932,In_515);
nand U793 (N_793,In_1392,In_1591);
nand U794 (N_794,In_404,In_1599);
or U795 (N_795,In_1926,In_1106);
xnor U796 (N_796,In_1831,In_615);
nor U797 (N_797,In_187,In_1299);
nand U798 (N_798,In_108,In_1342);
and U799 (N_799,In_1878,In_25);
and U800 (N_800,N_280,In_1059);
or U801 (N_801,N_795,N_574);
and U802 (N_802,N_124,N_113);
or U803 (N_803,N_545,N_207);
xnor U804 (N_804,N_72,In_662);
nor U805 (N_805,N_410,N_705);
or U806 (N_806,N_231,In_984);
or U807 (N_807,In_27,N_390);
nand U808 (N_808,N_402,N_797);
or U809 (N_809,In_1829,In_926);
xor U810 (N_810,N_378,N_301);
and U811 (N_811,N_631,In_1841);
or U812 (N_812,N_74,N_125);
and U813 (N_813,In_1366,In_96);
nor U814 (N_814,N_381,N_152);
and U815 (N_815,N_311,In_1307);
and U816 (N_816,N_541,N_44);
nor U817 (N_817,In_1159,N_588);
and U818 (N_818,N_189,N_341);
and U819 (N_819,N_165,N_518);
and U820 (N_820,N_772,N_23);
and U821 (N_821,N_391,N_676);
and U822 (N_822,N_211,N_289);
and U823 (N_823,In_66,In_174);
nand U824 (N_824,N_149,N_208);
nor U825 (N_825,N_548,N_491);
or U826 (N_826,N_375,N_363);
or U827 (N_827,N_210,In_1404);
xnor U828 (N_828,In_1265,N_270);
and U829 (N_829,In_504,N_203);
or U830 (N_830,N_786,N_53);
xor U831 (N_831,N_420,N_720);
nand U832 (N_832,N_340,N_319);
nor U833 (N_833,N_285,N_19);
and U834 (N_834,N_568,In_828);
xnor U835 (N_835,N_334,N_40);
or U836 (N_836,N_130,In_1068);
and U837 (N_837,N_546,N_489);
nor U838 (N_838,N_513,N_724);
nand U839 (N_839,N_741,N_443);
nand U840 (N_840,In_827,N_694);
nor U841 (N_841,N_729,In_1594);
and U842 (N_842,N_217,N_10);
nand U843 (N_843,N_182,In_893);
nor U844 (N_844,N_672,N_653);
or U845 (N_845,N_734,In_1048);
or U846 (N_846,N_793,In_1358);
or U847 (N_847,In_1867,N_121);
or U848 (N_848,N_241,N_179);
or U849 (N_849,In_548,N_542);
and U850 (N_850,N_445,N_364);
or U851 (N_851,In_594,N_214);
nor U852 (N_852,N_138,N_582);
nand U853 (N_853,N_222,N_605);
nor U854 (N_854,In_543,N_232);
and U855 (N_855,In_11,N_302);
and U856 (N_856,N_461,N_630);
nor U857 (N_857,In_1329,In_1007);
nand U858 (N_858,N_181,N_209);
nor U859 (N_859,In_1438,N_100);
or U860 (N_860,N_481,In_1804);
xor U861 (N_861,N_749,In_1174);
or U862 (N_862,N_354,In_1902);
nand U863 (N_863,N_62,In_1072);
nand U864 (N_864,N_350,N_34);
or U865 (N_865,N_712,N_487);
or U866 (N_866,N_530,N_661);
or U867 (N_867,N_384,N_106);
or U868 (N_868,N_246,In_1211);
and U869 (N_869,N_145,In_1314);
nor U870 (N_870,In_1537,N_187);
nand U871 (N_871,N_117,In_1103);
xor U872 (N_872,N_348,In_1562);
nor U873 (N_873,N_33,In_1897);
and U874 (N_874,N_439,N_306);
nor U875 (N_875,N_460,In_205);
xnor U876 (N_876,N_502,In_1532);
and U877 (N_877,In_200,In_1795);
xor U878 (N_878,N_769,In_866);
xor U879 (N_879,N_13,In_211);
nor U880 (N_880,N_477,In_376);
and U881 (N_881,N_110,N_14);
or U882 (N_882,In_760,In_924);
xor U883 (N_883,N_66,N_333);
or U884 (N_884,N_26,In_1603);
and U885 (N_885,N_36,N_560);
xor U886 (N_886,N_421,In_1655);
nor U887 (N_887,In_395,In_1970);
xnor U888 (N_888,N_466,N_558);
and U889 (N_889,In_1889,N_139);
or U890 (N_890,N_90,N_383);
xnor U891 (N_891,N_673,In_1858);
nand U892 (N_892,N_35,N_514);
nor U893 (N_893,In_735,N_433);
and U894 (N_894,N_748,N_611);
and U895 (N_895,N_59,N_308);
and U896 (N_896,In_710,In_1564);
and U897 (N_897,N_483,N_414);
and U898 (N_898,In_739,N_595);
nor U899 (N_899,In_1304,In_632);
nor U900 (N_900,N_604,N_430);
nand U901 (N_901,N_455,In_915);
or U902 (N_902,N_18,In_1997);
or U903 (N_903,N_282,N_409);
and U904 (N_904,N_96,In_900);
nor U905 (N_905,N_213,In_1870);
and U906 (N_906,N_654,In_1671);
xor U907 (N_907,N_664,In_1628);
or U908 (N_908,N_55,N_642);
or U909 (N_909,N_95,In_1251);
nor U910 (N_910,In_905,In_782);
nor U911 (N_911,In_1065,N_407);
nand U912 (N_912,In_837,N_474);
nor U913 (N_913,N_718,In_985);
or U914 (N_914,N_256,In_811);
nand U915 (N_915,N_767,N_320);
nor U916 (N_916,N_756,N_1);
nand U917 (N_917,In_97,N_388);
or U918 (N_918,N_504,N_198);
and U919 (N_919,In_1653,N_269);
nor U920 (N_920,In_1127,N_501);
and U921 (N_921,N_295,In_194);
or U922 (N_922,In_1541,N_12);
xnor U923 (N_923,N_730,In_30);
or U924 (N_924,In_1444,N_665);
nor U925 (N_925,In_159,N_0);
nor U926 (N_926,N_658,In_1505);
nand U927 (N_927,N_326,N_297);
and U928 (N_928,N_669,N_431);
xor U929 (N_929,N_580,In_1750);
nor U930 (N_930,In_1951,N_5);
nand U931 (N_931,In_1142,In_1656);
and U932 (N_932,N_190,N_250);
xor U933 (N_933,N_399,In_1851);
nand U934 (N_934,In_56,In_1710);
xnor U935 (N_935,N_111,N_359);
xnor U936 (N_936,In_359,In_1228);
nand U937 (N_937,N_163,N_16);
nand U938 (N_938,N_238,N_509);
nand U939 (N_939,N_778,N_37);
nand U940 (N_940,In_163,N_277);
nand U941 (N_941,N_54,N_395);
or U942 (N_942,N_463,N_162);
nor U943 (N_943,In_344,N_361);
and U944 (N_944,N_294,In_361);
and U945 (N_945,In_1283,N_393);
nand U946 (N_946,N_212,N_325);
or U947 (N_947,N_742,N_87);
nand U948 (N_948,N_651,N_98);
nor U949 (N_949,N_794,N_257);
nor U950 (N_950,In_614,N_752);
nand U951 (N_951,In_1277,In_37);
or U952 (N_952,N_147,In_1739);
nor U953 (N_953,N_740,N_493);
xnor U954 (N_954,In_579,In_948);
and U955 (N_955,N_609,N_271);
nand U956 (N_956,N_382,In_1498);
nor U957 (N_957,In_1296,N_726);
and U958 (N_958,In_1557,N_183);
nand U959 (N_959,In_15,In_1757);
nand U960 (N_960,N_150,In_1661);
xor U961 (N_961,N_429,N_775);
nand U962 (N_962,N_578,N_615);
nor U963 (N_963,In_1230,N_400);
nand U964 (N_964,N_456,N_178);
and U965 (N_965,N_692,N_68);
nor U966 (N_966,N_397,In_401);
nand U967 (N_967,N_567,In_1325);
and U968 (N_968,N_312,In_546);
xnor U969 (N_969,In_1451,N_675);
nand U970 (N_970,N_143,In_279);
nor U971 (N_971,In_676,N_529);
and U972 (N_972,In_1155,In_1149);
or U973 (N_973,N_172,N_127);
nand U974 (N_974,N_99,In_1736);
nand U975 (N_975,In_1344,In_681);
nand U976 (N_976,N_368,N_589);
and U977 (N_977,In_1077,In_962);
nand U978 (N_978,N_685,N_176);
and U979 (N_979,N_787,In_712);
or U980 (N_980,N_571,N_188);
and U981 (N_981,N_649,In_1874);
nand U982 (N_982,N_781,N_531);
or U983 (N_983,N_374,In_1608);
nor U984 (N_984,In_1182,In_1911);
nor U985 (N_985,N_744,In_1168);
xor U986 (N_986,In_1884,N_251);
or U987 (N_987,N_660,N_423);
and U988 (N_988,In_387,N_97);
or U989 (N_989,In_1468,N_335);
xor U990 (N_990,N_782,N_362);
and U991 (N_991,In_626,N_373);
nand U992 (N_992,N_617,N_329);
or U993 (N_993,In_247,N_69);
xnor U994 (N_994,N_495,N_677);
xor U995 (N_995,In_1722,In_1986);
and U996 (N_996,N_556,N_314);
xnor U997 (N_997,In_82,N_655);
xor U998 (N_998,N_620,In_1967);
nor U999 (N_999,N_750,N_614);
nor U1000 (N_1000,N_528,N_695);
or U1001 (N_1001,In_1447,N_161);
nor U1002 (N_1002,N_602,N_291);
nand U1003 (N_1003,N_102,In_1172);
nor U1004 (N_1004,In_1716,N_634);
nand U1005 (N_1005,In_110,In_1194);
and U1006 (N_1006,N_703,N_237);
or U1007 (N_1007,N_20,In_957);
and U1008 (N_1008,N_79,N_169);
nand U1009 (N_1009,In_264,N_129);
nor U1010 (N_1010,N_324,In_1961);
xor U1011 (N_1011,N_27,N_157);
and U1012 (N_1012,N_6,N_56);
nand U1013 (N_1013,N_643,N_435);
and U1014 (N_1014,In_98,N_520);
and U1015 (N_1015,In_57,N_592);
nand U1016 (N_1016,In_1950,N_698);
nor U1017 (N_1017,In_1472,N_245);
or U1018 (N_1018,In_1933,N_64);
nor U1019 (N_1019,In_613,In_920);
xor U1020 (N_1020,In_1339,In_1539);
xnor U1021 (N_1021,N_472,In_490);
nor U1022 (N_1022,In_186,In_929);
xor U1023 (N_1023,N_349,In_1615);
or U1024 (N_1024,N_31,In_876);
and U1025 (N_1025,N_77,In_904);
and U1026 (N_1026,In_1607,N_753);
xor U1027 (N_1027,N_141,N_638);
xor U1028 (N_1028,In_1506,In_1021);
xnor U1029 (N_1029,N_315,In_1353);
or U1030 (N_1030,N_156,In_1901);
and U1031 (N_1031,N_597,N_136);
nor U1032 (N_1032,In_1419,In_1223);
or U1033 (N_1033,In_624,In_217);
and U1034 (N_1034,In_1497,In_651);
xnor U1035 (N_1035,In_131,In_1082);
xor U1036 (N_1036,N_464,N_151);
or U1037 (N_1037,N_667,N_709);
or U1038 (N_1038,In_471,N_777);
xor U1039 (N_1039,N_173,N_690);
or U1040 (N_1040,In_1246,N_764);
nor U1041 (N_1041,In_1790,In_1773);
and U1042 (N_1042,In_600,N_264);
nand U1043 (N_1043,N_446,N_158);
nor U1044 (N_1044,N_401,N_467);
and U1045 (N_1045,N_674,In_1094);
nand U1046 (N_1046,N_263,N_790);
nor U1047 (N_1047,In_1275,N_680);
or U1048 (N_1048,N_532,In_1688);
nand U1049 (N_1049,N_688,N_339);
and U1050 (N_1050,In_1384,N_784);
nor U1051 (N_1051,N_716,In_1117);
and U1052 (N_1052,N_259,N_248);
nand U1053 (N_1053,In_1545,N_155);
and U1054 (N_1054,In_1840,In_52);
or U1055 (N_1055,N_755,N_229);
nand U1056 (N_1056,In_434,N_305);
nor U1057 (N_1057,N_197,N_475);
nor U1058 (N_1058,N_91,N_547);
xnor U1059 (N_1059,N_357,N_253);
nor U1060 (N_1060,In_832,N_450);
nor U1061 (N_1061,In_845,N_613);
xnor U1062 (N_1062,In_1894,In_533);
or U1063 (N_1063,N_22,N_17);
and U1064 (N_1064,In_183,In_1558);
xnor U1065 (N_1065,N_70,N_544);
nor U1066 (N_1066,N_449,In_1429);
nand U1067 (N_1067,In_1905,N_134);
or U1068 (N_1068,N_180,N_83);
and U1069 (N_1069,N_496,N_606);
nor U1070 (N_1070,In_1010,N_171);
nor U1071 (N_1071,In_842,In_752);
xnor U1072 (N_1072,N_583,N_780);
nor U1073 (N_1073,N_488,N_243);
or U1074 (N_1074,N_219,N_590);
xnor U1075 (N_1075,N_337,In_728);
and U1076 (N_1076,N_132,N_550);
nor U1077 (N_1077,N_510,N_133);
nor U1078 (N_1078,In_945,N_57);
nand U1079 (N_1079,In_1160,N_566);
xnor U1080 (N_1080,In_765,N_476);
or U1081 (N_1081,N_385,In_1476);
and U1082 (N_1082,N_516,N_771);
and U1083 (N_1083,In_1398,In_1484);
and U1084 (N_1084,N_146,N_426);
and U1085 (N_1085,N_494,N_697);
or U1086 (N_1086,In_580,N_785);
xnor U1087 (N_1087,N_153,N_32);
nand U1088 (N_1088,N_81,In_892);
or U1089 (N_1089,In_500,In_85);
nor U1090 (N_1090,In_1492,In_1225);
nand U1091 (N_1091,N_46,In_1632);
and U1092 (N_1092,N_168,N_45);
nand U1093 (N_1093,In_453,N_118);
and U1094 (N_1094,N_108,N_268);
nand U1095 (N_1095,N_733,N_265);
nor U1096 (N_1096,In_753,N_338);
and U1097 (N_1097,N_540,N_63);
nor U1098 (N_1098,In_839,In_1574);
nand U1099 (N_1099,In_1085,N_766);
or U1100 (N_1100,N_300,N_612);
or U1101 (N_1101,N_38,N_668);
xnor U1102 (N_1102,N_278,N_227);
and U1103 (N_1103,In_1066,In_585);
and U1104 (N_1104,N_763,N_292);
xnor U1105 (N_1105,N_367,N_369);
or U1106 (N_1106,N_313,In_1235);
or U1107 (N_1107,N_506,In_1087);
nand U1108 (N_1108,N_719,In_958);
nor U1109 (N_1109,N_714,N_48);
xnor U1110 (N_1110,In_225,N_629);
xor U1111 (N_1111,N_663,In_277);
nand U1112 (N_1112,N_737,N_296);
xnor U1113 (N_1113,N_204,In_584);
xor U1114 (N_1114,N_577,In_1657);
nand U1115 (N_1115,N_279,In_1937);
xnor U1116 (N_1116,In_1559,N_93);
xnor U1117 (N_1117,N_184,N_115);
nand U1118 (N_1118,In_1877,In_1135);
nand U1119 (N_1119,In_1242,In_275);
nand U1120 (N_1120,N_307,N_576);
nand U1121 (N_1121,N_86,N_343);
xor U1122 (N_1122,N_418,N_538);
nand U1123 (N_1123,In_1400,N_281);
xnor U1124 (N_1124,In_393,N_225);
nand U1125 (N_1125,In_697,In_1027);
or U1126 (N_1126,N_42,In_2);
xnor U1127 (N_1127,N_796,N_174);
nor U1128 (N_1128,In_221,N_600);
nand U1129 (N_1129,N_41,In_512);
nor U1130 (N_1130,N_406,N_75);
xor U1131 (N_1131,N_377,N_262);
nor U1132 (N_1132,N_164,N_621);
xnor U1133 (N_1133,In_1787,N_193);
xor U1134 (N_1134,N_486,N_167);
and U1135 (N_1135,N_536,In_1301);
nor U1136 (N_1136,In_17,N_273);
and U1137 (N_1137,In_786,N_671);
nor U1138 (N_1138,In_1844,N_773);
and U1139 (N_1139,In_1936,In_1658);
nor U1140 (N_1140,N_128,N_109);
nor U1141 (N_1141,In_690,In_373);
nand U1142 (N_1142,N_727,N_747);
nor U1143 (N_1143,N_116,N_586);
xnor U1144 (N_1144,In_1925,In_942);
xor U1145 (N_1145,N_230,N_266);
nor U1146 (N_1146,N_682,N_559);
nor U1147 (N_1147,N_735,N_71);
xnor U1148 (N_1148,In_1368,N_473);
and U1149 (N_1149,N_721,N_618);
and U1150 (N_1150,N_637,N_347);
nor U1151 (N_1151,N_411,N_686);
nand U1152 (N_1152,N_699,N_394);
nor U1153 (N_1153,N_601,N_523);
xor U1154 (N_1154,N_7,In_1234);
nand U1155 (N_1155,N_799,In_122);
xnor U1156 (N_1156,N_783,N_126);
and U1157 (N_1157,N_492,N_666);
and U1158 (N_1158,N_84,N_711);
nor U1159 (N_1159,N_417,N_224);
and U1160 (N_1160,N_317,N_706);
or U1161 (N_1161,N_500,N_353);
and U1162 (N_1162,N_105,N_759);
nor U1163 (N_1163,In_124,N_459);
xor U1164 (N_1164,In_869,In_607);
nand U1165 (N_1165,N_356,N_687);
nor U1166 (N_1166,In_1192,N_607);
or U1167 (N_1167,N_206,N_85);
xor U1168 (N_1168,N_635,N_441);
xor U1169 (N_1169,In_189,In_1005);
and U1170 (N_1170,N_387,In_747);
nor U1171 (N_1171,N_471,N_434);
nand U1172 (N_1172,N_205,In_1084);
nand U1173 (N_1173,In_422,N_585);
nand U1174 (N_1174,In_1711,In_81);
and U1175 (N_1175,N_30,N_526);
and U1176 (N_1176,N_322,N_452);
nor U1177 (N_1177,N_398,N_745);
and U1178 (N_1178,In_1271,N_551);
or U1179 (N_1179,In_1356,N_760);
nand U1180 (N_1180,N_332,In_634);
or U1181 (N_1181,N_424,In_959);
nor U1182 (N_1182,N_776,N_573);
and U1183 (N_1183,N_365,N_379);
or U1184 (N_1184,In_553,N_587);
and U1185 (N_1185,N_581,N_754);
or U1186 (N_1186,N_515,In_1751);
and U1187 (N_1187,N_233,N_372);
xor U1188 (N_1188,N_58,N_564);
xor U1189 (N_1189,In_671,N_195);
or U1190 (N_1190,N_440,N_722);
xnor U1191 (N_1191,N_342,N_235);
nand U1192 (N_1192,In_158,In_91);
nor U1193 (N_1193,N_683,N_226);
and U1194 (N_1194,N_554,N_521);
and U1195 (N_1195,In_1499,In_1208);
xnor U1196 (N_1196,N_624,N_318);
or U1197 (N_1197,N_49,N_701);
or U1198 (N_1198,N_533,N_380);
nor U1199 (N_1199,In_1477,N_287);
or U1200 (N_1200,In_1297,N_249);
or U1201 (N_1201,In_718,N_284);
or U1202 (N_1202,N_689,N_28);
xor U1203 (N_1203,In_202,N_330);
or U1204 (N_1204,N_625,N_267);
nand U1205 (N_1205,N_107,N_479);
or U1206 (N_1206,N_645,In_1491);
and U1207 (N_1207,N_484,N_360);
nor U1208 (N_1208,N_779,N_82);
nand U1209 (N_1209,N_24,N_275);
nor U1210 (N_1210,N_469,In_109);
and U1211 (N_1211,N_221,N_9);
and U1212 (N_1212,In_419,In_406);
nand U1213 (N_1213,N_331,In_859);
nand U1214 (N_1214,In_1639,N_623);
or U1215 (N_1215,N_639,N_732);
nor U1216 (N_1216,N_371,In_1215);
nor U1217 (N_1217,N_696,In_830);
nor U1218 (N_1218,N_29,N_8);
or U1219 (N_1219,N_681,N_572);
xnor U1220 (N_1220,N_298,N_316);
nand U1221 (N_1221,N_557,N_52);
nor U1222 (N_1222,N_261,N_490);
and U1223 (N_1223,N_344,N_199);
or U1224 (N_1224,In_1070,N_154);
nor U1225 (N_1225,In_967,In_826);
or U1226 (N_1226,N_355,N_43);
nor U1227 (N_1227,In_1090,N_196);
or U1228 (N_1228,N_700,In_385);
nand U1229 (N_1229,In_1733,In_528);
nand U1230 (N_1230,In_1335,N_140);
and U1231 (N_1231,N_370,N_525);
and U1232 (N_1232,N_562,N_608);
and U1233 (N_1233,N_186,In_882);
nand U1234 (N_1234,N_470,N_148);
nand U1235 (N_1235,N_101,In_1689);
xnor U1236 (N_1236,In_333,N_254);
nor U1237 (N_1237,N_765,N_413);
and U1238 (N_1238,N_236,N_462);
xor U1239 (N_1239,In_1637,N_570);
or U1240 (N_1240,In_1962,N_239);
xor U1241 (N_1241,In_1701,N_553);
or U1242 (N_1242,In_1332,N_404);
nand U1243 (N_1243,In_1931,N_192);
and U1244 (N_1244,N_142,N_626);
and U1245 (N_1245,In_1272,N_392);
nand U1246 (N_1246,N_216,N_499);
and U1247 (N_1247,N_537,N_603);
and U1248 (N_1248,N_512,In_425);
or U1249 (N_1249,N_438,N_622);
and U1250 (N_1250,N_112,N_791);
and U1251 (N_1251,N_647,In_1365);
nand U1252 (N_1252,N_67,In_1253);
nor U1253 (N_1253,N_761,In_572);
nor U1254 (N_1254,N_223,N_628);
xor U1255 (N_1255,In_1791,N_166);
and U1256 (N_1256,N_274,In_1092);
nand U1257 (N_1257,N_323,In_232);
nor U1258 (N_1258,N_757,N_276);
nor U1259 (N_1259,N_565,N_480);
and U1260 (N_1260,In_883,N_684);
or U1261 (N_1261,In_1128,N_122);
nand U1262 (N_1262,N_746,N_92);
or U1263 (N_1263,In_970,N_774);
or U1264 (N_1264,N_743,In_1249);
xor U1265 (N_1265,In_154,N_412);
and U1266 (N_1266,In_321,N_731);
or U1267 (N_1267,In_716,N_691);
xnor U1268 (N_1268,N_498,N_534);
nor U1269 (N_1269,N_713,N_228);
or U1270 (N_1270,N_220,N_563);
nand U1271 (N_1271,N_524,N_200);
or U1272 (N_1272,In_1979,N_159);
nand U1273 (N_1273,In_1992,N_648);
or U1274 (N_1274,N_15,In_841);
and U1275 (N_1275,In_1929,In_93);
nor U1276 (N_1276,N_457,N_652);
or U1277 (N_1277,In_1236,N_619);
xnor U1278 (N_1278,In_246,N_448);
nand U1279 (N_1279,In_100,N_60);
xnor U1280 (N_1280,In_795,N_792);
xor U1281 (N_1281,In_176,N_61);
or U1282 (N_1282,N_3,N_288);
xnor U1283 (N_1283,N_662,N_610);
nor U1284 (N_1284,N_328,N_427);
nor U1285 (N_1285,N_65,N_594);
or U1286 (N_1286,N_646,N_717);
nor U1287 (N_1287,N_693,In_1617);
and U1288 (N_1288,In_1912,N_505);
or U1289 (N_1289,In_593,N_657);
nor U1290 (N_1290,N_591,N_454);
nor U1291 (N_1291,N_405,N_584);
or U1292 (N_1292,N_644,In_370);
xnor U1293 (N_1293,In_1528,N_707);
nand U1294 (N_1294,In_1529,In_940);
xnor U1295 (N_1295,N_656,In_1351);
or U1296 (N_1296,In_1076,N_788);
or U1297 (N_1297,In_136,N_458);
nor U1298 (N_1298,N_659,N_710);
nand U1299 (N_1299,N_389,N_453);
nor U1300 (N_1300,In_358,In_0);
and U1301 (N_1301,N_447,N_194);
and U1302 (N_1302,In_26,N_114);
nand U1303 (N_1303,N_708,In_570);
and U1304 (N_1304,N_599,N_444);
and U1305 (N_1305,In_429,N_4);
or U1306 (N_1306,N_478,N_403);
or U1307 (N_1307,N_352,In_271);
nand U1308 (N_1308,N_511,N_503);
nor U1309 (N_1309,In_780,N_321);
nand U1310 (N_1310,N_351,N_386);
xor U1311 (N_1311,In_1759,In_451);
nand U1312 (N_1312,N_247,In_1430);
nor U1313 (N_1313,In_751,N_73);
or U1314 (N_1314,N_552,N_627);
nor U1315 (N_1315,N_535,N_739);
nand U1316 (N_1316,N_76,N_422);
xnor U1317 (N_1317,In_1462,N_728);
nor U1318 (N_1318,N_290,N_89);
or U1319 (N_1319,In_1227,N_252);
nor U1320 (N_1320,In_206,N_283);
xnor U1321 (N_1321,N_723,N_120);
nand U1322 (N_1322,In_1340,N_650);
nand U1323 (N_1323,N_240,N_2);
nor U1324 (N_1324,In_748,In_1752);
or U1325 (N_1325,N_336,N_497);
and U1326 (N_1326,In_745,In_927);
and U1327 (N_1327,N_346,N_144);
nor U1328 (N_1328,N_303,In_1887);
and U1329 (N_1329,N_215,N_679);
nor U1330 (N_1330,N_242,N_517);
xor U1331 (N_1331,N_451,N_633);
nand U1332 (N_1332,In_168,N_366);
nand U1333 (N_1333,In_1853,In_1408);
and U1334 (N_1334,In_1971,N_80);
nor U1335 (N_1335,In_1212,N_598);
xnor U1336 (N_1336,N_408,In_1337);
nand U1337 (N_1337,N_104,N_304);
xnor U1338 (N_1338,N_425,N_135);
nand U1339 (N_1339,N_636,In_717);
nor U1340 (N_1340,In_1675,N_561);
nor U1341 (N_1341,N_47,N_376);
and U1342 (N_1342,N_555,N_78);
and U1343 (N_1343,N_482,In_693);
or U1344 (N_1344,N_432,N_507);
nor U1345 (N_1345,N_286,N_39);
or U1346 (N_1346,N_640,N_11);
nor U1347 (N_1347,N_575,N_768);
or U1348 (N_1348,N_160,N_272);
xnor U1349 (N_1349,N_468,In_1930);
and U1350 (N_1350,N_770,In_1842);
nand U1351 (N_1351,N_798,In_1044);
nand U1352 (N_1352,N_244,In_1659);
nor U1353 (N_1353,In_467,In_1237);
or U1354 (N_1354,N_442,N_437);
or U1355 (N_1355,N_50,N_201);
xnor U1356 (N_1356,In_1868,N_543);
xor U1357 (N_1357,N_485,In_541);
nand U1358 (N_1358,N_396,In_1612);
xor U1359 (N_1359,N_131,N_51);
and U1360 (N_1360,N_416,In_574);
and U1361 (N_1361,N_345,N_255);
xnor U1362 (N_1362,N_119,N_519);
nand U1363 (N_1363,In_416,N_185);
and U1364 (N_1364,N_202,N_549);
nand U1365 (N_1365,In_1179,N_309);
and U1366 (N_1366,N_704,In_1596);
nand U1367 (N_1367,N_758,In_1834);
xnor U1368 (N_1368,In_1560,In_1664);
and U1369 (N_1369,In_1482,N_88);
nor U1370 (N_1370,N_123,N_299);
xor U1371 (N_1371,N_593,N_736);
nor U1372 (N_1372,In_655,In_746);
or U1373 (N_1373,N_358,N_569);
nand U1374 (N_1374,In_578,In_1989);
nand U1375 (N_1375,In_683,N_137);
xor U1376 (N_1376,N_327,In_1189);
nor U1377 (N_1377,N_170,N_175);
xnor U1378 (N_1378,N_177,N_428);
nand U1379 (N_1379,N_260,N_539);
or U1380 (N_1380,N_596,In_1996);
nand U1381 (N_1381,N_641,N_94);
xnor U1382 (N_1382,N_191,N_527);
and U1383 (N_1383,N_218,N_522);
and U1384 (N_1384,N_508,In_431);
nor U1385 (N_1385,N_21,N_103);
or U1386 (N_1386,N_632,N_234);
nand U1387 (N_1387,In_1515,N_293);
xnor U1388 (N_1388,N_310,N_465);
and U1389 (N_1389,N_25,N_725);
nor U1390 (N_1390,In_476,In_1713);
and U1391 (N_1391,N_670,In_1974);
and U1392 (N_1392,N_738,In_695);
nor U1393 (N_1393,N_762,N_436);
nor U1394 (N_1394,N_415,N_789);
or U1395 (N_1395,N_751,In_1156);
nand U1396 (N_1396,N_715,N_616);
or U1397 (N_1397,N_678,N_419);
nand U1398 (N_1398,N_579,In_1920);
or U1399 (N_1399,N_702,N_258);
xor U1400 (N_1400,N_246,N_274);
nor U1401 (N_1401,N_43,N_71);
nand U1402 (N_1402,In_1246,N_785);
and U1403 (N_1403,N_667,N_455);
or U1404 (N_1404,N_776,In_194);
or U1405 (N_1405,N_289,N_626);
or U1406 (N_1406,N_533,N_449);
xor U1407 (N_1407,N_278,In_1212);
xor U1408 (N_1408,In_159,In_1368);
or U1409 (N_1409,N_6,N_555);
or U1410 (N_1410,N_368,In_574);
and U1411 (N_1411,N_261,N_2);
nor U1412 (N_1412,N_669,In_1713);
nor U1413 (N_1413,N_81,N_258);
and U1414 (N_1414,In_745,N_510);
nor U1415 (N_1415,In_1351,N_657);
nand U1416 (N_1416,In_1149,In_614);
or U1417 (N_1417,In_395,N_199);
and U1418 (N_1418,In_232,N_706);
xor U1419 (N_1419,N_331,In_1253);
nor U1420 (N_1420,N_376,N_178);
nor U1421 (N_1421,In_1419,N_81);
or U1422 (N_1422,In_866,N_11);
nor U1423 (N_1423,N_387,N_2);
nand U1424 (N_1424,N_422,In_52);
or U1425 (N_1425,N_213,N_238);
nor U1426 (N_1426,N_587,N_427);
xnor U1427 (N_1427,In_271,N_623);
nand U1428 (N_1428,N_474,In_37);
or U1429 (N_1429,N_496,N_533);
xor U1430 (N_1430,N_784,N_471);
nand U1431 (N_1431,N_582,N_328);
or U1432 (N_1432,N_173,N_721);
xnor U1433 (N_1433,N_490,N_227);
nand U1434 (N_1434,N_274,N_748);
or U1435 (N_1435,N_129,N_476);
or U1436 (N_1436,In_206,N_165);
and U1437 (N_1437,In_26,N_86);
nand U1438 (N_1438,N_293,In_1688);
nor U1439 (N_1439,N_263,N_422);
nand U1440 (N_1440,N_30,In_1834);
and U1441 (N_1441,N_355,N_387);
xor U1442 (N_1442,N_659,In_1048);
nor U1443 (N_1443,N_470,N_162);
nand U1444 (N_1444,In_584,N_777);
nand U1445 (N_1445,N_648,In_1773);
xnor U1446 (N_1446,In_1353,In_1937);
nor U1447 (N_1447,In_1858,N_686);
or U1448 (N_1448,N_580,N_280);
or U1449 (N_1449,N_204,N_284);
xnor U1450 (N_1450,In_1237,In_26);
nand U1451 (N_1451,N_675,In_1841);
xor U1452 (N_1452,In_543,In_1066);
nor U1453 (N_1453,In_98,In_970);
nor U1454 (N_1454,N_129,In_1066);
xnor U1455 (N_1455,N_236,N_363);
or U1456 (N_1456,In_811,N_59);
xor U1457 (N_1457,N_241,N_605);
xor U1458 (N_1458,In_358,In_1408);
and U1459 (N_1459,In_1332,In_651);
xnor U1460 (N_1460,In_748,In_948);
and U1461 (N_1461,N_568,N_232);
nand U1462 (N_1462,N_761,N_264);
or U1463 (N_1463,In_716,N_312);
nor U1464 (N_1464,N_47,In_546);
and U1465 (N_1465,In_655,In_1658);
or U1466 (N_1466,N_441,In_1297);
nand U1467 (N_1467,N_514,N_629);
or U1468 (N_1468,N_505,N_194);
xor U1469 (N_1469,N_670,In_1007);
xor U1470 (N_1470,N_741,N_129);
nor U1471 (N_1471,N_534,N_701);
nor U1472 (N_1472,N_490,N_668);
nand U1473 (N_1473,In_189,N_311);
nand U1474 (N_1474,N_630,N_583);
nor U1475 (N_1475,In_1751,N_737);
nor U1476 (N_1476,N_463,In_543);
or U1477 (N_1477,N_258,N_294);
nor U1478 (N_1478,N_573,N_211);
nor U1479 (N_1479,N_669,N_214);
or U1480 (N_1480,N_739,In_1182);
xnor U1481 (N_1481,N_477,N_507);
nand U1482 (N_1482,N_541,In_624);
and U1483 (N_1483,In_1558,N_771);
and U1484 (N_1484,In_780,N_251);
xor U1485 (N_1485,In_1979,N_711);
or U1486 (N_1486,N_599,N_350);
and U1487 (N_1487,N_679,N_584);
nand U1488 (N_1488,N_31,N_433);
nor U1489 (N_1489,N_338,N_486);
nor U1490 (N_1490,In_832,In_585);
xor U1491 (N_1491,N_570,In_1325);
or U1492 (N_1492,N_227,N_689);
nand U1493 (N_1493,N_658,N_513);
nor U1494 (N_1494,N_242,In_1759);
nand U1495 (N_1495,N_71,In_940);
nand U1496 (N_1496,N_324,N_566);
and U1497 (N_1497,In_782,N_324);
and U1498 (N_1498,N_333,N_445);
xnor U1499 (N_1499,In_422,N_274);
nor U1500 (N_1500,N_688,N_114);
xor U1501 (N_1501,N_472,In_1242);
or U1502 (N_1502,N_50,N_662);
nand U1503 (N_1503,In_614,In_710);
nand U1504 (N_1504,N_374,N_180);
nor U1505 (N_1505,In_683,N_255);
and U1506 (N_1506,N_24,N_436);
and U1507 (N_1507,N_225,N_610);
nor U1508 (N_1508,In_1297,N_759);
or U1509 (N_1509,N_664,In_1757);
and U1510 (N_1510,N_605,N_229);
or U1511 (N_1511,N_424,N_620);
and U1512 (N_1512,N_615,N_372);
and U1513 (N_1513,N_59,N_781);
nand U1514 (N_1514,N_694,N_418);
nor U1515 (N_1515,N_314,N_692);
nand U1516 (N_1516,N_422,N_736);
and U1517 (N_1517,In_344,N_538);
nand U1518 (N_1518,N_372,In_962);
and U1519 (N_1519,N_624,N_686);
xor U1520 (N_1520,In_1773,N_535);
or U1521 (N_1521,In_984,N_48);
or U1522 (N_1522,N_201,In_1068);
nand U1523 (N_1523,N_398,N_26);
nand U1524 (N_1524,N_402,In_1332);
xor U1525 (N_1525,N_729,N_551);
xor U1526 (N_1526,N_295,N_334);
and U1527 (N_1527,In_1962,N_444);
nand U1528 (N_1528,In_693,N_569);
nor U1529 (N_1529,N_571,N_179);
nor U1530 (N_1530,N_739,N_532);
nand U1531 (N_1531,N_727,In_401);
nor U1532 (N_1532,N_575,N_1);
xor U1533 (N_1533,In_1497,N_256);
nor U1534 (N_1534,N_285,N_436);
or U1535 (N_1535,In_1902,N_110);
xnor U1536 (N_1536,N_510,In_1560);
nand U1537 (N_1537,N_55,In_1841);
xor U1538 (N_1538,N_340,N_741);
and U1539 (N_1539,In_1272,N_585);
xor U1540 (N_1540,N_697,In_97);
nor U1541 (N_1541,N_209,N_704);
or U1542 (N_1542,N_190,N_730);
xnor U1543 (N_1543,N_206,In_1048);
or U1544 (N_1544,N_359,N_198);
and U1545 (N_1545,In_1545,N_298);
or U1546 (N_1546,N_777,N_535);
xor U1547 (N_1547,N_629,N_326);
nand U1548 (N_1548,N_185,N_47);
or U1549 (N_1549,In_1419,N_493);
nor U1550 (N_1550,In_1277,N_325);
or U1551 (N_1551,N_732,N_315);
nor U1552 (N_1552,In_1215,N_323);
xnor U1553 (N_1553,N_634,N_131);
nand U1554 (N_1554,N_779,N_554);
xnor U1555 (N_1555,N_551,In_752);
xnor U1556 (N_1556,N_285,N_530);
nor U1557 (N_1557,N_23,In_795);
and U1558 (N_1558,In_174,In_739);
nand U1559 (N_1559,N_610,N_31);
nand U1560 (N_1560,N_286,N_715);
or U1561 (N_1561,In_1007,In_434);
nor U1562 (N_1562,In_225,In_859);
xnor U1563 (N_1563,N_64,N_90);
or U1564 (N_1564,N_631,N_785);
nand U1565 (N_1565,N_99,In_747);
nand U1566 (N_1566,N_271,N_448);
xnor U1567 (N_1567,N_334,N_73);
or U1568 (N_1568,N_546,N_66);
xnor U1569 (N_1569,N_186,N_103);
nor U1570 (N_1570,In_467,N_659);
nor U1571 (N_1571,N_432,In_904);
nor U1572 (N_1572,In_1076,N_300);
nor U1573 (N_1573,N_420,N_785);
or U1574 (N_1574,N_217,N_466);
and U1575 (N_1575,In_1506,N_162);
nor U1576 (N_1576,N_531,N_682);
nor U1577 (N_1577,N_594,N_278);
or U1578 (N_1578,N_247,N_192);
nor U1579 (N_1579,In_416,N_177);
and U1580 (N_1580,N_196,N_653);
or U1581 (N_1581,In_416,N_40);
and U1582 (N_1582,N_275,In_1661);
and U1583 (N_1583,N_273,N_60);
and U1584 (N_1584,N_380,In_1398);
or U1585 (N_1585,N_594,N_631);
and U1586 (N_1586,In_82,In_929);
and U1587 (N_1587,N_636,In_1477);
or U1588 (N_1588,N_792,N_660);
and U1589 (N_1589,N_124,N_357);
or U1590 (N_1590,N_14,N_499);
and U1591 (N_1591,In_1142,In_613);
or U1592 (N_1592,In_826,N_100);
nor U1593 (N_1593,N_766,N_507);
nor U1594 (N_1594,N_119,N_725);
and U1595 (N_1595,N_664,N_287);
nand U1596 (N_1596,N_333,N_52);
xnor U1597 (N_1597,N_524,N_673);
xor U1598 (N_1598,N_48,N_44);
nor U1599 (N_1599,In_1498,N_624);
nor U1600 (N_1600,N_1587,N_1477);
nand U1601 (N_1601,N_1363,N_1485);
nand U1602 (N_1602,N_1349,N_1436);
and U1603 (N_1603,N_1005,N_1410);
nand U1604 (N_1604,N_1521,N_844);
and U1605 (N_1605,N_1007,N_1448);
or U1606 (N_1606,N_1472,N_1104);
and U1607 (N_1607,N_1434,N_1532);
or U1608 (N_1608,N_952,N_1562);
or U1609 (N_1609,N_1474,N_802);
nand U1610 (N_1610,N_1105,N_1245);
and U1611 (N_1611,N_1298,N_1133);
or U1612 (N_1612,N_1130,N_1328);
xor U1613 (N_1613,N_980,N_833);
and U1614 (N_1614,N_1218,N_1152);
and U1615 (N_1615,N_1422,N_1077);
or U1616 (N_1616,N_1376,N_1356);
and U1617 (N_1617,N_1172,N_1572);
nor U1618 (N_1618,N_1259,N_989);
and U1619 (N_1619,N_843,N_1519);
and U1620 (N_1620,N_1284,N_839);
nand U1621 (N_1621,N_1462,N_1101);
xnor U1622 (N_1622,N_1553,N_870);
or U1623 (N_1623,N_1453,N_1237);
nand U1624 (N_1624,N_1203,N_949);
and U1625 (N_1625,N_907,N_1306);
and U1626 (N_1626,N_1093,N_1407);
nor U1627 (N_1627,N_1252,N_1289);
or U1628 (N_1628,N_1234,N_1095);
and U1629 (N_1629,N_1489,N_1327);
or U1630 (N_1630,N_1466,N_1382);
nor U1631 (N_1631,N_1146,N_1364);
nand U1632 (N_1632,N_937,N_1272);
or U1633 (N_1633,N_1323,N_1311);
nand U1634 (N_1634,N_1182,N_935);
or U1635 (N_1635,N_1230,N_1255);
nor U1636 (N_1636,N_930,N_1401);
xnor U1637 (N_1637,N_1303,N_1269);
and U1638 (N_1638,N_1540,N_1208);
and U1639 (N_1639,N_852,N_1546);
and U1640 (N_1640,N_1568,N_1511);
nor U1641 (N_1641,N_1261,N_938);
or U1642 (N_1642,N_1052,N_982);
nand U1643 (N_1643,N_1174,N_1515);
xnor U1644 (N_1644,N_1461,N_805);
or U1645 (N_1645,N_1342,N_1508);
or U1646 (N_1646,N_1417,N_1447);
nor U1647 (N_1647,N_1374,N_1022);
or U1648 (N_1648,N_1192,N_1025);
or U1649 (N_1649,N_1078,N_1247);
and U1650 (N_1650,N_1340,N_1277);
nor U1651 (N_1651,N_1278,N_1391);
xor U1652 (N_1652,N_979,N_1274);
nor U1653 (N_1653,N_1556,N_943);
or U1654 (N_1654,N_1488,N_871);
or U1655 (N_1655,N_841,N_1563);
or U1656 (N_1656,N_1249,N_1299);
nor U1657 (N_1657,N_1367,N_1501);
xor U1658 (N_1658,N_823,N_940);
nand U1659 (N_1659,N_906,N_1227);
and U1660 (N_1660,N_1313,N_1525);
xor U1661 (N_1661,N_1020,N_1383);
nand U1662 (N_1662,N_1350,N_1431);
or U1663 (N_1663,N_1395,N_969);
and U1664 (N_1664,N_908,N_836);
nor U1665 (N_1665,N_1512,N_1564);
or U1666 (N_1666,N_1074,N_916);
nand U1667 (N_1667,N_1281,N_1111);
and U1668 (N_1668,N_978,N_1345);
xnor U1669 (N_1669,N_992,N_1034);
and U1670 (N_1670,N_1004,N_1045);
or U1671 (N_1671,N_951,N_1483);
xor U1672 (N_1672,N_1221,N_1468);
xnor U1673 (N_1673,N_990,N_1549);
nand U1674 (N_1674,N_1292,N_911);
nand U1675 (N_1675,N_1075,N_1557);
and U1676 (N_1676,N_910,N_1390);
xnor U1677 (N_1677,N_1148,N_876);
and U1678 (N_1678,N_909,N_1479);
nor U1679 (N_1679,N_803,N_1404);
xor U1680 (N_1680,N_882,N_1056);
xnor U1681 (N_1681,N_1484,N_864);
nand U1682 (N_1682,N_1341,N_1150);
nor U1683 (N_1683,N_950,N_1589);
or U1684 (N_1684,N_1571,N_996);
nor U1685 (N_1685,N_1517,N_1217);
xnor U1686 (N_1686,N_945,N_1055);
xor U1687 (N_1687,N_1082,N_1051);
xnor U1688 (N_1688,N_1403,N_1015);
nor U1689 (N_1689,N_1362,N_1091);
xnor U1690 (N_1690,N_1533,N_971);
and U1691 (N_1691,N_821,N_1033);
or U1692 (N_1692,N_1251,N_1547);
and U1693 (N_1693,N_1087,N_1331);
and U1694 (N_1694,N_927,N_1180);
and U1695 (N_1695,N_1348,N_1316);
and U1696 (N_1696,N_1337,N_1595);
nor U1697 (N_1697,N_1302,N_1548);
xor U1698 (N_1698,N_883,N_1239);
xor U1699 (N_1699,N_1165,N_856);
xor U1700 (N_1700,N_1329,N_1013);
nor U1701 (N_1701,N_1469,N_1365);
or U1702 (N_1702,N_1442,N_1144);
nor U1703 (N_1703,N_1042,N_1076);
xor U1704 (N_1704,N_1314,N_1481);
and U1705 (N_1705,N_947,N_923);
nand U1706 (N_1706,N_1153,N_1392);
nor U1707 (N_1707,N_1393,N_926);
xor U1708 (N_1708,N_964,N_1223);
xor U1709 (N_1709,N_1206,N_1565);
nand U1710 (N_1710,N_1355,N_1145);
nand U1711 (N_1711,N_977,N_875);
nand U1712 (N_1712,N_1044,N_1119);
xnor U1713 (N_1713,N_1186,N_1063);
nor U1714 (N_1714,N_1232,N_1072);
or U1715 (N_1715,N_1283,N_1019);
or U1716 (N_1716,N_1575,N_1086);
or U1717 (N_1717,N_965,N_1188);
nand U1718 (N_1718,N_1419,N_1509);
nand U1719 (N_1719,N_1199,N_1377);
nand U1720 (N_1720,N_924,N_1287);
xor U1721 (N_1721,N_1271,N_878);
xnor U1722 (N_1722,N_986,N_970);
xnor U1723 (N_1723,N_958,N_1193);
or U1724 (N_1724,N_1092,N_1071);
nand U1725 (N_1725,N_1433,N_1200);
nor U1726 (N_1726,N_1409,N_860);
nor U1727 (N_1727,N_1372,N_1233);
nand U1728 (N_1728,N_1301,N_1163);
nor U1729 (N_1729,N_1586,N_1458);
nor U1730 (N_1730,N_999,N_810);
and U1731 (N_1731,N_913,N_955);
or U1732 (N_1732,N_1368,N_1369);
and U1733 (N_1733,N_988,N_1324);
nand U1734 (N_1734,N_1585,N_1432);
and U1735 (N_1735,N_894,N_861);
or U1736 (N_1736,N_1495,N_1122);
and U1737 (N_1737,N_942,N_824);
nor U1738 (N_1738,N_1579,N_1094);
nor U1739 (N_1739,N_1293,N_807);
nor U1740 (N_1740,N_1507,N_1260);
or U1741 (N_1741,N_1475,N_1097);
nor U1742 (N_1742,N_1347,N_1225);
xor U1743 (N_1743,N_1139,N_1136);
nand U1744 (N_1744,N_1318,N_892);
and U1745 (N_1745,N_1116,N_1228);
or U1746 (N_1746,N_1574,N_826);
or U1747 (N_1747,N_1543,N_1213);
or U1748 (N_1748,N_983,N_885);
or U1749 (N_1749,N_1142,N_1598);
xnor U1750 (N_1750,N_1351,N_1421);
and U1751 (N_1751,N_1167,N_1343);
nand U1752 (N_1752,N_1229,N_1524);
and U1753 (N_1753,N_1244,N_954);
xnor U1754 (N_1754,N_1099,N_809);
nand U1755 (N_1755,N_1505,N_1439);
xnor U1756 (N_1756,N_1235,N_1427);
nor U1757 (N_1757,N_960,N_1581);
or U1758 (N_1758,N_1336,N_1184);
nor U1759 (N_1759,N_1081,N_828);
or U1760 (N_1760,N_873,N_1420);
or U1761 (N_1761,N_1067,N_936);
xor U1762 (N_1762,N_1147,N_917);
or U1763 (N_1763,N_1242,N_1179);
nor U1764 (N_1764,N_931,N_1010);
nand U1765 (N_1765,N_1268,N_1175);
xnor U1766 (N_1766,N_1236,N_1106);
and U1767 (N_1767,N_1493,N_1135);
or U1768 (N_1768,N_874,N_1330);
nand U1769 (N_1769,N_898,N_1338);
and U1770 (N_1770,N_1522,N_896);
xor U1771 (N_1771,N_1499,N_1513);
and U1772 (N_1772,N_1154,N_1588);
and U1773 (N_1773,N_1321,N_1370);
nor U1774 (N_1774,N_816,N_1064);
nand U1775 (N_1775,N_1123,N_957);
and U1776 (N_1776,N_1412,N_1248);
xnor U1777 (N_1777,N_1118,N_1189);
nand U1778 (N_1778,N_1423,N_1191);
nor U1779 (N_1779,N_1584,N_1357);
or U1780 (N_1780,N_1538,N_1280);
nor U1781 (N_1781,N_1276,N_1240);
and U1782 (N_1782,N_1117,N_974);
and U1783 (N_1783,N_1264,N_1219);
nand U1784 (N_1784,N_1467,N_1109);
xnor U1785 (N_1785,N_1429,N_963);
xor U1786 (N_1786,N_1487,N_1492);
and U1787 (N_1787,N_1541,N_975);
nand U1788 (N_1788,N_877,N_842);
and U1789 (N_1789,N_1202,N_1291);
nor U1790 (N_1790,N_995,N_1282);
nand U1791 (N_1791,N_1378,N_1437);
or U1792 (N_1792,N_1120,N_1465);
xor U1793 (N_1793,N_1576,N_879);
or U1794 (N_1794,N_1346,N_933);
and U1795 (N_1795,N_1426,N_887);
xor U1796 (N_1796,N_1275,N_890);
nor U1797 (N_1797,N_1577,N_1344);
xor U1798 (N_1798,N_1596,N_800);
and U1799 (N_1799,N_1173,N_1195);
xnor U1800 (N_1800,N_1267,N_929);
nand U1801 (N_1801,N_1542,N_1387);
nand U1802 (N_1802,N_811,N_1121);
or U1803 (N_1803,N_851,N_1325);
nor U1804 (N_1804,N_925,N_1161);
nor U1805 (N_1805,N_1386,N_1138);
nor U1806 (N_1806,N_1384,N_1058);
and U1807 (N_1807,N_1534,N_1373);
nand U1808 (N_1808,N_1494,N_1220);
and U1809 (N_1809,N_904,N_1049);
nor U1810 (N_1810,N_1128,N_1100);
or U1811 (N_1811,N_813,N_1389);
xnor U1812 (N_1812,N_1243,N_919);
or U1813 (N_1813,N_862,N_854);
and U1814 (N_1814,N_1198,N_1171);
and U1815 (N_1815,N_1021,N_829);
and U1816 (N_1816,N_1250,N_1226);
and U1817 (N_1817,N_1295,N_899);
and U1818 (N_1818,N_1496,N_1441);
nand U1819 (N_1819,N_900,N_946);
nand U1820 (N_1820,N_1454,N_948);
nand U1821 (N_1821,N_845,N_1204);
xnor U1822 (N_1822,N_1084,N_1270);
or U1823 (N_1823,N_1039,N_1023);
or U1824 (N_1824,N_1594,N_840);
nand U1825 (N_1825,N_1569,N_994);
and U1826 (N_1826,N_1418,N_1523);
and U1827 (N_1827,N_1444,N_959);
xor U1828 (N_1828,N_1134,N_1307);
nand U1829 (N_1829,N_1177,N_944);
xnor U1830 (N_1830,N_1497,N_847);
nand U1831 (N_1831,N_1215,N_1285);
and U1832 (N_1832,N_1408,N_1471);
nor U1833 (N_1833,N_1551,N_1560);
nor U1834 (N_1834,N_1253,N_1246);
nor U1835 (N_1835,N_1539,N_973);
or U1836 (N_1836,N_812,N_855);
xnor U1837 (N_1837,N_1108,N_1416);
and U1838 (N_1838,N_859,N_1405);
nand U1839 (N_1839,N_1222,N_953);
or U1840 (N_1840,N_1414,N_1151);
and U1841 (N_1841,N_1238,N_1181);
xnor U1842 (N_1842,N_1452,N_1070);
nor U1843 (N_1843,N_1290,N_1381);
nor U1844 (N_1844,N_1411,N_1085);
nand U1845 (N_1845,N_1506,N_962);
nand U1846 (N_1846,N_1201,N_1380);
xnor U1847 (N_1847,N_1090,N_1046);
nand U1848 (N_1848,N_991,N_1455);
nand U1849 (N_1849,N_848,N_1354);
and U1850 (N_1850,N_1319,N_1583);
xor U1851 (N_1851,N_1024,N_822);
nand U1852 (N_1852,N_1265,N_1486);
and U1853 (N_1853,N_1555,N_1040);
nand U1854 (N_1854,N_1504,N_1043);
xnor U1855 (N_1855,N_1332,N_1279);
nand U1856 (N_1856,N_997,N_1257);
or U1857 (N_1857,N_1402,N_967);
xor U1858 (N_1858,N_1209,N_830);
nand U1859 (N_1859,N_872,N_1320);
nor U1860 (N_1860,N_1582,N_1141);
and U1861 (N_1861,N_1162,N_1187);
xnor U1862 (N_1862,N_897,N_857);
nor U1863 (N_1863,N_1166,N_1001);
or U1864 (N_1864,N_849,N_1003);
xnor U1865 (N_1865,N_1088,N_1456);
or U1866 (N_1866,N_1322,N_838);
or U1867 (N_1867,N_1176,N_1359);
nor U1868 (N_1868,N_1224,N_1593);
nand U1869 (N_1869,N_934,N_1125);
nand U1870 (N_1870,N_1096,N_1379);
or U1871 (N_1871,N_1459,N_1190);
nor U1872 (N_1872,N_1537,N_1559);
nor U1873 (N_1873,N_1573,N_976);
nand U1874 (N_1874,N_1566,N_1169);
and U1875 (N_1875,N_868,N_1503);
or U1876 (N_1876,N_1527,N_834);
nand U1877 (N_1877,N_837,N_1529);
nand U1878 (N_1878,N_1544,N_1273);
xor U1879 (N_1879,N_1068,N_1254);
and U1880 (N_1880,N_884,N_1413);
and U1881 (N_1881,N_1062,N_1300);
and U1882 (N_1882,N_1490,N_1438);
nor U1883 (N_1883,N_932,N_1590);
or U1884 (N_1884,N_1157,N_1041);
and U1885 (N_1885,N_961,N_972);
nand U1886 (N_1886,N_1140,N_1371);
xor U1887 (N_1887,N_1425,N_1516);
or U1888 (N_1888,N_1578,N_1170);
and U1889 (N_1889,N_1032,N_863);
nor U1890 (N_1890,N_998,N_1388);
xnor U1891 (N_1891,N_1263,N_869);
and U1892 (N_1892,N_1591,N_1057);
or U1893 (N_1893,N_1194,N_1258);
xor U1894 (N_1894,N_956,N_1498);
and U1895 (N_1895,N_1476,N_1183);
nand U1896 (N_1896,N_1478,N_1114);
or U1897 (N_1897,N_914,N_1011);
and U1898 (N_1898,N_1463,N_1143);
and U1899 (N_1899,N_985,N_1210);
xor U1900 (N_1900,N_1335,N_1297);
nand U1901 (N_1901,N_1470,N_818);
and U1902 (N_1902,N_1396,N_920);
nor U1903 (N_1903,N_1031,N_1502);
nand U1904 (N_1904,N_1531,N_1028);
or U1905 (N_1905,N_1030,N_891);
xor U1906 (N_1906,N_1266,N_1443);
xor U1907 (N_1907,N_1083,N_1334);
nor U1908 (N_1908,N_1399,N_1262);
xnor U1909 (N_1909,N_1016,N_1110);
or U1910 (N_1910,N_1164,N_1530);
xnor U1911 (N_1911,N_1103,N_1137);
xor U1912 (N_1912,N_1536,N_1400);
nor U1913 (N_1913,N_902,N_968);
and U1914 (N_1914,N_1149,N_889);
nand U1915 (N_1915,N_1567,N_1446);
or U1916 (N_1916,N_1288,N_1514);
or U1917 (N_1917,N_1286,N_804);
and U1918 (N_1918,N_966,N_939);
nor U1919 (N_1919,N_1445,N_1061);
and U1920 (N_1920,N_1000,N_1113);
or U1921 (N_1921,N_1027,N_1535);
nand U1922 (N_1922,N_1102,N_1360);
nor U1923 (N_1923,N_1552,N_1006);
or U1924 (N_1924,N_1500,N_867);
nor U1925 (N_1925,N_827,N_1449);
nand U1926 (N_1926,N_993,N_1518);
xor U1927 (N_1927,N_928,N_1231);
xor U1928 (N_1928,N_865,N_1214);
nor U1929 (N_1929,N_1066,N_1014);
xnor U1930 (N_1930,N_1304,N_817);
and U1931 (N_1931,N_1440,N_825);
and U1932 (N_1932,N_1385,N_1089);
nor U1933 (N_1933,N_987,N_918);
and U1934 (N_1934,N_1570,N_1333);
nand U1935 (N_1935,N_1315,N_1296);
nand U1936 (N_1936,N_1358,N_886);
xnor U1937 (N_1937,N_1353,N_1361);
nand U1938 (N_1938,N_1415,N_1480);
or U1939 (N_1939,N_881,N_1550);
nand U1940 (N_1940,N_1435,N_1080);
nor U1941 (N_1941,N_1036,N_1491);
xor U1942 (N_1942,N_1129,N_1107);
xnor U1943 (N_1943,N_1178,N_1394);
and U1944 (N_1944,N_1047,N_806);
and U1945 (N_1945,N_808,N_853);
nor U1946 (N_1946,N_1450,N_1305);
or U1947 (N_1947,N_866,N_984);
nand U1948 (N_1948,N_1207,N_1132);
xor U1949 (N_1949,N_1561,N_1256);
or U1950 (N_1950,N_1185,N_1160);
xnor U1951 (N_1951,N_1029,N_1326);
nand U1952 (N_1952,N_1079,N_1464);
and U1953 (N_1953,N_1580,N_1197);
xor U1954 (N_1954,N_1599,N_1060);
nand U1955 (N_1955,N_981,N_915);
and U1956 (N_1956,N_1339,N_1558);
and U1957 (N_1957,N_819,N_1460);
and U1958 (N_1958,N_1430,N_1398);
xnor U1959 (N_1959,N_835,N_801);
nand U1960 (N_1960,N_1312,N_1526);
and U1961 (N_1961,N_912,N_815);
nor U1962 (N_1962,N_1310,N_903);
nand U1963 (N_1963,N_1158,N_1037);
nor U1964 (N_1964,N_1352,N_1159);
nor U1965 (N_1965,N_1196,N_1406);
nor U1966 (N_1966,N_1451,N_1069);
nor U1967 (N_1967,N_1155,N_1592);
and U1968 (N_1968,N_1424,N_1127);
nor U1969 (N_1969,N_888,N_1098);
and U1970 (N_1970,N_1308,N_1012);
nand U1971 (N_1971,N_1126,N_1050);
and U1972 (N_1972,N_1124,N_1241);
or U1973 (N_1973,N_1309,N_858);
or U1974 (N_1974,N_1009,N_831);
nor U1975 (N_1975,N_832,N_1366);
nor U1976 (N_1976,N_1212,N_1375);
nand U1977 (N_1977,N_1317,N_1035);
and U1978 (N_1978,N_1008,N_1002);
xor U1979 (N_1979,N_1073,N_1054);
xor U1980 (N_1980,N_1397,N_1294);
or U1981 (N_1981,N_941,N_905);
or U1982 (N_1982,N_1038,N_1211);
nand U1983 (N_1983,N_1048,N_1428);
or U1984 (N_1984,N_895,N_846);
and U1985 (N_1985,N_1112,N_1059);
and U1986 (N_1986,N_893,N_1018);
or U1987 (N_1987,N_820,N_1205);
or U1988 (N_1988,N_1520,N_1156);
xor U1989 (N_1989,N_1528,N_880);
nor U1990 (N_1990,N_850,N_1115);
xor U1991 (N_1991,N_1053,N_1017);
nand U1992 (N_1992,N_1473,N_1216);
nand U1993 (N_1993,N_1131,N_1510);
nor U1994 (N_1994,N_1554,N_1482);
nor U1995 (N_1995,N_1597,N_1545);
nand U1996 (N_1996,N_1168,N_1457);
or U1997 (N_1997,N_921,N_1065);
xor U1998 (N_1998,N_901,N_1026);
nand U1999 (N_1999,N_814,N_922);
nor U2000 (N_2000,N_1256,N_1407);
and U2001 (N_2001,N_1417,N_964);
and U2002 (N_2002,N_1572,N_884);
or U2003 (N_2003,N_834,N_1041);
or U2004 (N_2004,N_1533,N_1387);
nor U2005 (N_2005,N_973,N_844);
nor U2006 (N_2006,N_1460,N_1044);
or U2007 (N_2007,N_1285,N_1532);
nor U2008 (N_2008,N_949,N_885);
or U2009 (N_2009,N_1095,N_1394);
xnor U2010 (N_2010,N_1226,N_881);
nand U2011 (N_2011,N_1423,N_1208);
nor U2012 (N_2012,N_1556,N_1206);
and U2013 (N_2013,N_1007,N_941);
and U2014 (N_2014,N_1077,N_1466);
nand U2015 (N_2015,N_1564,N_1268);
nor U2016 (N_2016,N_1035,N_1320);
and U2017 (N_2017,N_1526,N_850);
nand U2018 (N_2018,N_944,N_1506);
or U2019 (N_2019,N_1591,N_1215);
xnor U2020 (N_2020,N_1443,N_1403);
or U2021 (N_2021,N_1160,N_1432);
nor U2022 (N_2022,N_1024,N_1392);
and U2023 (N_2023,N_1281,N_960);
xnor U2024 (N_2024,N_950,N_1199);
xnor U2025 (N_2025,N_1098,N_962);
nand U2026 (N_2026,N_1080,N_1410);
xor U2027 (N_2027,N_1233,N_1368);
or U2028 (N_2028,N_918,N_1066);
and U2029 (N_2029,N_1244,N_1327);
nor U2030 (N_2030,N_1359,N_800);
nor U2031 (N_2031,N_1230,N_1527);
nor U2032 (N_2032,N_1405,N_1445);
and U2033 (N_2033,N_1220,N_930);
xor U2034 (N_2034,N_1597,N_887);
and U2035 (N_2035,N_1521,N_1073);
and U2036 (N_2036,N_1218,N_826);
nor U2037 (N_2037,N_1318,N_1280);
nand U2038 (N_2038,N_1505,N_1583);
xor U2039 (N_2039,N_1438,N_1235);
nor U2040 (N_2040,N_1426,N_976);
nor U2041 (N_2041,N_874,N_1063);
and U2042 (N_2042,N_1559,N_1494);
nor U2043 (N_2043,N_1390,N_1343);
xnor U2044 (N_2044,N_1023,N_818);
or U2045 (N_2045,N_1010,N_904);
xor U2046 (N_2046,N_993,N_1507);
or U2047 (N_2047,N_1469,N_1375);
or U2048 (N_2048,N_1143,N_1384);
and U2049 (N_2049,N_1443,N_1200);
nand U2050 (N_2050,N_1292,N_1453);
nor U2051 (N_2051,N_1275,N_1355);
nor U2052 (N_2052,N_1265,N_992);
xnor U2053 (N_2053,N_1314,N_1003);
and U2054 (N_2054,N_927,N_1328);
nand U2055 (N_2055,N_1232,N_1010);
xnor U2056 (N_2056,N_1531,N_1326);
xor U2057 (N_2057,N_1224,N_1197);
and U2058 (N_2058,N_1059,N_1080);
nand U2059 (N_2059,N_1047,N_917);
nor U2060 (N_2060,N_1173,N_1240);
and U2061 (N_2061,N_1457,N_1217);
nor U2062 (N_2062,N_911,N_1228);
nor U2063 (N_2063,N_1169,N_1589);
xnor U2064 (N_2064,N_831,N_1150);
or U2065 (N_2065,N_1198,N_1126);
xnor U2066 (N_2066,N_1103,N_888);
xnor U2067 (N_2067,N_975,N_1200);
and U2068 (N_2068,N_1004,N_1214);
or U2069 (N_2069,N_1599,N_1312);
nor U2070 (N_2070,N_1536,N_985);
and U2071 (N_2071,N_1069,N_1225);
or U2072 (N_2072,N_1552,N_1227);
and U2073 (N_2073,N_1341,N_1190);
or U2074 (N_2074,N_1592,N_1034);
nand U2075 (N_2075,N_1008,N_1294);
or U2076 (N_2076,N_1554,N_1178);
nand U2077 (N_2077,N_966,N_1575);
and U2078 (N_2078,N_1401,N_1475);
nor U2079 (N_2079,N_808,N_1585);
and U2080 (N_2080,N_1055,N_1039);
nor U2081 (N_2081,N_1164,N_835);
and U2082 (N_2082,N_1312,N_1053);
nor U2083 (N_2083,N_1176,N_843);
nor U2084 (N_2084,N_1253,N_1156);
and U2085 (N_2085,N_1044,N_1163);
xnor U2086 (N_2086,N_1315,N_1573);
and U2087 (N_2087,N_1270,N_1307);
xor U2088 (N_2088,N_1440,N_1133);
nor U2089 (N_2089,N_895,N_1353);
nor U2090 (N_2090,N_1167,N_891);
or U2091 (N_2091,N_1588,N_946);
or U2092 (N_2092,N_1022,N_907);
and U2093 (N_2093,N_1134,N_1147);
nor U2094 (N_2094,N_912,N_1174);
nand U2095 (N_2095,N_1228,N_1160);
nor U2096 (N_2096,N_853,N_804);
or U2097 (N_2097,N_973,N_1212);
or U2098 (N_2098,N_949,N_1280);
xor U2099 (N_2099,N_1152,N_961);
and U2100 (N_2100,N_1535,N_1309);
xor U2101 (N_2101,N_1474,N_1188);
nand U2102 (N_2102,N_1317,N_867);
nand U2103 (N_2103,N_1227,N_1107);
or U2104 (N_2104,N_1227,N_1443);
nor U2105 (N_2105,N_1098,N_866);
or U2106 (N_2106,N_1517,N_1390);
xor U2107 (N_2107,N_1185,N_1444);
nand U2108 (N_2108,N_1044,N_963);
and U2109 (N_2109,N_1323,N_1410);
and U2110 (N_2110,N_1581,N_1387);
xor U2111 (N_2111,N_1200,N_1145);
xnor U2112 (N_2112,N_1321,N_1228);
nand U2113 (N_2113,N_1182,N_1009);
nand U2114 (N_2114,N_1366,N_853);
nand U2115 (N_2115,N_1399,N_1555);
nor U2116 (N_2116,N_1192,N_1539);
nand U2117 (N_2117,N_1357,N_1462);
nor U2118 (N_2118,N_1365,N_851);
or U2119 (N_2119,N_1545,N_1252);
nand U2120 (N_2120,N_1153,N_1305);
nor U2121 (N_2121,N_1243,N_933);
and U2122 (N_2122,N_955,N_934);
nand U2123 (N_2123,N_1275,N_910);
or U2124 (N_2124,N_1338,N_997);
and U2125 (N_2125,N_1424,N_801);
and U2126 (N_2126,N_877,N_1145);
nor U2127 (N_2127,N_1363,N_1127);
or U2128 (N_2128,N_961,N_1440);
xnor U2129 (N_2129,N_830,N_1193);
xor U2130 (N_2130,N_1170,N_1253);
nand U2131 (N_2131,N_849,N_1504);
nor U2132 (N_2132,N_1470,N_1269);
and U2133 (N_2133,N_1526,N_1231);
or U2134 (N_2134,N_1422,N_851);
and U2135 (N_2135,N_1587,N_1351);
xnor U2136 (N_2136,N_1026,N_1279);
nand U2137 (N_2137,N_1436,N_1221);
nand U2138 (N_2138,N_1058,N_1302);
xnor U2139 (N_2139,N_970,N_1555);
xor U2140 (N_2140,N_878,N_1097);
and U2141 (N_2141,N_1233,N_1489);
nand U2142 (N_2142,N_1189,N_1454);
and U2143 (N_2143,N_1282,N_1384);
nor U2144 (N_2144,N_1269,N_1007);
xnor U2145 (N_2145,N_812,N_1329);
nor U2146 (N_2146,N_1136,N_1356);
or U2147 (N_2147,N_1111,N_1541);
xnor U2148 (N_2148,N_832,N_1367);
nor U2149 (N_2149,N_1564,N_1186);
xor U2150 (N_2150,N_970,N_1105);
nand U2151 (N_2151,N_1063,N_1196);
or U2152 (N_2152,N_1421,N_1331);
xor U2153 (N_2153,N_1472,N_1175);
and U2154 (N_2154,N_1398,N_1157);
or U2155 (N_2155,N_1033,N_1086);
or U2156 (N_2156,N_903,N_1102);
and U2157 (N_2157,N_1066,N_897);
nor U2158 (N_2158,N_1455,N_1416);
xnor U2159 (N_2159,N_891,N_1473);
nand U2160 (N_2160,N_817,N_1373);
xnor U2161 (N_2161,N_1558,N_1375);
and U2162 (N_2162,N_1541,N_1559);
xnor U2163 (N_2163,N_1472,N_961);
or U2164 (N_2164,N_1400,N_1448);
or U2165 (N_2165,N_979,N_1097);
or U2166 (N_2166,N_1288,N_818);
nand U2167 (N_2167,N_1574,N_1256);
nor U2168 (N_2168,N_1502,N_1450);
or U2169 (N_2169,N_906,N_1314);
and U2170 (N_2170,N_1190,N_885);
nor U2171 (N_2171,N_806,N_1519);
and U2172 (N_2172,N_1157,N_837);
and U2173 (N_2173,N_1590,N_1412);
xnor U2174 (N_2174,N_922,N_1283);
nor U2175 (N_2175,N_1160,N_865);
and U2176 (N_2176,N_1117,N_1110);
nand U2177 (N_2177,N_1181,N_1460);
or U2178 (N_2178,N_1137,N_1576);
nand U2179 (N_2179,N_879,N_974);
xnor U2180 (N_2180,N_1228,N_1177);
nor U2181 (N_2181,N_1374,N_1035);
nor U2182 (N_2182,N_1354,N_892);
and U2183 (N_2183,N_1051,N_1080);
or U2184 (N_2184,N_1372,N_849);
nand U2185 (N_2185,N_904,N_1430);
xor U2186 (N_2186,N_1305,N_1286);
or U2187 (N_2187,N_1556,N_1290);
nand U2188 (N_2188,N_1397,N_998);
or U2189 (N_2189,N_1051,N_904);
and U2190 (N_2190,N_1408,N_1125);
or U2191 (N_2191,N_1100,N_980);
xnor U2192 (N_2192,N_1290,N_1362);
nor U2193 (N_2193,N_1542,N_1088);
and U2194 (N_2194,N_868,N_824);
nor U2195 (N_2195,N_939,N_843);
nand U2196 (N_2196,N_809,N_1413);
nor U2197 (N_2197,N_1306,N_1384);
nand U2198 (N_2198,N_902,N_802);
nor U2199 (N_2199,N_957,N_1476);
xnor U2200 (N_2200,N_1527,N_1344);
or U2201 (N_2201,N_878,N_1329);
nand U2202 (N_2202,N_1135,N_1514);
nand U2203 (N_2203,N_1146,N_1018);
xor U2204 (N_2204,N_926,N_1560);
and U2205 (N_2205,N_1438,N_1559);
xor U2206 (N_2206,N_1547,N_1513);
nor U2207 (N_2207,N_911,N_1588);
nor U2208 (N_2208,N_843,N_1086);
and U2209 (N_2209,N_1112,N_1224);
nor U2210 (N_2210,N_1315,N_1003);
nor U2211 (N_2211,N_1421,N_1136);
and U2212 (N_2212,N_1204,N_1348);
nor U2213 (N_2213,N_833,N_1018);
nor U2214 (N_2214,N_1056,N_1296);
nand U2215 (N_2215,N_1481,N_1455);
or U2216 (N_2216,N_1559,N_1319);
xor U2217 (N_2217,N_1474,N_1334);
and U2218 (N_2218,N_1460,N_1146);
nor U2219 (N_2219,N_1161,N_1320);
nand U2220 (N_2220,N_977,N_1125);
or U2221 (N_2221,N_1220,N_1495);
xor U2222 (N_2222,N_1225,N_1457);
nand U2223 (N_2223,N_1259,N_1144);
or U2224 (N_2224,N_1349,N_1157);
nor U2225 (N_2225,N_1338,N_1354);
nor U2226 (N_2226,N_1222,N_1339);
and U2227 (N_2227,N_932,N_1320);
nand U2228 (N_2228,N_1491,N_1001);
or U2229 (N_2229,N_1183,N_1428);
nor U2230 (N_2230,N_1408,N_828);
or U2231 (N_2231,N_1303,N_983);
nand U2232 (N_2232,N_1094,N_1317);
nand U2233 (N_2233,N_1514,N_1346);
nor U2234 (N_2234,N_1093,N_1329);
nor U2235 (N_2235,N_882,N_1218);
or U2236 (N_2236,N_914,N_1186);
and U2237 (N_2237,N_1274,N_1513);
nor U2238 (N_2238,N_1131,N_831);
nor U2239 (N_2239,N_1563,N_1150);
and U2240 (N_2240,N_1328,N_946);
or U2241 (N_2241,N_964,N_1479);
or U2242 (N_2242,N_1106,N_854);
xnor U2243 (N_2243,N_1279,N_860);
or U2244 (N_2244,N_905,N_1308);
or U2245 (N_2245,N_1516,N_1594);
or U2246 (N_2246,N_1388,N_1103);
xnor U2247 (N_2247,N_1493,N_1074);
nand U2248 (N_2248,N_1090,N_1330);
or U2249 (N_2249,N_1353,N_1418);
nor U2250 (N_2250,N_912,N_1309);
nor U2251 (N_2251,N_973,N_1335);
xor U2252 (N_2252,N_1552,N_1282);
or U2253 (N_2253,N_1107,N_994);
or U2254 (N_2254,N_1067,N_848);
or U2255 (N_2255,N_1049,N_852);
nor U2256 (N_2256,N_948,N_1194);
nand U2257 (N_2257,N_825,N_1520);
xnor U2258 (N_2258,N_883,N_1511);
or U2259 (N_2259,N_1334,N_1507);
or U2260 (N_2260,N_1472,N_932);
and U2261 (N_2261,N_1286,N_1147);
and U2262 (N_2262,N_1308,N_1293);
or U2263 (N_2263,N_1437,N_1432);
nor U2264 (N_2264,N_1100,N_898);
xnor U2265 (N_2265,N_1360,N_1218);
xor U2266 (N_2266,N_1157,N_1590);
or U2267 (N_2267,N_1542,N_1439);
and U2268 (N_2268,N_1252,N_1188);
nand U2269 (N_2269,N_1173,N_1180);
xnor U2270 (N_2270,N_1037,N_807);
and U2271 (N_2271,N_1174,N_1307);
nor U2272 (N_2272,N_1297,N_1275);
xor U2273 (N_2273,N_1391,N_1180);
or U2274 (N_2274,N_1156,N_834);
and U2275 (N_2275,N_1059,N_1356);
nand U2276 (N_2276,N_1533,N_1312);
or U2277 (N_2277,N_1593,N_1079);
xnor U2278 (N_2278,N_1124,N_1582);
nor U2279 (N_2279,N_977,N_881);
or U2280 (N_2280,N_1007,N_1487);
nor U2281 (N_2281,N_1086,N_1040);
nor U2282 (N_2282,N_1492,N_1076);
or U2283 (N_2283,N_1432,N_1384);
nand U2284 (N_2284,N_1472,N_944);
nor U2285 (N_2285,N_1561,N_1066);
or U2286 (N_2286,N_1298,N_1296);
nand U2287 (N_2287,N_825,N_1123);
nand U2288 (N_2288,N_1136,N_1002);
and U2289 (N_2289,N_1384,N_837);
nand U2290 (N_2290,N_839,N_970);
nor U2291 (N_2291,N_1240,N_1256);
and U2292 (N_2292,N_1261,N_1341);
nor U2293 (N_2293,N_1088,N_1293);
and U2294 (N_2294,N_1280,N_865);
or U2295 (N_2295,N_1002,N_1076);
nor U2296 (N_2296,N_839,N_1243);
and U2297 (N_2297,N_1580,N_949);
nor U2298 (N_2298,N_892,N_957);
or U2299 (N_2299,N_1377,N_1284);
nor U2300 (N_2300,N_996,N_1261);
nor U2301 (N_2301,N_1168,N_1263);
xnor U2302 (N_2302,N_1540,N_1328);
nand U2303 (N_2303,N_1227,N_1043);
nor U2304 (N_2304,N_947,N_1496);
xnor U2305 (N_2305,N_1128,N_1163);
xnor U2306 (N_2306,N_914,N_892);
or U2307 (N_2307,N_861,N_1023);
or U2308 (N_2308,N_1154,N_1313);
nor U2309 (N_2309,N_940,N_1452);
and U2310 (N_2310,N_1537,N_852);
nor U2311 (N_2311,N_1006,N_1401);
nand U2312 (N_2312,N_1526,N_1585);
xnor U2313 (N_2313,N_1036,N_834);
nor U2314 (N_2314,N_1193,N_1429);
nand U2315 (N_2315,N_1150,N_1200);
and U2316 (N_2316,N_1025,N_1007);
nor U2317 (N_2317,N_1443,N_1267);
and U2318 (N_2318,N_814,N_1525);
nand U2319 (N_2319,N_923,N_1419);
nor U2320 (N_2320,N_1302,N_1236);
nand U2321 (N_2321,N_912,N_1015);
and U2322 (N_2322,N_1489,N_1586);
nor U2323 (N_2323,N_1572,N_1105);
and U2324 (N_2324,N_1053,N_846);
nand U2325 (N_2325,N_1059,N_1368);
xor U2326 (N_2326,N_1287,N_896);
xnor U2327 (N_2327,N_1352,N_827);
nand U2328 (N_2328,N_1293,N_832);
xnor U2329 (N_2329,N_1556,N_1596);
nor U2330 (N_2330,N_1090,N_858);
nand U2331 (N_2331,N_1080,N_1533);
nand U2332 (N_2332,N_1135,N_1143);
xor U2333 (N_2333,N_1402,N_1444);
nand U2334 (N_2334,N_1146,N_1017);
and U2335 (N_2335,N_1354,N_1306);
xnor U2336 (N_2336,N_1282,N_1292);
nand U2337 (N_2337,N_1137,N_1205);
or U2338 (N_2338,N_1083,N_929);
and U2339 (N_2339,N_1063,N_1326);
and U2340 (N_2340,N_1279,N_1042);
nand U2341 (N_2341,N_994,N_840);
xnor U2342 (N_2342,N_1285,N_818);
and U2343 (N_2343,N_1433,N_1368);
and U2344 (N_2344,N_905,N_1128);
nand U2345 (N_2345,N_1549,N_1160);
nand U2346 (N_2346,N_1361,N_1446);
and U2347 (N_2347,N_1495,N_865);
or U2348 (N_2348,N_1476,N_1215);
nand U2349 (N_2349,N_995,N_1091);
xnor U2350 (N_2350,N_924,N_912);
and U2351 (N_2351,N_911,N_846);
xor U2352 (N_2352,N_1577,N_1346);
nor U2353 (N_2353,N_1282,N_1373);
or U2354 (N_2354,N_1201,N_958);
nand U2355 (N_2355,N_1064,N_1059);
and U2356 (N_2356,N_1073,N_972);
nand U2357 (N_2357,N_928,N_819);
nor U2358 (N_2358,N_1189,N_1164);
nor U2359 (N_2359,N_1523,N_818);
nor U2360 (N_2360,N_1393,N_1017);
nor U2361 (N_2361,N_917,N_1223);
xnor U2362 (N_2362,N_1517,N_1444);
nor U2363 (N_2363,N_872,N_1409);
nand U2364 (N_2364,N_1144,N_1111);
nor U2365 (N_2365,N_860,N_1139);
or U2366 (N_2366,N_1403,N_1346);
nor U2367 (N_2367,N_1322,N_1187);
xnor U2368 (N_2368,N_880,N_853);
and U2369 (N_2369,N_1018,N_1507);
or U2370 (N_2370,N_1242,N_1129);
nor U2371 (N_2371,N_812,N_1188);
or U2372 (N_2372,N_1392,N_1246);
and U2373 (N_2373,N_905,N_1278);
xor U2374 (N_2374,N_1295,N_1153);
xnor U2375 (N_2375,N_1414,N_1015);
nor U2376 (N_2376,N_1298,N_1479);
xor U2377 (N_2377,N_1565,N_959);
and U2378 (N_2378,N_878,N_845);
and U2379 (N_2379,N_1124,N_1205);
and U2380 (N_2380,N_1207,N_1040);
xor U2381 (N_2381,N_845,N_1019);
and U2382 (N_2382,N_1089,N_900);
xnor U2383 (N_2383,N_1394,N_913);
xnor U2384 (N_2384,N_1584,N_1445);
xor U2385 (N_2385,N_1042,N_1470);
xnor U2386 (N_2386,N_1414,N_1428);
or U2387 (N_2387,N_1202,N_956);
nor U2388 (N_2388,N_1124,N_834);
and U2389 (N_2389,N_1579,N_1110);
nand U2390 (N_2390,N_992,N_1569);
and U2391 (N_2391,N_1386,N_941);
and U2392 (N_2392,N_946,N_905);
nand U2393 (N_2393,N_828,N_1267);
nand U2394 (N_2394,N_966,N_1543);
nor U2395 (N_2395,N_900,N_1084);
and U2396 (N_2396,N_1341,N_1138);
or U2397 (N_2397,N_1412,N_1522);
and U2398 (N_2398,N_1073,N_1589);
or U2399 (N_2399,N_918,N_1590);
nor U2400 (N_2400,N_2054,N_2329);
and U2401 (N_2401,N_2361,N_2064);
or U2402 (N_2402,N_2227,N_2123);
nand U2403 (N_2403,N_1900,N_1622);
and U2404 (N_2404,N_2339,N_2039);
or U2405 (N_2405,N_2033,N_2210);
or U2406 (N_2406,N_2344,N_2258);
or U2407 (N_2407,N_2201,N_1672);
xnor U2408 (N_2408,N_1769,N_1984);
xnor U2409 (N_2409,N_1709,N_2379);
or U2410 (N_2410,N_2251,N_1616);
nand U2411 (N_2411,N_1704,N_2074);
or U2412 (N_2412,N_1848,N_1806);
xor U2413 (N_2413,N_2300,N_1665);
and U2414 (N_2414,N_1954,N_1803);
and U2415 (N_2415,N_2101,N_2085);
xnor U2416 (N_2416,N_1706,N_1661);
or U2417 (N_2417,N_2208,N_1750);
nor U2418 (N_2418,N_1705,N_1938);
nand U2419 (N_2419,N_2096,N_2268);
and U2420 (N_2420,N_1965,N_2030);
or U2421 (N_2421,N_1896,N_1825);
or U2422 (N_2422,N_2021,N_1720);
nand U2423 (N_2423,N_2367,N_2051);
and U2424 (N_2424,N_2116,N_2248);
or U2425 (N_2425,N_2285,N_2071);
and U2426 (N_2426,N_2386,N_1810);
or U2427 (N_2427,N_1689,N_1939);
and U2428 (N_2428,N_2372,N_1666);
nand U2429 (N_2429,N_1785,N_2387);
nand U2430 (N_2430,N_1717,N_2115);
nor U2431 (N_2431,N_2345,N_2356);
xnor U2432 (N_2432,N_1787,N_2390);
nor U2433 (N_2433,N_2183,N_1950);
or U2434 (N_2434,N_2257,N_2266);
and U2435 (N_2435,N_2079,N_2126);
nand U2436 (N_2436,N_2037,N_1885);
xnor U2437 (N_2437,N_1962,N_1707);
xor U2438 (N_2438,N_1636,N_1923);
or U2439 (N_2439,N_1768,N_2172);
or U2440 (N_2440,N_1654,N_1735);
or U2441 (N_2441,N_1739,N_1851);
and U2442 (N_2442,N_2306,N_1731);
and U2443 (N_2443,N_1692,N_1872);
nand U2444 (N_2444,N_1862,N_1745);
nand U2445 (N_2445,N_2003,N_1747);
xnor U2446 (N_2446,N_2331,N_1817);
xor U2447 (N_2447,N_1897,N_1725);
xor U2448 (N_2448,N_1643,N_1601);
nand U2449 (N_2449,N_2236,N_1829);
xor U2450 (N_2450,N_1813,N_2063);
xnor U2451 (N_2451,N_1767,N_1873);
and U2452 (N_2452,N_2217,N_2380);
xor U2453 (N_2453,N_2006,N_1920);
nand U2454 (N_2454,N_2381,N_2125);
nor U2455 (N_2455,N_2360,N_1975);
nand U2456 (N_2456,N_2001,N_1853);
nor U2457 (N_2457,N_2168,N_1884);
nand U2458 (N_2458,N_2137,N_1635);
and U2459 (N_2459,N_1909,N_1964);
nor U2460 (N_2460,N_2288,N_1657);
nor U2461 (N_2461,N_1949,N_1934);
nand U2462 (N_2462,N_1634,N_1763);
nor U2463 (N_2463,N_1760,N_1606);
or U2464 (N_2464,N_2365,N_1611);
nor U2465 (N_2465,N_2272,N_2199);
or U2466 (N_2466,N_2271,N_2034);
xnor U2467 (N_2467,N_2351,N_2298);
xor U2468 (N_2468,N_2154,N_2082);
or U2469 (N_2469,N_2309,N_2289);
xor U2470 (N_2470,N_2225,N_2165);
xnor U2471 (N_2471,N_2273,N_1935);
nand U2472 (N_2472,N_1960,N_2252);
xnor U2473 (N_2473,N_2099,N_2226);
nor U2474 (N_2474,N_1815,N_2015);
or U2475 (N_2475,N_1662,N_1898);
or U2476 (N_2476,N_1926,N_1904);
nand U2477 (N_2477,N_2335,N_2221);
nor U2478 (N_2478,N_2169,N_1757);
xnor U2479 (N_2479,N_2263,N_1660);
xor U2480 (N_2480,N_2004,N_2173);
nand U2481 (N_2481,N_1795,N_2355);
and U2482 (N_2482,N_2105,N_2358);
xnor U2483 (N_2483,N_2328,N_1983);
xnor U2484 (N_2484,N_1740,N_1959);
and U2485 (N_2485,N_1880,N_1866);
or U2486 (N_2486,N_2188,N_2133);
nor U2487 (N_2487,N_2167,N_2277);
nand U2488 (N_2488,N_1834,N_1821);
nor U2489 (N_2489,N_1697,N_2012);
nand U2490 (N_2490,N_1742,N_2291);
or U2491 (N_2491,N_2028,N_2233);
nor U2492 (N_2492,N_1857,N_1933);
or U2493 (N_2493,N_2066,N_2073);
nand U2494 (N_2494,N_2293,N_1868);
or U2495 (N_2495,N_1694,N_2060);
or U2496 (N_2496,N_2260,N_1708);
nand U2497 (N_2497,N_2363,N_1685);
and U2498 (N_2498,N_1711,N_1681);
nor U2499 (N_2499,N_2136,N_2232);
nor U2500 (N_2500,N_2052,N_1889);
and U2501 (N_2501,N_2196,N_2254);
or U2502 (N_2502,N_2162,N_1713);
nor U2503 (N_2503,N_2193,N_2156);
nand U2504 (N_2504,N_2385,N_2398);
xnor U2505 (N_2505,N_2202,N_2212);
or U2506 (N_2506,N_2124,N_2264);
xor U2507 (N_2507,N_2005,N_2297);
nor U2508 (N_2508,N_1921,N_2131);
nand U2509 (N_2509,N_1625,N_1819);
nor U2510 (N_2510,N_1756,N_1780);
and U2511 (N_2511,N_1907,N_2171);
or U2512 (N_2512,N_2159,N_1727);
nand U2513 (N_2513,N_2336,N_2370);
xor U2514 (N_2514,N_1976,N_2278);
or U2515 (N_2515,N_2206,N_1618);
nand U2516 (N_2516,N_1746,N_2035);
nand U2517 (N_2517,N_2118,N_1721);
and U2518 (N_2518,N_2397,N_2055);
and U2519 (N_2519,N_1928,N_2102);
or U2520 (N_2520,N_2150,N_2223);
nor U2521 (N_2521,N_1628,N_1836);
and U2522 (N_2522,N_1640,N_1605);
or U2523 (N_2523,N_2230,N_2182);
xnor U2524 (N_2524,N_1980,N_2100);
and U2525 (N_2525,N_2145,N_1734);
or U2526 (N_2526,N_2368,N_2235);
xnor U2527 (N_2527,N_1793,N_1609);
nor U2528 (N_2528,N_2093,N_1841);
and U2529 (N_2529,N_1905,N_1649);
xor U2530 (N_2530,N_1641,N_1676);
nand U2531 (N_2531,N_2058,N_1936);
nor U2532 (N_2532,N_2138,N_1675);
and U2533 (N_2533,N_2312,N_1632);
nor U2534 (N_2534,N_2245,N_1818);
xor U2535 (N_2535,N_1869,N_2249);
xor U2536 (N_2536,N_2255,N_2200);
nor U2537 (N_2537,N_1948,N_1807);
and U2538 (N_2538,N_2092,N_1703);
nor U2539 (N_2539,N_1722,N_2149);
nand U2540 (N_2540,N_2106,N_1630);
and U2541 (N_2541,N_1922,N_1974);
nand U2542 (N_2542,N_1881,N_2184);
and U2543 (N_2543,N_1982,N_1970);
xor U2544 (N_2544,N_1919,N_1981);
and U2545 (N_2545,N_2177,N_2211);
nand U2546 (N_2546,N_2049,N_1973);
nor U2547 (N_2547,N_1623,N_2274);
and U2548 (N_2548,N_2152,N_1751);
nand U2549 (N_2549,N_2238,N_1668);
and U2550 (N_2550,N_2341,N_1781);
or U2551 (N_2551,N_2376,N_2394);
nor U2552 (N_2552,N_2319,N_1762);
nand U2553 (N_2553,N_1682,N_2283);
nor U2554 (N_2554,N_2280,N_2275);
xnor U2555 (N_2555,N_1842,N_1990);
xor U2556 (N_2556,N_2347,N_1658);
and U2557 (N_2557,N_1797,N_2259);
and U2558 (N_2558,N_1669,N_2242);
nor U2559 (N_2559,N_2010,N_2359);
nand U2560 (N_2560,N_2067,N_1858);
xnor U2561 (N_2561,N_1995,N_1788);
or U2562 (N_2562,N_2192,N_1929);
nand U2563 (N_2563,N_1695,N_2190);
or U2564 (N_2564,N_2218,N_2186);
nand U2565 (N_2565,N_2295,N_1651);
nor U2566 (N_2566,N_2086,N_1833);
xor U2567 (N_2567,N_1883,N_2127);
and U2568 (N_2568,N_1794,N_1892);
nor U2569 (N_2569,N_2326,N_1847);
or U2570 (N_2570,N_2237,N_2229);
or U2571 (N_2571,N_1816,N_1996);
or U2572 (N_2572,N_2377,N_2378);
or U2573 (N_2573,N_1613,N_2155);
and U2574 (N_2574,N_2296,N_1765);
nand U2575 (N_2575,N_1968,N_1719);
nand U2576 (N_2576,N_1792,N_1871);
xor U2577 (N_2577,N_1927,N_1716);
or U2578 (N_2578,N_1867,N_1958);
or U2579 (N_2579,N_1683,N_1997);
xor U2580 (N_2580,N_1728,N_2097);
or U2581 (N_2581,N_1966,N_2213);
xor U2582 (N_2582,N_2017,N_2044);
xnor U2583 (N_2583,N_1701,N_1778);
xor U2584 (N_2584,N_2181,N_1998);
nand U2585 (N_2585,N_1930,N_2318);
nor U2586 (N_2586,N_2382,N_1838);
or U2587 (N_2587,N_1631,N_1808);
and U2588 (N_2588,N_2014,N_2391);
or U2589 (N_2589,N_2323,N_2352);
and U2590 (N_2590,N_2038,N_1863);
or U2591 (N_2591,N_1820,N_2354);
and U2592 (N_2592,N_1771,N_2027);
nand U2593 (N_2593,N_2143,N_1911);
xor U2594 (N_2594,N_1673,N_1835);
xnor U2595 (N_2595,N_2164,N_2239);
nor U2596 (N_2596,N_1865,N_1830);
xnor U2597 (N_2597,N_2147,N_1678);
nand U2598 (N_2598,N_2139,N_1967);
nor U2599 (N_2599,N_1754,N_1809);
and U2600 (N_2600,N_1844,N_1684);
nor U2601 (N_2601,N_2179,N_1796);
and U2602 (N_2602,N_1969,N_2163);
nand U2603 (N_2603,N_2000,N_2151);
xnor U2604 (N_2604,N_2216,N_1633);
xnor U2605 (N_2605,N_1743,N_2089);
xnor U2606 (N_2606,N_2045,N_2234);
nand U2607 (N_2607,N_1648,N_2393);
or U2608 (N_2608,N_2310,N_1859);
xor U2609 (N_2609,N_1688,N_2317);
xnor U2610 (N_2610,N_2036,N_2069);
or U2611 (N_2611,N_2357,N_1991);
nor U2612 (N_2612,N_2141,N_2088);
nand U2613 (N_2613,N_1843,N_1952);
and U2614 (N_2614,N_2203,N_1639);
nor U2615 (N_2615,N_2029,N_1822);
or U2616 (N_2616,N_1789,N_2120);
and U2617 (N_2617,N_1947,N_1617);
or U2618 (N_2618,N_1744,N_2343);
or U2619 (N_2619,N_1702,N_2094);
xnor U2620 (N_2620,N_1963,N_2135);
xnor U2621 (N_2621,N_1840,N_1615);
nand U2622 (N_2622,N_1993,N_1864);
nor U2623 (N_2623,N_2128,N_1908);
nor U2624 (N_2624,N_2311,N_2170);
nor U2625 (N_2625,N_1612,N_1645);
nand U2626 (N_2626,N_1946,N_1753);
nand U2627 (N_2627,N_1729,N_2122);
nor U2628 (N_2628,N_1999,N_2353);
and U2629 (N_2629,N_1801,N_1893);
and U2630 (N_2630,N_1749,N_1989);
or U2631 (N_2631,N_2068,N_2207);
or U2632 (N_2632,N_1839,N_1931);
nor U2633 (N_2633,N_1887,N_2107);
xor U2634 (N_2634,N_2046,N_1957);
or U2635 (N_2635,N_1626,N_2025);
nand U2636 (N_2636,N_2132,N_1755);
or U2637 (N_2637,N_1903,N_1775);
nand U2638 (N_2638,N_2020,N_1770);
or U2639 (N_2639,N_2090,N_2292);
nor U2640 (N_2640,N_1691,N_2140);
xnor U2641 (N_2641,N_1764,N_2321);
nor U2642 (N_2642,N_1942,N_2198);
xor U2643 (N_2643,N_2110,N_2290);
xnor U2644 (N_2644,N_1953,N_2187);
nor U2645 (N_2645,N_1619,N_2314);
nand U2646 (N_2646,N_1971,N_1659);
or U2647 (N_2647,N_2080,N_1901);
and U2648 (N_2648,N_2346,N_2322);
xor U2649 (N_2649,N_2325,N_2384);
and U2650 (N_2650,N_2270,N_1629);
or U2651 (N_2651,N_1894,N_2399);
nor U2652 (N_2652,N_1891,N_1978);
and U2653 (N_2653,N_1696,N_1824);
nor U2654 (N_2654,N_2303,N_2224);
nor U2655 (N_2655,N_2267,N_2209);
or U2656 (N_2656,N_2134,N_2304);
and U2657 (N_2657,N_1642,N_1943);
xnor U2658 (N_2658,N_1724,N_1610);
nand U2659 (N_2659,N_1888,N_1917);
nand U2660 (N_2660,N_1644,N_2109);
xor U2661 (N_2661,N_1812,N_1603);
or U2662 (N_2662,N_1786,N_2011);
or U2663 (N_2663,N_1832,N_2175);
nand U2664 (N_2664,N_1876,N_1798);
xor U2665 (N_2665,N_2059,N_2294);
xor U2666 (N_2666,N_1621,N_1600);
nor U2667 (N_2667,N_2219,N_1604);
or U2668 (N_2668,N_2305,N_1860);
or U2669 (N_2669,N_1992,N_2327);
or U2670 (N_2670,N_2215,N_2315);
nor U2671 (N_2671,N_2158,N_1680);
and U2672 (N_2672,N_2042,N_1723);
nand U2673 (N_2673,N_1945,N_1886);
nor U2674 (N_2674,N_1916,N_2308);
nor U2675 (N_2675,N_1726,N_1693);
or U2676 (N_2676,N_1773,N_1977);
and U2677 (N_2677,N_1667,N_1653);
nand U2678 (N_2678,N_2176,N_1624);
nor U2679 (N_2679,N_1674,N_2180);
nor U2680 (N_2680,N_2253,N_2389);
and U2681 (N_2681,N_1782,N_1655);
and U2682 (N_2682,N_1986,N_1766);
and U2683 (N_2683,N_1846,N_1955);
nor U2684 (N_2684,N_1870,N_2032);
nor U2685 (N_2685,N_1761,N_1718);
nor U2686 (N_2686,N_2338,N_2084);
nor U2687 (N_2687,N_2195,N_2392);
or U2688 (N_2688,N_1855,N_1712);
nand U2689 (N_2689,N_1698,N_1687);
or U2690 (N_2690,N_2286,N_2349);
nand U2691 (N_2691,N_1814,N_2129);
nand U2692 (N_2692,N_2364,N_2061);
nand U2693 (N_2693,N_1679,N_1856);
and U2694 (N_2694,N_1805,N_2075);
and U2695 (N_2695,N_2383,N_1906);
xnor U2696 (N_2696,N_2050,N_1602);
nand U2697 (N_2697,N_2031,N_2191);
nand U2698 (N_2698,N_2009,N_1831);
and U2699 (N_2699,N_2161,N_1845);
and U2700 (N_2700,N_2316,N_2048);
nor U2701 (N_2701,N_1972,N_1944);
and U2702 (N_2702,N_1710,N_2016);
nor U2703 (N_2703,N_2396,N_1987);
or U2704 (N_2704,N_2369,N_1850);
or U2705 (N_2705,N_1647,N_2284);
xnor U2706 (N_2706,N_2250,N_1837);
and U2707 (N_2707,N_2007,N_1784);
nor U2708 (N_2708,N_2374,N_1854);
nand U2709 (N_2709,N_2301,N_2204);
nand U2710 (N_2710,N_1925,N_1924);
nor U2711 (N_2711,N_1902,N_1890);
nor U2712 (N_2712,N_2130,N_1776);
nor U2713 (N_2713,N_1811,N_2078);
nand U2714 (N_2714,N_2340,N_2040);
nand U2715 (N_2715,N_2324,N_2062);
or U2716 (N_2716,N_2395,N_1759);
xor U2717 (N_2717,N_2222,N_2178);
and U2718 (N_2718,N_1912,N_1874);
or U2719 (N_2719,N_2166,N_1656);
nand U2720 (N_2720,N_2189,N_2026);
xor U2721 (N_2721,N_2350,N_1878);
xnor U2722 (N_2722,N_2065,N_1700);
or U2723 (N_2723,N_2111,N_2330);
or U2724 (N_2724,N_2081,N_2146);
xnor U2725 (N_2725,N_2153,N_1741);
or U2726 (N_2726,N_2269,N_2279);
nand U2727 (N_2727,N_2243,N_1879);
nand U2728 (N_2728,N_1671,N_1979);
xnor U2729 (N_2729,N_2121,N_2282);
nand U2730 (N_2730,N_1882,N_2197);
nand U2731 (N_2731,N_2320,N_2261);
nand U2732 (N_2732,N_2119,N_2307);
nor U2733 (N_2733,N_1915,N_1748);
xor U2734 (N_2734,N_1774,N_2098);
nor U2735 (N_2735,N_1985,N_2041);
and U2736 (N_2736,N_1637,N_2246);
and U2737 (N_2737,N_1828,N_1646);
nand U2738 (N_2738,N_2302,N_2205);
and U2739 (N_2739,N_1714,N_2241);
or U2740 (N_2740,N_2070,N_2194);
nand U2741 (N_2741,N_1961,N_1910);
nand U2742 (N_2742,N_1690,N_2281);
or U2743 (N_2743,N_2371,N_2019);
nand U2744 (N_2744,N_1802,N_2112);
or U2745 (N_2745,N_1737,N_1790);
nor U2746 (N_2746,N_1686,N_2114);
or U2747 (N_2747,N_1826,N_2018);
xnor U2748 (N_2748,N_2256,N_2056);
nor U2749 (N_2749,N_1663,N_2342);
or U2750 (N_2750,N_2231,N_1918);
and U2751 (N_2751,N_2262,N_2095);
xor U2752 (N_2752,N_2087,N_1988);
nand U2753 (N_2753,N_1664,N_2333);
xnor U2754 (N_2754,N_1677,N_1804);
and U2755 (N_2755,N_2348,N_2091);
nand U2756 (N_2756,N_2117,N_2023);
and U2757 (N_2757,N_1732,N_1758);
and U2758 (N_2758,N_1932,N_1827);
or U2759 (N_2759,N_2337,N_1823);
nand U2760 (N_2760,N_2024,N_1733);
and U2761 (N_2761,N_2142,N_1799);
nor U2762 (N_2762,N_2057,N_1620);
xor U2763 (N_2763,N_2287,N_1627);
nor U2764 (N_2764,N_1895,N_2299);
xor U2765 (N_2765,N_1940,N_2072);
xnor U2766 (N_2766,N_2002,N_2148);
and U2767 (N_2767,N_2388,N_2008);
and U2768 (N_2768,N_2174,N_1899);
or U2769 (N_2769,N_1607,N_2375);
and U2770 (N_2770,N_1913,N_2334);
or U2771 (N_2771,N_2247,N_2077);
nand U2772 (N_2772,N_1670,N_2108);
xor U2773 (N_2773,N_1638,N_1779);
or U2774 (N_2774,N_2214,N_2362);
nand U2775 (N_2775,N_1914,N_1777);
and U2776 (N_2776,N_1861,N_1800);
nor U2777 (N_2777,N_2160,N_1994);
nor U2778 (N_2778,N_1608,N_1650);
nor U2779 (N_2779,N_2103,N_2083);
xnor U2780 (N_2780,N_1937,N_2228);
nor U2781 (N_2781,N_2244,N_1614);
and U2782 (N_2782,N_2185,N_1951);
nor U2783 (N_2783,N_2240,N_2373);
xor U2784 (N_2784,N_2013,N_2053);
nand U2785 (N_2785,N_2076,N_1652);
xor U2786 (N_2786,N_1877,N_1738);
or U2787 (N_2787,N_2113,N_2104);
nor U2788 (N_2788,N_2265,N_2047);
nand U2789 (N_2789,N_2313,N_1852);
or U2790 (N_2790,N_2220,N_2043);
or U2791 (N_2791,N_1699,N_2366);
xnor U2792 (N_2792,N_1783,N_2276);
and U2793 (N_2793,N_1791,N_2332);
nand U2794 (N_2794,N_2022,N_1715);
xor U2795 (N_2795,N_1956,N_1736);
xor U2796 (N_2796,N_1941,N_2144);
nor U2797 (N_2797,N_1730,N_1752);
or U2798 (N_2798,N_1772,N_2157);
and U2799 (N_2799,N_1849,N_1875);
or U2800 (N_2800,N_1812,N_1860);
and U2801 (N_2801,N_2190,N_1845);
and U2802 (N_2802,N_2117,N_2042);
xor U2803 (N_2803,N_2018,N_1614);
nand U2804 (N_2804,N_1647,N_1980);
and U2805 (N_2805,N_1612,N_2194);
xor U2806 (N_2806,N_2201,N_2177);
xnor U2807 (N_2807,N_1760,N_2305);
and U2808 (N_2808,N_2011,N_2236);
or U2809 (N_2809,N_2217,N_1753);
and U2810 (N_2810,N_2112,N_2329);
nor U2811 (N_2811,N_2208,N_2332);
and U2812 (N_2812,N_2089,N_1779);
and U2813 (N_2813,N_2285,N_2230);
and U2814 (N_2814,N_1627,N_1906);
nand U2815 (N_2815,N_1665,N_1617);
nand U2816 (N_2816,N_1805,N_1825);
or U2817 (N_2817,N_1982,N_1896);
xnor U2818 (N_2818,N_1645,N_2058);
or U2819 (N_2819,N_2367,N_1923);
nand U2820 (N_2820,N_2297,N_2242);
and U2821 (N_2821,N_1720,N_1841);
and U2822 (N_2822,N_2137,N_2236);
xnor U2823 (N_2823,N_1843,N_1728);
nand U2824 (N_2824,N_1614,N_1850);
and U2825 (N_2825,N_2194,N_2167);
xor U2826 (N_2826,N_1678,N_1970);
and U2827 (N_2827,N_1940,N_1605);
nor U2828 (N_2828,N_2281,N_1743);
nand U2829 (N_2829,N_2334,N_2273);
nor U2830 (N_2830,N_2274,N_1695);
nand U2831 (N_2831,N_2351,N_1683);
or U2832 (N_2832,N_1738,N_2166);
xor U2833 (N_2833,N_2172,N_2376);
xnor U2834 (N_2834,N_1794,N_1623);
or U2835 (N_2835,N_2273,N_1852);
xor U2836 (N_2836,N_2291,N_2265);
nand U2837 (N_2837,N_1862,N_1661);
and U2838 (N_2838,N_1864,N_2351);
and U2839 (N_2839,N_2131,N_2223);
nand U2840 (N_2840,N_2375,N_2034);
xnor U2841 (N_2841,N_1877,N_2353);
xor U2842 (N_2842,N_2205,N_2165);
and U2843 (N_2843,N_2037,N_1774);
and U2844 (N_2844,N_1726,N_1790);
or U2845 (N_2845,N_2006,N_2352);
xor U2846 (N_2846,N_2292,N_2217);
nand U2847 (N_2847,N_1628,N_2304);
or U2848 (N_2848,N_2094,N_2119);
or U2849 (N_2849,N_1755,N_2115);
nor U2850 (N_2850,N_2199,N_1796);
nor U2851 (N_2851,N_1839,N_1801);
nand U2852 (N_2852,N_1688,N_2211);
xor U2853 (N_2853,N_1632,N_1980);
nand U2854 (N_2854,N_1774,N_1610);
or U2855 (N_2855,N_2286,N_1937);
and U2856 (N_2856,N_1774,N_1941);
or U2857 (N_2857,N_2025,N_1825);
or U2858 (N_2858,N_2127,N_1712);
xor U2859 (N_2859,N_1856,N_1717);
and U2860 (N_2860,N_2161,N_1999);
nand U2861 (N_2861,N_2378,N_2391);
xnor U2862 (N_2862,N_2074,N_2214);
or U2863 (N_2863,N_2326,N_1804);
nor U2864 (N_2864,N_2317,N_1667);
and U2865 (N_2865,N_2093,N_2071);
xor U2866 (N_2866,N_2360,N_2108);
nor U2867 (N_2867,N_2044,N_1622);
or U2868 (N_2868,N_2170,N_2101);
nand U2869 (N_2869,N_1634,N_2246);
nor U2870 (N_2870,N_1825,N_1935);
nand U2871 (N_2871,N_1615,N_2099);
xnor U2872 (N_2872,N_2005,N_1616);
and U2873 (N_2873,N_2321,N_2371);
nor U2874 (N_2874,N_1682,N_1827);
nor U2875 (N_2875,N_1609,N_1840);
xor U2876 (N_2876,N_2385,N_2248);
or U2877 (N_2877,N_2184,N_2110);
nor U2878 (N_2878,N_1639,N_1755);
nand U2879 (N_2879,N_2298,N_2130);
and U2880 (N_2880,N_1760,N_2040);
xor U2881 (N_2881,N_1666,N_2047);
nor U2882 (N_2882,N_1971,N_2311);
and U2883 (N_2883,N_1990,N_1797);
and U2884 (N_2884,N_2062,N_2020);
and U2885 (N_2885,N_1741,N_2279);
nor U2886 (N_2886,N_2299,N_1921);
nor U2887 (N_2887,N_2144,N_2327);
or U2888 (N_2888,N_1873,N_1848);
and U2889 (N_2889,N_2311,N_1743);
or U2890 (N_2890,N_1805,N_1879);
xor U2891 (N_2891,N_1953,N_1802);
nor U2892 (N_2892,N_1913,N_1737);
xor U2893 (N_2893,N_1758,N_2080);
xor U2894 (N_2894,N_1712,N_1985);
or U2895 (N_2895,N_2132,N_2306);
xnor U2896 (N_2896,N_1717,N_2085);
and U2897 (N_2897,N_2342,N_1650);
nor U2898 (N_2898,N_2361,N_1826);
nor U2899 (N_2899,N_1621,N_2205);
or U2900 (N_2900,N_2366,N_1963);
nor U2901 (N_2901,N_2354,N_1656);
nand U2902 (N_2902,N_1958,N_2208);
or U2903 (N_2903,N_2229,N_1949);
and U2904 (N_2904,N_2323,N_1900);
and U2905 (N_2905,N_1642,N_1605);
nand U2906 (N_2906,N_2031,N_2192);
nand U2907 (N_2907,N_2026,N_1718);
nor U2908 (N_2908,N_1987,N_1626);
or U2909 (N_2909,N_1844,N_2387);
and U2910 (N_2910,N_2293,N_1615);
xnor U2911 (N_2911,N_1981,N_2336);
nand U2912 (N_2912,N_1934,N_1804);
or U2913 (N_2913,N_1897,N_2338);
nand U2914 (N_2914,N_1765,N_1823);
xnor U2915 (N_2915,N_1979,N_1976);
or U2916 (N_2916,N_2129,N_2333);
or U2917 (N_2917,N_1833,N_1620);
nand U2918 (N_2918,N_2258,N_2026);
nand U2919 (N_2919,N_1669,N_1821);
and U2920 (N_2920,N_1963,N_1973);
xnor U2921 (N_2921,N_1972,N_2114);
nand U2922 (N_2922,N_1751,N_2270);
nor U2923 (N_2923,N_1717,N_2150);
xnor U2924 (N_2924,N_1865,N_2380);
nor U2925 (N_2925,N_1911,N_2315);
and U2926 (N_2926,N_2010,N_2358);
and U2927 (N_2927,N_2360,N_1800);
xnor U2928 (N_2928,N_1778,N_1682);
and U2929 (N_2929,N_1600,N_1790);
or U2930 (N_2930,N_1836,N_2384);
nand U2931 (N_2931,N_2109,N_2244);
nor U2932 (N_2932,N_1747,N_1940);
nand U2933 (N_2933,N_2282,N_1916);
and U2934 (N_2934,N_1823,N_2194);
xor U2935 (N_2935,N_1900,N_1652);
nor U2936 (N_2936,N_1724,N_1762);
nor U2937 (N_2937,N_1696,N_2360);
nand U2938 (N_2938,N_2395,N_2236);
nand U2939 (N_2939,N_1752,N_2110);
nor U2940 (N_2940,N_2143,N_2090);
and U2941 (N_2941,N_1702,N_1963);
or U2942 (N_2942,N_1602,N_1656);
nand U2943 (N_2943,N_2070,N_1757);
xnor U2944 (N_2944,N_2063,N_2252);
nor U2945 (N_2945,N_2155,N_2092);
xnor U2946 (N_2946,N_2367,N_2395);
or U2947 (N_2947,N_2168,N_2339);
xnor U2948 (N_2948,N_1721,N_1987);
or U2949 (N_2949,N_1780,N_2140);
and U2950 (N_2950,N_1894,N_2311);
xnor U2951 (N_2951,N_1623,N_2086);
nor U2952 (N_2952,N_1927,N_2261);
or U2953 (N_2953,N_2023,N_1725);
nor U2954 (N_2954,N_2204,N_1935);
nor U2955 (N_2955,N_2051,N_2055);
nor U2956 (N_2956,N_2130,N_1714);
nor U2957 (N_2957,N_1982,N_1861);
nor U2958 (N_2958,N_2220,N_2366);
xor U2959 (N_2959,N_1829,N_1743);
and U2960 (N_2960,N_1625,N_2261);
xnor U2961 (N_2961,N_1809,N_2112);
nand U2962 (N_2962,N_1823,N_1977);
xnor U2963 (N_2963,N_1720,N_1879);
nor U2964 (N_2964,N_1649,N_2080);
xnor U2965 (N_2965,N_2247,N_2190);
xor U2966 (N_2966,N_2135,N_1617);
or U2967 (N_2967,N_1920,N_1843);
xnor U2968 (N_2968,N_1700,N_2396);
nor U2969 (N_2969,N_2035,N_2285);
xor U2970 (N_2970,N_2041,N_2072);
nand U2971 (N_2971,N_1786,N_1607);
nand U2972 (N_2972,N_2166,N_2165);
or U2973 (N_2973,N_1618,N_2084);
or U2974 (N_2974,N_1956,N_2338);
and U2975 (N_2975,N_2288,N_1734);
nand U2976 (N_2976,N_2264,N_1680);
nand U2977 (N_2977,N_2089,N_1696);
xor U2978 (N_2978,N_1727,N_1627);
or U2979 (N_2979,N_1923,N_1995);
nand U2980 (N_2980,N_1800,N_1822);
nand U2981 (N_2981,N_1835,N_1677);
or U2982 (N_2982,N_1792,N_1699);
nor U2983 (N_2983,N_1937,N_2377);
or U2984 (N_2984,N_1908,N_1757);
and U2985 (N_2985,N_1811,N_2156);
and U2986 (N_2986,N_1680,N_2268);
and U2987 (N_2987,N_2043,N_2097);
or U2988 (N_2988,N_1942,N_2266);
nor U2989 (N_2989,N_2127,N_2172);
or U2990 (N_2990,N_1728,N_1688);
nand U2991 (N_2991,N_2328,N_2368);
xnor U2992 (N_2992,N_1758,N_1656);
or U2993 (N_2993,N_2315,N_1896);
or U2994 (N_2994,N_2392,N_1798);
and U2995 (N_2995,N_1939,N_1908);
xor U2996 (N_2996,N_2136,N_2095);
and U2997 (N_2997,N_1775,N_1772);
and U2998 (N_2998,N_2305,N_2119);
nand U2999 (N_2999,N_2125,N_2256);
nand U3000 (N_3000,N_2273,N_1798);
and U3001 (N_3001,N_2164,N_1796);
or U3002 (N_3002,N_2383,N_2389);
nor U3003 (N_3003,N_1989,N_1660);
nand U3004 (N_3004,N_2199,N_2208);
xnor U3005 (N_3005,N_1788,N_2015);
and U3006 (N_3006,N_1771,N_1901);
or U3007 (N_3007,N_2192,N_1784);
nand U3008 (N_3008,N_2113,N_1769);
xnor U3009 (N_3009,N_1963,N_2175);
or U3010 (N_3010,N_1602,N_2037);
nor U3011 (N_3011,N_2187,N_1666);
nand U3012 (N_3012,N_1864,N_2180);
nand U3013 (N_3013,N_1687,N_2129);
xnor U3014 (N_3014,N_2368,N_1917);
or U3015 (N_3015,N_2180,N_2034);
and U3016 (N_3016,N_2268,N_2213);
or U3017 (N_3017,N_2067,N_1622);
or U3018 (N_3018,N_2199,N_2132);
nand U3019 (N_3019,N_2298,N_1795);
nand U3020 (N_3020,N_1704,N_2064);
or U3021 (N_3021,N_1805,N_1757);
nor U3022 (N_3022,N_2285,N_2051);
xnor U3023 (N_3023,N_1600,N_2274);
nand U3024 (N_3024,N_1628,N_2345);
nor U3025 (N_3025,N_2130,N_2338);
nor U3026 (N_3026,N_1910,N_1826);
nor U3027 (N_3027,N_2325,N_2164);
nor U3028 (N_3028,N_2200,N_1863);
nor U3029 (N_3029,N_1720,N_2215);
nand U3030 (N_3030,N_1911,N_1645);
xnor U3031 (N_3031,N_1871,N_1684);
xor U3032 (N_3032,N_1778,N_2044);
nand U3033 (N_3033,N_1891,N_1777);
xor U3034 (N_3034,N_1618,N_1641);
or U3035 (N_3035,N_1773,N_2235);
nor U3036 (N_3036,N_2149,N_2261);
xor U3037 (N_3037,N_2315,N_1611);
xnor U3038 (N_3038,N_1752,N_1879);
nor U3039 (N_3039,N_1945,N_1828);
or U3040 (N_3040,N_1662,N_1791);
and U3041 (N_3041,N_2207,N_2192);
xnor U3042 (N_3042,N_1832,N_1899);
and U3043 (N_3043,N_1991,N_2222);
nor U3044 (N_3044,N_2022,N_1754);
and U3045 (N_3045,N_1659,N_2062);
and U3046 (N_3046,N_1835,N_2176);
and U3047 (N_3047,N_1754,N_2059);
and U3048 (N_3048,N_2348,N_2173);
or U3049 (N_3049,N_1673,N_1853);
or U3050 (N_3050,N_1763,N_1920);
or U3051 (N_3051,N_1874,N_1988);
nor U3052 (N_3052,N_2241,N_1921);
and U3053 (N_3053,N_1666,N_1668);
nand U3054 (N_3054,N_2359,N_2237);
and U3055 (N_3055,N_1773,N_1994);
nor U3056 (N_3056,N_2155,N_2223);
nand U3057 (N_3057,N_2133,N_1783);
or U3058 (N_3058,N_2148,N_2212);
nand U3059 (N_3059,N_2124,N_1801);
xnor U3060 (N_3060,N_1676,N_2208);
nor U3061 (N_3061,N_2104,N_1853);
or U3062 (N_3062,N_1977,N_1787);
xor U3063 (N_3063,N_2009,N_2225);
and U3064 (N_3064,N_1618,N_2120);
xor U3065 (N_3065,N_2384,N_2024);
xor U3066 (N_3066,N_2051,N_1691);
nor U3067 (N_3067,N_1892,N_2268);
xnor U3068 (N_3068,N_2344,N_1980);
or U3069 (N_3069,N_2394,N_2054);
nor U3070 (N_3070,N_2244,N_1848);
xnor U3071 (N_3071,N_1826,N_1832);
nor U3072 (N_3072,N_1759,N_2389);
xnor U3073 (N_3073,N_1997,N_2390);
xor U3074 (N_3074,N_2132,N_2119);
xor U3075 (N_3075,N_1818,N_1794);
xnor U3076 (N_3076,N_2117,N_2394);
nand U3077 (N_3077,N_1671,N_1950);
and U3078 (N_3078,N_1959,N_2140);
xor U3079 (N_3079,N_1748,N_1643);
or U3080 (N_3080,N_1795,N_2011);
nand U3081 (N_3081,N_1618,N_1854);
nor U3082 (N_3082,N_1801,N_2120);
and U3083 (N_3083,N_2061,N_1751);
nor U3084 (N_3084,N_1947,N_2066);
nor U3085 (N_3085,N_1608,N_1667);
nand U3086 (N_3086,N_1746,N_1745);
nand U3087 (N_3087,N_1957,N_1791);
xnor U3088 (N_3088,N_1647,N_2026);
or U3089 (N_3089,N_2209,N_2185);
or U3090 (N_3090,N_1842,N_2334);
xnor U3091 (N_3091,N_1854,N_2193);
and U3092 (N_3092,N_2360,N_1813);
nor U3093 (N_3093,N_1925,N_2200);
nand U3094 (N_3094,N_1900,N_2328);
and U3095 (N_3095,N_2328,N_1907);
nor U3096 (N_3096,N_1636,N_1675);
nand U3097 (N_3097,N_2115,N_2071);
and U3098 (N_3098,N_1827,N_2149);
nand U3099 (N_3099,N_2127,N_2051);
and U3100 (N_3100,N_1893,N_1984);
or U3101 (N_3101,N_1627,N_2211);
nand U3102 (N_3102,N_2160,N_1777);
and U3103 (N_3103,N_1908,N_1730);
nand U3104 (N_3104,N_1995,N_1736);
nand U3105 (N_3105,N_1856,N_2240);
or U3106 (N_3106,N_2054,N_1601);
or U3107 (N_3107,N_2161,N_1917);
xnor U3108 (N_3108,N_2094,N_1656);
and U3109 (N_3109,N_1990,N_1655);
or U3110 (N_3110,N_1837,N_1939);
nor U3111 (N_3111,N_1739,N_2228);
or U3112 (N_3112,N_2145,N_1641);
xnor U3113 (N_3113,N_2010,N_2273);
xor U3114 (N_3114,N_2355,N_2011);
xor U3115 (N_3115,N_2095,N_1614);
nor U3116 (N_3116,N_2211,N_2142);
nor U3117 (N_3117,N_2312,N_1834);
or U3118 (N_3118,N_1747,N_1982);
and U3119 (N_3119,N_1983,N_1923);
nor U3120 (N_3120,N_1886,N_1996);
nor U3121 (N_3121,N_2336,N_2319);
nor U3122 (N_3122,N_1795,N_1609);
or U3123 (N_3123,N_2003,N_1799);
or U3124 (N_3124,N_1887,N_2207);
nand U3125 (N_3125,N_1925,N_2351);
xnor U3126 (N_3126,N_1619,N_2189);
or U3127 (N_3127,N_1909,N_1997);
nand U3128 (N_3128,N_1968,N_2298);
nand U3129 (N_3129,N_1774,N_1872);
xnor U3130 (N_3130,N_2160,N_1603);
xnor U3131 (N_3131,N_1880,N_1988);
xnor U3132 (N_3132,N_1734,N_2023);
or U3133 (N_3133,N_1805,N_2194);
xor U3134 (N_3134,N_2281,N_2188);
or U3135 (N_3135,N_2039,N_1617);
xnor U3136 (N_3136,N_1689,N_2034);
or U3137 (N_3137,N_1882,N_2366);
nand U3138 (N_3138,N_2397,N_2142);
or U3139 (N_3139,N_1828,N_1900);
xnor U3140 (N_3140,N_2035,N_1925);
xor U3141 (N_3141,N_2058,N_1983);
nand U3142 (N_3142,N_1962,N_1719);
nor U3143 (N_3143,N_2025,N_2056);
xor U3144 (N_3144,N_2216,N_2121);
xor U3145 (N_3145,N_2166,N_1647);
nand U3146 (N_3146,N_1644,N_2172);
nand U3147 (N_3147,N_2029,N_2275);
or U3148 (N_3148,N_2291,N_1608);
nor U3149 (N_3149,N_2224,N_2222);
xnor U3150 (N_3150,N_1684,N_1731);
or U3151 (N_3151,N_1608,N_1868);
or U3152 (N_3152,N_2172,N_2178);
nand U3153 (N_3153,N_2192,N_1647);
and U3154 (N_3154,N_1923,N_2000);
or U3155 (N_3155,N_2194,N_1625);
or U3156 (N_3156,N_1602,N_2100);
nor U3157 (N_3157,N_1972,N_2277);
xor U3158 (N_3158,N_1865,N_2363);
or U3159 (N_3159,N_1626,N_1922);
xor U3160 (N_3160,N_1937,N_2101);
nand U3161 (N_3161,N_1734,N_1911);
and U3162 (N_3162,N_1856,N_2349);
or U3163 (N_3163,N_2046,N_1885);
xnor U3164 (N_3164,N_1643,N_1958);
nor U3165 (N_3165,N_1751,N_1790);
and U3166 (N_3166,N_1970,N_1603);
or U3167 (N_3167,N_2351,N_2191);
or U3168 (N_3168,N_1641,N_1801);
and U3169 (N_3169,N_1647,N_1676);
and U3170 (N_3170,N_1864,N_1810);
nor U3171 (N_3171,N_2186,N_2005);
xnor U3172 (N_3172,N_1623,N_1734);
nor U3173 (N_3173,N_2334,N_1914);
and U3174 (N_3174,N_2217,N_1670);
xnor U3175 (N_3175,N_1979,N_1941);
and U3176 (N_3176,N_1660,N_1933);
and U3177 (N_3177,N_1636,N_1626);
xnor U3178 (N_3178,N_2155,N_2291);
and U3179 (N_3179,N_2237,N_1931);
and U3180 (N_3180,N_1782,N_2234);
xnor U3181 (N_3181,N_2092,N_1944);
nand U3182 (N_3182,N_1854,N_2015);
xor U3183 (N_3183,N_2225,N_1674);
and U3184 (N_3184,N_2109,N_2285);
and U3185 (N_3185,N_2302,N_2311);
or U3186 (N_3186,N_2331,N_2361);
xor U3187 (N_3187,N_1871,N_1726);
xnor U3188 (N_3188,N_2291,N_2373);
xnor U3189 (N_3189,N_2069,N_2207);
and U3190 (N_3190,N_1851,N_2303);
nand U3191 (N_3191,N_2249,N_1980);
nor U3192 (N_3192,N_1833,N_2198);
xnor U3193 (N_3193,N_2245,N_2048);
or U3194 (N_3194,N_1626,N_1801);
or U3195 (N_3195,N_1943,N_2365);
or U3196 (N_3196,N_2000,N_2005);
and U3197 (N_3197,N_2051,N_1662);
nor U3198 (N_3198,N_1661,N_2393);
or U3199 (N_3199,N_2195,N_1883);
nor U3200 (N_3200,N_2425,N_3095);
or U3201 (N_3201,N_3054,N_2843);
nor U3202 (N_3202,N_3107,N_3125);
or U3203 (N_3203,N_3070,N_2516);
nand U3204 (N_3204,N_3089,N_3061);
nand U3205 (N_3205,N_2649,N_2565);
xnor U3206 (N_3206,N_2519,N_2821);
and U3207 (N_3207,N_2995,N_3157);
nor U3208 (N_3208,N_2677,N_2596);
nor U3209 (N_3209,N_2695,N_2772);
nand U3210 (N_3210,N_3092,N_3074);
nor U3211 (N_3211,N_2422,N_2631);
nand U3212 (N_3212,N_2952,N_3028);
and U3213 (N_3213,N_2652,N_3072);
nand U3214 (N_3214,N_2598,N_2826);
xnor U3215 (N_3215,N_3088,N_2432);
xor U3216 (N_3216,N_2840,N_3140);
xnor U3217 (N_3217,N_3009,N_3039);
nor U3218 (N_3218,N_2650,N_3014);
nor U3219 (N_3219,N_3026,N_2403);
nor U3220 (N_3220,N_2878,N_2480);
or U3221 (N_3221,N_2756,N_2497);
and U3222 (N_3222,N_3106,N_2586);
nor U3223 (N_3223,N_2564,N_2767);
nor U3224 (N_3224,N_2965,N_3192);
xnor U3225 (N_3225,N_2656,N_2887);
or U3226 (N_3226,N_3045,N_2799);
nand U3227 (N_3227,N_3082,N_2646);
nor U3228 (N_3228,N_2701,N_2980);
nand U3229 (N_3229,N_2414,N_2934);
xor U3230 (N_3230,N_2825,N_3042);
nor U3231 (N_3231,N_2522,N_2736);
nand U3232 (N_3232,N_2713,N_3069);
nor U3233 (N_3233,N_3123,N_2809);
xor U3234 (N_3234,N_3118,N_2563);
or U3235 (N_3235,N_2890,N_2907);
and U3236 (N_3236,N_2600,N_2764);
and U3237 (N_3237,N_2913,N_3098);
or U3238 (N_3238,N_2437,N_2456);
nor U3239 (N_3239,N_2739,N_2629);
or U3240 (N_3240,N_2939,N_3030);
nand U3241 (N_3241,N_2711,N_2828);
nand U3242 (N_3242,N_2839,N_2618);
nand U3243 (N_3243,N_2542,N_2611);
and U3244 (N_3244,N_3182,N_2568);
or U3245 (N_3245,N_3141,N_3068);
and U3246 (N_3246,N_2694,N_3010);
nand U3247 (N_3247,N_2751,N_3184);
or U3248 (N_3248,N_2663,N_2836);
xor U3249 (N_3249,N_2576,N_2612);
and U3250 (N_3250,N_2477,N_2640);
xor U3251 (N_3251,N_2962,N_3119);
xor U3252 (N_3252,N_3195,N_3162);
xor U3253 (N_3253,N_2945,N_2816);
nand U3254 (N_3254,N_2651,N_2472);
or U3255 (N_3255,N_2408,N_3059);
or U3256 (N_3256,N_2879,N_2909);
xor U3257 (N_3257,N_2720,N_2538);
xnor U3258 (N_3258,N_2637,N_2513);
nor U3259 (N_3259,N_2504,N_2998);
and U3260 (N_3260,N_2871,N_2850);
nor U3261 (N_3261,N_2492,N_2754);
and U3262 (N_3262,N_2536,N_2426);
and U3263 (N_3263,N_3078,N_2628);
xor U3264 (N_3264,N_3019,N_2876);
nand U3265 (N_3265,N_2479,N_2758);
nor U3266 (N_3266,N_3036,N_2963);
xnor U3267 (N_3267,N_2654,N_2874);
or U3268 (N_3268,N_2558,N_2891);
nand U3269 (N_3269,N_3115,N_2419);
and U3270 (N_3270,N_2551,N_2853);
xnor U3271 (N_3271,N_2901,N_2657);
or U3272 (N_3272,N_2931,N_2421);
or U3273 (N_3273,N_2499,N_2732);
and U3274 (N_3274,N_2888,N_2814);
nand U3275 (N_3275,N_2620,N_2418);
and U3276 (N_3276,N_2495,N_2520);
and U3277 (N_3277,N_2793,N_2979);
and U3278 (N_3278,N_2482,N_3194);
xor U3279 (N_3279,N_2737,N_2703);
and U3280 (N_3280,N_2669,N_2606);
and U3281 (N_3281,N_3016,N_2777);
xnor U3282 (N_3282,N_2983,N_3071);
and U3283 (N_3283,N_2433,N_3170);
xor U3284 (N_3284,N_3056,N_2447);
nand U3285 (N_3285,N_2765,N_2916);
xor U3286 (N_3286,N_2429,N_2986);
nor U3287 (N_3287,N_2784,N_2993);
and U3288 (N_3288,N_2857,N_3165);
or U3289 (N_3289,N_2743,N_2817);
or U3290 (N_3290,N_2506,N_2942);
xor U3291 (N_3291,N_2543,N_2760);
xor U3292 (N_3292,N_2574,N_3117);
or U3293 (N_3293,N_2645,N_3155);
xnor U3294 (N_3294,N_3049,N_2729);
xor U3295 (N_3295,N_2678,N_3132);
nor U3296 (N_3296,N_3159,N_2577);
xor U3297 (N_3297,N_2607,N_3024);
or U3298 (N_3298,N_2539,N_2666);
nand U3299 (N_3299,N_2885,N_3094);
xor U3300 (N_3300,N_2977,N_2725);
xor U3301 (N_3301,N_2929,N_2978);
nand U3302 (N_3302,N_2483,N_2500);
nand U3303 (N_3303,N_2575,N_2768);
and U3304 (N_3304,N_2683,N_2707);
and U3305 (N_3305,N_2485,N_2440);
xor U3306 (N_3306,N_2400,N_2859);
nand U3307 (N_3307,N_2451,N_2560);
nand U3308 (N_3308,N_2445,N_2959);
or U3309 (N_3309,N_2687,N_2493);
xor U3310 (N_3310,N_2863,N_3080);
and U3311 (N_3311,N_3047,N_2727);
nand U3312 (N_3312,N_2582,N_2795);
nand U3313 (N_3313,N_2921,N_2638);
xnor U3314 (N_3314,N_2868,N_2904);
nand U3315 (N_3315,N_2601,N_3005);
xnor U3316 (N_3316,N_2439,N_2923);
and U3317 (N_3317,N_2593,N_2409);
and U3318 (N_3318,N_2416,N_3096);
nor U3319 (N_3319,N_2566,N_2441);
xor U3320 (N_3320,N_3146,N_3137);
nor U3321 (N_3321,N_3189,N_2761);
nand U3322 (N_3322,N_2436,N_2639);
xnor U3323 (N_3323,N_2546,N_3066);
or U3324 (N_3324,N_2412,N_2501);
and U3325 (N_3325,N_3179,N_3062);
and U3326 (N_3326,N_3169,N_3081);
nand U3327 (N_3327,N_2824,N_2991);
and U3328 (N_3328,N_2625,N_2918);
nor U3329 (N_3329,N_3167,N_2442);
nor U3330 (N_3330,N_2457,N_3037);
and U3331 (N_3331,N_2689,N_2877);
or U3332 (N_3332,N_2498,N_2590);
and U3333 (N_3333,N_2829,N_2721);
and U3334 (N_3334,N_2599,N_2886);
and U3335 (N_3335,N_3105,N_2982);
nor U3336 (N_3336,N_2967,N_2800);
and U3337 (N_3337,N_2641,N_2933);
nor U3338 (N_3338,N_2510,N_2774);
and U3339 (N_3339,N_2700,N_3160);
xnor U3340 (N_3340,N_3143,N_3032);
and U3341 (N_3341,N_2884,N_2699);
xnor U3342 (N_3342,N_2692,N_2435);
xnor U3343 (N_3343,N_2420,N_2849);
xor U3344 (N_3344,N_2449,N_2405);
xor U3345 (N_3345,N_2697,N_2917);
or U3346 (N_3346,N_2752,N_3128);
nor U3347 (N_3347,N_2734,N_2935);
or U3348 (N_3348,N_2941,N_3158);
nand U3349 (N_3349,N_2984,N_2526);
nor U3350 (N_3350,N_2806,N_2897);
nand U3351 (N_3351,N_2922,N_2655);
and U3352 (N_3352,N_2659,N_3110);
and U3353 (N_3353,N_3191,N_3156);
xnor U3354 (N_3354,N_2402,N_3171);
or U3355 (N_3355,N_2555,N_3154);
xnor U3356 (N_3356,N_2759,N_2423);
nand U3357 (N_3357,N_2410,N_3175);
or U3358 (N_3358,N_2708,N_2748);
and U3359 (N_3359,N_3147,N_2512);
nor U3360 (N_3360,N_2723,N_3002);
nor U3361 (N_3361,N_2804,N_2446);
nor U3362 (N_3362,N_3161,N_2910);
nand U3363 (N_3363,N_2893,N_2667);
nor U3364 (N_3364,N_2511,N_2844);
and U3365 (N_3365,N_2514,N_2838);
and U3366 (N_3366,N_3058,N_2744);
nand U3367 (N_3367,N_2489,N_2448);
nor U3368 (N_3368,N_3178,N_3104);
and U3369 (N_3369,N_3011,N_2573);
nor U3370 (N_3370,N_2580,N_2609);
xor U3371 (N_3371,N_2679,N_2930);
or U3372 (N_3372,N_3187,N_2515);
or U3373 (N_3373,N_2894,N_2726);
nor U3374 (N_3374,N_2818,N_2675);
nand U3375 (N_3375,N_2668,N_2658);
xor U3376 (N_3376,N_2534,N_2985);
nand U3377 (N_3377,N_2788,N_2858);
xor U3378 (N_3378,N_2633,N_2428);
or U3379 (N_3379,N_2594,N_2680);
nor U3380 (N_3380,N_2938,N_2462);
and U3381 (N_3381,N_2898,N_2584);
nand U3382 (N_3382,N_3087,N_2460);
and U3383 (N_3383,N_2769,N_3017);
or U3384 (N_3384,N_2535,N_3057);
or U3385 (N_3385,N_2530,N_2610);
or U3386 (N_3386,N_2947,N_2578);
nand U3387 (N_3387,N_2411,N_2648);
nor U3388 (N_3388,N_2808,N_2773);
nor U3389 (N_3389,N_2592,N_2827);
and U3390 (N_3390,N_3112,N_2527);
nor U3391 (N_3391,N_3084,N_3018);
or U3392 (N_3392,N_3109,N_2822);
nor U3393 (N_3393,N_2617,N_2523);
nand U3394 (N_3394,N_2554,N_3197);
and U3395 (N_3395,N_2624,N_3079);
or U3396 (N_3396,N_2789,N_2796);
nand U3397 (N_3397,N_3000,N_2770);
nor U3398 (N_3398,N_2819,N_2763);
or U3399 (N_3399,N_3097,N_2518);
nand U3400 (N_3400,N_2621,N_3035);
nor U3401 (N_3401,N_2541,N_2927);
and U3402 (N_3402,N_2453,N_2973);
nand U3403 (N_3403,N_2999,N_2745);
and U3404 (N_3404,N_2717,N_3124);
nand U3405 (N_3405,N_2988,N_3073);
or U3406 (N_3406,N_2908,N_2567);
xnor U3407 (N_3407,N_2873,N_2940);
xor U3408 (N_3408,N_2968,N_2803);
nand U3409 (N_3409,N_2686,N_3183);
nor U3410 (N_3410,N_3043,N_3145);
xor U3411 (N_3411,N_2684,N_2889);
and U3412 (N_3412,N_2488,N_3193);
xnor U3413 (N_3413,N_2544,N_3100);
nor U3414 (N_3414,N_3065,N_2862);
xnor U3415 (N_3415,N_2994,N_2895);
xor U3416 (N_3416,N_3060,N_2545);
nor U3417 (N_3417,N_2807,N_2430);
and U3418 (N_3418,N_2996,N_2562);
and U3419 (N_3419,N_2509,N_2473);
and U3420 (N_3420,N_2989,N_2602);
and U3421 (N_3421,N_2470,N_2757);
xnor U3422 (N_3422,N_3034,N_2531);
xnor U3423 (N_3423,N_2549,N_2802);
nor U3424 (N_3424,N_3113,N_2956);
xor U3425 (N_3425,N_2966,N_2834);
or U3426 (N_3426,N_2925,N_2883);
nand U3427 (N_3427,N_2688,N_2466);
nor U3428 (N_3428,N_2860,N_3173);
nor U3429 (N_3429,N_2791,N_2861);
nand U3430 (N_3430,N_2899,N_2661);
xnor U3431 (N_3431,N_3055,N_2815);
nor U3432 (N_3432,N_3199,N_3083);
and U3433 (N_3433,N_2997,N_3122);
xnor U3434 (N_3434,N_2676,N_2969);
or U3435 (N_3435,N_2992,N_3085);
xnor U3436 (N_3436,N_2719,N_2949);
or U3437 (N_3437,N_3181,N_2914);
or U3438 (N_3438,N_2714,N_2948);
or U3439 (N_3439,N_2557,N_2778);
nand U3440 (N_3440,N_2797,N_3185);
or U3441 (N_3441,N_2468,N_2615);
nand U3442 (N_3442,N_2706,N_3022);
nand U3443 (N_3443,N_2529,N_2681);
nor U3444 (N_3444,N_2932,N_2981);
and U3445 (N_3445,N_3135,N_2912);
or U3446 (N_3446,N_2845,N_2444);
nand U3447 (N_3447,N_3126,N_3013);
or U3448 (N_3448,N_3004,N_3027);
xnor U3449 (N_3449,N_2842,N_2953);
or U3450 (N_3450,N_2704,N_3196);
nand U3451 (N_3451,N_2835,N_2792);
nand U3452 (N_3452,N_3150,N_2605);
xor U3453 (N_3453,N_3142,N_2944);
nand U3454 (N_3454,N_3099,N_2823);
nor U3455 (N_3455,N_2670,N_2943);
nor U3456 (N_3456,N_3186,N_2766);
and U3457 (N_3457,N_2569,N_2787);
nor U3458 (N_3458,N_2958,N_3006);
or U3459 (N_3459,N_2852,N_2902);
xnor U3460 (N_3460,N_3108,N_3101);
nor U3461 (N_3461,N_2532,N_2798);
or U3462 (N_3462,N_2710,N_2865);
xnor U3463 (N_3463,N_2730,N_2762);
nand U3464 (N_3464,N_2525,N_2459);
or U3465 (N_3465,N_2870,N_2785);
or U3466 (N_3466,N_3075,N_3031);
or U3467 (N_3467,N_3077,N_2603);
or U3468 (N_3468,N_2464,N_2434);
nor U3469 (N_3469,N_2552,N_2954);
and U3470 (N_3470,N_2961,N_3076);
xor U3471 (N_3471,N_2790,N_3180);
nor U3472 (N_3472,N_2415,N_2753);
or U3473 (N_3473,N_3051,N_2452);
nor U3474 (N_3474,N_3103,N_2589);
or U3475 (N_3475,N_2846,N_2653);
xor U3476 (N_3476,N_2467,N_2747);
or U3477 (N_3477,N_3138,N_2928);
nand U3478 (N_3478,N_3046,N_3048);
xnor U3479 (N_3479,N_2465,N_3023);
nor U3480 (N_3480,N_2682,N_3064);
or U3481 (N_3481,N_2484,N_2964);
and U3482 (N_3482,N_2749,N_2705);
and U3483 (N_3483,N_2672,N_3149);
nand U3484 (N_3484,N_3041,N_3090);
nor U3485 (N_3485,N_2561,N_2851);
nor U3486 (N_3486,N_2841,N_2696);
nor U3487 (N_3487,N_3190,N_2623);
and U3488 (N_3488,N_2476,N_2443);
xnor U3489 (N_3489,N_2698,N_2946);
or U3490 (N_3490,N_2693,N_2794);
nor U3491 (N_3491,N_3116,N_3144);
or U3492 (N_3492,N_2671,N_2524);
or U3493 (N_3493,N_2716,N_2626);
nand U3494 (N_3494,N_3003,N_2583);
nor U3495 (N_3495,N_2553,N_2556);
or U3496 (N_3496,N_2937,N_2970);
nor U3497 (N_3497,N_2820,N_3063);
and U3498 (N_3498,N_2587,N_2974);
xnor U3499 (N_3499,N_2722,N_2801);
xnor U3500 (N_3500,N_2627,N_3102);
nor U3501 (N_3501,N_2571,N_2882);
nor U3502 (N_3502,N_2951,N_3152);
nand U3503 (N_3503,N_2735,N_3134);
and U3504 (N_3504,N_2957,N_2608);
nand U3505 (N_3505,N_3029,N_2588);
xnor U3506 (N_3506,N_2741,N_2634);
xor U3507 (N_3507,N_2481,N_3164);
xnor U3508 (N_3508,N_2496,N_3093);
nand U3509 (N_3509,N_3130,N_3050);
or U3510 (N_3510,N_2597,N_2550);
xnor U3511 (N_3511,N_2810,N_2503);
and U3512 (N_3512,N_2406,N_3021);
nor U3513 (N_3513,N_2872,N_2643);
nand U3514 (N_3514,N_2517,N_2647);
and U3515 (N_3515,N_2781,N_3038);
xor U3516 (N_3516,N_2662,N_2673);
xnor U3517 (N_3517,N_2417,N_2595);
xnor U3518 (N_3518,N_2461,N_2502);
nand U3519 (N_3519,N_2664,N_2740);
nor U3520 (N_3520,N_2869,N_2854);
nand U3521 (N_3521,N_2960,N_2616);
or U3522 (N_3522,N_2955,N_2471);
or U3523 (N_3523,N_2614,N_2507);
xor U3524 (N_3524,N_2490,N_3025);
or U3525 (N_3525,N_3121,N_2478);
or U3526 (N_3526,N_2926,N_2585);
nor U3527 (N_3527,N_2642,N_2572);
nand U3528 (N_3528,N_2867,N_3120);
and U3529 (N_3529,N_2474,N_3052);
nor U3530 (N_3530,N_2724,N_2491);
nor U3531 (N_3531,N_3136,N_2548);
nor U3532 (N_3532,N_2559,N_2454);
xor U3533 (N_3533,N_2537,N_3133);
or U3534 (N_3534,N_2463,N_2487);
nor U3535 (N_3535,N_2805,N_3153);
nor U3536 (N_3536,N_2830,N_3007);
and U3537 (N_3537,N_2903,N_2950);
xor U3538 (N_3538,N_3166,N_2469);
nor U3539 (N_3539,N_3148,N_2728);
xor U3540 (N_3540,N_3111,N_2712);
nor U3541 (N_3541,N_2579,N_2738);
nand U3542 (N_3542,N_2866,N_2709);
nand U3543 (N_3543,N_3001,N_2864);
xor U3544 (N_3544,N_2831,N_3151);
or U3545 (N_3545,N_2972,N_3174);
nor U3546 (N_3546,N_3127,N_2505);
and U3547 (N_3547,N_3020,N_3053);
and U3548 (N_3548,N_2832,N_2905);
or U3549 (N_3549,N_2750,N_2775);
and U3550 (N_3550,N_2855,N_2880);
nor U3551 (N_3551,N_3067,N_2811);
or U3552 (N_3552,N_2733,N_2779);
and U3553 (N_3553,N_2665,N_3188);
nor U3554 (N_3554,N_3012,N_2427);
nand U3555 (N_3555,N_2521,N_2540);
nor U3556 (N_3556,N_2976,N_2674);
nor U3557 (N_3557,N_2570,N_2475);
and U3558 (N_3558,N_2780,N_2630);
xnor U3559 (N_3559,N_2875,N_2848);
xnor U3560 (N_3560,N_2782,N_2746);
or U3561 (N_3561,N_2581,N_2896);
nor U3562 (N_3562,N_2690,N_3040);
and U3563 (N_3563,N_2776,N_3114);
nand U3564 (N_3564,N_2881,N_2783);
or U3565 (N_3565,N_2401,N_2936);
and U3566 (N_3566,N_2892,N_3129);
and U3567 (N_3567,N_2486,N_3015);
and U3568 (N_3568,N_2715,N_2833);
or U3569 (N_3569,N_2533,N_2702);
nor U3570 (N_3570,N_2494,N_2906);
or U3571 (N_3571,N_2619,N_2431);
or U3572 (N_3572,N_3033,N_2742);
nor U3573 (N_3573,N_2660,N_2547);
nand U3574 (N_3574,N_2990,N_3086);
nand U3575 (N_3575,N_2812,N_2900);
and U3576 (N_3576,N_2438,N_2591);
nor U3577 (N_3577,N_2755,N_3176);
nand U3578 (N_3578,N_3163,N_2632);
nor U3579 (N_3579,N_2856,N_2458);
and U3580 (N_3580,N_3091,N_2975);
nor U3581 (N_3581,N_2731,N_3139);
nand U3582 (N_3582,N_2455,N_2920);
or U3583 (N_3583,N_2636,N_2924);
and U3584 (N_3584,N_3168,N_2691);
nand U3585 (N_3585,N_2644,N_3172);
and U3586 (N_3586,N_3044,N_2424);
xnor U3587 (N_3587,N_2407,N_2635);
nand U3588 (N_3588,N_2613,N_2528);
nor U3589 (N_3589,N_2987,N_2622);
or U3590 (N_3590,N_2604,N_2915);
and U3591 (N_3591,N_3008,N_2718);
nand U3592 (N_3592,N_3198,N_2847);
or U3593 (N_3593,N_2786,N_2837);
nor U3594 (N_3594,N_2911,N_2919);
nand U3595 (N_3595,N_2404,N_2771);
or U3596 (N_3596,N_2971,N_3177);
and U3597 (N_3597,N_2685,N_2450);
nand U3598 (N_3598,N_2508,N_2413);
nor U3599 (N_3599,N_2813,N_3131);
xnor U3600 (N_3600,N_2597,N_2722);
and U3601 (N_3601,N_2454,N_3186);
xor U3602 (N_3602,N_3003,N_2977);
and U3603 (N_3603,N_3098,N_2785);
xor U3604 (N_3604,N_3041,N_2789);
or U3605 (N_3605,N_2694,N_2624);
nand U3606 (N_3606,N_2944,N_2741);
nand U3607 (N_3607,N_3105,N_2758);
or U3608 (N_3608,N_2927,N_2865);
nor U3609 (N_3609,N_2549,N_2586);
and U3610 (N_3610,N_2523,N_2483);
or U3611 (N_3611,N_2463,N_2855);
nor U3612 (N_3612,N_2426,N_2438);
xnor U3613 (N_3613,N_2537,N_3151);
or U3614 (N_3614,N_2854,N_2573);
xnor U3615 (N_3615,N_2784,N_2531);
and U3616 (N_3616,N_2816,N_2454);
xnor U3617 (N_3617,N_3133,N_3086);
nor U3618 (N_3618,N_2876,N_2871);
xor U3619 (N_3619,N_2549,N_2675);
nand U3620 (N_3620,N_2667,N_2689);
and U3621 (N_3621,N_2834,N_2414);
xnor U3622 (N_3622,N_2704,N_2849);
nor U3623 (N_3623,N_2552,N_2695);
nand U3624 (N_3624,N_3063,N_2750);
xor U3625 (N_3625,N_3008,N_3003);
and U3626 (N_3626,N_2473,N_2996);
and U3627 (N_3627,N_2458,N_2954);
nand U3628 (N_3628,N_2648,N_2445);
nor U3629 (N_3629,N_2460,N_2939);
nor U3630 (N_3630,N_3113,N_3177);
or U3631 (N_3631,N_2818,N_2420);
and U3632 (N_3632,N_3058,N_2502);
or U3633 (N_3633,N_3194,N_3187);
nor U3634 (N_3634,N_2776,N_3054);
and U3635 (N_3635,N_2570,N_2684);
xnor U3636 (N_3636,N_2682,N_2564);
xor U3637 (N_3637,N_3188,N_2597);
and U3638 (N_3638,N_2404,N_3152);
or U3639 (N_3639,N_3164,N_2935);
and U3640 (N_3640,N_2976,N_2849);
xor U3641 (N_3641,N_2776,N_2677);
nor U3642 (N_3642,N_3100,N_2763);
xnor U3643 (N_3643,N_2954,N_2651);
and U3644 (N_3644,N_2981,N_2681);
and U3645 (N_3645,N_2861,N_2827);
and U3646 (N_3646,N_2817,N_2556);
and U3647 (N_3647,N_2968,N_2990);
and U3648 (N_3648,N_3023,N_2686);
or U3649 (N_3649,N_3108,N_2562);
or U3650 (N_3650,N_2525,N_2813);
nor U3651 (N_3651,N_2576,N_2937);
and U3652 (N_3652,N_2863,N_2623);
and U3653 (N_3653,N_2459,N_2787);
nor U3654 (N_3654,N_2472,N_2646);
xnor U3655 (N_3655,N_2624,N_2882);
nor U3656 (N_3656,N_2956,N_2906);
or U3657 (N_3657,N_2647,N_3135);
or U3658 (N_3658,N_2965,N_3196);
or U3659 (N_3659,N_2759,N_2740);
or U3660 (N_3660,N_2709,N_2465);
or U3661 (N_3661,N_2779,N_2948);
and U3662 (N_3662,N_3086,N_2519);
nor U3663 (N_3663,N_2736,N_2859);
xnor U3664 (N_3664,N_2625,N_2531);
xnor U3665 (N_3665,N_2604,N_3063);
and U3666 (N_3666,N_2774,N_2677);
nor U3667 (N_3667,N_3048,N_2739);
nor U3668 (N_3668,N_2913,N_2639);
xnor U3669 (N_3669,N_2656,N_3118);
nand U3670 (N_3670,N_2472,N_3023);
xnor U3671 (N_3671,N_2842,N_2745);
xnor U3672 (N_3672,N_2659,N_3196);
xor U3673 (N_3673,N_3020,N_2513);
or U3674 (N_3674,N_2662,N_2872);
or U3675 (N_3675,N_3134,N_2603);
nor U3676 (N_3676,N_2916,N_2823);
and U3677 (N_3677,N_2970,N_2525);
nand U3678 (N_3678,N_3054,N_2718);
and U3679 (N_3679,N_2420,N_3009);
and U3680 (N_3680,N_3015,N_2600);
nand U3681 (N_3681,N_2785,N_2823);
or U3682 (N_3682,N_2773,N_2606);
or U3683 (N_3683,N_2932,N_2407);
xor U3684 (N_3684,N_2946,N_2522);
nor U3685 (N_3685,N_2632,N_2816);
nand U3686 (N_3686,N_3183,N_2960);
and U3687 (N_3687,N_2465,N_3158);
nand U3688 (N_3688,N_2889,N_2569);
nand U3689 (N_3689,N_3052,N_2686);
nor U3690 (N_3690,N_3091,N_3182);
nor U3691 (N_3691,N_2558,N_2685);
nor U3692 (N_3692,N_3058,N_3167);
and U3693 (N_3693,N_3046,N_2634);
nand U3694 (N_3694,N_2618,N_2407);
xor U3695 (N_3695,N_3016,N_2440);
xnor U3696 (N_3696,N_3109,N_2746);
and U3697 (N_3697,N_2489,N_2955);
or U3698 (N_3698,N_2581,N_2650);
nor U3699 (N_3699,N_2631,N_2566);
and U3700 (N_3700,N_3179,N_2697);
nand U3701 (N_3701,N_2635,N_2682);
nand U3702 (N_3702,N_3053,N_3174);
and U3703 (N_3703,N_2753,N_2471);
xor U3704 (N_3704,N_2527,N_2623);
or U3705 (N_3705,N_3077,N_2692);
or U3706 (N_3706,N_2674,N_3035);
and U3707 (N_3707,N_2630,N_2731);
nor U3708 (N_3708,N_2928,N_2596);
or U3709 (N_3709,N_2778,N_2811);
or U3710 (N_3710,N_2766,N_2637);
and U3711 (N_3711,N_2590,N_2428);
and U3712 (N_3712,N_2585,N_2470);
or U3713 (N_3713,N_2637,N_2747);
or U3714 (N_3714,N_3096,N_2636);
xor U3715 (N_3715,N_2665,N_2492);
and U3716 (N_3716,N_2643,N_2781);
nand U3717 (N_3717,N_2798,N_2454);
or U3718 (N_3718,N_2536,N_3048);
or U3719 (N_3719,N_2506,N_3064);
xor U3720 (N_3720,N_2447,N_2964);
and U3721 (N_3721,N_3141,N_2482);
xor U3722 (N_3722,N_3016,N_2997);
and U3723 (N_3723,N_2820,N_3058);
nor U3724 (N_3724,N_3011,N_2818);
nor U3725 (N_3725,N_2449,N_2740);
and U3726 (N_3726,N_2614,N_2587);
nor U3727 (N_3727,N_2852,N_3068);
and U3728 (N_3728,N_3096,N_3063);
and U3729 (N_3729,N_3190,N_2552);
or U3730 (N_3730,N_2934,N_2906);
nand U3731 (N_3731,N_2767,N_3116);
xnor U3732 (N_3732,N_2924,N_2537);
or U3733 (N_3733,N_2874,N_2805);
or U3734 (N_3734,N_2678,N_2632);
nand U3735 (N_3735,N_2570,N_3129);
nor U3736 (N_3736,N_2512,N_2972);
xnor U3737 (N_3737,N_2805,N_2413);
nor U3738 (N_3738,N_2877,N_2970);
xnor U3739 (N_3739,N_2543,N_2991);
nand U3740 (N_3740,N_2799,N_2602);
xnor U3741 (N_3741,N_3186,N_2885);
xnor U3742 (N_3742,N_2567,N_2732);
and U3743 (N_3743,N_2758,N_2636);
or U3744 (N_3744,N_2627,N_2968);
xnor U3745 (N_3745,N_2452,N_2688);
nand U3746 (N_3746,N_3081,N_2453);
xor U3747 (N_3747,N_3143,N_3030);
and U3748 (N_3748,N_2607,N_2701);
xor U3749 (N_3749,N_3035,N_2704);
nand U3750 (N_3750,N_2893,N_2532);
and U3751 (N_3751,N_2885,N_3147);
nand U3752 (N_3752,N_2686,N_2700);
nand U3753 (N_3753,N_2758,N_2645);
or U3754 (N_3754,N_3139,N_2422);
or U3755 (N_3755,N_2738,N_2899);
xor U3756 (N_3756,N_2557,N_3008);
nor U3757 (N_3757,N_2973,N_2958);
nand U3758 (N_3758,N_3021,N_2473);
nand U3759 (N_3759,N_2790,N_3089);
and U3760 (N_3760,N_2545,N_2435);
nor U3761 (N_3761,N_2558,N_3172);
and U3762 (N_3762,N_2923,N_2527);
or U3763 (N_3763,N_2471,N_3096);
or U3764 (N_3764,N_2958,N_2431);
xor U3765 (N_3765,N_2703,N_2634);
xnor U3766 (N_3766,N_2917,N_2716);
nand U3767 (N_3767,N_2503,N_2421);
or U3768 (N_3768,N_2594,N_2463);
or U3769 (N_3769,N_3083,N_3026);
or U3770 (N_3770,N_3173,N_2905);
or U3771 (N_3771,N_3100,N_3109);
xnor U3772 (N_3772,N_2512,N_2652);
nand U3773 (N_3773,N_2688,N_3139);
nand U3774 (N_3774,N_3020,N_2443);
and U3775 (N_3775,N_2951,N_3001);
or U3776 (N_3776,N_2543,N_2577);
or U3777 (N_3777,N_2614,N_3040);
xor U3778 (N_3778,N_3176,N_2566);
nand U3779 (N_3779,N_2613,N_2966);
or U3780 (N_3780,N_2951,N_2683);
and U3781 (N_3781,N_3076,N_2583);
and U3782 (N_3782,N_2932,N_3092);
nor U3783 (N_3783,N_2707,N_2789);
xor U3784 (N_3784,N_2428,N_2943);
or U3785 (N_3785,N_2566,N_2973);
nor U3786 (N_3786,N_2965,N_2812);
nor U3787 (N_3787,N_2766,N_2900);
nor U3788 (N_3788,N_2977,N_3140);
nand U3789 (N_3789,N_2690,N_2613);
nand U3790 (N_3790,N_2974,N_2580);
or U3791 (N_3791,N_2611,N_2495);
nor U3792 (N_3792,N_3100,N_2506);
nand U3793 (N_3793,N_2482,N_3012);
xnor U3794 (N_3794,N_2937,N_3160);
and U3795 (N_3795,N_2692,N_2426);
or U3796 (N_3796,N_2561,N_2684);
nand U3797 (N_3797,N_3144,N_3093);
nor U3798 (N_3798,N_3015,N_3198);
and U3799 (N_3799,N_2955,N_2666);
nor U3800 (N_3800,N_3008,N_2777);
nand U3801 (N_3801,N_3199,N_3194);
nor U3802 (N_3802,N_2563,N_3104);
xnor U3803 (N_3803,N_3016,N_2757);
nor U3804 (N_3804,N_2433,N_2957);
and U3805 (N_3805,N_2960,N_2516);
nor U3806 (N_3806,N_2849,N_2654);
or U3807 (N_3807,N_3063,N_2959);
nor U3808 (N_3808,N_2808,N_2475);
nor U3809 (N_3809,N_2493,N_2576);
nor U3810 (N_3810,N_2790,N_3021);
nand U3811 (N_3811,N_2524,N_3085);
and U3812 (N_3812,N_2412,N_2820);
nand U3813 (N_3813,N_2949,N_2763);
and U3814 (N_3814,N_2726,N_2751);
xor U3815 (N_3815,N_2645,N_2859);
nand U3816 (N_3816,N_2683,N_2785);
and U3817 (N_3817,N_2906,N_3026);
nor U3818 (N_3818,N_2507,N_2599);
nor U3819 (N_3819,N_2444,N_3014);
nand U3820 (N_3820,N_3102,N_2576);
nor U3821 (N_3821,N_3144,N_2784);
nor U3822 (N_3822,N_2767,N_2673);
nor U3823 (N_3823,N_2772,N_2812);
or U3824 (N_3824,N_3000,N_2845);
nor U3825 (N_3825,N_2518,N_2936);
nor U3826 (N_3826,N_2958,N_2636);
and U3827 (N_3827,N_2627,N_3119);
xnor U3828 (N_3828,N_2445,N_2498);
xnor U3829 (N_3829,N_2624,N_2622);
nor U3830 (N_3830,N_2632,N_2704);
nand U3831 (N_3831,N_2956,N_2585);
nand U3832 (N_3832,N_2805,N_2808);
nor U3833 (N_3833,N_2589,N_2577);
xnor U3834 (N_3834,N_2493,N_2435);
xor U3835 (N_3835,N_2666,N_3042);
and U3836 (N_3836,N_3180,N_2946);
xnor U3837 (N_3837,N_3101,N_3086);
nand U3838 (N_3838,N_2810,N_2795);
nor U3839 (N_3839,N_2751,N_3152);
nor U3840 (N_3840,N_2788,N_3012);
nor U3841 (N_3841,N_2935,N_2484);
and U3842 (N_3842,N_2545,N_2827);
nand U3843 (N_3843,N_2747,N_2923);
nand U3844 (N_3844,N_2428,N_2927);
nand U3845 (N_3845,N_2486,N_2958);
xnor U3846 (N_3846,N_3127,N_2844);
or U3847 (N_3847,N_2970,N_3026);
nor U3848 (N_3848,N_3069,N_2534);
and U3849 (N_3849,N_3142,N_2508);
nor U3850 (N_3850,N_2908,N_2510);
and U3851 (N_3851,N_3065,N_2794);
or U3852 (N_3852,N_3140,N_2778);
and U3853 (N_3853,N_2747,N_2483);
nand U3854 (N_3854,N_2695,N_2612);
nor U3855 (N_3855,N_2632,N_3156);
nand U3856 (N_3856,N_2856,N_2905);
nor U3857 (N_3857,N_2947,N_2484);
nor U3858 (N_3858,N_2538,N_2549);
nand U3859 (N_3859,N_2997,N_2895);
and U3860 (N_3860,N_3116,N_3042);
nand U3861 (N_3861,N_3091,N_2711);
or U3862 (N_3862,N_2612,N_2867);
nor U3863 (N_3863,N_2796,N_2647);
nand U3864 (N_3864,N_2467,N_2862);
and U3865 (N_3865,N_2838,N_3124);
or U3866 (N_3866,N_2726,N_2838);
or U3867 (N_3867,N_3146,N_2697);
or U3868 (N_3868,N_2456,N_3076);
and U3869 (N_3869,N_2922,N_2499);
xnor U3870 (N_3870,N_2787,N_3095);
or U3871 (N_3871,N_2939,N_3071);
and U3872 (N_3872,N_3050,N_2743);
and U3873 (N_3873,N_2837,N_2778);
and U3874 (N_3874,N_3100,N_3015);
nand U3875 (N_3875,N_2890,N_3070);
and U3876 (N_3876,N_2690,N_3111);
nand U3877 (N_3877,N_2615,N_2427);
nand U3878 (N_3878,N_2911,N_3181);
and U3879 (N_3879,N_2542,N_2645);
and U3880 (N_3880,N_2429,N_2623);
nand U3881 (N_3881,N_2404,N_3062);
or U3882 (N_3882,N_2954,N_2885);
nand U3883 (N_3883,N_2930,N_2611);
nor U3884 (N_3884,N_2606,N_2498);
xor U3885 (N_3885,N_2421,N_2646);
nor U3886 (N_3886,N_2441,N_2806);
nor U3887 (N_3887,N_3143,N_2486);
and U3888 (N_3888,N_2517,N_2566);
or U3889 (N_3889,N_2658,N_2455);
xnor U3890 (N_3890,N_2719,N_2925);
and U3891 (N_3891,N_2855,N_2508);
or U3892 (N_3892,N_2865,N_2561);
and U3893 (N_3893,N_2947,N_2588);
nand U3894 (N_3894,N_2618,N_3140);
nand U3895 (N_3895,N_2770,N_2981);
or U3896 (N_3896,N_3143,N_2581);
and U3897 (N_3897,N_3099,N_2722);
nor U3898 (N_3898,N_3082,N_3122);
nand U3899 (N_3899,N_2494,N_3129);
nand U3900 (N_3900,N_3043,N_2808);
nor U3901 (N_3901,N_2786,N_2769);
nor U3902 (N_3902,N_2813,N_2549);
nor U3903 (N_3903,N_3078,N_2662);
nand U3904 (N_3904,N_2508,N_3076);
xor U3905 (N_3905,N_2512,N_2775);
nand U3906 (N_3906,N_2684,N_2820);
or U3907 (N_3907,N_2575,N_3107);
or U3908 (N_3908,N_2803,N_2689);
and U3909 (N_3909,N_2895,N_3015);
and U3910 (N_3910,N_2774,N_2876);
xor U3911 (N_3911,N_2713,N_2807);
nor U3912 (N_3912,N_2561,N_3071);
or U3913 (N_3913,N_3005,N_2895);
nand U3914 (N_3914,N_2766,N_2675);
nor U3915 (N_3915,N_2942,N_2773);
and U3916 (N_3916,N_2592,N_2611);
xnor U3917 (N_3917,N_3187,N_2945);
or U3918 (N_3918,N_2692,N_2500);
nor U3919 (N_3919,N_2462,N_3145);
nor U3920 (N_3920,N_2920,N_3158);
nor U3921 (N_3921,N_2639,N_3198);
nor U3922 (N_3922,N_2755,N_2559);
or U3923 (N_3923,N_2706,N_2651);
nand U3924 (N_3924,N_2716,N_2764);
nor U3925 (N_3925,N_2870,N_3052);
xnor U3926 (N_3926,N_2722,N_2488);
nand U3927 (N_3927,N_3159,N_2917);
nor U3928 (N_3928,N_2487,N_2501);
and U3929 (N_3929,N_2845,N_2668);
xor U3930 (N_3930,N_2798,N_3115);
xor U3931 (N_3931,N_2885,N_2902);
and U3932 (N_3932,N_2581,N_2448);
and U3933 (N_3933,N_2782,N_3003);
or U3934 (N_3934,N_2596,N_2649);
nand U3935 (N_3935,N_2730,N_2543);
nor U3936 (N_3936,N_2593,N_2945);
and U3937 (N_3937,N_2580,N_2964);
or U3938 (N_3938,N_3061,N_3046);
and U3939 (N_3939,N_2506,N_2477);
nand U3940 (N_3940,N_2509,N_2579);
nor U3941 (N_3941,N_2896,N_2907);
or U3942 (N_3942,N_2438,N_2952);
or U3943 (N_3943,N_2522,N_2534);
nor U3944 (N_3944,N_2420,N_2793);
nor U3945 (N_3945,N_2666,N_3015);
nor U3946 (N_3946,N_2729,N_3055);
xor U3947 (N_3947,N_2618,N_3183);
or U3948 (N_3948,N_2537,N_2672);
nor U3949 (N_3949,N_2892,N_2654);
and U3950 (N_3950,N_2833,N_2523);
or U3951 (N_3951,N_2631,N_3036);
and U3952 (N_3952,N_2657,N_2613);
and U3953 (N_3953,N_2755,N_2818);
nor U3954 (N_3954,N_2765,N_2927);
nand U3955 (N_3955,N_2796,N_3187);
nand U3956 (N_3956,N_2611,N_2548);
xor U3957 (N_3957,N_2700,N_2590);
or U3958 (N_3958,N_2577,N_2422);
or U3959 (N_3959,N_2931,N_2965);
nor U3960 (N_3960,N_3106,N_2476);
xnor U3961 (N_3961,N_3114,N_3017);
nor U3962 (N_3962,N_2997,N_3110);
and U3963 (N_3963,N_2712,N_3083);
nand U3964 (N_3964,N_3004,N_2861);
or U3965 (N_3965,N_2411,N_2525);
and U3966 (N_3966,N_3040,N_2798);
nor U3967 (N_3967,N_3185,N_2595);
and U3968 (N_3968,N_2775,N_2746);
nor U3969 (N_3969,N_2838,N_2526);
nor U3970 (N_3970,N_2872,N_2664);
or U3971 (N_3971,N_2817,N_2697);
xnor U3972 (N_3972,N_2718,N_2623);
xnor U3973 (N_3973,N_2620,N_2559);
nand U3974 (N_3974,N_2461,N_2633);
nand U3975 (N_3975,N_2659,N_3058);
xnor U3976 (N_3976,N_2515,N_2865);
or U3977 (N_3977,N_2925,N_2773);
or U3978 (N_3978,N_2467,N_2571);
nor U3979 (N_3979,N_3107,N_3120);
xnor U3980 (N_3980,N_2518,N_3081);
or U3981 (N_3981,N_2993,N_2761);
xnor U3982 (N_3982,N_2733,N_2735);
and U3983 (N_3983,N_2946,N_3094);
nand U3984 (N_3984,N_2705,N_3036);
or U3985 (N_3985,N_2641,N_3092);
or U3986 (N_3986,N_2751,N_2953);
xnor U3987 (N_3987,N_3028,N_3092);
nor U3988 (N_3988,N_2981,N_2746);
xor U3989 (N_3989,N_3166,N_2941);
xnor U3990 (N_3990,N_2665,N_2733);
nand U3991 (N_3991,N_3010,N_3068);
nor U3992 (N_3992,N_2942,N_2726);
and U3993 (N_3993,N_2511,N_3055);
xnor U3994 (N_3994,N_3136,N_2771);
nand U3995 (N_3995,N_2572,N_2723);
and U3996 (N_3996,N_2745,N_2585);
or U3997 (N_3997,N_3082,N_2580);
nand U3998 (N_3998,N_2514,N_2625);
and U3999 (N_3999,N_2715,N_2970);
nand U4000 (N_4000,N_3285,N_3694);
or U4001 (N_4001,N_3782,N_3678);
and U4002 (N_4002,N_3809,N_3721);
nand U4003 (N_4003,N_3723,N_3507);
nor U4004 (N_4004,N_3778,N_3235);
xor U4005 (N_4005,N_3747,N_3556);
and U4006 (N_4006,N_3211,N_3319);
and U4007 (N_4007,N_3299,N_3934);
or U4008 (N_4008,N_3866,N_3518);
nor U4009 (N_4009,N_3442,N_3832);
and U4010 (N_4010,N_3440,N_3743);
and U4011 (N_4011,N_3535,N_3687);
nand U4012 (N_4012,N_3595,N_3589);
or U4013 (N_4013,N_3824,N_3246);
or U4014 (N_4014,N_3660,N_3405);
and U4015 (N_4015,N_3690,N_3281);
xor U4016 (N_4016,N_3975,N_3466);
and U4017 (N_4017,N_3280,N_3762);
nor U4018 (N_4018,N_3392,N_3910);
xnor U4019 (N_4019,N_3909,N_3839);
nor U4020 (N_4020,N_3879,N_3653);
xor U4021 (N_4021,N_3978,N_3963);
nor U4022 (N_4022,N_3401,N_3689);
or U4023 (N_4023,N_3645,N_3306);
or U4024 (N_4024,N_3383,N_3302);
and U4025 (N_4025,N_3863,N_3918);
xor U4026 (N_4026,N_3759,N_3977);
and U4027 (N_4027,N_3756,N_3477);
and U4028 (N_4028,N_3525,N_3711);
or U4029 (N_4029,N_3993,N_3467);
nor U4030 (N_4030,N_3336,N_3633);
xor U4031 (N_4031,N_3382,N_3958);
nor U4032 (N_4032,N_3643,N_3966);
nor U4033 (N_4033,N_3287,N_3601);
xor U4034 (N_4034,N_3305,N_3991);
or U4035 (N_4035,N_3376,N_3635);
nor U4036 (N_4036,N_3321,N_3438);
nand U4037 (N_4037,N_3845,N_3668);
nor U4038 (N_4038,N_3770,N_3929);
xnor U4039 (N_4039,N_3823,N_3219);
xnor U4040 (N_4040,N_3881,N_3834);
or U4041 (N_4041,N_3730,N_3524);
nor U4042 (N_4042,N_3533,N_3250);
and U4043 (N_4043,N_3223,N_3421);
nand U4044 (N_4044,N_3844,N_3362);
nand U4045 (N_4045,N_3781,N_3527);
and U4046 (N_4046,N_3444,N_3840);
nand U4047 (N_4047,N_3658,N_3649);
xnor U4048 (N_4048,N_3373,N_3509);
nand U4049 (N_4049,N_3921,N_3487);
nand U4050 (N_4050,N_3818,N_3346);
xnor U4051 (N_4051,N_3473,N_3957);
xnor U4052 (N_4052,N_3245,N_3899);
xnor U4053 (N_4053,N_3741,N_3684);
or U4054 (N_4054,N_3697,N_3399);
or U4055 (N_4055,N_3669,N_3430);
xnor U4056 (N_4056,N_3544,N_3365);
nor U4057 (N_4057,N_3941,N_3768);
and U4058 (N_4058,N_3853,N_3644);
or U4059 (N_4059,N_3386,N_3790);
and U4060 (N_4060,N_3271,N_3751);
and U4061 (N_4061,N_3474,N_3354);
nand U4062 (N_4062,N_3590,N_3608);
and U4063 (N_4063,N_3923,N_3462);
and U4064 (N_4064,N_3422,N_3693);
xor U4065 (N_4065,N_3406,N_3709);
nand U4066 (N_4066,N_3603,N_3883);
and U4067 (N_4067,N_3279,N_3969);
and U4068 (N_4068,N_3855,N_3682);
or U4069 (N_4069,N_3695,N_3380);
nor U4070 (N_4070,N_3638,N_3291);
and U4071 (N_4071,N_3418,N_3565);
or U4072 (N_4072,N_3309,N_3979);
nand U4073 (N_4073,N_3901,N_3785);
and U4074 (N_4074,N_3715,N_3911);
and U4075 (N_4075,N_3688,N_3630);
nor U4076 (N_4076,N_3404,N_3596);
xnor U4077 (N_4077,N_3940,N_3893);
nor U4078 (N_4078,N_3435,N_3240);
xor U4079 (N_4079,N_3862,N_3582);
nor U4080 (N_4080,N_3870,N_3588);
xnor U4081 (N_4081,N_3976,N_3642);
nand U4082 (N_4082,N_3522,N_3787);
or U4083 (N_4083,N_3258,N_3446);
or U4084 (N_4084,N_3998,N_3740);
nand U4085 (N_4085,N_3935,N_3463);
or U4086 (N_4086,N_3683,N_3924);
nor U4087 (N_4087,N_3858,N_3915);
xnor U4088 (N_4088,N_3411,N_3772);
nor U4089 (N_4089,N_3414,N_3361);
nand U4090 (N_4090,N_3810,N_3625);
or U4091 (N_4091,N_3852,N_3699);
or U4092 (N_4092,N_3674,N_3433);
or U4093 (N_4093,N_3311,N_3805);
or U4094 (N_4094,N_3746,N_3803);
nor U4095 (N_4095,N_3583,N_3381);
xor U4096 (N_4096,N_3260,N_3586);
nor U4097 (N_4097,N_3303,N_3322);
xor U4098 (N_4098,N_3946,N_3367);
xnor U4099 (N_4099,N_3618,N_3729);
and U4100 (N_4100,N_3542,N_3454);
xor U4101 (N_4101,N_3835,N_3552);
or U4102 (N_4102,N_3791,N_3428);
nor U4103 (N_4103,N_3480,N_3594);
nand U4104 (N_4104,N_3988,N_3591);
nor U4105 (N_4105,N_3974,N_3263);
and U4106 (N_4106,N_3502,N_3310);
xnor U4107 (N_4107,N_3248,N_3256);
nor U4108 (N_4108,N_3388,N_3953);
nor U4109 (N_4109,N_3575,N_3308);
and U4110 (N_4110,N_3553,N_3985);
xor U4111 (N_4111,N_3597,N_3707);
or U4112 (N_4112,N_3842,N_3478);
nand U4113 (N_4113,N_3857,N_3609);
or U4114 (N_4114,N_3402,N_3528);
nor U4115 (N_4115,N_3249,N_3584);
nand U4116 (N_4116,N_3698,N_3836);
xor U4117 (N_4117,N_3812,N_3926);
nor U4118 (N_4118,N_3754,N_3821);
nand U4119 (N_4119,N_3794,N_3387);
nand U4120 (N_4120,N_3573,N_3622);
or U4121 (N_4121,N_3702,N_3546);
xnor U4122 (N_4122,N_3341,N_3403);
or U4123 (N_4123,N_3548,N_3936);
xor U4124 (N_4124,N_3885,N_3728);
or U4125 (N_4125,N_3676,N_3592);
nor U4126 (N_4126,N_3445,N_3201);
and U4127 (N_4127,N_3566,N_3726);
or U4128 (N_4128,N_3615,N_3491);
nor U4129 (N_4129,N_3357,N_3878);
nand U4130 (N_4130,N_3973,N_3300);
nor U4131 (N_4131,N_3580,N_3710);
xnor U4132 (N_4132,N_3620,N_3833);
and U4133 (N_4133,N_3352,N_3904);
and U4134 (N_4134,N_3780,N_3817);
or U4135 (N_4135,N_3455,N_3202);
or U4136 (N_4136,N_3345,N_3242);
xnor U4137 (N_4137,N_3505,N_3465);
nor U4138 (N_4138,N_3912,N_3907);
nand U4139 (N_4139,N_3439,N_3708);
xnor U4140 (N_4140,N_3512,N_3364);
xnor U4141 (N_4141,N_3587,N_3892);
and U4142 (N_4142,N_3247,N_3931);
or U4143 (N_4143,N_3236,N_3757);
nor U4144 (N_4144,N_3788,N_3232);
and U4145 (N_4145,N_3513,N_3875);
and U4146 (N_4146,N_3297,N_3578);
or U4147 (N_4147,N_3469,N_3207);
xnor U4148 (N_4148,N_3717,N_3749);
nand U4149 (N_4149,N_3771,N_3971);
or U4150 (N_4150,N_3860,N_3825);
nand U4151 (N_4151,N_3396,N_3680);
nand U4152 (N_4152,N_3972,N_3511);
and U4153 (N_4153,N_3324,N_3316);
nand U4154 (N_4154,N_3523,N_3335);
and U4155 (N_4155,N_3704,N_3673);
nor U4156 (N_4156,N_3970,N_3342);
nor U4157 (N_4157,N_3943,N_3610);
nand U4158 (N_4158,N_3654,N_3779);
and U4159 (N_4159,N_3983,N_3871);
or U4160 (N_4160,N_3994,N_3363);
nor U4161 (N_4161,N_3488,N_3278);
xnor U4162 (N_4162,N_3337,N_3604);
xor U4163 (N_4163,N_3431,N_3323);
nand U4164 (N_4164,N_3774,N_3626);
xor U4165 (N_4165,N_3510,N_3407);
nor U4166 (N_4166,N_3358,N_3298);
xor U4167 (N_4167,N_3508,N_3456);
nand U4168 (N_4168,N_3877,N_3200);
xor U4169 (N_4169,N_3284,N_3270);
xor U4170 (N_4170,N_3896,N_3636);
nor U4171 (N_4171,N_3783,N_3732);
xnor U4172 (N_4172,N_3962,N_3868);
and U4173 (N_4173,N_3629,N_3558);
nor U4174 (N_4174,N_3951,N_3313);
and U4175 (N_4175,N_3797,N_3549);
and U4176 (N_4176,N_3360,N_3887);
and U4177 (N_4177,N_3882,N_3811);
nand U4178 (N_4178,N_3916,N_3713);
nand U4179 (N_4179,N_3332,N_3716);
nand U4180 (N_4180,N_3777,N_3696);
xnor U4181 (N_4181,N_3437,N_3205);
nor U4182 (N_4182,N_3218,N_3449);
xnor U4183 (N_4183,N_3492,N_3353);
or U4184 (N_4184,N_3600,N_3476);
xor U4185 (N_4185,N_3925,N_3990);
nor U4186 (N_4186,N_3920,N_3413);
xor U4187 (N_4187,N_3334,N_3217);
nor U4188 (N_4188,N_3801,N_3914);
or U4189 (N_4189,N_3289,N_3350);
xnor U4190 (N_4190,N_3420,N_3656);
and U4191 (N_4191,N_3233,N_3226);
nand U4192 (N_4192,N_3900,N_3532);
nor U4193 (N_4193,N_3616,N_3400);
nor U4194 (N_4194,N_3631,N_3927);
xor U4195 (N_4195,N_3451,N_3489);
or U4196 (N_4196,N_3841,N_3331);
xnor U4197 (N_4197,N_3724,N_3624);
xnor U4198 (N_4198,N_3355,N_3763);
xnor U4199 (N_4199,N_3908,N_3955);
or U4200 (N_4200,N_3889,N_3436);
nor U4201 (N_4201,N_3786,N_3798);
nand U4202 (N_4202,N_3939,N_3867);
or U4203 (N_4203,N_3898,N_3735);
nand U4204 (N_4204,N_3415,N_3826);
or U4205 (N_4205,N_3423,N_3458);
or U4206 (N_4206,N_3733,N_3734);
or U4207 (N_4207,N_3275,N_3210);
nand U4208 (N_4208,N_3228,N_3831);
nor U4209 (N_4209,N_3767,N_3390);
nor U4210 (N_4210,N_3292,N_3813);
and U4211 (N_4211,N_3214,N_3829);
xor U4212 (N_4212,N_3419,N_3526);
or U4213 (N_4213,N_3338,N_3706);
or U4214 (N_4214,N_3581,N_3425);
and U4215 (N_4215,N_3417,N_3937);
nand U4216 (N_4216,N_3808,N_3662);
nand U4217 (N_4217,N_3238,N_3320);
nand U4218 (N_4218,N_3956,N_3452);
nor U4219 (N_4219,N_3393,N_3718);
xor U4220 (N_4220,N_3448,N_3574);
nand U4221 (N_4221,N_3257,N_3495);
or U4222 (N_4222,N_3391,N_3277);
and U4223 (N_4223,N_3989,N_3517);
or U4224 (N_4224,N_3529,N_3369);
xor U4225 (N_4225,N_3619,N_3269);
nand U4226 (N_4226,N_3816,N_3274);
nor U4227 (N_4227,N_3579,N_3340);
or U4228 (N_4228,N_3384,N_3377);
nor U4229 (N_4229,N_3426,N_3252);
nand U4230 (N_4230,N_3560,N_3276);
nand U4231 (N_4231,N_3986,N_3992);
xor U4232 (N_4232,N_3234,N_3820);
xnor U4233 (N_4233,N_3472,N_3379);
and U4234 (N_4234,N_3577,N_3551);
nor U4235 (N_4235,N_3216,N_3550);
or U4236 (N_4236,N_3765,N_3731);
or U4237 (N_4237,N_3325,N_3344);
nor U4238 (N_4238,N_3224,N_3888);
and U4239 (N_4239,N_3627,N_3776);
or U4240 (N_4240,N_3959,N_3459);
or U4241 (N_4241,N_3980,N_3482);
xnor U4242 (N_4242,N_3412,N_3846);
or U4243 (N_4243,N_3521,N_3481);
and U4244 (N_4244,N_3851,N_3906);
and U4245 (N_4245,N_3547,N_3461);
nand U4246 (N_4246,N_3330,N_3672);
or U4247 (N_4247,N_3997,N_3536);
and U4248 (N_4248,N_3231,N_3950);
nand U4249 (N_4249,N_3691,N_3944);
nand U4250 (N_4250,N_3539,N_3348);
xnor U4251 (N_4251,N_3891,N_3744);
or U4252 (N_4252,N_3960,N_3286);
or U4253 (N_4253,N_3204,N_3349);
and U4254 (N_4254,N_3515,N_3766);
nand U4255 (N_4255,N_3736,N_3819);
or U4256 (N_4256,N_3634,N_3516);
nand U4257 (N_4257,N_3827,N_3370);
xor U4258 (N_4258,N_3239,N_3244);
nor U4259 (N_4259,N_3475,N_3880);
nor U4260 (N_4260,N_3612,N_3623);
xor U4261 (N_4261,N_3666,N_3792);
nand U4262 (N_4262,N_3295,N_3470);
nand U4263 (N_4263,N_3203,N_3564);
and U4264 (N_4264,N_3947,N_3828);
or U4265 (N_4265,N_3995,N_3850);
and U4266 (N_4266,N_3395,N_3215);
or U4267 (N_4267,N_3640,N_3496);
nor U4268 (N_4268,N_3617,N_3967);
or U4269 (N_4269,N_3519,N_3290);
xnor U4270 (N_4270,N_3621,N_3922);
xnor U4271 (N_4271,N_3722,N_3847);
or U4272 (N_4272,N_3614,N_3639);
nor U4273 (N_4273,N_3351,N_3272);
nand U4274 (N_4274,N_3498,N_3543);
xor U4275 (N_4275,N_3429,N_3659);
and U4276 (N_4276,N_3865,N_3359);
nor U4277 (N_4277,N_3237,N_3784);
xor U4278 (N_4278,N_3987,N_3534);
and U4279 (N_4279,N_3576,N_3606);
or U4280 (N_4280,N_3737,N_3930);
nand U4281 (N_4281,N_3490,N_3854);
nor U4282 (N_4282,N_3514,N_3494);
and U4283 (N_4283,N_3651,N_3227);
and U4284 (N_4284,N_3796,N_3366);
nor U4285 (N_4285,N_3307,N_3830);
nand U4286 (N_4286,N_3241,N_3389);
or U4287 (N_4287,N_3856,N_3356);
nor U4288 (N_4288,N_3304,N_3264);
or U4289 (N_4289,N_3982,N_3876);
and U4290 (N_4290,N_3464,N_3919);
xor U4291 (N_4291,N_3965,N_3646);
and U4292 (N_4292,N_3685,N_3628);
nor U4293 (N_4293,N_3571,N_3679);
and U4294 (N_4294,N_3874,N_3554);
and U4295 (N_4295,N_3301,N_3869);
xor U4296 (N_4296,N_3692,N_3501);
nor U4297 (N_4297,N_3572,N_3329);
xor U4298 (N_4298,N_3569,N_3557);
and U4299 (N_4299,N_3681,N_3948);
and U4300 (N_4300,N_3984,N_3761);
and U4301 (N_4301,N_3486,N_3374);
nor U4302 (N_4302,N_3670,N_3282);
nor U4303 (N_4303,N_3570,N_3760);
and U4304 (N_4304,N_3409,N_3593);
xor U4305 (N_4305,N_3471,N_3312);
and U4306 (N_4306,N_3563,N_3714);
xnor U4307 (N_4307,N_3720,N_3945);
xnor U4308 (N_4308,N_3652,N_3917);
xnor U4309 (N_4309,N_3410,N_3849);
or U4310 (N_4310,N_3611,N_3637);
and U4311 (N_4311,N_3567,N_3333);
nand U4312 (N_4312,N_3665,N_3408);
xor U4313 (N_4313,N_3802,N_3253);
xor U4314 (N_4314,N_3657,N_3378);
or U4315 (N_4315,N_3913,N_3251);
and U4316 (N_4316,N_3457,N_3686);
and U4317 (N_4317,N_3799,N_3326);
xor U4318 (N_4318,N_3795,N_3942);
or U4319 (N_4319,N_3859,N_3755);
xnor U4320 (N_4320,N_3450,N_3460);
nor U4321 (N_4321,N_3894,N_3703);
nand U4322 (N_4322,N_3999,N_3328);
and U4323 (N_4323,N_3398,N_3933);
nand U4324 (N_4324,N_3753,N_3647);
xor U4325 (N_4325,N_3664,N_3314);
and U4326 (N_4326,N_3424,N_3468);
and U4327 (N_4327,N_3255,N_3837);
xnor U4328 (N_4328,N_3520,N_3769);
nor U4329 (N_4329,N_3745,N_3206);
or U4330 (N_4330,N_3208,N_3559);
and U4331 (N_4331,N_3229,N_3266);
or U4332 (N_4332,N_3375,N_3432);
and U4333 (N_4333,N_3928,N_3758);
nor U4334 (N_4334,N_3775,N_3738);
nand U4335 (N_4335,N_3905,N_3562);
nor U4336 (N_4336,N_3497,N_3750);
and U4337 (N_4337,N_3773,N_3602);
or U4338 (N_4338,N_3561,N_3372);
and U4339 (N_4339,N_3212,N_3895);
nand U4340 (N_4340,N_3954,N_3537);
nand U4341 (N_4341,N_3864,N_3221);
nand U4342 (N_4342,N_3964,N_3479);
and U4343 (N_4343,N_3952,N_3222);
nor U4344 (N_4344,N_3434,N_3800);
and U4345 (N_4345,N_3873,N_3555);
nor U4346 (N_4346,N_3296,N_3506);
nand U4347 (N_4347,N_3283,N_3230);
and U4348 (N_4348,N_3262,N_3504);
xnor U4349 (N_4349,N_3394,N_3371);
nand U4350 (N_4350,N_3485,N_3822);
nand U4351 (N_4351,N_3725,N_3872);
and U4352 (N_4352,N_3568,N_3938);
nand U4353 (N_4353,N_3447,N_3339);
xor U4354 (N_4354,N_3397,N_3343);
nand U4355 (N_4355,N_3949,N_3667);
and U4356 (N_4356,N_3503,N_3453);
nor U4357 (N_4357,N_3294,N_3317);
and U4358 (N_4358,N_3605,N_3661);
nand U4359 (N_4359,N_3500,N_3752);
xor U4360 (N_4360,N_3427,N_3385);
and U4361 (N_4361,N_3902,N_3499);
or U4362 (N_4362,N_3789,N_3804);
nor U4363 (N_4363,N_3968,N_3265);
nand U4364 (N_4364,N_3650,N_3632);
and U4365 (N_4365,N_3607,N_3268);
xor U4366 (N_4366,N_3961,N_3648);
nand U4367 (N_4367,N_3932,N_3318);
nand U4368 (N_4368,N_3742,N_3261);
nor U4369 (N_4369,N_3981,N_3897);
or U4370 (N_4370,N_3599,N_3288);
and U4371 (N_4371,N_3838,N_3727);
nor U4372 (N_4372,N_3764,N_3598);
nand U4373 (N_4373,N_3493,N_3484);
xnor U4374 (N_4374,N_3443,N_3719);
and U4375 (N_4375,N_3541,N_3675);
nor U4376 (N_4376,N_3677,N_3814);
nor U4377 (N_4377,N_3225,N_3531);
or U4378 (N_4378,N_3848,N_3538);
and U4379 (N_4379,N_3712,N_3441);
xor U4380 (N_4380,N_3807,N_3613);
or U4381 (N_4381,N_3213,N_3843);
xnor U4382 (N_4382,N_3903,N_3545);
nand U4383 (N_4383,N_3641,N_3793);
nor U4384 (N_4384,N_3267,N_3861);
nor U4385 (N_4385,N_3663,N_3886);
nor U4386 (N_4386,N_3209,N_3327);
or U4387 (N_4387,N_3890,N_3700);
and U4388 (N_4388,N_3254,N_3259);
nor U4389 (N_4389,N_3220,N_3273);
nor U4390 (N_4390,N_3884,N_3701);
or U4391 (N_4391,N_3705,N_3368);
nand U4392 (N_4392,N_3671,N_3416);
nor U4393 (N_4393,N_3585,N_3540);
nor U4394 (N_4394,N_3655,N_3530);
nand U4395 (N_4395,N_3748,N_3996);
xnor U4396 (N_4396,N_3293,N_3315);
or U4397 (N_4397,N_3739,N_3815);
nand U4398 (N_4398,N_3347,N_3483);
xor U4399 (N_4399,N_3806,N_3243);
and U4400 (N_4400,N_3873,N_3297);
or U4401 (N_4401,N_3704,N_3510);
nand U4402 (N_4402,N_3506,N_3983);
or U4403 (N_4403,N_3993,N_3847);
and U4404 (N_4404,N_3391,N_3626);
or U4405 (N_4405,N_3682,N_3605);
and U4406 (N_4406,N_3568,N_3711);
nand U4407 (N_4407,N_3615,N_3318);
nor U4408 (N_4408,N_3718,N_3430);
nand U4409 (N_4409,N_3232,N_3382);
nand U4410 (N_4410,N_3667,N_3749);
and U4411 (N_4411,N_3891,N_3521);
or U4412 (N_4412,N_3214,N_3481);
nor U4413 (N_4413,N_3779,N_3863);
or U4414 (N_4414,N_3722,N_3935);
or U4415 (N_4415,N_3597,N_3283);
xor U4416 (N_4416,N_3484,N_3765);
and U4417 (N_4417,N_3527,N_3517);
xor U4418 (N_4418,N_3846,N_3879);
xnor U4419 (N_4419,N_3921,N_3888);
nor U4420 (N_4420,N_3776,N_3745);
nor U4421 (N_4421,N_3803,N_3887);
or U4422 (N_4422,N_3945,N_3232);
and U4423 (N_4423,N_3436,N_3649);
nand U4424 (N_4424,N_3499,N_3985);
nor U4425 (N_4425,N_3250,N_3723);
nand U4426 (N_4426,N_3923,N_3402);
or U4427 (N_4427,N_3588,N_3670);
nor U4428 (N_4428,N_3531,N_3842);
or U4429 (N_4429,N_3522,N_3706);
nand U4430 (N_4430,N_3841,N_3451);
nor U4431 (N_4431,N_3649,N_3512);
xnor U4432 (N_4432,N_3785,N_3551);
nor U4433 (N_4433,N_3899,N_3233);
and U4434 (N_4434,N_3232,N_3874);
or U4435 (N_4435,N_3516,N_3285);
and U4436 (N_4436,N_3985,N_3948);
xnor U4437 (N_4437,N_3744,N_3428);
nand U4438 (N_4438,N_3666,N_3730);
nand U4439 (N_4439,N_3239,N_3780);
nand U4440 (N_4440,N_3512,N_3748);
nand U4441 (N_4441,N_3801,N_3792);
nor U4442 (N_4442,N_3729,N_3730);
and U4443 (N_4443,N_3546,N_3831);
and U4444 (N_4444,N_3449,N_3462);
nand U4445 (N_4445,N_3829,N_3565);
and U4446 (N_4446,N_3221,N_3483);
xor U4447 (N_4447,N_3711,N_3312);
or U4448 (N_4448,N_3430,N_3234);
xor U4449 (N_4449,N_3883,N_3647);
or U4450 (N_4450,N_3825,N_3200);
and U4451 (N_4451,N_3531,N_3775);
nand U4452 (N_4452,N_3827,N_3458);
nand U4453 (N_4453,N_3861,N_3923);
xnor U4454 (N_4454,N_3798,N_3523);
or U4455 (N_4455,N_3706,N_3510);
xor U4456 (N_4456,N_3314,N_3434);
and U4457 (N_4457,N_3559,N_3229);
xor U4458 (N_4458,N_3555,N_3330);
xor U4459 (N_4459,N_3723,N_3392);
nand U4460 (N_4460,N_3482,N_3922);
nand U4461 (N_4461,N_3932,N_3381);
and U4462 (N_4462,N_3990,N_3404);
xor U4463 (N_4463,N_3695,N_3395);
nand U4464 (N_4464,N_3406,N_3928);
nor U4465 (N_4465,N_3231,N_3850);
or U4466 (N_4466,N_3359,N_3482);
xnor U4467 (N_4467,N_3602,N_3550);
nor U4468 (N_4468,N_3748,N_3669);
xnor U4469 (N_4469,N_3238,N_3580);
nor U4470 (N_4470,N_3769,N_3424);
xnor U4471 (N_4471,N_3515,N_3810);
nand U4472 (N_4472,N_3365,N_3505);
nand U4473 (N_4473,N_3615,N_3444);
or U4474 (N_4474,N_3885,N_3750);
and U4475 (N_4475,N_3725,N_3636);
and U4476 (N_4476,N_3254,N_3274);
and U4477 (N_4477,N_3354,N_3746);
nor U4478 (N_4478,N_3526,N_3843);
nand U4479 (N_4479,N_3625,N_3904);
or U4480 (N_4480,N_3589,N_3831);
nand U4481 (N_4481,N_3616,N_3814);
or U4482 (N_4482,N_3928,N_3344);
or U4483 (N_4483,N_3452,N_3793);
or U4484 (N_4484,N_3420,N_3266);
or U4485 (N_4485,N_3359,N_3388);
or U4486 (N_4486,N_3762,N_3894);
or U4487 (N_4487,N_3312,N_3601);
and U4488 (N_4488,N_3572,N_3761);
xnor U4489 (N_4489,N_3836,N_3817);
nand U4490 (N_4490,N_3899,N_3227);
nor U4491 (N_4491,N_3671,N_3545);
or U4492 (N_4492,N_3694,N_3578);
xor U4493 (N_4493,N_3785,N_3414);
xnor U4494 (N_4494,N_3841,N_3718);
or U4495 (N_4495,N_3575,N_3292);
and U4496 (N_4496,N_3868,N_3825);
nand U4497 (N_4497,N_3495,N_3700);
xnor U4498 (N_4498,N_3220,N_3432);
nor U4499 (N_4499,N_3452,N_3768);
and U4500 (N_4500,N_3860,N_3331);
and U4501 (N_4501,N_3233,N_3511);
xor U4502 (N_4502,N_3274,N_3728);
xnor U4503 (N_4503,N_3801,N_3749);
and U4504 (N_4504,N_3631,N_3486);
xnor U4505 (N_4505,N_3223,N_3734);
xor U4506 (N_4506,N_3262,N_3459);
and U4507 (N_4507,N_3526,N_3410);
nand U4508 (N_4508,N_3594,N_3741);
and U4509 (N_4509,N_3775,N_3410);
nor U4510 (N_4510,N_3893,N_3609);
xor U4511 (N_4511,N_3902,N_3970);
nand U4512 (N_4512,N_3791,N_3234);
xnor U4513 (N_4513,N_3536,N_3287);
and U4514 (N_4514,N_3244,N_3853);
xor U4515 (N_4515,N_3813,N_3357);
nand U4516 (N_4516,N_3259,N_3765);
and U4517 (N_4517,N_3293,N_3604);
and U4518 (N_4518,N_3292,N_3671);
and U4519 (N_4519,N_3399,N_3510);
xnor U4520 (N_4520,N_3208,N_3210);
or U4521 (N_4521,N_3384,N_3556);
or U4522 (N_4522,N_3866,N_3520);
nand U4523 (N_4523,N_3910,N_3518);
nor U4524 (N_4524,N_3546,N_3695);
nand U4525 (N_4525,N_3780,N_3480);
nor U4526 (N_4526,N_3627,N_3877);
xnor U4527 (N_4527,N_3776,N_3291);
xor U4528 (N_4528,N_3809,N_3865);
nor U4529 (N_4529,N_3776,N_3895);
and U4530 (N_4530,N_3356,N_3422);
nor U4531 (N_4531,N_3202,N_3663);
and U4532 (N_4532,N_3920,N_3755);
nor U4533 (N_4533,N_3720,N_3317);
or U4534 (N_4534,N_3604,N_3888);
xnor U4535 (N_4535,N_3210,N_3860);
xnor U4536 (N_4536,N_3350,N_3974);
xor U4537 (N_4537,N_3253,N_3599);
nor U4538 (N_4538,N_3473,N_3819);
nand U4539 (N_4539,N_3925,N_3758);
or U4540 (N_4540,N_3854,N_3266);
xnor U4541 (N_4541,N_3976,N_3296);
nor U4542 (N_4542,N_3599,N_3862);
xnor U4543 (N_4543,N_3898,N_3496);
nor U4544 (N_4544,N_3975,N_3236);
nor U4545 (N_4545,N_3769,N_3736);
and U4546 (N_4546,N_3396,N_3703);
nand U4547 (N_4547,N_3363,N_3208);
and U4548 (N_4548,N_3438,N_3582);
xor U4549 (N_4549,N_3734,N_3780);
and U4550 (N_4550,N_3673,N_3943);
nor U4551 (N_4551,N_3953,N_3344);
or U4552 (N_4552,N_3276,N_3770);
nand U4553 (N_4553,N_3613,N_3610);
nor U4554 (N_4554,N_3542,N_3641);
nor U4555 (N_4555,N_3554,N_3838);
and U4556 (N_4556,N_3875,N_3508);
xnor U4557 (N_4557,N_3211,N_3232);
or U4558 (N_4558,N_3719,N_3664);
nand U4559 (N_4559,N_3741,N_3618);
xnor U4560 (N_4560,N_3529,N_3913);
xnor U4561 (N_4561,N_3607,N_3427);
nand U4562 (N_4562,N_3639,N_3997);
or U4563 (N_4563,N_3948,N_3763);
and U4564 (N_4564,N_3838,N_3259);
nand U4565 (N_4565,N_3656,N_3941);
xnor U4566 (N_4566,N_3608,N_3399);
or U4567 (N_4567,N_3815,N_3429);
or U4568 (N_4568,N_3434,N_3685);
nor U4569 (N_4569,N_3812,N_3264);
nor U4570 (N_4570,N_3595,N_3638);
nor U4571 (N_4571,N_3486,N_3555);
or U4572 (N_4572,N_3754,N_3226);
and U4573 (N_4573,N_3568,N_3983);
nor U4574 (N_4574,N_3533,N_3456);
or U4575 (N_4575,N_3707,N_3666);
nor U4576 (N_4576,N_3713,N_3213);
or U4577 (N_4577,N_3534,N_3765);
nand U4578 (N_4578,N_3469,N_3667);
nand U4579 (N_4579,N_3901,N_3826);
nand U4580 (N_4580,N_3691,N_3592);
nand U4581 (N_4581,N_3290,N_3588);
and U4582 (N_4582,N_3506,N_3351);
and U4583 (N_4583,N_3935,N_3720);
nand U4584 (N_4584,N_3209,N_3991);
and U4585 (N_4585,N_3261,N_3595);
nand U4586 (N_4586,N_3706,N_3328);
nor U4587 (N_4587,N_3357,N_3703);
nand U4588 (N_4588,N_3432,N_3900);
nand U4589 (N_4589,N_3732,N_3630);
or U4590 (N_4590,N_3881,N_3214);
nor U4591 (N_4591,N_3453,N_3429);
nor U4592 (N_4592,N_3751,N_3231);
nand U4593 (N_4593,N_3882,N_3688);
or U4594 (N_4594,N_3344,N_3713);
or U4595 (N_4595,N_3636,N_3222);
nand U4596 (N_4596,N_3999,N_3425);
nor U4597 (N_4597,N_3506,N_3857);
and U4598 (N_4598,N_3803,N_3304);
xnor U4599 (N_4599,N_3942,N_3869);
nor U4600 (N_4600,N_3894,N_3691);
and U4601 (N_4601,N_3599,N_3290);
or U4602 (N_4602,N_3255,N_3893);
or U4603 (N_4603,N_3399,N_3971);
xor U4604 (N_4604,N_3895,N_3572);
xor U4605 (N_4605,N_3928,N_3933);
or U4606 (N_4606,N_3334,N_3624);
nand U4607 (N_4607,N_3745,N_3816);
or U4608 (N_4608,N_3886,N_3915);
nand U4609 (N_4609,N_3860,N_3409);
nand U4610 (N_4610,N_3935,N_3472);
or U4611 (N_4611,N_3366,N_3290);
and U4612 (N_4612,N_3946,N_3737);
xor U4613 (N_4613,N_3461,N_3541);
or U4614 (N_4614,N_3652,N_3200);
nor U4615 (N_4615,N_3628,N_3727);
and U4616 (N_4616,N_3810,N_3285);
xor U4617 (N_4617,N_3231,N_3243);
and U4618 (N_4618,N_3358,N_3609);
and U4619 (N_4619,N_3584,N_3424);
or U4620 (N_4620,N_3946,N_3472);
and U4621 (N_4621,N_3974,N_3699);
nand U4622 (N_4622,N_3550,N_3391);
nor U4623 (N_4623,N_3474,N_3883);
and U4624 (N_4624,N_3486,N_3581);
xnor U4625 (N_4625,N_3826,N_3717);
and U4626 (N_4626,N_3444,N_3297);
and U4627 (N_4627,N_3375,N_3269);
and U4628 (N_4628,N_3377,N_3213);
xor U4629 (N_4629,N_3869,N_3244);
or U4630 (N_4630,N_3903,N_3998);
nor U4631 (N_4631,N_3812,N_3248);
or U4632 (N_4632,N_3789,N_3572);
xnor U4633 (N_4633,N_3394,N_3277);
nand U4634 (N_4634,N_3746,N_3862);
xor U4635 (N_4635,N_3233,N_3379);
xnor U4636 (N_4636,N_3759,N_3768);
xor U4637 (N_4637,N_3960,N_3449);
nand U4638 (N_4638,N_3851,N_3579);
nor U4639 (N_4639,N_3814,N_3286);
xor U4640 (N_4640,N_3238,N_3662);
xnor U4641 (N_4641,N_3555,N_3923);
and U4642 (N_4642,N_3458,N_3631);
and U4643 (N_4643,N_3925,N_3464);
and U4644 (N_4644,N_3373,N_3335);
nor U4645 (N_4645,N_3236,N_3821);
and U4646 (N_4646,N_3710,N_3757);
nand U4647 (N_4647,N_3359,N_3724);
xnor U4648 (N_4648,N_3421,N_3680);
nand U4649 (N_4649,N_3294,N_3865);
or U4650 (N_4650,N_3794,N_3478);
nor U4651 (N_4651,N_3412,N_3557);
nand U4652 (N_4652,N_3820,N_3266);
xnor U4653 (N_4653,N_3495,N_3845);
or U4654 (N_4654,N_3714,N_3977);
or U4655 (N_4655,N_3405,N_3829);
nor U4656 (N_4656,N_3243,N_3272);
and U4657 (N_4657,N_3725,N_3292);
nand U4658 (N_4658,N_3592,N_3633);
nor U4659 (N_4659,N_3981,N_3378);
or U4660 (N_4660,N_3363,N_3346);
xnor U4661 (N_4661,N_3533,N_3803);
or U4662 (N_4662,N_3969,N_3600);
or U4663 (N_4663,N_3594,N_3200);
nor U4664 (N_4664,N_3797,N_3225);
or U4665 (N_4665,N_3386,N_3417);
xnor U4666 (N_4666,N_3580,N_3348);
or U4667 (N_4667,N_3896,N_3376);
and U4668 (N_4668,N_3780,N_3909);
nor U4669 (N_4669,N_3377,N_3456);
nor U4670 (N_4670,N_3611,N_3247);
nand U4671 (N_4671,N_3987,N_3962);
or U4672 (N_4672,N_3389,N_3990);
or U4673 (N_4673,N_3464,N_3714);
or U4674 (N_4674,N_3664,N_3980);
and U4675 (N_4675,N_3499,N_3935);
nor U4676 (N_4676,N_3834,N_3967);
xnor U4677 (N_4677,N_3263,N_3261);
xnor U4678 (N_4678,N_3358,N_3281);
xnor U4679 (N_4679,N_3403,N_3379);
and U4680 (N_4680,N_3391,N_3574);
xnor U4681 (N_4681,N_3906,N_3695);
or U4682 (N_4682,N_3943,N_3502);
and U4683 (N_4683,N_3626,N_3203);
nor U4684 (N_4684,N_3353,N_3468);
or U4685 (N_4685,N_3687,N_3652);
and U4686 (N_4686,N_3931,N_3717);
nor U4687 (N_4687,N_3418,N_3551);
nor U4688 (N_4688,N_3567,N_3341);
nor U4689 (N_4689,N_3323,N_3866);
nand U4690 (N_4690,N_3899,N_3939);
xor U4691 (N_4691,N_3787,N_3935);
and U4692 (N_4692,N_3542,N_3231);
or U4693 (N_4693,N_3427,N_3634);
nand U4694 (N_4694,N_3984,N_3553);
or U4695 (N_4695,N_3264,N_3923);
xor U4696 (N_4696,N_3229,N_3998);
or U4697 (N_4697,N_3380,N_3574);
and U4698 (N_4698,N_3827,N_3669);
nand U4699 (N_4699,N_3970,N_3310);
nand U4700 (N_4700,N_3491,N_3768);
or U4701 (N_4701,N_3332,N_3526);
nor U4702 (N_4702,N_3356,N_3658);
xnor U4703 (N_4703,N_3408,N_3813);
and U4704 (N_4704,N_3868,N_3870);
nor U4705 (N_4705,N_3403,N_3254);
xor U4706 (N_4706,N_3625,N_3524);
or U4707 (N_4707,N_3805,N_3318);
xor U4708 (N_4708,N_3729,N_3689);
nor U4709 (N_4709,N_3314,N_3737);
and U4710 (N_4710,N_3370,N_3355);
nor U4711 (N_4711,N_3313,N_3941);
and U4712 (N_4712,N_3735,N_3599);
xor U4713 (N_4713,N_3600,N_3762);
and U4714 (N_4714,N_3958,N_3202);
or U4715 (N_4715,N_3263,N_3891);
and U4716 (N_4716,N_3416,N_3623);
and U4717 (N_4717,N_3999,N_3993);
nor U4718 (N_4718,N_3527,N_3634);
and U4719 (N_4719,N_3966,N_3803);
and U4720 (N_4720,N_3534,N_3215);
nor U4721 (N_4721,N_3749,N_3448);
xnor U4722 (N_4722,N_3670,N_3358);
or U4723 (N_4723,N_3464,N_3902);
and U4724 (N_4724,N_3780,N_3697);
and U4725 (N_4725,N_3246,N_3790);
xnor U4726 (N_4726,N_3963,N_3918);
nand U4727 (N_4727,N_3637,N_3368);
or U4728 (N_4728,N_3503,N_3336);
xor U4729 (N_4729,N_3663,N_3962);
and U4730 (N_4730,N_3814,N_3447);
and U4731 (N_4731,N_3769,N_3837);
and U4732 (N_4732,N_3459,N_3360);
and U4733 (N_4733,N_3665,N_3719);
and U4734 (N_4734,N_3341,N_3222);
or U4735 (N_4735,N_3434,N_3788);
or U4736 (N_4736,N_3366,N_3751);
nand U4737 (N_4737,N_3901,N_3825);
xor U4738 (N_4738,N_3373,N_3521);
xor U4739 (N_4739,N_3925,N_3940);
and U4740 (N_4740,N_3537,N_3508);
xor U4741 (N_4741,N_3770,N_3841);
nor U4742 (N_4742,N_3492,N_3571);
nand U4743 (N_4743,N_3547,N_3622);
nor U4744 (N_4744,N_3340,N_3680);
or U4745 (N_4745,N_3583,N_3429);
and U4746 (N_4746,N_3490,N_3461);
nand U4747 (N_4747,N_3527,N_3393);
or U4748 (N_4748,N_3250,N_3970);
xnor U4749 (N_4749,N_3706,N_3705);
nand U4750 (N_4750,N_3516,N_3733);
xor U4751 (N_4751,N_3692,N_3864);
and U4752 (N_4752,N_3751,N_3545);
nand U4753 (N_4753,N_3847,N_3554);
nand U4754 (N_4754,N_3797,N_3741);
and U4755 (N_4755,N_3226,N_3749);
nand U4756 (N_4756,N_3950,N_3401);
xnor U4757 (N_4757,N_3359,N_3869);
nand U4758 (N_4758,N_3676,N_3564);
nor U4759 (N_4759,N_3462,N_3539);
or U4760 (N_4760,N_3580,N_3895);
nor U4761 (N_4761,N_3515,N_3687);
and U4762 (N_4762,N_3666,N_3804);
nor U4763 (N_4763,N_3998,N_3314);
or U4764 (N_4764,N_3733,N_3936);
and U4765 (N_4765,N_3395,N_3739);
or U4766 (N_4766,N_3671,N_3738);
nor U4767 (N_4767,N_3977,N_3621);
or U4768 (N_4768,N_3581,N_3759);
or U4769 (N_4769,N_3503,N_3557);
and U4770 (N_4770,N_3636,N_3248);
or U4771 (N_4771,N_3201,N_3271);
and U4772 (N_4772,N_3536,N_3943);
nor U4773 (N_4773,N_3573,N_3503);
nor U4774 (N_4774,N_3980,N_3265);
nor U4775 (N_4775,N_3442,N_3568);
nor U4776 (N_4776,N_3657,N_3902);
nand U4777 (N_4777,N_3991,N_3512);
or U4778 (N_4778,N_3671,N_3505);
xnor U4779 (N_4779,N_3736,N_3468);
xor U4780 (N_4780,N_3517,N_3879);
nand U4781 (N_4781,N_3767,N_3757);
and U4782 (N_4782,N_3512,N_3293);
nor U4783 (N_4783,N_3875,N_3337);
and U4784 (N_4784,N_3223,N_3745);
xor U4785 (N_4785,N_3264,N_3747);
nor U4786 (N_4786,N_3945,N_3552);
nor U4787 (N_4787,N_3876,N_3349);
nor U4788 (N_4788,N_3914,N_3282);
nand U4789 (N_4789,N_3525,N_3505);
and U4790 (N_4790,N_3667,N_3511);
nor U4791 (N_4791,N_3335,N_3831);
xnor U4792 (N_4792,N_3356,N_3994);
nand U4793 (N_4793,N_3706,N_3350);
and U4794 (N_4794,N_3642,N_3563);
nand U4795 (N_4795,N_3711,N_3976);
or U4796 (N_4796,N_3695,N_3475);
and U4797 (N_4797,N_3794,N_3958);
and U4798 (N_4798,N_3995,N_3369);
and U4799 (N_4799,N_3668,N_3710);
nor U4800 (N_4800,N_4794,N_4729);
xnor U4801 (N_4801,N_4439,N_4627);
and U4802 (N_4802,N_4248,N_4123);
nor U4803 (N_4803,N_4149,N_4027);
xor U4804 (N_4804,N_4402,N_4060);
nand U4805 (N_4805,N_4131,N_4358);
nor U4806 (N_4806,N_4089,N_4718);
xnor U4807 (N_4807,N_4314,N_4421);
and U4808 (N_4808,N_4492,N_4604);
xor U4809 (N_4809,N_4649,N_4447);
and U4810 (N_4810,N_4217,N_4650);
or U4811 (N_4811,N_4449,N_4504);
nor U4812 (N_4812,N_4619,N_4456);
xnor U4813 (N_4813,N_4130,N_4352);
xor U4814 (N_4814,N_4667,N_4674);
and U4815 (N_4815,N_4574,N_4680);
xor U4816 (N_4816,N_4632,N_4422);
xor U4817 (N_4817,N_4068,N_4158);
xor U4818 (N_4818,N_4730,N_4350);
nor U4819 (N_4819,N_4359,N_4142);
nor U4820 (N_4820,N_4624,N_4625);
xnor U4821 (N_4821,N_4773,N_4768);
and U4822 (N_4822,N_4086,N_4761);
nand U4823 (N_4823,N_4030,N_4668);
and U4824 (N_4824,N_4677,N_4382);
or U4825 (N_4825,N_4072,N_4782);
or U4826 (N_4826,N_4398,N_4695);
nor U4827 (N_4827,N_4496,N_4375);
and U4828 (N_4828,N_4615,N_4361);
nand U4829 (N_4829,N_4512,N_4503);
xor U4830 (N_4830,N_4155,N_4393);
and U4831 (N_4831,N_4058,N_4021);
xnor U4832 (N_4832,N_4013,N_4454);
nor U4833 (N_4833,N_4357,N_4560);
nor U4834 (N_4834,N_4283,N_4328);
nand U4835 (N_4835,N_4047,N_4691);
and U4836 (N_4836,N_4128,N_4073);
and U4837 (N_4837,N_4090,N_4573);
nand U4838 (N_4838,N_4260,N_4211);
or U4839 (N_4839,N_4309,N_4440);
nand U4840 (N_4840,N_4708,N_4420);
or U4841 (N_4841,N_4025,N_4316);
xor U4842 (N_4842,N_4431,N_4475);
xnor U4843 (N_4843,N_4596,N_4381);
nand U4844 (N_4844,N_4009,N_4436);
nor U4845 (N_4845,N_4722,N_4781);
and U4846 (N_4846,N_4061,N_4687);
and U4847 (N_4847,N_4480,N_4719);
nand U4848 (N_4848,N_4701,N_4497);
or U4849 (N_4849,N_4714,N_4276);
xor U4850 (N_4850,N_4799,N_4105);
xnor U4851 (N_4851,N_4124,N_4723);
nor U4852 (N_4852,N_4502,N_4172);
nand U4853 (N_4853,N_4593,N_4100);
xnor U4854 (N_4854,N_4499,N_4786);
or U4855 (N_4855,N_4157,N_4366);
or U4856 (N_4856,N_4379,N_4261);
nor U4857 (N_4857,N_4783,N_4281);
xor U4858 (N_4858,N_4132,N_4648);
nand U4859 (N_4859,N_4050,N_4616);
and U4860 (N_4860,N_4653,N_4081);
nand U4861 (N_4861,N_4034,N_4195);
and U4862 (N_4862,N_4642,N_4666);
nand U4863 (N_4863,N_4269,N_4535);
or U4864 (N_4864,N_4312,N_4553);
nand U4865 (N_4865,N_4111,N_4519);
nand U4866 (N_4866,N_4255,N_4310);
and U4867 (N_4867,N_4663,N_4394);
nand U4868 (N_4868,N_4004,N_4167);
or U4869 (N_4869,N_4197,N_4360);
nand U4870 (N_4870,N_4715,N_4640);
nand U4871 (N_4871,N_4607,N_4003);
xor U4872 (N_4872,N_4726,N_4661);
and U4873 (N_4873,N_4230,N_4411);
or U4874 (N_4874,N_4139,N_4313);
nor U4875 (N_4875,N_4654,N_4057);
and U4876 (N_4876,N_4184,N_4622);
or U4877 (N_4877,N_4041,N_4389);
nand U4878 (N_4878,N_4481,N_4019);
nor U4879 (N_4879,N_4369,N_4007);
nor U4880 (N_4880,N_4231,N_4554);
nor U4881 (N_4881,N_4024,N_4750);
or U4882 (N_4882,N_4017,N_4305);
and U4883 (N_4883,N_4662,N_4270);
and U4884 (N_4884,N_4699,N_4777);
nor U4885 (N_4885,N_4603,N_4612);
nand U4886 (N_4886,N_4159,N_4724);
nor U4887 (N_4887,N_4566,N_4344);
or U4888 (N_4888,N_4678,N_4216);
and U4889 (N_4889,N_4247,N_4169);
nand U4890 (N_4890,N_4378,N_4706);
nor U4891 (N_4891,N_4153,N_4367);
xnor U4892 (N_4892,N_4785,N_4215);
or U4893 (N_4893,N_4442,N_4537);
xnor U4894 (N_4894,N_4323,N_4075);
nor U4895 (N_4895,N_4183,N_4513);
or U4896 (N_4896,N_4403,N_4225);
nor U4897 (N_4897,N_4235,N_4698);
or U4898 (N_4898,N_4737,N_4336);
nand U4899 (N_4899,N_4087,N_4505);
and U4900 (N_4900,N_4372,N_4459);
nor U4901 (N_4901,N_4646,N_4052);
nor U4902 (N_4902,N_4441,N_4580);
or U4903 (N_4903,N_4204,N_4088);
nand U4904 (N_4904,N_4126,N_4765);
nor U4905 (N_4905,N_4268,N_4322);
nor U4906 (N_4906,N_4080,N_4735);
or U4907 (N_4907,N_4177,N_4584);
or U4908 (N_4908,N_4078,N_4220);
xnor U4909 (N_4909,N_4239,N_4386);
nor U4910 (N_4910,N_4570,N_4536);
nor U4911 (N_4911,N_4747,N_4498);
xnor U4912 (N_4912,N_4115,N_4334);
nor U4913 (N_4913,N_4067,N_4355);
or U4914 (N_4914,N_4005,N_4198);
xnor U4915 (N_4915,N_4464,N_4438);
nand U4916 (N_4916,N_4410,N_4201);
nand U4917 (N_4917,N_4577,N_4285);
or U4918 (N_4918,N_4252,N_4134);
and U4919 (N_4919,N_4397,N_4018);
xnor U4920 (N_4920,N_4745,N_4094);
xnor U4921 (N_4921,N_4462,N_4401);
and U4922 (N_4922,N_4032,N_4483);
nand U4923 (N_4923,N_4154,N_4308);
nand U4924 (N_4924,N_4685,N_4544);
or U4925 (N_4925,N_4563,N_4364);
nand U4926 (N_4926,N_4277,N_4222);
nand U4927 (N_4927,N_4213,N_4766);
or U4928 (N_4928,N_4414,N_4404);
or U4929 (N_4929,N_4598,N_4302);
or U4930 (N_4930,N_4788,N_4053);
or U4931 (N_4931,N_4156,N_4099);
nand U4932 (N_4932,N_4258,N_4575);
and U4933 (N_4933,N_4145,N_4428);
or U4934 (N_4934,N_4092,N_4340);
xnor U4935 (N_4935,N_4348,N_4753);
nand U4936 (N_4936,N_4317,N_4510);
nand U4937 (N_4937,N_4793,N_4406);
or U4938 (N_4938,N_4259,N_4614);
and U4939 (N_4939,N_4203,N_4174);
nor U4940 (N_4940,N_4748,N_4494);
or U4941 (N_4941,N_4689,N_4085);
nand U4942 (N_4942,N_4096,N_4567);
or U4943 (N_4943,N_4486,N_4409);
or U4944 (N_4944,N_4795,N_4109);
nand U4945 (N_4945,N_4339,N_4547);
xor U4946 (N_4946,N_4545,N_4621);
or U4947 (N_4947,N_4071,N_4610);
xor U4948 (N_4948,N_4186,N_4733);
nor U4949 (N_4949,N_4396,N_4168);
or U4950 (N_4950,N_4415,N_4098);
nor U4951 (N_4951,N_4446,N_4083);
nor U4952 (N_4952,N_4688,N_4368);
or U4953 (N_4953,N_4370,N_4743);
nand U4954 (N_4954,N_4137,N_4295);
nand U4955 (N_4955,N_4026,N_4246);
and U4956 (N_4956,N_4338,N_4669);
and U4957 (N_4957,N_4709,N_4407);
and U4958 (N_4958,N_4552,N_4046);
xor U4959 (N_4959,N_4635,N_4636);
or U4960 (N_4960,N_4304,N_4187);
xnor U4961 (N_4961,N_4602,N_4644);
xnor U4962 (N_4962,N_4490,N_4558);
nand U4963 (N_4963,N_4556,N_4125);
nor U4964 (N_4964,N_4417,N_4694);
xor U4965 (N_4965,N_4233,N_4327);
and U4966 (N_4966,N_4790,N_4194);
xor U4967 (N_4967,N_4265,N_4645);
or U4968 (N_4968,N_4051,N_4144);
or U4969 (N_4969,N_4416,N_4728);
nand U4970 (N_4970,N_4597,N_4116);
nor U4971 (N_4971,N_4263,N_4541);
nand U4972 (N_4972,N_4683,N_4031);
nand U4973 (N_4973,N_4564,N_4345);
or U4974 (N_4974,N_4569,N_4444);
nand U4975 (N_4975,N_4756,N_4101);
or U4976 (N_4976,N_4509,N_4571);
or U4977 (N_4977,N_4329,N_4387);
nand U4978 (N_4978,N_4595,N_4084);
nand U4979 (N_4979,N_4725,N_4507);
or U4980 (N_4980,N_4696,N_4453);
xor U4981 (N_4981,N_4193,N_4228);
nor U4982 (N_4982,N_4559,N_4141);
or U4983 (N_4983,N_4792,N_4214);
nor U4984 (N_4984,N_4738,N_4609);
nor U4985 (N_4985,N_4136,N_4717);
or U4986 (N_4986,N_4478,N_4572);
nor U4987 (N_4987,N_4757,N_4672);
nor U4988 (N_4988,N_4097,N_4471);
or U4989 (N_4989,N_4008,N_4022);
or U4990 (N_4990,N_4010,N_4237);
nand U4991 (N_4991,N_4550,N_4710);
xor U4992 (N_4992,N_4165,N_4755);
and U4993 (N_4993,N_4079,N_4796);
nand U4994 (N_4994,N_4122,N_4301);
nand U4995 (N_4995,N_4207,N_4495);
nor U4996 (N_4996,N_4658,N_4266);
nand U4997 (N_4997,N_4767,N_4095);
nor U4998 (N_4998,N_4484,N_4180);
nor U4999 (N_4999,N_4659,N_4190);
or U5000 (N_5000,N_4226,N_4298);
xor U5001 (N_5001,N_4555,N_4307);
xnor U5002 (N_5002,N_4742,N_4690);
and U5003 (N_5003,N_4206,N_4399);
xnor U5004 (N_5004,N_4133,N_4530);
xnor U5005 (N_5005,N_4641,N_4290);
nand U5006 (N_5006,N_4349,N_4630);
nand U5007 (N_5007,N_4430,N_4435);
nand U5008 (N_5008,N_4129,N_4294);
nor U5009 (N_5009,N_4582,N_4288);
xnor U5010 (N_5010,N_4458,N_4039);
xor U5011 (N_5011,N_4063,N_4043);
xnor U5012 (N_5012,N_4380,N_4476);
and U5013 (N_5013,N_4526,N_4353);
xor U5014 (N_5014,N_4011,N_4146);
nand U5015 (N_5015,N_4160,N_4171);
nor U5016 (N_5016,N_4200,N_4532);
xor U5017 (N_5017,N_4751,N_4205);
xor U5018 (N_5018,N_4511,N_4245);
nand U5019 (N_5019,N_4676,N_4055);
and U5020 (N_5020,N_4373,N_4589);
or U5021 (N_5021,N_4351,N_4267);
or U5022 (N_5022,N_4749,N_4427);
nand U5023 (N_5023,N_4601,N_4271);
nor U5024 (N_5024,N_4529,N_4395);
or U5025 (N_5025,N_4721,N_4272);
and U5026 (N_5026,N_4371,N_4059);
xnor U5027 (N_5027,N_4346,N_4716);
xor U5028 (N_5028,N_4113,N_4482);
and U5029 (N_5029,N_4196,N_4287);
or U5030 (N_5030,N_4434,N_4289);
nor U5031 (N_5031,N_4606,N_4682);
nand U5032 (N_5032,N_4250,N_4551);
and U5033 (N_5033,N_4639,N_4209);
xor U5034 (N_5034,N_4769,N_4363);
nor U5035 (N_5035,N_4771,N_4508);
nand U5036 (N_5036,N_4776,N_4107);
nor U5037 (N_5037,N_4221,N_4588);
xnor U5038 (N_5038,N_4631,N_4229);
xor U5039 (N_5039,N_4091,N_4332);
or U5040 (N_5040,N_4450,N_4684);
or U5041 (N_5041,N_4712,N_4347);
or U5042 (N_5042,N_4188,N_4383);
xor U5043 (N_5043,N_4705,N_4741);
nand U5044 (N_5044,N_4489,N_4686);
xnor U5045 (N_5045,N_4292,N_4493);
or U5046 (N_5046,N_4320,N_4506);
or U5047 (N_5047,N_4054,N_4652);
and U5048 (N_5048,N_4585,N_4150);
or U5049 (N_5049,N_4224,N_4121);
or U5050 (N_5050,N_4590,N_4576);
nor U5051 (N_5051,N_4335,N_4423);
xor U5052 (N_5052,N_4759,N_4744);
nand U5053 (N_5053,N_4711,N_4102);
xor U5054 (N_5054,N_4070,N_4693);
nand U5055 (N_5055,N_4049,N_4176);
nor U5056 (N_5056,N_4538,N_4628);
and U5057 (N_5057,N_4119,N_4178);
nand U5058 (N_5058,N_4181,N_4219);
nand U5059 (N_5059,N_4212,N_4179);
nand U5060 (N_5060,N_4056,N_4135);
nand U5061 (N_5061,N_4704,N_4779);
and U5062 (N_5062,N_4605,N_4736);
and U5063 (N_5063,N_4152,N_4223);
nor U5064 (N_5064,N_4429,N_4477);
or U5065 (N_5065,N_4425,N_4400);
or U5066 (N_5066,N_4740,N_4539);
nand U5067 (N_5067,N_4557,N_4643);
xnor U5068 (N_5068,N_4048,N_4020);
and U5069 (N_5069,N_4293,N_4012);
and U5070 (N_5070,N_4789,N_4664);
and U5071 (N_5071,N_4463,N_4657);
or U5072 (N_5072,N_4093,N_4419);
nor U5073 (N_5073,N_4273,N_4148);
xnor U5074 (N_5074,N_4045,N_4611);
xnor U5075 (N_5075,N_4465,N_4426);
xor U5076 (N_5076,N_4077,N_4700);
nand U5077 (N_5077,N_4791,N_4384);
nand U5078 (N_5078,N_4501,N_4437);
nand U5079 (N_5079,N_4412,N_4586);
and U5080 (N_5080,N_4433,N_4548);
xnor U5081 (N_5081,N_4208,N_4166);
nor U5082 (N_5082,N_4164,N_4066);
and U5083 (N_5083,N_4354,N_4562);
or U5084 (N_5084,N_4254,N_4234);
nor U5085 (N_5085,N_4278,N_4330);
and U5086 (N_5086,N_4210,N_4479);
and U5087 (N_5087,N_4637,N_4044);
and U5088 (N_5088,N_4028,N_4533);
xnor U5089 (N_5089,N_4182,N_4731);
and U5090 (N_5090,N_4117,N_4065);
xor U5091 (N_5091,N_4001,N_4306);
xnor U5092 (N_5092,N_4487,N_4634);
nand U5093 (N_5093,N_4485,N_4326);
nand U5094 (N_5094,N_4798,N_4524);
and U5095 (N_5095,N_4325,N_4517);
nor U5096 (N_5096,N_4408,N_4448);
nand U5097 (N_5097,N_4284,N_4762);
nor U5098 (N_5098,N_4540,N_4734);
nor U5099 (N_5099,N_4774,N_4418);
and U5100 (N_5100,N_4467,N_4282);
nor U5101 (N_5101,N_4042,N_4752);
or U5102 (N_5102,N_4623,N_4170);
nor U5103 (N_5103,N_4673,N_4500);
and U5104 (N_5104,N_4191,N_4445);
nor U5105 (N_5105,N_4527,N_4778);
nor U5106 (N_5106,N_4120,N_4062);
nand U5107 (N_5107,N_4703,N_4275);
xnor U5108 (N_5108,N_4561,N_4660);
xor U5109 (N_5109,N_4787,N_4138);
nor U5110 (N_5110,N_4746,N_4469);
nand U5111 (N_5111,N_4472,N_4488);
nand U5112 (N_5112,N_4280,N_4702);
and U5113 (N_5113,N_4587,N_4618);
nand U5114 (N_5114,N_4390,N_4432);
nand U5115 (N_5115,N_4739,N_4036);
or U5116 (N_5116,N_4770,N_4473);
xnor U5117 (N_5117,N_4000,N_4175);
nor U5118 (N_5118,N_4474,N_4238);
or U5119 (N_5119,N_4015,N_4424);
and U5120 (N_5120,N_4232,N_4377);
and U5121 (N_5121,N_4274,N_4104);
nand U5122 (N_5122,N_4002,N_4405);
nand U5123 (N_5123,N_4006,N_4376);
and U5124 (N_5124,N_4331,N_4118);
nor U5125 (N_5125,N_4244,N_4392);
nand U5126 (N_5126,N_4035,N_4029);
nand U5127 (N_5127,N_4675,N_4681);
nand U5128 (N_5128,N_4784,N_4256);
nor U5129 (N_5129,N_4037,N_4491);
nor U5130 (N_5130,N_4249,N_4754);
nor U5131 (N_5131,N_4218,N_4106);
nor U5132 (N_5132,N_4362,N_4279);
nand U5133 (N_5133,N_4516,N_4594);
nor U5134 (N_5134,N_4656,N_4599);
nor U5135 (N_5135,N_4525,N_4023);
or U5136 (N_5136,N_4633,N_4568);
and U5137 (N_5137,N_4592,N_4546);
and U5138 (N_5138,N_4651,N_4460);
nand U5139 (N_5139,N_4522,N_4227);
xnor U5140 (N_5140,N_4720,N_4162);
nand U5141 (N_5141,N_4240,N_4758);
xnor U5142 (N_5142,N_4443,N_4518);
nor U5143 (N_5143,N_4679,N_4665);
nand U5144 (N_5144,N_4670,N_4775);
or U5145 (N_5145,N_4760,N_4707);
nand U5146 (N_5146,N_4253,N_4189);
nand U5147 (N_5147,N_4655,N_4543);
xnor U5148 (N_5148,N_4147,N_4626);
or U5149 (N_5149,N_4727,N_4365);
or U5150 (N_5150,N_4413,N_4033);
nor U5151 (N_5151,N_4192,N_4242);
and U5152 (N_5152,N_4385,N_4613);
xnor U5153 (N_5153,N_4515,N_4534);
and U5154 (N_5154,N_4581,N_4297);
nor U5155 (N_5155,N_4151,N_4583);
or U5156 (N_5156,N_4671,N_4251);
and U5157 (N_5157,N_4243,N_4457);
nor U5158 (N_5158,N_4466,N_4236);
nand U5159 (N_5159,N_4324,N_4199);
xnor U5160 (N_5160,N_4161,N_4514);
or U5161 (N_5161,N_4531,N_4311);
or U5162 (N_5162,N_4797,N_4074);
nor U5163 (N_5163,N_4040,N_4103);
xnor U5164 (N_5164,N_4600,N_4319);
nand U5165 (N_5165,N_4391,N_4647);
nor U5166 (N_5166,N_4713,N_4523);
nand U5167 (N_5167,N_4455,N_4470);
and U5168 (N_5168,N_4638,N_4076);
or U5169 (N_5169,N_4374,N_4356);
or U5170 (N_5170,N_4296,N_4697);
or U5171 (N_5171,N_4764,N_4333);
nand U5172 (N_5172,N_4451,N_4064);
and U5173 (N_5173,N_4341,N_4608);
or U5174 (N_5174,N_4114,N_4014);
and U5175 (N_5175,N_4772,N_4140);
or U5176 (N_5176,N_4016,N_4112);
nand U5177 (N_5177,N_4300,N_4591);
xor U5178 (N_5178,N_4264,N_4528);
and U5179 (N_5179,N_4579,N_4542);
nand U5180 (N_5180,N_4549,N_4692);
nand U5181 (N_5181,N_4763,N_4082);
and U5182 (N_5182,N_4241,N_4318);
or U5183 (N_5183,N_4520,N_4286);
or U5184 (N_5184,N_4343,N_4163);
or U5185 (N_5185,N_4291,N_4173);
or U5186 (N_5186,N_4337,N_4303);
nor U5187 (N_5187,N_4732,N_4342);
or U5188 (N_5188,N_4069,N_4110);
nor U5189 (N_5189,N_4299,N_4108);
nor U5190 (N_5190,N_4468,N_4127);
and U5191 (N_5191,N_4315,N_4202);
or U5192 (N_5192,N_4578,N_4629);
nor U5193 (N_5193,N_4038,N_4262);
xor U5194 (N_5194,N_4521,N_4185);
and U5195 (N_5195,N_4321,N_4565);
or U5196 (N_5196,N_4452,N_4461);
and U5197 (N_5197,N_4617,N_4388);
and U5198 (N_5198,N_4143,N_4257);
or U5199 (N_5199,N_4780,N_4620);
nor U5200 (N_5200,N_4377,N_4733);
nor U5201 (N_5201,N_4114,N_4348);
nand U5202 (N_5202,N_4433,N_4358);
and U5203 (N_5203,N_4185,N_4600);
xnor U5204 (N_5204,N_4452,N_4022);
and U5205 (N_5205,N_4356,N_4265);
and U5206 (N_5206,N_4014,N_4646);
or U5207 (N_5207,N_4666,N_4286);
or U5208 (N_5208,N_4190,N_4424);
or U5209 (N_5209,N_4210,N_4038);
or U5210 (N_5210,N_4570,N_4658);
nand U5211 (N_5211,N_4281,N_4660);
and U5212 (N_5212,N_4297,N_4179);
nor U5213 (N_5213,N_4654,N_4510);
and U5214 (N_5214,N_4661,N_4610);
and U5215 (N_5215,N_4255,N_4373);
nor U5216 (N_5216,N_4020,N_4539);
or U5217 (N_5217,N_4076,N_4202);
nor U5218 (N_5218,N_4468,N_4029);
or U5219 (N_5219,N_4370,N_4685);
nor U5220 (N_5220,N_4372,N_4356);
and U5221 (N_5221,N_4222,N_4711);
or U5222 (N_5222,N_4220,N_4623);
nor U5223 (N_5223,N_4286,N_4532);
and U5224 (N_5224,N_4341,N_4122);
nor U5225 (N_5225,N_4267,N_4261);
nand U5226 (N_5226,N_4349,N_4799);
and U5227 (N_5227,N_4105,N_4543);
nor U5228 (N_5228,N_4781,N_4482);
or U5229 (N_5229,N_4050,N_4434);
xnor U5230 (N_5230,N_4484,N_4490);
nor U5231 (N_5231,N_4588,N_4554);
xor U5232 (N_5232,N_4422,N_4327);
nor U5233 (N_5233,N_4650,N_4176);
nand U5234 (N_5234,N_4225,N_4667);
and U5235 (N_5235,N_4128,N_4189);
xnor U5236 (N_5236,N_4105,N_4690);
nor U5237 (N_5237,N_4642,N_4362);
nand U5238 (N_5238,N_4180,N_4674);
and U5239 (N_5239,N_4294,N_4669);
and U5240 (N_5240,N_4299,N_4030);
nor U5241 (N_5241,N_4701,N_4428);
or U5242 (N_5242,N_4642,N_4439);
or U5243 (N_5243,N_4035,N_4349);
or U5244 (N_5244,N_4147,N_4470);
nor U5245 (N_5245,N_4390,N_4761);
or U5246 (N_5246,N_4474,N_4480);
nor U5247 (N_5247,N_4492,N_4407);
xor U5248 (N_5248,N_4426,N_4142);
nor U5249 (N_5249,N_4269,N_4096);
xnor U5250 (N_5250,N_4460,N_4562);
or U5251 (N_5251,N_4410,N_4766);
nor U5252 (N_5252,N_4752,N_4513);
nand U5253 (N_5253,N_4426,N_4329);
nand U5254 (N_5254,N_4568,N_4593);
nand U5255 (N_5255,N_4726,N_4434);
and U5256 (N_5256,N_4473,N_4724);
nor U5257 (N_5257,N_4381,N_4257);
xor U5258 (N_5258,N_4351,N_4104);
and U5259 (N_5259,N_4202,N_4207);
and U5260 (N_5260,N_4347,N_4483);
nand U5261 (N_5261,N_4005,N_4264);
and U5262 (N_5262,N_4386,N_4201);
nor U5263 (N_5263,N_4292,N_4549);
or U5264 (N_5264,N_4079,N_4239);
or U5265 (N_5265,N_4617,N_4467);
and U5266 (N_5266,N_4198,N_4062);
xor U5267 (N_5267,N_4381,N_4129);
or U5268 (N_5268,N_4634,N_4410);
nor U5269 (N_5269,N_4759,N_4221);
nand U5270 (N_5270,N_4098,N_4665);
and U5271 (N_5271,N_4541,N_4756);
and U5272 (N_5272,N_4252,N_4739);
nor U5273 (N_5273,N_4667,N_4370);
or U5274 (N_5274,N_4329,N_4635);
or U5275 (N_5275,N_4342,N_4691);
nand U5276 (N_5276,N_4721,N_4638);
or U5277 (N_5277,N_4372,N_4450);
nand U5278 (N_5278,N_4150,N_4554);
or U5279 (N_5279,N_4592,N_4130);
nor U5280 (N_5280,N_4304,N_4616);
or U5281 (N_5281,N_4389,N_4613);
nand U5282 (N_5282,N_4191,N_4420);
nor U5283 (N_5283,N_4688,N_4789);
nand U5284 (N_5284,N_4408,N_4016);
xor U5285 (N_5285,N_4310,N_4793);
nor U5286 (N_5286,N_4094,N_4535);
xnor U5287 (N_5287,N_4669,N_4036);
or U5288 (N_5288,N_4007,N_4376);
nor U5289 (N_5289,N_4097,N_4069);
xor U5290 (N_5290,N_4678,N_4599);
or U5291 (N_5291,N_4316,N_4777);
and U5292 (N_5292,N_4339,N_4548);
nand U5293 (N_5293,N_4449,N_4580);
xor U5294 (N_5294,N_4698,N_4709);
nor U5295 (N_5295,N_4575,N_4198);
xnor U5296 (N_5296,N_4015,N_4614);
or U5297 (N_5297,N_4755,N_4203);
and U5298 (N_5298,N_4743,N_4778);
nor U5299 (N_5299,N_4299,N_4775);
or U5300 (N_5300,N_4460,N_4279);
nand U5301 (N_5301,N_4659,N_4048);
and U5302 (N_5302,N_4781,N_4149);
nand U5303 (N_5303,N_4451,N_4766);
or U5304 (N_5304,N_4726,N_4540);
nor U5305 (N_5305,N_4603,N_4604);
and U5306 (N_5306,N_4150,N_4413);
nor U5307 (N_5307,N_4604,N_4389);
xor U5308 (N_5308,N_4774,N_4056);
nand U5309 (N_5309,N_4730,N_4501);
or U5310 (N_5310,N_4498,N_4682);
nand U5311 (N_5311,N_4002,N_4384);
nor U5312 (N_5312,N_4204,N_4442);
nand U5313 (N_5313,N_4371,N_4623);
nor U5314 (N_5314,N_4686,N_4302);
or U5315 (N_5315,N_4505,N_4048);
or U5316 (N_5316,N_4130,N_4673);
xor U5317 (N_5317,N_4269,N_4473);
nor U5318 (N_5318,N_4418,N_4684);
nand U5319 (N_5319,N_4008,N_4397);
xor U5320 (N_5320,N_4251,N_4191);
xor U5321 (N_5321,N_4496,N_4440);
xor U5322 (N_5322,N_4448,N_4343);
nand U5323 (N_5323,N_4773,N_4060);
or U5324 (N_5324,N_4706,N_4099);
nand U5325 (N_5325,N_4097,N_4578);
or U5326 (N_5326,N_4543,N_4600);
and U5327 (N_5327,N_4715,N_4534);
xnor U5328 (N_5328,N_4760,N_4202);
nand U5329 (N_5329,N_4275,N_4230);
xor U5330 (N_5330,N_4678,N_4795);
xor U5331 (N_5331,N_4430,N_4773);
nand U5332 (N_5332,N_4127,N_4750);
xor U5333 (N_5333,N_4150,N_4632);
or U5334 (N_5334,N_4683,N_4127);
and U5335 (N_5335,N_4082,N_4109);
xor U5336 (N_5336,N_4326,N_4447);
nand U5337 (N_5337,N_4369,N_4604);
xnor U5338 (N_5338,N_4309,N_4022);
nand U5339 (N_5339,N_4449,N_4041);
and U5340 (N_5340,N_4044,N_4625);
and U5341 (N_5341,N_4176,N_4336);
or U5342 (N_5342,N_4068,N_4277);
and U5343 (N_5343,N_4580,N_4664);
nand U5344 (N_5344,N_4273,N_4655);
nor U5345 (N_5345,N_4136,N_4567);
and U5346 (N_5346,N_4775,N_4681);
nor U5347 (N_5347,N_4048,N_4451);
xor U5348 (N_5348,N_4085,N_4653);
xor U5349 (N_5349,N_4464,N_4133);
and U5350 (N_5350,N_4724,N_4503);
xor U5351 (N_5351,N_4499,N_4648);
and U5352 (N_5352,N_4218,N_4369);
or U5353 (N_5353,N_4310,N_4130);
and U5354 (N_5354,N_4452,N_4381);
nor U5355 (N_5355,N_4705,N_4611);
and U5356 (N_5356,N_4479,N_4503);
and U5357 (N_5357,N_4328,N_4772);
nand U5358 (N_5358,N_4312,N_4575);
xnor U5359 (N_5359,N_4191,N_4048);
xnor U5360 (N_5360,N_4078,N_4671);
nand U5361 (N_5361,N_4080,N_4542);
nand U5362 (N_5362,N_4253,N_4217);
and U5363 (N_5363,N_4281,N_4579);
nand U5364 (N_5364,N_4493,N_4564);
or U5365 (N_5365,N_4653,N_4203);
or U5366 (N_5366,N_4677,N_4792);
nand U5367 (N_5367,N_4604,N_4329);
and U5368 (N_5368,N_4671,N_4783);
nand U5369 (N_5369,N_4701,N_4732);
or U5370 (N_5370,N_4176,N_4474);
and U5371 (N_5371,N_4172,N_4651);
and U5372 (N_5372,N_4612,N_4796);
xor U5373 (N_5373,N_4515,N_4386);
xor U5374 (N_5374,N_4718,N_4525);
nand U5375 (N_5375,N_4111,N_4040);
and U5376 (N_5376,N_4793,N_4754);
nand U5377 (N_5377,N_4791,N_4502);
or U5378 (N_5378,N_4319,N_4052);
and U5379 (N_5379,N_4535,N_4448);
xnor U5380 (N_5380,N_4084,N_4359);
nor U5381 (N_5381,N_4584,N_4273);
or U5382 (N_5382,N_4027,N_4010);
and U5383 (N_5383,N_4277,N_4696);
xor U5384 (N_5384,N_4274,N_4003);
xnor U5385 (N_5385,N_4181,N_4669);
or U5386 (N_5386,N_4675,N_4190);
nand U5387 (N_5387,N_4115,N_4314);
nor U5388 (N_5388,N_4711,N_4034);
and U5389 (N_5389,N_4140,N_4047);
nand U5390 (N_5390,N_4320,N_4186);
nor U5391 (N_5391,N_4046,N_4699);
and U5392 (N_5392,N_4096,N_4235);
xor U5393 (N_5393,N_4537,N_4205);
xor U5394 (N_5394,N_4306,N_4497);
or U5395 (N_5395,N_4441,N_4445);
and U5396 (N_5396,N_4765,N_4045);
or U5397 (N_5397,N_4723,N_4245);
nor U5398 (N_5398,N_4673,N_4699);
xnor U5399 (N_5399,N_4448,N_4120);
or U5400 (N_5400,N_4540,N_4003);
xor U5401 (N_5401,N_4074,N_4693);
nand U5402 (N_5402,N_4101,N_4086);
nor U5403 (N_5403,N_4736,N_4307);
and U5404 (N_5404,N_4648,N_4382);
and U5405 (N_5405,N_4327,N_4710);
nor U5406 (N_5406,N_4588,N_4771);
nor U5407 (N_5407,N_4137,N_4451);
nand U5408 (N_5408,N_4709,N_4271);
nor U5409 (N_5409,N_4583,N_4621);
xor U5410 (N_5410,N_4513,N_4382);
nor U5411 (N_5411,N_4758,N_4195);
nor U5412 (N_5412,N_4656,N_4593);
nor U5413 (N_5413,N_4309,N_4406);
xnor U5414 (N_5414,N_4230,N_4055);
or U5415 (N_5415,N_4694,N_4347);
xnor U5416 (N_5416,N_4384,N_4313);
nand U5417 (N_5417,N_4136,N_4100);
xnor U5418 (N_5418,N_4304,N_4429);
or U5419 (N_5419,N_4291,N_4743);
or U5420 (N_5420,N_4370,N_4227);
xnor U5421 (N_5421,N_4169,N_4071);
nand U5422 (N_5422,N_4548,N_4785);
nor U5423 (N_5423,N_4604,N_4065);
and U5424 (N_5424,N_4433,N_4460);
nor U5425 (N_5425,N_4284,N_4631);
or U5426 (N_5426,N_4556,N_4495);
or U5427 (N_5427,N_4350,N_4218);
and U5428 (N_5428,N_4428,N_4218);
nand U5429 (N_5429,N_4040,N_4018);
nand U5430 (N_5430,N_4037,N_4338);
nor U5431 (N_5431,N_4168,N_4725);
nand U5432 (N_5432,N_4035,N_4667);
nand U5433 (N_5433,N_4518,N_4625);
nor U5434 (N_5434,N_4290,N_4541);
nor U5435 (N_5435,N_4085,N_4321);
and U5436 (N_5436,N_4000,N_4078);
xor U5437 (N_5437,N_4756,N_4399);
xnor U5438 (N_5438,N_4064,N_4370);
and U5439 (N_5439,N_4278,N_4186);
xor U5440 (N_5440,N_4407,N_4493);
nor U5441 (N_5441,N_4301,N_4583);
nor U5442 (N_5442,N_4785,N_4515);
nor U5443 (N_5443,N_4372,N_4040);
nor U5444 (N_5444,N_4297,N_4336);
xor U5445 (N_5445,N_4116,N_4776);
or U5446 (N_5446,N_4574,N_4398);
nand U5447 (N_5447,N_4657,N_4507);
nand U5448 (N_5448,N_4409,N_4043);
nand U5449 (N_5449,N_4581,N_4325);
nand U5450 (N_5450,N_4243,N_4472);
or U5451 (N_5451,N_4319,N_4607);
nand U5452 (N_5452,N_4078,N_4604);
or U5453 (N_5453,N_4458,N_4426);
xnor U5454 (N_5454,N_4739,N_4576);
and U5455 (N_5455,N_4698,N_4359);
nor U5456 (N_5456,N_4532,N_4158);
nor U5457 (N_5457,N_4064,N_4028);
nor U5458 (N_5458,N_4396,N_4355);
and U5459 (N_5459,N_4205,N_4283);
nor U5460 (N_5460,N_4039,N_4792);
and U5461 (N_5461,N_4509,N_4155);
nand U5462 (N_5462,N_4370,N_4421);
nand U5463 (N_5463,N_4174,N_4237);
or U5464 (N_5464,N_4188,N_4099);
or U5465 (N_5465,N_4024,N_4799);
nand U5466 (N_5466,N_4459,N_4013);
and U5467 (N_5467,N_4297,N_4449);
nand U5468 (N_5468,N_4763,N_4354);
or U5469 (N_5469,N_4024,N_4585);
and U5470 (N_5470,N_4750,N_4484);
nand U5471 (N_5471,N_4562,N_4557);
or U5472 (N_5472,N_4487,N_4762);
and U5473 (N_5473,N_4575,N_4713);
and U5474 (N_5474,N_4611,N_4590);
nand U5475 (N_5475,N_4080,N_4570);
nor U5476 (N_5476,N_4270,N_4426);
nand U5477 (N_5477,N_4774,N_4039);
nand U5478 (N_5478,N_4454,N_4410);
or U5479 (N_5479,N_4681,N_4187);
xnor U5480 (N_5480,N_4630,N_4367);
nand U5481 (N_5481,N_4176,N_4271);
nand U5482 (N_5482,N_4697,N_4528);
nor U5483 (N_5483,N_4562,N_4059);
nor U5484 (N_5484,N_4014,N_4071);
xnor U5485 (N_5485,N_4598,N_4699);
xor U5486 (N_5486,N_4282,N_4716);
nand U5487 (N_5487,N_4509,N_4181);
or U5488 (N_5488,N_4506,N_4416);
or U5489 (N_5489,N_4521,N_4046);
and U5490 (N_5490,N_4213,N_4496);
and U5491 (N_5491,N_4145,N_4706);
and U5492 (N_5492,N_4797,N_4362);
or U5493 (N_5493,N_4507,N_4155);
xor U5494 (N_5494,N_4099,N_4006);
xnor U5495 (N_5495,N_4051,N_4262);
or U5496 (N_5496,N_4265,N_4623);
or U5497 (N_5497,N_4004,N_4744);
or U5498 (N_5498,N_4028,N_4282);
nand U5499 (N_5499,N_4045,N_4269);
and U5500 (N_5500,N_4793,N_4607);
and U5501 (N_5501,N_4024,N_4607);
nand U5502 (N_5502,N_4566,N_4696);
nor U5503 (N_5503,N_4070,N_4704);
nor U5504 (N_5504,N_4033,N_4502);
xor U5505 (N_5505,N_4085,N_4197);
xor U5506 (N_5506,N_4398,N_4779);
or U5507 (N_5507,N_4583,N_4121);
or U5508 (N_5508,N_4700,N_4474);
or U5509 (N_5509,N_4188,N_4196);
nor U5510 (N_5510,N_4001,N_4555);
nor U5511 (N_5511,N_4519,N_4771);
nand U5512 (N_5512,N_4134,N_4472);
xor U5513 (N_5513,N_4500,N_4418);
or U5514 (N_5514,N_4235,N_4213);
or U5515 (N_5515,N_4157,N_4535);
xnor U5516 (N_5516,N_4768,N_4656);
xor U5517 (N_5517,N_4357,N_4012);
xor U5518 (N_5518,N_4359,N_4053);
or U5519 (N_5519,N_4562,N_4086);
nor U5520 (N_5520,N_4683,N_4611);
nand U5521 (N_5521,N_4582,N_4157);
and U5522 (N_5522,N_4200,N_4061);
xor U5523 (N_5523,N_4749,N_4285);
and U5524 (N_5524,N_4038,N_4551);
nor U5525 (N_5525,N_4276,N_4205);
nor U5526 (N_5526,N_4027,N_4424);
nor U5527 (N_5527,N_4739,N_4287);
nor U5528 (N_5528,N_4115,N_4368);
and U5529 (N_5529,N_4495,N_4063);
xor U5530 (N_5530,N_4076,N_4328);
nand U5531 (N_5531,N_4555,N_4178);
and U5532 (N_5532,N_4613,N_4465);
nor U5533 (N_5533,N_4349,N_4369);
nor U5534 (N_5534,N_4505,N_4280);
xor U5535 (N_5535,N_4026,N_4675);
nor U5536 (N_5536,N_4685,N_4614);
and U5537 (N_5537,N_4766,N_4096);
nor U5538 (N_5538,N_4307,N_4007);
xnor U5539 (N_5539,N_4760,N_4347);
nand U5540 (N_5540,N_4611,N_4262);
nor U5541 (N_5541,N_4795,N_4461);
or U5542 (N_5542,N_4418,N_4654);
and U5543 (N_5543,N_4283,N_4471);
nand U5544 (N_5544,N_4775,N_4018);
xor U5545 (N_5545,N_4020,N_4426);
nand U5546 (N_5546,N_4638,N_4336);
nand U5547 (N_5547,N_4415,N_4251);
and U5548 (N_5548,N_4299,N_4448);
xnor U5549 (N_5549,N_4471,N_4642);
xor U5550 (N_5550,N_4298,N_4290);
and U5551 (N_5551,N_4525,N_4395);
and U5552 (N_5552,N_4444,N_4184);
and U5553 (N_5553,N_4575,N_4438);
xnor U5554 (N_5554,N_4441,N_4493);
nand U5555 (N_5555,N_4206,N_4572);
xor U5556 (N_5556,N_4562,N_4318);
nor U5557 (N_5557,N_4185,N_4622);
and U5558 (N_5558,N_4529,N_4103);
nand U5559 (N_5559,N_4459,N_4427);
nor U5560 (N_5560,N_4323,N_4288);
and U5561 (N_5561,N_4644,N_4789);
and U5562 (N_5562,N_4696,N_4493);
nor U5563 (N_5563,N_4463,N_4205);
xor U5564 (N_5564,N_4039,N_4693);
nor U5565 (N_5565,N_4693,N_4772);
and U5566 (N_5566,N_4193,N_4387);
or U5567 (N_5567,N_4587,N_4271);
and U5568 (N_5568,N_4573,N_4359);
and U5569 (N_5569,N_4291,N_4517);
xnor U5570 (N_5570,N_4388,N_4253);
nand U5571 (N_5571,N_4353,N_4485);
xnor U5572 (N_5572,N_4695,N_4342);
or U5573 (N_5573,N_4301,N_4400);
or U5574 (N_5574,N_4345,N_4089);
and U5575 (N_5575,N_4640,N_4632);
nand U5576 (N_5576,N_4385,N_4458);
xor U5577 (N_5577,N_4587,N_4288);
nand U5578 (N_5578,N_4000,N_4469);
or U5579 (N_5579,N_4596,N_4312);
nor U5580 (N_5580,N_4794,N_4552);
or U5581 (N_5581,N_4531,N_4597);
or U5582 (N_5582,N_4614,N_4424);
xnor U5583 (N_5583,N_4556,N_4680);
nor U5584 (N_5584,N_4469,N_4722);
or U5585 (N_5585,N_4543,N_4476);
or U5586 (N_5586,N_4414,N_4499);
xnor U5587 (N_5587,N_4409,N_4673);
nor U5588 (N_5588,N_4173,N_4193);
or U5589 (N_5589,N_4708,N_4459);
and U5590 (N_5590,N_4536,N_4534);
nor U5591 (N_5591,N_4378,N_4024);
and U5592 (N_5592,N_4332,N_4650);
xor U5593 (N_5593,N_4587,N_4674);
and U5594 (N_5594,N_4321,N_4793);
nand U5595 (N_5595,N_4543,N_4205);
nand U5596 (N_5596,N_4106,N_4189);
nand U5597 (N_5597,N_4428,N_4227);
or U5598 (N_5598,N_4000,N_4109);
or U5599 (N_5599,N_4552,N_4619);
nand U5600 (N_5600,N_5493,N_5498);
xnor U5601 (N_5601,N_5518,N_4900);
xnor U5602 (N_5602,N_4837,N_5239);
nand U5603 (N_5603,N_5220,N_5261);
nor U5604 (N_5604,N_5533,N_4915);
xor U5605 (N_5605,N_4805,N_5043);
xnor U5606 (N_5606,N_5328,N_5171);
nor U5607 (N_5607,N_5262,N_5151);
xnor U5608 (N_5608,N_5044,N_5318);
and U5609 (N_5609,N_5197,N_5434);
nand U5610 (N_5610,N_5460,N_4980);
nand U5611 (N_5611,N_4959,N_5126);
or U5612 (N_5612,N_5010,N_5119);
and U5613 (N_5613,N_5167,N_5224);
nor U5614 (N_5614,N_5316,N_5065);
or U5615 (N_5615,N_4840,N_5441);
nor U5616 (N_5616,N_5557,N_5101);
and U5617 (N_5617,N_5323,N_5428);
nand U5618 (N_5618,N_5061,N_5464);
xor U5619 (N_5619,N_4942,N_5025);
and U5620 (N_5620,N_5280,N_5144);
nand U5621 (N_5621,N_4993,N_4896);
nor U5622 (N_5622,N_5391,N_5185);
nor U5623 (N_5623,N_5283,N_4892);
nand U5624 (N_5624,N_5034,N_5582);
nor U5625 (N_5625,N_4812,N_4862);
nor U5626 (N_5626,N_5045,N_5544);
or U5627 (N_5627,N_5535,N_5115);
xor U5628 (N_5628,N_4893,N_4841);
xor U5629 (N_5629,N_4887,N_5108);
nor U5630 (N_5630,N_4803,N_5068);
nor U5631 (N_5631,N_5430,N_4952);
and U5632 (N_5632,N_5335,N_5306);
nand U5633 (N_5633,N_4801,N_4999);
or U5634 (N_5634,N_5103,N_5522);
and U5635 (N_5635,N_4804,N_5500);
xnor U5636 (N_5636,N_4859,N_5507);
xor U5637 (N_5637,N_5122,N_5146);
xor U5638 (N_5638,N_5514,N_4904);
or U5639 (N_5639,N_5424,N_4964);
or U5640 (N_5640,N_5150,N_5540);
nor U5641 (N_5641,N_5375,N_5593);
or U5642 (N_5642,N_5282,N_4890);
nand U5643 (N_5643,N_5267,N_5290);
nand U5644 (N_5644,N_4869,N_5003);
or U5645 (N_5645,N_5259,N_5455);
nor U5646 (N_5646,N_5551,N_5016);
xnor U5647 (N_5647,N_5104,N_5447);
and U5648 (N_5648,N_4923,N_5134);
nand U5649 (N_5649,N_5199,N_4830);
and U5650 (N_5650,N_5212,N_5577);
or U5651 (N_5651,N_5338,N_5058);
nor U5652 (N_5652,N_5450,N_5260);
nand U5653 (N_5653,N_4948,N_4907);
nand U5654 (N_5654,N_4976,N_4932);
xnor U5655 (N_5655,N_5344,N_5189);
or U5656 (N_5656,N_5164,N_5550);
xor U5657 (N_5657,N_4858,N_5091);
nor U5658 (N_5658,N_5399,N_5117);
or U5659 (N_5659,N_5148,N_5305);
or U5660 (N_5660,N_4977,N_5321);
xor U5661 (N_5661,N_5573,N_5243);
nand U5662 (N_5662,N_5439,N_5071);
nand U5663 (N_5663,N_5308,N_5476);
nor U5664 (N_5664,N_5165,N_5405);
or U5665 (N_5665,N_5511,N_5599);
xnor U5666 (N_5666,N_4941,N_5192);
or U5667 (N_5667,N_5254,N_5423);
and U5668 (N_5668,N_4916,N_5039);
nand U5669 (N_5669,N_5408,N_5118);
and U5670 (N_5670,N_4960,N_5594);
or U5671 (N_5671,N_4950,N_5247);
nand U5672 (N_5672,N_5370,N_5504);
and U5673 (N_5673,N_5334,N_5386);
or U5674 (N_5674,N_5143,N_5555);
xnor U5675 (N_5675,N_4845,N_5092);
and U5676 (N_5676,N_5495,N_4940);
xor U5677 (N_5677,N_5549,N_5036);
nor U5678 (N_5678,N_4894,N_5017);
and U5679 (N_5679,N_4963,N_5079);
nor U5680 (N_5680,N_4835,N_5240);
or U5681 (N_5681,N_5309,N_5049);
nand U5682 (N_5682,N_5516,N_4946);
nand U5683 (N_5683,N_5138,N_5057);
and U5684 (N_5684,N_5166,N_5411);
and U5685 (N_5685,N_4990,N_5054);
nor U5686 (N_5686,N_5575,N_5461);
and U5687 (N_5687,N_5481,N_4899);
or U5688 (N_5688,N_4992,N_5128);
nor U5689 (N_5689,N_5011,N_5510);
xor U5690 (N_5690,N_5513,N_5395);
xor U5691 (N_5691,N_4895,N_5085);
xnor U5692 (N_5692,N_5176,N_5287);
nand U5693 (N_5693,N_5569,N_5404);
or U5694 (N_5694,N_5041,N_5178);
and U5695 (N_5695,N_4975,N_5113);
nand U5696 (N_5696,N_5515,N_5018);
nor U5697 (N_5697,N_5420,N_5517);
or U5698 (N_5698,N_5040,N_5547);
xnor U5699 (N_5699,N_5250,N_5022);
xor U5700 (N_5700,N_4868,N_5561);
xor U5701 (N_5701,N_4857,N_4860);
or U5702 (N_5702,N_5362,N_4938);
and U5703 (N_5703,N_5466,N_5401);
xnor U5704 (N_5704,N_5210,N_5278);
or U5705 (N_5705,N_5374,N_5028);
nand U5706 (N_5706,N_5312,N_4842);
or U5707 (N_5707,N_5292,N_5353);
nor U5708 (N_5708,N_4861,N_4818);
and U5709 (N_5709,N_5494,N_4831);
nand U5710 (N_5710,N_4852,N_5440);
xor U5711 (N_5711,N_4807,N_4881);
nand U5712 (N_5712,N_5426,N_5421);
nor U5713 (N_5713,N_5565,N_5233);
or U5714 (N_5714,N_5135,N_5311);
xor U5715 (N_5715,N_5572,N_4829);
nand U5716 (N_5716,N_5392,N_5453);
nand U5717 (N_5717,N_5067,N_4867);
xnor U5718 (N_5718,N_5145,N_4880);
nor U5719 (N_5719,N_5444,N_5348);
xor U5720 (N_5720,N_5400,N_4956);
and U5721 (N_5721,N_5449,N_5443);
nor U5722 (N_5722,N_5106,N_5203);
and U5723 (N_5723,N_5592,N_5172);
and U5724 (N_5724,N_5284,N_5096);
xnor U5725 (N_5725,N_5160,N_5505);
nand U5726 (N_5726,N_4988,N_5258);
xnor U5727 (N_5727,N_4995,N_4951);
nand U5728 (N_5728,N_5448,N_4920);
and U5729 (N_5729,N_5088,N_5351);
or U5730 (N_5730,N_5075,N_5452);
nor U5731 (N_5731,N_5116,N_5469);
nand U5732 (N_5732,N_5310,N_5536);
nand U5733 (N_5733,N_5163,N_4871);
nor U5734 (N_5734,N_5340,N_5445);
or U5735 (N_5735,N_5286,N_5070);
or U5736 (N_5736,N_5207,N_5398);
or U5737 (N_5737,N_5030,N_5064);
and U5738 (N_5738,N_4879,N_5142);
nand U5739 (N_5739,N_4806,N_4848);
and U5740 (N_5740,N_4989,N_5086);
nand U5741 (N_5741,N_5154,N_5479);
xnor U5742 (N_5742,N_5325,N_4906);
xnor U5743 (N_5743,N_4833,N_4800);
nand U5744 (N_5744,N_5059,N_4935);
xor U5745 (N_5745,N_4839,N_5007);
xor U5746 (N_5746,N_5066,N_5158);
xnor U5747 (N_5747,N_5277,N_5174);
or U5748 (N_5748,N_4936,N_4969);
nor U5749 (N_5749,N_4973,N_5161);
nand U5750 (N_5750,N_5581,N_5585);
nand U5751 (N_5751,N_5074,N_4821);
nand U5752 (N_5752,N_5201,N_5035);
and U5753 (N_5753,N_5417,N_5105);
and U5754 (N_5754,N_5379,N_5433);
and U5755 (N_5755,N_5098,N_5179);
nand U5756 (N_5756,N_5237,N_5038);
xor U5757 (N_5757,N_4918,N_5390);
and U5758 (N_5758,N_5406,N_5214);
nand U5759 (N_5759,N_4824,N_5056);
nor U5760 (N_5760,N_5188,N_5191);
and U5761 (N_5761,N_5205,N_4828);
nor U5762 (N_5762,N_4864,N_5598);
nor U5763 (N_5763,N_5322,N_5442);
and U5764 (N_5764,N_5006,N_5491);
and U5765 (N_5765,N_4844,N_5396);
and U5766 (N_5766,N_4825,N_5490);
xnor U5767 (N_5767,N_5190,N_4886);
nor U5768 (N_5768,N_4849,N_5000);
nor U5769 (N_5769,N_5459,N_5365);
or U5770 (N_5770,N_5545,N_5590);
nand U5771 (N_5771,N_5266,N_5489);
and U5772 (N_5772,N_5388,N_5526);
or U5773 (N_5773,N_5350,N_4930);
and U5774 (N_5774,N_5271,N_5378);
nand U5775 (N_5775,N_5554,N_5520);
xnor U5776 (N_5776,N_5078,N_5478);
xnor U5777 (N_5777,N_5298,N_5413);
xor U5778 (N_5778,N_5027,N_5169);
or U5779 (N_5779,N_4877,N_4985);
nor U5780 (N_5780,N_5275,N_5072);
nand U5781 (N_5781,N_5576,N_5299);
xnor U5782 (N_5782,N_5596,N_5465);
and U5783 (N_5783,N_4820,N_5241);
nand U5784 (N_5784,N_4961,N_5217);
or U5785 (N_5785,N_5242,N_5488);
nand U5786 (N_5786,N_5208,N_5288);
and U5787 (N_5787,N_5228,N_4929);
xnor U5788 (N_5788,N_5111,N_5177);
nand U5789 (N_5789,N_5457,N_5087);
and U5790 (N_5790,N_5032,N_5425);
and U5791 (N_5791,N_5530,N_5415);
xor U5792 (N_5792,N_5324,N_5361);
nand U5793 (N_5793,N_4926,N_5485);
nor U5794 (N_5794,N_5120,N_4802);
or U5795 (N_5795,N_4836,N_5437);
and U5796 (N_5796,N_5355,N_5436);
nor U5797 (N_5797,N_4846,N_4974);
or U5798 (N_5798,N_5496,N_5230);
nor U5799 (N_5799,N_5371,N_5053);
and U5800 (N_5800,N_5213,N_5559);
xnor U5801 (N_5801,N_5089,N_5281);
and U5802 (N_5802,N_4937,N_5588);
or U5803 (N_5803,N_5130,N_5245);
nor U5804 (N_5804,N_5337,N_4965);
and U5805 (N_5805,N_5473,N_4986);
nor U5806 (N_5806,N_5184,N_4968);
or U5807 (N_5807,N_5276,N_4813);
xnor U5808 (N_5808,N_5069,N_5410);
and U5809 (N_5809,N_5499,N_5004);
or U5810 (N_5810,N_5564,N_5364);
nor U5811 (N_5811,N_5471,N_5023);
and U5812 (N_5812,N_5357,N_5380);
nand U5813 (N_5813,N_5005,N_5194);
xnor U5814 (N_5814,N_4897,N_5541);
and U5815 (N_5815,N_5238,N_5249);
nand U5816 (N_5816,N_5571,N_5216);
or U5817 (N_5817,N_5029,N_4826);
and U5818 (N_5818,N_5232,N_5492);
nand U5819 (N_5819,N_5257,N_5497);
xnor U5820 (N_5820,N_4889,N_5556);
and U5821 (N_5821,N_4922,N_5209);
nor U5822 (N_5822,N_4875,N_5501);
xor U5823 (N_5823,N_5048,N_5367);
and U5824 (N_5824,N_4850,N_5578);
and U5825 (N_5825,N_5315,N_5094);
nand U5826 (N_5826,N_5539,N_4809);
or U5827 (N_5827,N_5427,N_4905);
nand U5828 (N_5828,N_5269,N_5270);
and U5829 (N_5829,N_5253,N_5302);
nand U5830 (N_5830,N_5402,N_5397);
and U5831 (N_5831,N_5055,N_4882);
and U5832 (N_5832,N_5429,N_5236);
nor U5833 (N_5833,N_5506,N_5552);
nand U5834 (N_5834,N_5435,N_5330);
or U5835 (N_5835,N_4984,N_5475);
or U5836 (N_5836,N_5393,N_5314);
nand U5837 (N_5837,N_5597,N_5063);
nand U5838 (N_5838,N_5422,N_5508);
and U5839 (N_5839,N_5407,N_5273);
and U5840 (N_5840,N_5102,N_5204);
or U5841 (N_5841,N_5123,N_5432);
and U5842 (N_5842,N_5317,N_5026);
xnor U5843 (N_5843,N_5431,N_5538);
xnor U5844 (N_5844,N_4945,N_5409);
or U5845 (N_5845,N_4921,N_5046);
nor U5846 (N_5846,N_5595,N_5438);
or U5847 (N_5847,N_5587,N_5186);
or U5848 (N_5848,N_5419,N_5339);
and U5849 (N_5849,N_5519,N_5131);
xor U5850 (N_5850,N_4884,N_5296);
nand U5851 (N_5851,N_4832,N_4856);
xnor U5852 (N_5852,N_4908,N_4885);
nand U5853 (N_5853,N_5215,N_5454);
nand U5854 (N_5854,N_5525,N_4972);
xnor U5855 (N_5855,N_5195,N_4817);
xnor U5856 (N_5856,N_5418,N_5531);
nand U5857 (N_5857,N_4934,N_5121);
and U5858 (N_5858,N_5295,N_4814);
or U5859 (N_5859,N_5524,N_5196);
nand U5860 (N_5860,N_5182,N_4851);
nand U5861 (N_5861,N_5156,N_5385);
or U5862 (N_5862,N_5414,N_5081);
nand U5863 (N_5863,N_5542,N_4954);
nor U5864 (N_5864,N_5532,N_5366);
and U5865 (N_5865,N_5358,N_4943);
nand U5866 (N_5866,N_5368,N_5009);
xor U5867 (N_5867,N_5175,N_4996);
xor U5868 (N_5868,N_5133,N_5080);
nand U5869 (N_5869,N_5170,N_5042);
or U5870 (N_5870,N_5301,N_5248);
or U5871 (N_5871,N_5246,N_4981);
or U5872 (N_5872,N_5137,N_5579);
xnor U5873 (N_5873,N_5206,N_4914);
or U5874 (N_5874,N_5095,N_5187);
nor U5875 (N_5875,N_5279,N_5155);
nand U5876 (N_5876,N_5180,N_5487);
and U5877 (N_5877,N_5077,N_5183);
nand U5878 (N_5878,N_5019,N_5008);
nand U5879 (N_5879,N_4967,N_5583);
xnor U5880 (N_5880,N_5162,N_5014);
and U5881 (N_5881,N_5384,N_5200);
or U5882 (N_5882,N_5580,N_5093);
and U5883 (N_5883,N_4847,N_5149);
nand U5884 (N_5884,N_5377,N_4997);
or U5885 (N_5885,N_4987,N_5002);
or U5886 (N_5886,N_5193,N_4822);
or U5887 (N_5887,N_5264,N_4909);
xnor U5888 (N_5888,N_5467,N_5293);
nor U5889 (N_5889,N_5319,N_5231);
nand U5890 (N_5890,N_4827,N_4903);
nand U5891 (N_5891,N_4811,N_5484);
or U5892 (N_5892,N_4955,N_5589);
or U5893 (N_5893,N_5219,N_4810);
or U5894 (N_5894,N_5256,N_4854);
xnor U5895 (N_5895,N_5221,N_5218);
or U5896 (N_5896,N_4898,N_5568);
nand U5897 (N_5897,N_5387,N_5354);
xor U5898 (N_5898,N_5463,N_5147);
xnor U5899 (N_5899,N_5528,N_4933);
and U5900 (N_5900,N_5502,N_5382);
xor U5901 (N_5901,N_5486,N_5047);
or U5902 (N_5902,N_5225,N_5020);
and U5903 (N_5903,N_5403,N_5458);
and U5904 (N_5904,N_5509,N_4878);
and U5905 (N_5905,N_4970,N_4874);
and U5906 (N_5906,N_5474,N_5252);
and U5907 (N_5907,N_5050,N_4978);
xnor U5908 (N_5908,N_5263,N_4910);
and U5909 (N_5909,N_5125,N_4808);
and U5910 (N_5910,N_5446,N_5132);
or U5911 (N_5911,N_5234,N_5110);
or U5912 (N_5912,N_5255,N_5168);
or U5913 (N_5913,N_5558,N_5124);
nor U5914 (N_5914,N_5015,N_4953);
and U5915 (N_5915,N_5332,N_5229);
xnor U5916 (N_5916,N_5251,N_4991);
or U5917 (N_5917,N_5303,N_4982);
or U5918 (N_5918,N_5326,N_5001);
nand U5919 (N_5919,N_5416,N_5320);
nand U5920 (N_5920,N_5372,N_5562);
xnor U5921 (N_5921,N_5470,N_4855);
nor U5922 (N_5922,N_5352,N_5294);
nor U5923 (N_5923,N_4888,N_5127);
nor U5924 (N_5924,N_4815,N_5462);
and U5925 (N_5925,N_5553,N_5451);
nand U5926 (N_5926,N_4912,N_5383);
or U5927 (N_5927,N_5345,N_5527);
nand U5928 (N_5928,N_5534,N_5483);
xor U5929 (N_5929,N_5341,N_5181);
nand U5930 (N_5930,N_4853,N_4865);
or U5931 (N_5931,N_5477,N_4924);
nor U5932 (N_5932,N_5369,N_5331);
nand U5933 (N_5933,N_5272,N_4971);
or U5934 (N_5934,N_5211,N_5346);
nor U5935 (N_5935,N_5356,N_5073);
xor U5936 (N_5936,N_5376,N_4902);
nor U5937 (N_5937,N_4979,N_5297);
xnor U5938 (N_5938,N_5394,N_5548);
nand U5939 (N_5939,N_5084,N_4873);
xor U5940 (N_5940,N_4823,N_5347);
nor U5941 (N_5941,N_5265,N_5329);
xnor U5942 (N_5942,N_5360,N_5342);
or U5943 (N_5943,N_4962,N_5512);
and U5944 (N_5944,N_5304,N_5567);
and U5945 (N_5945,N_5523,N_5159);
or U5946 (N_5946,N_5097,N_5244);
nor U5947 (N_5947,N_4870,N_4957);
or U5948 (N_5948,N_5153,N_5521);
xor U5949 (N_5949,N_5136,N_5107);
nand U5950 (N_5950,N_4872,N_4838);
nand U5951 (N_5951,N_5031,N_5373);
xor U5952 (N_5952,N_5051,N_5152);
xor U5953 (N_5953,N_5291,N_5574);
nor U5954 (N_5954,N_5099,N_5198);
and U5955 (N_5955,N_5591,N_5389);
xnor U5956 (N_5956,N_5060,N_5336);
and U5957 (N_5957,N_5381,N_5503);
nor U5958 (N_5958,N_5307,N_4939);
and U5959 (N_5959,N_5033,N_5082);
or U5960 (N_5960,N_4925,N_4876);
or U5961 (N_5961,N_5560,N_5139);
and U5962 (N_5962,N_5090,N_5480);
nor U5963 (N_5963,N_5083,N_5012);
xor U5964 (N_5964,N_5300,N_5223);
nand U5965 (N_5965,N_4927,N_5141);
xor U5966 (N_5966,N_5021,N_5202);
nand U5967 (N_5967,N_4883,N_5584);
nand U5968 (N_5968,N_4901,N_5285);
nor U5969 (N_5969,N_4966,N_5349);
nand U5970 (N_5970,N_4816,N_5343);
xnor U5971 (N_5971,N_4843,N_5566);
xnor U5972 (N_5972,N_5570,N_5235);
nand U5973 (N_5973,N_5173,N_4863);
and U5974 (N_5974,N_4944,N_5586);
or U5975 (N_5975,N_5112,N_5359);
nand U5976 (N_5976,N_5227,N_5140);
xnor U5977 (N_5977,N_4958,N_5157);
or U5978 (N_5978,N_4866,N_5226);
or U5979 (N_5979,N_4994,N_4819);
nand U5980 (N_5980,N_4919,N_5289);
xor U5981 (N_5981,N_5563,N_5222);
or U5982 (N_5982,N_4891,N_5013);
or U5983 (N_5983,N_4917,N_4928);
nor U5984 (N_5984,N_5333,N_4911);
nand U5985 (N_5985,N_5327,N_5062);
and U5986 (N_5986,N_5268,N_5274);
nor U5987 (N_5987,N_5076,N_5537);
nor U5988 (N_5988,N_5037,N_5109);
or U5989 (N_5989,N_5129,N_5313);
nand U5990 (N_5990,N_5412,N_4834);
xnor U5991 (N_5991,N_5024,N_5363);
and U5992 (N_5992,N_5472,N_4983);
nor U5993 (N_5993,N_4949,N_5468);
xor U5994 (N_5994,N_5529,N_5482);
nand U5995 (N_5995,N_5543,N_4913);
nor U5996 (N_5996,N_4931,N_5546);
nor U5997 (N_5997,N_5456,N_4947);
or U5998 (N_5998,N_5052,N_5114);
nand U5999 (N_5999,N_4998,N_5100);
nand U6000 (N_6000,N_5384,N_5533);
nor U6001 (N_6001,N_5087,N_5434);
or U6002 (N_6002,N_5050,N_5020);
or U6003 (N_6003,N_5324,N_4849);
nand U6004 (N_6004,N_5077,N_4923);
and U6005 (N_6005,N_5183,N_5579);
xor U6006 (N_6006,N_5250,N_5490);
nand U6007 (N_6007,N_5066,N_5314);
xor U6008 (N_6008,N_5118,N_5052);
xor U6009 (N_6009,N_5101,N_5507);
or U6010 (N_6010,N_5060,N_5133);
nor U6011 (N_6011,N_4987,N_4908);
nor U6012 (N_6012,N_4987,N_4963);
or U6013 (N_6013,N_5238,N_5121);
and U6014 (N_6014,N_5497,N_5017);
xnor U6015 (N_6015,N_5555,N_5458);
nand U6016 (N_6016,N_4891,N_5045);
and U6017 (N_6017,N_5402,N_5125);
or U6018 (N_6018,N_5369,N_5031);
or U6019 (N_6019,N_4809,N_5463);
nor U6020 (N_6020,N_4822,N_5326);
or U6021 (N_6021,N_5219,N_4943);
xor U6022 (N_6022,N_5228,N_5160);
nand U6023 (N_6023,N_5054,N_5160);
xnor U6024 (N_6024,N_5054,N_4856);
or U6025 (N_6025,N_5337,N_5460);
nand U6026 (N_6026,N_5417,N_4960);
xor U6027 (N_6027,N_5591,N_5303);
xor U6028 (N_6028,N_4839,N_4887);
nor U6029 (N_6029,N_5167,N_5488);
and U6030 (N_6030,N_5292,N_5397);
nand U6031 (N_6031,N_5241,N_5201);
nor U6032 (N_6032,N_5146,N_5152);
or U6033 (N_6033,N_4918,N_4893);
and U6034 (N_6034,N_5190,N_4875);
and U6035 (N_6035,N_5053,N_5329);
nor U6036 (N_6036,N_4902,N_5286);
or U6037 (N_6037,N_5419,N_5495);
nand U6038 (N_6038,N_5231,N_4941);
xor U6039 (N_6039,N_4986,N_5130);
nand U6040 (N_6040,N_5288,N_5381);
xor U6041 (N_6041,N_5567,N_4852);
xor U6042 (N_6042,N_5263,N_4894);
nor U6043 (N_6043,N_4906,N_5547);
nor U6044 (N_6044,N_5315,N_5369);
and U6045 (N_6045,N_5295,N_5015);
nand U6046 (N_6046,N_5100,N_5440);
or U6047 (N_6047,N_5319,N_5078);
nand U6048 (N_6048,N_4942,N_5585);
and U6049 (N_6049,N_5584,N_5454);
nand U6050 (N_6050,N_4945,N_5170);
xnor U6051 (N_6051,N_5552,N_5533);
nor U6052 (N_6052,N_5104,N_5402);
or U6053 (N_6053,N_5492,N_5315);
nand U6054 (N_6054,N_5323,N_5202);
nand U6055 (N_6055,N_4928,N_5584);
nor U6056 (N_6056,N_5364,N_5395);
nor U6057 (N_6057,N_5281,N_5498);
nand U6058 (N_6058,N_5378,N_5114);
nand U6059 (N_6059,N_5226,N_5515);
nand U6060 (N_6060,N_5070,N_5514);
xnor U6061 (N_6061,N_5196,N_5296);
nor U6062 (N_6062,N_5591,N_4828);
nand U6063 (N_6063,N_5137,N_5099);
nand U6064 (N_6064,N_5501,N_5059);
nor U6065 (N_6065,N_5183,N_4821);
and U6066 (N_6066,N_5403,N_5244);
and U6067 (N_6067,N_5287,N_5557);
nand U6068 (N_6068,N_5136,N_4854);
nand U6069 (N_6069,N_5303,N_4881);
and U6070 (N_6070,N_5447,N_4851);
nand U6071 (N_6071,N_5585,N_4904);
xnor U6072 (N_6072,N_4808,N_5331);
xnor U6073 (N_6073,N_5514,N_5431);
or U6074 (N_6074,N_5103,N_5129);
and U6075 (N_6075,N_4956,N_5033);
nand U6076 (N_6076,N_5505,N_5257);
or U6077 (N_6077,N_5227,N_5366);
nand U6078 (N_6078,N_5135,N_5497);
nand U6079 (N_6079,N_5136,N_5085);
nor U6080 (N_6080,N_5149,N_4837);
xnor U6081 (N_6081,N_5448,N_5319);
or U6082 (N_6082,N_5319,N_4940);
nor U6083 (N_6083,N_5183,N_4956);
nor U6084 (N_6084,N_4932,N_4850);
nor U6085 (N_6085,N_5244,N_5521);
or U6086 (N_6086,N_5458,N_5166);
nand U6087 (N_6087,N_5267,N_4898);
nor U6088 (N_6088,N_5026,N_5396);
and U6089 (N_6089,N_5153,N_5037);
nand U6090 (N_6090,N_5542,N_5385);
nand U6091 (N_6091,N_5428,N_4933);
and U6092 (N_6092,N_5227,N_5278);
xor U6093 (N_6093,N_5408,N_5474);
or U6094 (N_6094,N_5596,N_5272);
xor U6095 (N_6095,N_5128,N_4998);
and U6096 (N_6096,N_5284,N_5588);
or U6097 (N_6097,N_5072,N_5429);
and U6098 (N_6098,N_5158,N_5025);
xor U6099 (N_6099,N_4917,N_5357);
and U6100 (N_6100,N_5587,N_5019);
and U6101 (N_6101,N_5174,N_5085);
or U6102 (N_6102,N_5068,N_5543);
xor U6103 (N_6103,N_4879,N_5180);
xor U6104 (N_6104,N_4873,N_5211);
nor U6105 (N_6105,N_5372,N_5390);
nand U6106 (N_6106,N_4982,N_5086);
or U6107 (N_6107,N_5598,N_5005);
xnor U6108 (N_6108,N_5565,N_5239);
xor U6109 (N_6109,N_4911,N_5268);
nor U6110 (N_6110,N_4961,N_5546);
nor U6111 (N_6111,N_5477,N_5172);
nor U6112 (N_6112,N_5413,N_5235);
xnor U6113 (N_6113,N_5157,N_5476);
or U6114 (N_6114,N_5587,N_4996);
nor U6115 (N_6115,N_5321,N_5009);
or U6116 (N_6116,N_5463,N_5497);
nor U6117 (N_6117,N_4914,N_5419);
or U6118 (N_6118,N_5281,N_5027);
nand U6119 (N_6119,N_5333,N_4978);
xor U6120 (N_6120,N_5023,N_4801);
xor U6121 (N_6121,N_5046,N_5134);
and U6122 (N_6122,N_5114,N_4807);
and U6123 (N_6123,N_5443,N_5114);
nor U6124 (N_6124,N_5316,N_5156);
nor U6125 (N_6125,N_5004,N_4883);
and U6126 (N_6126,N_5582,N_4806);
nand U6127 (N_6127,N_5306,N_4975);
nor U6128 (N_6128,N_5566,N_5175);
nor U6129 (N_6129,N_5318,N_5510);
and U6130 (N_6130,N_5012,N_5512);
nand U6131 (N_6131,N_4903,N_5346);
nand U6132 (N_6132,N_5054,N_4932);
and U6133 (N_6133,N_5096,N_5584);
or U6134 (N_6134,N_5330,N_4902);
nor U6135 (N_6135,N_4805,N_4838);
nor U6136 (N_6136,N_4984,N_4976);
and U6137 (N_6137,N_5046,N_5071);
or U6138 (N_6138,N_5201,N_5190);
and U6139 (N_6139,N_5077,N_4851);
nand U6140 (N_6140,N_4843,N_5322);
nor U6141 (N_6141,N_4859,N_5420);
xor U6142 (N_6142,N_5451,N_4998);
nand U6143 (N_6143,N_5369,N_4800);
or U6144 (N_6144,N_5165,N_4950);
or U6145 (N_6145,N_5525,N_4961);
xor U6146 (N_6146,N_4964,N_4841);
and U6147 (N_6147,N_5093,N_5137);
xor U6148 (N_6148,N_5536,N_5462);
xor U6149 (N_6149,N_5258,N_4892);
and U6150 (N_6150,N_4838,N_5052);
nand U6151 (N_6151,N_5524,N_5024);
xnor U6152 (N_6152,N_5053,N_4844);
xnor U6153 (N_6153,N_4965,N_5529);
nand U6154 (N_6154,N_5305,N_4978);
xnor U6155 (N_6155,N_5434,N_4822);
and U6156 (N_6156,N_5169,N_5580);
xor U6157 (N_6157,N_4881,N_4981);
xnor U6158 (N_6158,N_5381,N_5374);
nor U6159 (N_6159,N_5296,N_5310);
and U6160 (N_6160,N_5201,N_5395);
nor U6161 (N_6161,N_5231,N_5143);
or U6162 (N_6162,N_5417,N_5083);
or U6163 (N_6163,N_5126,N_5338);
or U6164 (N_6164,N_5018,N_5093);
or U6165 (N_6165,N_5096,N_5391);
or U6166 (N_6166,N_5142,N_5059);
xnor U6167 (N_6167,N_5265,N_4854);
and U6168 (N_6168,N_4972,N_5129);
xnor U6169 (N_6169,N_5311,N_5532);
or U6170 (N_6170,N_4874,N_5501);
nor U6171 (N_6171,N_5460,N_5576);
and U6172 (N_6172,N_4936,N_5432);
nor U6173 (N_6173,N_4805,N_5229);
nand U6174 (N_6174,N_4886,N_5105);
nor U6175 (N_6175,N_5354,N_5025);
or U6176 (N_6176,N_5354,N_4820);
xor U6177 (N_6177,N_4817,N_4998);
or U6178 (N_6178,N_5530,N_5503);
nor U6179 (N_6179,N_5593,N_5090);
xnor U6180 (N_6180,N_5307,N_5275);
nor U6181 (N_6181,N_5317,N_5444);
and U6182 (N_6182,N_4952,N_5057);
nor U6183 (N_6183,N_5584,N_5592);
or U6184 (N_6184,N_5358,N_5392);
nand U6185 (N_6185,N_5277,N_5444);
xnor U6186 (N_6186,N_5114,N_5112);
xnor U6187 (N_6187,N_5456,N_5216);
nand U6188 (N_6188,N_5348,N_4813);
xor U6189 (N_6189,N_5316,N_5154);
nand U6190 (N_6190,N_5031,N_5275);
nand U6191 (N_6191,N_4966,N_5565);
nand U6192 (N_6192,N_5108,N_4872);
or U6193 (N_6193,N_4994,N_5235);
xor U6194 (N_6194,N_4867,N_5069);
nand U6195 (N_6195,N_5122,N_5044);
or U6196 (N_6196,N_5388,N_5482);
and U6197 (N_6197,N_4974,N_5314);
and U6198 (N_6198,N_5343,N_5105);
or U6199 (N_6199,N_5474,N_5337);
and U6200 (N_6200,N_5165,N_5250);
or U6201 (N_6201,N_5243,N_5496);
xnor U6202 (N_6202,N_5021,N_5463);
nor U6203 (N_6203,N_4909,N_5517);
nand U6204 (N_6204,N_4807,N_5338);
or U6205 (N_6205,N_4818,N_4919);
nor U6206 (N_6206,N_5389,N_5366);
or U6207 (N_6207,N_5072,N_5568);
nand U6208 (N_6208,N_5044,N_5483);
nor U6209 (N_6209,N_5389,N_5133);
xor U6210 (N_6210,N_4833,N_5282);
and U6211 (N_6211,N_5430,N_5090);
and U6212 (N_6212,N_5065,N_4997);
nor U6213 (N_6213,N_5165,N_5437);
or U6214 (N_6214,N_5129,N_5100);
xor U6215 (N_6215,N_5326,N_4996);
xnor U6216 (N_6216,N_5489,N_5196);
and U6217 (N_6217,N_5304,N_4816);
nand U6218 (N_6218,N_4876,N_5470);
nor U6219 (N_6219,N_5084,N_5511);
nor U6220 (N_6220,N_5365,N_5558);
and U6221 (N_6221,N_5183,N_5487);
and U6222 (N_6222,N_4932,N_5086);
nand U6223 (N_6223,N_5222,N_5292);
and U6224 (N_6224,N_5291,N_5236);
or U6225 (N_6225,N_5090,N_5431);
or U6226 (N_6226,N_5432,N_5372);
or U6227 (N_6227,N_5243,N_4941);
or U6228 (N_6228,N_4863,N_4948);
and U6229 (N_6229,N_5396,N_5045);
nor U6230 (N_6230,N_5585,N_5191);
xor U6231 (N_6231,N_5082,N_4909);
xnor U6232 (N_6232,N_5360,N_5466);
nor U6233 (N_6233,N_4966,N_4932);
nand U6234 (N_6234,N_5414,N_5006);
nor U6235 (N_6235,N_5086,N_4809);
and U6236 (N_6236,N_5331,N_5261);
xnor U6237 (N_6237,N_4868,N_5015);
and U6238 (N_6238,N_5360,N_5067);
or U6239 (N_6239,N_5509,N_4865);
or U6240 (N_6240,N_5220,N_5066);
nand U6241 (N_6241,N_4879,N_5146);
nor U6242 (N_6242,N_5394,N_5132);
or U6243 (N_6243,N_5025,N_5473);
nor U6244 (N_6244,N_4953,N_5198);
or U6245 (N_6245,N_5370,N_4830);
xnor U6246 (N_6246,N_4872,N_5531);
xor U6247 (N_6247,N_4959,N_5001);
xnor U6248 (N_6248,N_5511,N_4951);
or U6249 (N_6249,N_5512,N_4977);
nor U6250 (N_6250,N_5150,N_5421);
nand U6251 (N_6251,N_5343,N_4862);
and U6252 (N_6252,N_4935,N_5275);
xor U6253 (N_6253,N_5201,N_4922);
and U6254 (N_6254,N_5018,N_5544);
and U6255 (N_6255,N_5422,N_4879);
or U6256 (N_6256,N_5172,N_4949);
xor U6257 (N_6257,N_5482,N_5206);
xnor U6258 (N_6258,N_4827,N_5158);
nand U6259 (N_6259,N_5110,N_5457);
or U6260 (N_6260,N_5235,N_5587);
nand U6261 (N_6261,N_5166,N_5220);
nand U6262 (N_6262,N_4884,N_4906);
xor U6263 (N_6263,N_4970,N_5101);
nand U6264 (N_6264,N_5553,N_4941);
or U6265 (N_6265,N_4951,N_5546);
nand U6266 (N_6266,N_4868,N_5203);
xor U6267 (N_6267,N_5401,N_4836);
or U6268 (N_6268,N_5169,N_5152);
xor U6269 (N_6269,N_5586,N_4823);
xor U6270 (N_6270,N_4884,N_4955);
or U6271 (N_6271,N_5109,N_5483);
nor U6272 (N_6272,N_5398,N_4910);
and U6273 (N_6273,N_5231,N_5094);
nand U6274 (N_6274,N_4970,N_4903);
xnor U6275 (N_6275,N_5397,N_5444);
and U6276 (N_6276,N_5137,N_5239);
and U6277 (N_6277,N_5168,N_4901);
or U6278 (N_6278,N_4978,N_5232);
or U6279 (N_6279,N_5187,N_4912);
nor U6280 (N_6280,N_5001,N_5011);
nand U6281 (N_6281,N_5490,N_5463);
and U6282 (N_6282,N_5265,N_5580);
nor U6283 (N_6283,N_5429,N_5111);
nor U6284 (N_6284,N_5579,N_5542);
or U6285 (N_6285,N_5552,N_4883);
and U6286 (N_6286,N_5462,N_5208);
xor U6287 (N_6287,N_5440,N_5160);
or U6288 (N_6288,N_5235,N_5424);
or U6289 (N_6289,N_5210,N_4913);
nor U6290 (N_6290,N_4919,N_5054);
nor U6291 (N_6291,N_5570,N_5415);
xor U6292 (N_6292,N_4896,N_5207);
or U6293 (N_6293,N_5424,N_5086);
nand U6294 (N_6294,N_4946,N_4941);
xnor U6295 (N_6295,N_5106,N_4837);
and U6296 (N_6296,N_4804,N_4949);
or U6297 (N_6297,N_4967,N_4985);
and U6298 (N_6298,N_4844,N_5337);
nor U6299 (N_6299,N_5555,N_5522);
and U6300 (N_6300,N_4855,N_5122);
or U6301 (N_6301,N_5221,N_5448);
nand U6302 (N_6302,N_4961,N_5362);
xor U6303 (N_6303,N_4910,N_5072);
or U6304 (N_6304,N_5393,N_4965);
nor U6305 (N_6305,N_5375,N_4851);
or U6306 (N_6306,N_5587,N_4947);
and U6307 (N_6307,N_5457,N_5422);
nand U6308 (N_6308,N_5127,N_5338);
nor U6309 (N_6309,N_5086,N_5462);
or U6310 (N_6310,N_5486,N_5472);
xnor U6311 (N_6311,N_4831,N_5569);
xnor U6312 (N_6312,N_5542,N_5052);
nand U6313 (N_6313,N_5111,N_5539);
xor U6314 (N_6314,N_5489,N_5299);
and U6315 (N_6315,N_5531,N_5511);
and U6316 (N_6316,N_5007,N_4924);
xnor U6317 (N_6317,N_5105,N_4912);
nand U6318 (N_6318,N_5567,N_4959);
or U6319 (N_6319,N_4960,N_4847);
nor U6320 (N_6320,N_5473,N_5059);
nor U6321 (N_6321,N_5017,N_4998);
nand U6322 (N_6322,N_5545,N_5029);
xor U6323 (N_6323,N_5164,N_4842);
or U6324 (N_6324,N_5257,N_5181);
nand U6325 (N_6325,N_5404,N_5271);
xor U6326 (N_6326,N_4887,N_5023);
nor U6327 (N_6327,N_5314,N_5411);
nand U6328 (N_6328,N_5434,N_4829);
nand U6329 (N_6329,N_5246,N_4891);
nand U6330 (N_6330,N_5573,N_4938);
or U6331 (N_6331,N_5024,N_5528);
xnor U6332 (N_6332,N_4802,N_5178);
nand U6333 (N_6333,N_5290,N_5493);
nor U6334 (N_6334,N_4969,N_5065);
and U6335 (N_6335,N_4828,N_5387);
or U6336 (N_6336,N_5274,N_5139);
xor U6337 (N_6337,N_5034,N_4950);
nor U6338 (N_6338,N_5195,N_5430);
or U6339 (N_6339,N_5561,N_5349);
nand U6340 (N_6340,N_5412,N_5170);
xnor U6341 (N_6341,N_5493,N_5090);
nand U6342 (N_6342,N_5429,N_5338);
and U6343 (N_6343,N_5090,N_4993);
nand U6344 (N_6344,N_5288,N_5262);
or U6345 (N_6345,N_5076,N_5496);
or U6346 (N_6346,N_4855,N_4831);
nor U6347 (N_6347,N_4953,N_4903);
and U6348 (N_6348,N_5228,N_5541);
xor U6349 (N_6349,N_5583,N_5105);
and U6350 (N_6350,N_5328,N_4810);
xnor U6351 (N_6351,N_5449,N_5444);
or U6352 (N_6352,N_4960,N_5245);
and U6353 (N_6353,N_5412,N_4867);
nand U6354 (N_6354,N_4854,N_4980);
xnor U6355 (N_6355,N_5133,N_5423);
or U6356 (N_6356,N_5475,N_5304);
nand U6357 (N_6357,N_4973,N_4950);
nor U6358 (N_6358,N_5599,N_4867);
nor U6359 (N_6359,N_4823,N_5496);
xor U6360 (N_6360,N_4943,N_4977);
xnor U6361 (N_6361,N_5080,N_4876);
or U6362 (N_6362,N_4843,N_5396);
xor U6363 (N_6363,N_5305,N_5144);
nand U6364 (N_6364,N_4861,N_4863);
or U6365 (N_6365,N_5447,N_5075);
xnor U6366 (N_6366,N_4871,N_5208);
or U6367 (N_6367,N_5270,N_4935);
nor U6368 (N_6368,N_4850,N_4944);
xnor U6369 (N_6369,N_5271,N_5081);
and U6370 (N_6370,N_4975,N_5338);
xnor U6371 (N_6371,N_5166,N_4857);
nor U6372 (N_6372,N_5029,N_4846);
or U6373 (N_6373,N_5105,N_5242);
or U6374 (N_6374,N_5250,N_4935);
nor U6375 (N_6375,N_5507,N_5234);
nor U6376 (N_6376,N_5021,N_4940);
xnor U6377 (N_6377,N_5386,N_5040);
xnor U6378 (N_6378,N_5537,N_5564);
or U6379 (N_6379,N_5298,N_5396);
or U6380 (N_6380,N_5116,N_4812);
or U6381 (N_6381,N_5240,N_5429);
xor U6382 (N_6382,N_4904,N_5450);
xor U6383 (N_6383,N_5599,N_5397);
or U6384 (N_6384,N_5161,N_4870);
nor U6385 (N_6385,N_5169,N_5456);
nand U6386 (N_6386,N_4936,N_4958);
and U6387 (N_6387,N_5379,N_5172);
xor U6388 (N_6388,N_4806,N_5029);
xnor U6389 (N_6389,N_5589,N_5426);
xnor U6390 (N_6390,N_5208,N_5369);
nor U6391 (N_6391,N_5136,N_5288);
xor U6392 (N_6392,N_4955,N_5585);
nand U6393 (N_6393,N_4978,N_5541);
and U6394 (N_6394,N_5337,N_5180);
or U6395 (N_6395,N_5575,N_4949);
nor U6396 (N_6396,N_4962,N_5380);
and U6397 (N_6397,N_5332,N_4952);
xnor U6398 (N_6398,N_5569,N_5290);
nor U6399 (N_6399,N_5028,N_4999);
and U6400 (N_6400,N_5705,N_6279);
nand U6401 (N_6401,N_5603,N_6055);
or U6402 (N_6402,N_6249,N_6372);
and U6403 (N_6403,N_5731,N_5871);
and U6404 (N_6404,N_6046,N_5861);
and U6405 (N_6405,N_5772,N_5972);
or U6406 (N_6406,N_6258,N_5804);
or U6407 (N_6407,N_6302,N_6362);
or U6408 (N_6408,N_5931,N_6301);
and U6409 (N_6409,N_5905,N_6032);
nand U6410 (N_6410,N_5870,N_5893);
or U6411 (N_6411,N_5835,N_6070);
and U6412 (N_6412,N_5950,N_5974);
nor U6413 (N_6413,N_6259,N_5612);
nor U6414 (N_6414,N_5765,N_5727);
nand U6415 (N_6415,N_5736,N_6242);
or U6416 (N_6416,N_5919,N_5933);
nor U6417 (N_6417,N_6061,N_5767);
xnor U6418 (N_6418,N_5797,N_6235);
xnor U6419 (N_6419,N_6311,N_5740);
nor U6420 (N_6420,N_5661,N_6024);
and U6421 (N_6421,N_6039,N_6113);
and U6422 (N_6422,N_6331,N_5730);
nand U6423 (N_6423,N_5602,N_5786);
and U6424 (N_6424,N_6236,N_5822);
nor U6425 (N_6425,N_6318,N_6391);
nand U6426 (N_6426,N_5640,N_5891);
nor U6427 (N_6427,N_6351,N_5794);
or U6428 (N_6428,N_5796,N_5968);
and U6429 (N_6429,N_5608,N_6095);
nor U6430 (N_6430,N_5660,N_6075);
nor U6431 (N_6431,N_5998,N_5915);
and U6432 (N_6432,N_5700,N_6117);
and U6433 (N_6433,N_6042,N_6197);
and U6434 (N_6434,N_6264,N_5724);
xnor U6435 (N_6435,N_6228,N_6299);
nand U6436 (N_6436,N_6066,N_5708);
and U6437 (N_6437,N_6270,N_6143);
and U6438 (N_6438,N_5795,N_6155);
or U6439 (N_6439,N_5646,N_5834);
and U6440 (N_6440,N_6247,N_5672);
nor U6441 (N_6441,N_6037,N_5890);
nand U6442 (N_6442,N_5941,N_5865);
and U6443 (N_6443,N_6102,N_6146);
nor U6444 (N_6444,N_6223,N_6166);
or U6445 (N_6445,N_5627,N_5840);
nand U6446 (N_6446,N_5799,N_5971);
or U6447 (N_6447,N_6163,N_6184);
nand U6448 (N_6448,N_5630,N_6380);
nor U6449 (N_6449,N_5788,N_5954);
or U6450 (N_6450,N_5889,N_6314);
and U6451 (N_6451,N_5956,N_6225);
and U6452 (N_6452,N_5748,N_6261);
or U6453 (N_6453,N_6052,N_5743);
nor U6454 (N_6454,N_6136,N_6110);
and U6455 (N_6455,N_5671,N_5802);
and U6456 (N_6456,N_6312,N_5645);
and U6457 (N_6457,N_6126,N_5668);
nor U6458 (N_6458,N_5754,N_5864);
nand U6459 (N_6459,N_6255,N_5658);
and U6460 (N_6460,N_5911,N_6149);
or U6461 (N_6461,N_5706,N_5914);
or U6462 (N_6462,N_5621,N_5981);
nand U6463 (N_6463,N_6229,N_5857);
nor U6464 (N_6464,N_5813,N_6240);
or U6465 (N_6465,N_5615,N_5841);
or U6466 (N_6466,N_6375,N_5928);
or U6467 (N_6467,N_5847,N_5644);
nor U6468 (N_6468,N_5854,N_6260);
xnor U6469 (N_6469,N_6142,N_6368);
or U6470 (N_6470,N_6180,N_6010);
or U6471 (N_6471,N_5780,N_5805);
or U6472 (N_6472,N_5641,N_6127);
nand U6473 (N_6473,N_6219,N_5634);
or U6474 (N_6474,N_6020,N_6073);
xnor U6475 (N_6475,N_5811,N_6334);
and U6476 (N_6476,N_5846,N_5701);
nor U6477 (N_6477,N_6332,N_5942);
nand U6478 (N_6478,N_5806,N_5878);
nand U6479 (N_6479,N_6144,N_5616);
nand U6480 (N_6480,N_5753,N_6213);
nor U6481 (N_6481,N_6088,N_6054);
nand U6482 (N_6482,N_5977,N_6145);
xnor U6483 (N_6483,N_5651,N_5939);
xor U6484 (N_6484,N_6252,N_5747);
xnor U6485 (N_6485,N_5844,N_5623);
nor U6486 (N_6486,N_5745,N_6385);
or U6487 (N_6487,N_5979,N_5978);
nand U6488 (N_6488,N_5716,N_5666);
and U6489 (N_6489,N_5965,N_6359);
xnor U6490 (N_6490,N_6370,N_6356);
xnor U6491 (N_6491,N_5992,N_6023);
nor U6492 (N_6492,N_5702,N_6273);
or U6493 (N_6493,N_5775,N_6369);
nand U6494 (N_6494,N_5960,N_6079);
and U6495 (N_6495,N_6243,N_5898);
xor U6496 (N_6496,N_6028,N_5924);
or U6497 (N_6497,N_5963,N_6305);
nand U6498 (N_6498,N_5613,N_6189);
or U6499 (N_6499,N_6014,N_6187);
or U6500 (N_6500,N_5899,N_6328);
nor U6501 (N_6501,N_6101,N_6103);
or U6502 (N_6502,N_5798,N_5885);
nor U6503 (N_6503,N_6390,N_5684);
xnor U6504 (N_6504,N_6324,N_5945);
nand U6505 (N_6505,N_5930,N_6220);
nor U6506 (N_6506,N_5638,N_6090);
and U6507 (N_6507,N_5962,N_6364);
nor U6508 (N_6508,N_6063,N_5860);
nand U6509 (N_6509,N_5696,N_6129);
and U6510 (N_6510,N_6160,N_6268);
or U6511 (N_6511,N_6076,N_6257);
or U6512 (N_6512,N_5738,N_6276);
and U6513 (N_6513,N_6360,N_6343);
or U6514 (N_6514,N_6285,N_5807);
or U6515 (N_6515,N_5699,N_6361);
or U6516 (N_6516,N_5784,N_5709);
or U6517 (N_6517,N_6043,N_5770);
nand U6518 (N_6518,N_5882,N_6005);
or U6519 (N_6519,N_5823,N_5764);
nand U6520 (N_6520,N_5869,N_5635);
nor U6521 (N_6521,N_6156,N_5663);
or U6522 (N_6522,N_6341,N_6111);
xnor U6523 (N_6523,N_5676,N_5987);
and U6524 (N_6524,N_6315,N_6135);
or U6525 (N_6525,N_5674,N_6104);
or U6526 (N_6526,N_6322,N_6122);
nor U6527 (N_6527,N_5734,N_5791);
nand U6528 (N_6528,N_6057,N_5852);
and U6529 (N_6529,N_6082,N_6224);
nor U6530 (N_6530,N_6137,N_6231);
or U6531 (N_6531,N_6041,N_6123);
or U6532 (N_6532,N_5913,N_6233);
and U6533 (N_6533,N_5717,N_5850);
nor U6534 (N_6534,N_5842,N_5648);
and U6535 (N_6535,N_5895,N_5925);
nor U6536 (N_6536,N_5779,N_6188);
xnor U6537 (N_6537,N_5703,N_5637);
xnor U6538 (N_6538,N_6193,N_6139);
or U6539 (N_6539,N_6350,N_6282);
nor U6540 (N_6540,N_5690,N_5848);
nand U6541 (N_6541,N_6326,N_6178);
nand U6542 (N_6542,N_5948,N_5910);
and U6543 (N_6543,N_6310,N_6033);
xor U6544 (N_6544,N_5995,N_5988);
or U6545 (N_6545,N_5722,N_5601);
nand U6546 (N_6546,N_6347,N_5920);
nor U6547 (N_6547,N_6296,N_6392);
nor U6548 (N_6548,N_6116,N_5946);
nand U6549 (N_6549,N_6298,N_6304);
or U6550 (N_6550,N_6294,N_5606);
xor U6551 (N_6551,N_5793,N_6287);
xnor U6552 (N_6552,N_5958,N_5940);
xor U6553 (N_6553,N_5994,N_6018);
and U6554 (N_6554,N_6140,N_6049);
or U6555 (N_6555,N_6256,N_5626);
nand U6556 (N_6556,N_6214,N_6040);
xnor U6557 (N_6557,N_6269,N_5952);
or U6558 (N_6558,N_6218,N_6281);
nand U6559 (N_6559,N_6093,N_5761);
nor U6560 (N_6560,N_5605,N_6044);
xor U6561 (N_6561,N_6297,N_5755);
nor U6562 (N_6562,N_6272,N_5787);
or U6563 (N_6563,N_6319,N_5728);
or U6564 (N_6564,N_5639,N_6004);
and U6565 (N_6565,N_5886,N_5636);
nor U6566 (N_6566,N_5888,N_6124);
nand U6567 (N_6567,N_5991,N_6118);
nor U6568 (N_6568,N_6352,N_6266);
nor U6569 (N_6569,N_6058,N_5678);
nor U6570 (N_6570,N_6340,N_6177);
or U6571 (N_6571,N_6141,N_5729);
or U6572 (N_6572,N_6098,N_6085);
xnor U6573 (N_6573,N_5820,N_5969);
and U6574 (N_6574,N_6164,N_5664);
nor U6575 (N_6575,N_6349,N_6196);
nor U6576 (N_6576,N_6363,N_6171);
and U6577 (N_6577,N_6115,N_5771);
xnor U6578 (N_6578,N_6374,N_6308);
or U6579 (N_6579,N_5725,N_6367);
nand U6580 (N_6580,N_6195,N_6176);
nand U6581 (N_6581,N_5762,N_5907);
or U6582 (N_6582,N_5826,N_5935);
nor U6583 (N_6583,N_5789,N_5611);
and U6584 (N_6584,N_6013,N_5906);
and U6585 (N_6585,N_6212,N_5752);
and U6586 (N_6586,N_5815,N_6207);
nand U6587 (N_6587,N_6080,N_6234);
nand U6588 (N_6588,N_5836,N_5726);
nand U6589 (N_6589,N_5733,N_6274);
nor U6590 (N_6590,N_6288,N_5961);
and U6591 (N_6591,N_5902,N_5713);
xnor U6592 (N_6592,N_6025,N_6353);
nand U6593 (N_6593,N_6151,N_6121);
nor U6594 (N_6594,N_5679,N_5629);
nor U6595 (N_6595,N_5973,N_5970);
and U6596 (N_6596,N_6377,N_5737);
and U6597 (N_6597,N_5916,N_6109);
nand U6598 (N_6598,N_6211,N_5883);
nor U6599 (N_6599,N_5665,N_6271);
nand U6600 (N_6600,N_5817,N_6064);
or U6601 (N_6601,N_5859,N_6344);
nand U6602 (N_6602,N_6148,N_5695);
nor U6603 (N_6603,N_5760,N_6008);
and U6604 (N_6604,N_6069,N_5633);
xnor U6605 (N_6605,N_6091,N_6190);
xor U6606 (N_6606,N_6208,N_6241);
or U6607 (N_6607,N_5845,N_5872);
nand U6608 (N_6608,N_6002,N_6333);
xnor U6609 (N_6609,N_6381,N_5758);
or U6610 (N_6610,N_5604,N_5909);
xnor U6611 (N_6611,N_6120,N_6267);
or U6612 (N_6612,N_6396,N_6316);
nand U6613 (N_6613,N_6003,N_5877);
nor U6614 (N_6614,N_5742,N_5618);
nor U6615 (N_6615,N_6017,N_6265);
xor U6616 (N_6616,N_6125,N_6194);
and U6617 (N_6617,N_6321,N_6339);
or U6618 (N_6618,N_5750,N_6048);
nand U6619 (N_6619,N_5715,N_5757);
xnor U6620 (N_6620,N_6320,N_6185);
xnor U6621 (N_6621,N_5620,N_5875);
nand U6622 (N_6622,N_5818,N_5964);
and U6623 (N_6623,N_5921,N_5918);
nor U6624 (N_6624,N_5783,N_5975);
nor U6625 (N_6625,N_6081,N_5867);
and U6626 (N_6626,N_6134,N_5862);
xor U6627 (N_6627,N_6210,N_6348);
nand U6628 (N_6628,N_5670,N_5986);
nand U6629 (N_6629,N_6153,N_5816);
and U6630 (N_6630,N_6071,N_5685);
nor U6631 (N_6631,N_6067,N_5934);
and U6632 (N_6632,N_6202,N_6289);
nand U6633 (N_6633,N_6376,N_6131);
xor U6634 (N_6634,N_6226,N_5617);
xnor U6635 (N_6635,N_5776,N_5989);
nor U6636 (N_6636,N_6152,N_5976);
nand U6637 (N_6637,N_6035,N_5751);
xnor U6638 (N_6638,N_5947,N_5686);
and U6639 (N_6639,N_5838,N_5720);
xor U6640 (N_6640,N_6133,N_5653);
nor U6641 (N_6641,N_6205,N_5614);
or U6642 (N_6642,N_5652,N_5773);
nand U6643 (N_6643,N_6387,N_5721);
or U6644 (N_6644,N_6337,N_6345);
and U6645 (N_6645,N_5829,N_5622);
or U6646 (N_6646,N_6161,N_6238);
nor U6647 (N_6647,N_6128,N_6206);
xor U6648 (N_6648,N_6094,N_6244);
nor U6649 (N_6649,N_5984,N_5719);
nand U6650 (N_6650,N_6378,N_6038);
nor U6651 (N_6651,N_6313,N_6277);
nor U6652 (N_6652,N_5607,N_6026);
xor U6653 (N_6653,N_6165,N_6373);
xor U6654 (N_6654,N_6114,N_5997);
and U6655 (N_6655,N_6072,N_6263);
xnor U6656 (N_6656,N_6130,N_5749);
xor U6657 (N_6657,N_5851,N_5959);
xnor U6658 (N_6658,N_6254,N_5936);
and U6659 (N_6659,N_6157,N_5812);
nor U6660 (N_6660,N_5853,N_6097);
nor U6661 (N_6661,N_6280,N_6059);
xnor U6662 (N_6662,N_5874,N_6016);
nand U6663 (N_6663,N_5912,N_5688);
xor U6664 (N_6664,N_6357,N_5632);
nand U6665 (N_6665,N_5662,N_5955);
nand U6666 (N_6666,N_5704,N_6087);
and U6667 (N_6667,N_6036,N_5832);
and U6668 (N_6668,N_6365,N_5763);
or U6669 (N_6669,N_5996,N_5903);
and U6670 (N_6670,N_5667,N_5609);
and U6671 (N_6671,N_5774,N_6275);
nor U6672 (N_6672,N_5675,N_6303);
or U6673 (N_6673,N_6031,N_5692);
nand U6674 (N_6674,N_6006,N_5766);
and U6675 (N_6675,N_5746,N_5693);
nand U6676 (N_6676,N_5687,N_5710);
and U6677 (N_6677,N_5863,N_5858);
nand U6678 (N_6678,N_6278,N_6245);
nor U6679 (N_6679,N_6317,N_6379);
and U6680 (N_6680,N_5677,N_6183);
nor U6681 (N_6681,N_5876,N_6366);
nor U6682 (N_6682,N_6009,N_5744);
or U6683 (N_6683,N_5792,N_5769);
nor U6684 (N_6684,N_6154,N_6012);
nor U6685 (N_6685,N_6216,N_5827);
xor U6686 (N_6686,N_5707,N_5610);
nand U6687 (N_6687,N_6394,N_5735);
and U6688 (N_6688,N_6092,N_6262);
nand U6689 (N_6689,N_6393,N_5654);
and U6690 (N_6690,N_5825,N_6181);
or U6691 (N_6691,N_6221,N_5982);
xor U6692 (N_6692,N_5628,N_6239);
nor U6693 (N_6693,N_6290,N_5781);
xor U6694 (N_6694,N_5682,N_5980);
nand U6695 (N_6695,N_5714,N_6172);
or U6696 (N_6696,N_5655,N_5814);
and U6697 (N_6697,N_5922,N_6253);
xor U6698 (N_6698,N_5689,N_6056);
xor U6699 (N_6699,N_5657,N_5741);
and U6700 (N_6700,N_6203,N_6011);
xnor U6701 (N_6701,N_6307,N_5723);
xnor U6702 (N_6702,N_5649,N_6293);
and U6703 (N_6703,N_6077,N_6100);
xor U6704 (N_6704,N_6291,N_6112);
nor U6705 (N_6705,N_6108,N_6295);
nand U6706 (N_6706,N_5839,N_6053);
nor U6707 (N_6707,N_6338,N_6179);
and U6708 (N_6708,N_5697,N_6045);
xnor U6709 (N_6709,N_5957,N_5868);
nand U6710 (N_6710,N_6167,N_5951);
and U6711 (N_6711,N_5999,N_5809);
nor U6712 (N_6712,N_6248,N_6034);
and U6713 (N_6713,N_6186,N_5831);
nor U6714 (N_6714,N_6099,N_6199);
nor U6715 (N_6715,N_6000,N_6105);
or U6716 (N_6716,N_5929,N_5949);
and U6717 (N_6717,N_6383,N_6162);
or U6718 (N_6718,N_5908,N_5647);
and U6719 (N_6719,N_5897,N_5953);
or U6720 (N_6720,N_5900,N_6106);
nand U6721 (N_6721,N_6062,N_6030);
or U6722 (N_6722,N_6201,N_6217);
nand U6723 (N_6723,N_5866,N_6089);
or U6724 (N_6724,N_5732,N_6138);
xnor U6725 (N_6725,N_5768,N_5739);
and U6726 (N_6726,N_5917,N_5937);
nor U6727 (N_6727,N_5698,N_6192);
xor U6728 (N_6728,N_5833,N_5892);
nor U6729 (N_6729,N_6222,N_6065);
nor U6730 (N_6730,N_6132,N_6060);
xnor U6731 (N_6731,N_5837,N_6251);
or U6732 (N_6732,N_5967,N_5887);
or U6733 (N_6733,N_6398,N_6386);
or U6734 (N_6734,N_5801,N_5966);
or U6735 (N_6735,N_6292,N_6169);
xnor U6736 (N_6736,N_6237,N_5691);
and U6737 (N_6737,N_6158,N_5923);
nor U6738 (N_6738,N_6204,N_5790);
or U6739 (N_6739,N_5873,N_5759);
and U6740 (N_6740,N_6084,N_6021);
and U6741 (N_6741,N_5927,N_6329);
nand U6742 (N_6742,N_5884,N_5694);
and U6743 (N_6743,N_6175,N_5856);
or U6744 (N_6744,N_6371,N_6286);
nand U6745 (N_6745,N_6330,N_6246);
nor U6746 (N_6746,N_5983,N_5643);
nor U6747 (N_6747,N_5600,N_5803);
or U6748 (N_6748,N_5824,N_6358);
xor U6749 (N_6749,N_5756,N_5843);
nor U6750 (N_6750,N_6159,N_6384);
nor U6751 (N_6751,N_6173,N_6083);
nor U6752 (N_6752,N_6029,N_6209);
or U6753 (N_6753,N_6323,N_5830);
nor U6754 (N_6754,N_5659,N_5828);
xnor U6755 (N_6755,N_5642,N_5619);
nand U6756 (N_6756,N_6346,N_6335);
and U6757 (N_6757,N_6047,N_6283);
and U6758 (N_6758,N_5625,N_5656);
and U6759 (N_6759,N_5879,N_6230);
nand U6760 (N_6760,N_5985,N_5932);
or U6761 (N_6761,N_6015,N_6232);
nor U6762 (N_6762,N_6336,N_6007);
or U6763 (N_6763,N_6001,N_6397);
and U6764 (N_6764,N_5673,N_6074);
and U6765 (N_6765,N_6174,N_5880);
and U6766 (N_6766,N_5938,N_5849);
and U6767 (N_6767,N_5624,N_6284);
or U6768 (N_6768,N_6022,N_6388);
or U6769 (N_6769,N_5894,N_5782);
and U6770 (N_6770,N_6227,N_6168);
nand U6771 (N_6771,N_5990,N_5810);
and U6772 (N_6772,N_6200,N_6150);
or U6773 (N_6773,N_6395,N_5808);
nand U6774 (N_6774,N_6215,N_6355);
nand U6775 (N_6775,N_5993,N_6250);
or U6776 (N_6776,N_5631,N_5926);
and U6777 (N_6777,N_6354,N_6198);
xnor U6778 (N_6778,N_5855,N_6300);
nand U6779 (N_6779,N_5712,N_6019);
xnor U6780 (N_6780,N_5901,N_6327);
nand U6781 (N_6781,N_5669,N_5819);
nand U6782 (N_6782,N_6325,N_5904);
nand U6783 (N_6783,N_5821,N_6399);
xnor U6784 (N_6784,N_5711,N_6096);
and U6785 (N_6785,N_6068,N_6191);
xor U6786 (N_6786,N_6147,N_5881);
and U6787 (N_6787,N_6078,N_6050);
or U6788 (N_6788,N_6051,N_6107);
xnor U6789 (N_6789,N_6306,N_6342);
xnor U6790 (N_6790,N_5800,N_5943);
nand U6791 (N_6791,N_5778,N_5777);
xor U6792 (N_6792,N_6382,N_6182);
nand U6793 (N_6793,N_5944,N_6119);
or U6794 (N_6794,N_5650,N_5680);
xnor U6795 (N_6795,N_6086,N_6309);
xnor U6796 (N_6796,N_6389,N_6027);
nand U6797 (N_6797,N_6170,N_5785);
and U6798 (N_6798,N_5896,N_5683);
nor U6799 (N_6799,N_5718,N_5681);
xor U6800 (N_6800,N_6150,N_5977);
nand U6801 (N_6801,N_5822,N_5890);
nand U6802 (N_6802,N_6313,N_6310);
nor U6803 (N_6803,N_5780,N_5952);
or U6804 (N_6804,N_5775,N_6255);
and U6805 (N_6805,N_6045,N_5801);
nand U6806 (N_6806,N_6160,N_5874);
or U6807 (N_6807,N_6023,N_5985);
nor U6808 (N_6808,N_5704,N_5622);
nand U6809 (N_6809,N_5919,N_5828);
or U6810 (N_6810,N_5723,N_5619);
nand U6811 (N_6811,N_6183,N_6033);
nand U6812 (N_6812,N_5833,N_6160);
nand U6813 (N_6813,N_5928,N_6389);
nand U6814 (N_6814,N_6345,N_5682);
xor U6815 (N_6815,N_6309,N_5728);
nand U6816 (N_6816,N_6208,N_5971);
nor U6817 (N_6817,N_5610,N_5711);
and U6818 (N_6818,N_6346,N_6001);
nand U6819 (N_6819,N_5918,N_6260);
and U6820 (N_6820,N_6298,N_6073);
xor U6821 (N_6821,N_5861,N_6382);
or U6822 (N_6822,N_6142,N_5890);
xnor U6823 (N_6823,N_5675,N_6259);
nand U6824 (N_6824,N_6295,N_5678);
or U6825 (N_6825,N_6236,N_5745);
xnor U6826 (N_6826,N_6160,N_6048);
and U6827 (N_6827,N_6030,N_5840);
xor U6828 (N_6828,N_5724,N_6256);
xnor U6829 (N_6829,N_6203,N_6212);
xnor U6830 (N_6830,N_5831,N_6361);
or U6831 (N_6831,N_5625,N_5818);
or U6832 (N_6832,N_5691,N_6073);
or U6833 (N_6833,N_5960,N_6082);
xor U6834 (N_6834,N_5618,N_6023);
nand U6835 (N_6835,N_5905,N_5841);
xnor U6836 (N_6836,N_5979,N_5981);
nor U6837 (N_6837,N_6111,N_6228);
or U6838 (N_6838,N_6375,N_5800);
and U6839 (N_6839,N_6248,N_6251);
xor U6840 (N_6840,N_6371,N_6229);
or U6841 (N_6841,N_6392,N_5616);
or U6842 (N_6842,N_6216,N_6293);
nand U6843 (N_6843,N_6171,N_6254);
xnor U6844 (N_6844,N_5756,N_6179);
nand U6845 (N_6845,N_6121,N_6264);
nand U6846 (N_6846,N_5638,N_6210);
xor U6847 (N_6847,N_6370,N_6024);
or U6848 (N_6848,N_6295,N_6385);
or U6849 (N_6849,N_5693,N_6026);
xnor U6850 (N_6850,N_6067,N_6269);
nor U6851 (N_6851,N_6369,N_6140);
xor U6852 (N_6852,N_5642,N_6264);
nor U6853 (N_6853,N_5959,N_5874);
nand U6854 (N_6854,N_6297,N_6301);
nand U6855 (N_6855,N_6215,N_5764);
nand U6856 (N_6856,N_6038,N_6142);
nor U6857 (N_6857,N_6168,N_6358);
or U6858 (N_6858,N_6006,N_6214);
or U6859 (N_6859,N_5628,N_6027);
xor U6860 (N_6860,N_5912,N_6226);
and U6861 (N_6861,N_5717,N_6133);
xnor U6862 (N_6862,N_6169,N_6063);
nand U6863 (N_6863,N_5795,N_6244);
xnor U6864 (N_6864,N_6322,N_6188);
or U6865 (N_6865,N_6215,N_5980);
or U6866 (N_6866,N_6383,N_5911);
and U6867 (N_6867,N_6034,N_5611);
nor U6868 (N_6868,N_5983,N_6059);
and U6869 (N_6869,N_6132,N_5677);
or U6870 (N_6870,N_5902,N_6292);
or U6871 (N_6871,N_5628,N_6083);
nor U6872 (N_6872,N_5629,N_5942);
nor U6873 (N_6873,N_5649,N_6371);
nand U6874 (N_6874,N_5654,N_6029);
nand U6875 (N_6875,N_6193,N_6099);
or U6876 (N_6876,N_5844,N_6016);
or U6877 (N_6877,N_6226,N_6004);
xnor U6878 (N_6878,N_6127,N_5625);
and U6879 (N_6879,N_6243,N_6359);
nor U6880 (N_6880,N_6050,N_5711);
xnor U6881 (N_6881,N_5847,N_5845);
nand U6882 (N_6882,N_6168,N_5778);
and U6883 (N_6883,N_6139,N_6088);
or U6884 (N_6884,N_5703,N_6131);
nor U6885 (N_6885,N_6143,N_6394);
or U6886 (N_6886,N_5677,N_5851);
or U6887 (N_6887,N_6362,N_6090);
nor U6888 (N_6888,N_6358,N_6076);
nor U6889 (N_6889,N_5885,N_5749);
nor U6890 (N_6890,N_5768,N_5730);
xor U6891 (N_6891,N_6258,N_5950);
or U6892 (N_6892,N_6207,N_6000);
nor U6893 (N_6893,N_5703,N_5931);
xnor U6894 (N_6894,N_5615,N_6294);
xnor U6895 (N_6895,N_6118,N_6184);
or U6896 (N_6896,N_6153,N_6145);
or U6897 (N_6897,N_6175,N_5838);
and U6898 (N_6898,N_5849,N_6207);
nor U6899 (N_6899,N_5912,N_5995);
and U6900 (N_6900,N_5969,N_6150);
xnor U6901 (N_6901,N_5738,N_5874);
nor U6902 (N_6902,N_6272,N_5677);
and U6903 (N_6903,N_5814,N_6075);
nor U6904 (N_6904,N_6296,N_6177);
nand U6905 (N_6905,N_5745,N_6304);
nor U6906 (N_6906,N_5748,N_5647);
or U6907 (N_6907,N_5960,N_5985);
xor U6908 (N_6908,N_5623,N_6067);
or U6909 (N_6909,N_6025,N_5643);
nor U6910 (N_6910,N_5760,N_6075);
nor U6911 (N_6911,N_6264,N_6148);
and U6912 (N_6912,N_5977,N_6241);
nor U6913 (N_6913,N_6150,N_6201);
or U6914 (N_6914,N_6178,N_5693);
or U6915 (N_6915,N_6289,N_5913);
and U6916 (N_6916,N_6252,N_6065);
xor U6917 (N_6917,N_5624,N_5626);
nor U6918 (N_6918,N_6202,N_5889);
nand U6919 (N_6919,N_5627,N_5734);
nand U6920 (N_6920,N_6006,N_5721);
xnor U6921 (N_6921,N_5952,N_5869);
and U6922 (N_6922,N_6157,N_5600);
nand U6923 (N_6923,N_5805,N_5912);
and U6924 (N_6924,N_6127,N_6363);
nand U6925 (N_6925,N_5711,N_5624);
or U6926 (N_6926,N_6311,N_6165);
nand U6927 (N_6927,N_6392,N_5724);
or U6928 (N_6928,N_6324,N_6245);
nand U6929 (N_6929,N_5602,N_5673);
and U6930 (N_6930,N_5613,N_5638);
and U6931 (N_6931,N_6331,N_5847);
xor U6932 (N_6932,N_5635,N_6245);
nand U6933 (N_6933,N_6046,N_6322);
nor U6934 (N_6934,N_6165,N_5790);
nand U6935 (N_6935,N_6302,N_6258);
xnor U6936 (N_6936,N_5777,N_5961);
or U6937 (N_6937,N_5790,N_6133);
nor U6938 (N_6938,N_5837,N_6271);
or U6939 (N_6939,N_6046,N_5987);
nand U6940 (N_6940,N_5694,N_5873);
xnor U6941 (N_6941,N_5855,N_6121);
nand U6942 (N_6942,N_6094,N_6366);
xor U6943 (N_6943,N_5933,N_5859);
nor U6944 (N_6944,N_6163,N_6274);
and U6945 (N_6945,N_6034,N_6209);
xnor U6946 (N_6946,N_6195,N_6378);
or U6947 (N_6947,N_6178,N_6279);
or U6948 (N_6948,N_6162,N_6258);
nand U6949 (N_6949,N_6116,N_6108);
xor U6950 (N_6950,N_5651,N_5662);
or U6951 (N_6951,N_5605,N_6082);
or U6952 (N_6952,N_6150,N_6313);
xnor U6953 (N_6953,N_5642,N_6116);
xor U6954 (N_6954,N_6061,N_6225);
and U6955 (N_6955,N_5820,N_5791);
and U6956 (N_6956,N_6270,N_6085);
or U6957 (N_6957,N_5761,N_5742);
and U6958 (N_6958,N_5727,N_6143);
nand U6959 (N_6959,N_6195,N_6010);
nand U6960 (N_6960,N_6371,N_5904);
nor U6961 (N_6961,N_6021,N_6097);
or U6962 (N_6962,N_5775,N_6175);
nor U6963 (N_6963,N_5993,N_5905);
and U6964 (N_6964,N_5894,N_6283);
nor U6965 (N_6965,N_6198,N_6011);
or U6966 (N_6966,N_6028,N_6143);
nor U6967 (N_6967,N_6056,N_5943);
nand U6968 (N_6968,N_6391,N_5997);
and U6969 (N_6969,N_6107,N_5837);
nor U6970 (N_6970,N_5788,N_6081);
and U6971 (N_6971,N_5733,N_5789);
or U6972 (N_6972,N_6364,N_6285);
or U6973 (N_6973,N_5884,N_6028);
and U6974 (N_6974,N_6056,N_5630);
nand U6975 (N_6975,N_5742,N_6295);
xnor U6976 (N_6976,N_5825,N_6190);
or U6977 (N_6977,N_6128,N_6324);
nor U6978 (N_6978,N_6088,N_5666);
and U6979 (N_6979,N_5771,N_5608);
xnor U6980 (N_6980,N_6140,N_5657);
nand U6981 (N_6981,N_6374,N_5898);
nand U6982 (N_6982,N_6295,N_5847);
nor U6983 (N_6983,N_6096,N_5884);
nor U6984 (N_6984,N_5670,N_6335);
xor U6985 (N_6985,N_6116,N_6151);
and U6986 (N_6986,N_5967,N_6167);
nor U6987 (N_6987,N_6199,N_5894);
nand U6988 (N_6988,N_5949,N_6262);
or U6989 (N_6989,N_5865,N_5849);
nand U6990 (N_6990,N_5758,N_5628);
nor U6991 (N_6991,N_6206,N_5937);
or U6992 (N_6992,N_5724,N_6356);
or U6993 (N_6993,N_5868,N_6080);
nor U6994 (N_6994,N_5602,N_5916);
and U6995 (N_6995,N_6107,N_6345);
xor U6996 (N_6996,N_6051,N_6335);
nor U6997 (N_6997,N_5612,N_5766);
nor U6998 (N_6998,N_5861,N_5663);
or U6999 (N_6999,N_6047,N_6326);
nor U7000 (N_7000,N_5846,N_6000);
xor U7001 (N_7001,N_6356,N_5725);
nor U7002 (N_7002,N_5613,N_5649);
or U7003 (N_7003,N_5988,N_6331);
nor U7004 (N_7004,N_5880,N_6143);
nand U7005 (N_7005,N_6029,N_6372);
and U7006 (N_7006,N_6259,N_6017);
or U7007 (N_7007,N_6028,N_6048);
and U7008 (N_7008,N_6291,N_6034);
or U7009 (N_7009,N_6396,N_6291);
nor U7010 (N_7010,N_6080,N_6309);
or U7011 (N_7011,N_5903,N_5666);
nand U7012 (N_7012,N_6165,N_5638);
and U7013 (N_7013,N_6238,N_6185);
xnor U7014 (N_7014,N_5752,N_6320);
and U7015 (N_7015,N_6057,N_5639);
nor U7016 (N_7016,N_5750,N_5941);
nand U7017 (N_7017,N_5737,N_6195);
nand U7018 (N_7018,N_6095,N_5842);
nor U7019 (N_7019,N_6028,N_6374);
nor U7020 (N_7020,N_5811,N_6134);
xor U7021 (N_7021,N_5927,N_6326);
nand U7022 (N_7022,N_6285,N_6042);
and U7023 (N_7023,N_5703,N_6135);
or U7024 (N_7024,N_6216,N_5658);
nand U7025 (N_7025,N_6073,N_5932);
xnor U7026 (N_7026,N_6143,N_5831);
nand U7027 (N_7027,N_6126,N_6076);
and U7028 (N_7028,N_5751,N_6119);
or U7029 (N_7029,N_6057,N_5904);
and U7030 (N_7030,N_5955,N_6050);
and U7031 (N_7031,N_5854,N_6055);
nor U7032 (N_7032,N_5827,N_5786);
or U7033 (N_7033,N_5646,N_5673);
nor U7034 (N_7034,N_5681,N_5816);
xor U7035 (N_7035,N_6108,N_6235);
nor U7036 (N_7036,N_5995,N_6082);
nor U7037 (N_7037,N_6309,N_6133);
nor U7038 (N_7038,N_5837,N_5746);
nor U7039 (N_7039,N_5699,N_5800);
nand U7040 (N_7040,N_6210,N_5602);
nand U7041 (N_7041,N_6185,N_5734);
and U7042 (N_7042,N_6168,N_6342);
and U7043 (N_7043,N_6227,N_6360);
nor U7044 (N_7044,N_6167,N_5979);
and U7045 (N_7045,N_6355,N_6398);
nor U7046 (N_7046,N_5998,N_5716);
xor U7047 (N_7047,N_6021,N_5665);
and U7048 (N_7048,N_5681,N_6336);
xnor U7049 (N_7049,N_5892,N_5746);
nor U7050 (N_7050,N_6172,N_6268);
or U7051 (N_7051,N_6128,N_6201);
nor U7052 (N_7052,N_5931,N_5812);
and U7053 (N_7053,N_6001,N_5794);
xnor U7054 (N_7054,N_6136,N_6326);
nor U7055 (N_7055,N_6168,N_5774);
and U7056 (N_7056,N_5851,N_5880);
nand U7057 (N_7057,N_5939,N_5749);
nor U7058 (N_7058,N_5789,N_5754);
xor U7059 (N_7059,N_6387,N_6207);
xnor U7060 (N_7060,N_6128,N_5727);
nor U7061 (N_7061,N_5987,N_5933);
nand U7062 (N_7062,N_5658,N_5739);
nand U7063 (N_7063,N_5675,N_5649);
xnor U7064 (N_7064,N_6192,N_5958);
and U7065 (N_7065,N_6022,N_5810);
nor U7066 (N_7066,N_5802,N_5635);
or U7067 (N_7067,N_6165,N_5729);
nor U7068 (N_7068,N_5997,N_5679);
or U7069 (N_7069,N_6046,N_6229);
and U7070 (N_7070,N_5904,N_6211);
and U7071 (N_7071,N_6320,N_5872);
xnor U7072 (N_7072,N_6299,N_6231);
xnor U7073 (N_7073,N_5751,N_6344);
and U7074 (N_7074,N_5814,N_6046);
and U7075 (N_7075,N_5954,N_6291);
and U7076 (N_7076,N_5967,N_5727);
nand U7077 (N_7077,N_6360,N_5665);
nor U7078 (N_7078,N_6215,N_6154);
nor U7079 (N_7079,N_6003,N_6072);
nor U7080 (N_7080,N_6383,N_6261);
nor U7081 (N_7081,N_5664,N_5926);
xor U7082 (N_7082,N_5807,N_5777);
xor U7083 (N_7083,N_6107,N_6372);
or U7084 (N_7084,N_5685,N_5871);
nor U7085 (N_7085,N_5708,N_6394);
xor U7086 (N_7086,N_6021,N_6207);
and U7087 (N_7087,N_5830,N_6243);
nand U7088 (N_7088,N_6386,N_6259);
xnor U7089 (N_7089,N_6198,N_6368);
xnor U7090 (N_7090,N_5944,N_6202);
xor U7091 (N_7091,N_6323,N_5996);
xnor U7092 (N_7092,N_6301,N_5901);
nand U7093 (N_7093,N_6112,N_5824);
xor U7094 (N_7094,N_5799,N_6395);
and U7095 (N_7095,N_6118,N_5836);
nor U7096 (N_7096,N_5936,N_6265);
nor U7097 (N_7097,N_5662,N_5785);
nand U7098 (N_7098,N_5766,N_5872);
xnor U7099 (N_7099,N_6319,N_6012);
nand U7100 (N_7100,N_6239,N_6061);
or U7101 (N_7101,N_6044,N_5687);
nand U7102 (N_7102,N_5770,N_6037);
nand U7103 (N_7103,N_6093,N_5926);
nand U7104 (N_7104,N_5644,N_6080);
xnor U7105 (N_7105,N_5629,N_6394);
nand U7106 (N_7106,N_5725,N_6273);
nand U7107 (N_7107,N_6126,N_6241);
and U7108 (N_7108,N_5754,N_6132);
nor U7109 (N_7109,N_5877,N_6073);
and U7110 (N_7110,N_5980,N_5616);
nor U7111 (N_7111,N_6124,N_6056);
nand U7112 (N_7112,N_5967,N_5680);
and U7113 (N_7113,N_6099,N_5714);
xor U7114 (N_7114,N_6153,N_5658);
nand U7115 (N_7115,N_5682,N_6315);
nand U7116 (N_7116,N_6136,N_5833);
or U7117 (N_7117,N_5899,N_6224);
and U7118 (N_7118,N_6342,N_6381);
and U7119 (N_7119,N_6397,N_5702);
nand U7120 (N_7120,N_5640,N_5639);
and U7121 (N_7121,N_5693,N_5630);
xnor U7122 (N_7122,N_6206,N_6361);
nand U7123 (N_7123,N_5765,N_6384);
or U7124 (N_7124,N_6369,N_5676);
xnor U7125 (N_7125,N_6174,N_5723);
nand U7126 (N_7126,N_6285,N_6188);
or U7127 (N_7127,N_5851,N_5755);
nor U7128 (N_7128,N_5851,N_5698);
xor U7129 (N_7129,N_6115,N_6347);
and U7130 (N_7130,N_5909,N_6259);
or U7131 (N_7131,N_5642,N_6102);
xnor U7132 (N_7132,N_6215,N_6390);
xnor U7133 (N_7133,N_6065,N_6040);
nand U7134 (N_7134,N_5641,N_6174);
and U7135 (N_7135,N_6242,N_5914);
and U7136 (N_7136,N_5974,N_5767);
xnor U7137 (N_7137,N_6015,N_6091);
and U7138 (N_7138,N_6066,N_6144);
xor U7139 (N_7139,N_6104,N_5852);
and U7140 (N_7140,N_6207,N_5684);
xor U7141 (N_7141,N_6327,N_5941);
nor U7142 (N_7142,N_5843,N_6231);
nand U7143 (N_7143,N_6017,N_5820);
and U7144 (N_7144,N_5606,N_6334);
nor U7145 (N_7145,N_5691,N_5976);
nor U7146 (N_7146,N_6264,N_6210);
or U7147 (N_7147,N_5690,N_5932);
nand U7148 (N_7148,N_5673,N_5984);
or U7149 (N_7149,N_5786,N_5880);
and U7150 (N_7150,N_6331,N_5710);
xor U7151 (N_7151,N_5933,N_5649);
and U7152 (N_7152,N_5724,N_6188);
nor U7153 (N_7153,N_6082,N_6015);
and U7154 (N_7154,N_6068,N_6176);
and U7155 (N_7155,N_5811,N_5802);
nor U7156 (N_7156,N_6006,N_5885);
xor U7157 (N_7157,N_5625,N_5700);
nand U7158 (N_7158,N_5888,N_6237);
nand U7159 (N_7159,N_5947,N_6334);
nand U7160 (N_7160,N_6173,N_5970);
or U7161 (N_7161,N_5665,N_5716);
nor U7162 (N_7162,N_5815,N_6355);
xnor U7163 (N_7163,N_6335,N_5701);
or U7164 (N_7164,N_5853,N_5722);
and U7165 (N_7165,N_5798,N_6100);
nor U7166 (N_7166,N_6049,N_5809);
or U7167 (N_7167,N_5888,N_6106);
xnor U7168 (N_7168,N_6237,N_5685);
nand U7169 (N_7169,N_5917,N_6142);
or U7170 (N_7170,N_6365,N_5607);
nor U7171 (N_7171,N_6079,N_5871);
nor U7172 (N_7172,N_5647,N_6102);
nor U7173 (N_7173,N_5654,N_5669);
or U7174 (N_7174,N_6265,N_6320);
nand U7175 (N_7175,N_5609,N_6311);
nor U7176 (N_7176,N_6026,N_6191);
or U7177 (N_7177,N_5689,N_5816);
or U7178 (N_7178,N_6158,N_5901);
xor U7179 (N_7179,N_5638,N_6298);
xor U7180 (N_7180,N_6160,N_6389);
xor U7181 (N_7181,N_5873,N_6305);
and U7182 (N_7182,N_6308,N_6340);
nor U7183 (N_7183,N_6132,N_6348);
nand U7184 (N_7184,N_5945,N_6020);
and U7185 (N_7185,N_5675,N_6354);
nor U7186 (N_7186,N_6379,N_5611);
or U7187 (N_7187,N_5805,N_6282);
xor U7188 (N_7188,N_5799,N_5646);
nand U7189 (N_7189,N_6311,N_6009);
or U7190 (N_7190,N_5996,N_6310);
nand U7191 (N_7191,N_5877,N_5815);
or U7192 (N_7192,N_5819,N_5968);
and U7193 (N_7193,N_5625,N_6398);
or U7194 (N_7194,N_6381,N_5990);
and U7195 (N_7195,N_5845,N_5631);
and U7196 (N_7196,N_5813,N_5881);
xnor U7197 (N_7197,N_5613,N_6207);
or U7198 (N_7198,N_5668,N_6041);
or U7199 (N_7199,N_6248,N_5815);
nand U7200 (N_7200,N_6628,N_6615);
nor U7201 (N_7201,N_7110,N_7191);
xnor U7202 (N_7202,N_6649,N_6881);
nor U7203 (N_7203,N_6608,N_6613);
xnor U7204 (N_7204,N_6620,N_6573);
xor U7205 (N_7205,N_7103,N_6859);
nor U7206 (N_7206,N_6557,N_6464);
xor U7207 (N_7207,N_6517,N_7144);
nand U7208 (N_7208,N_7097,N_6866);
nand U7209 (N_7209,N_7109,N_7112);
or U7210 (N_7210,N_6864,N_7133);
nand U7211 (N_7211,N_6463,N_6893);
nor U7212 (N_7212,N_7092,N_7107);
nor U7213 (N_7213,N_6883,N_6916);
xor U7214 (N_7214,N_6921,N_6880);
xnor U7215 (N_7215,N_6691,N_6872);
xnor U7216 (N_7216,N_6462,N_6721);
nor U7217 (N_7217,N_7094,N_7075);
or U7218 (N_7218,N_6842,N_6418);
or U7219 (N_7219,N_6946,N_6467);
nor U7220 (N_7220,N_6690,N_6824);
xor U7221 (N_7221,N_6572,N_6584);
nor U7222 (N_7222,N_6619,N_7132);
xnor U7223 (N_7223,N_6951,N_6475);
and U7224 (N_7224,N_6967,N_7083);
or U7225 (N_7225,N_6485,N_6840);
nor U7226 (N_7226,N_6739,N_6807);
or U7227 (N_7227,N_6993,N_7131);
and U7228 (N_7228,N_6565,N_6884);
or U7229 (N_7229,N_6830,N_6470);
and U7230 (N_7230,N_6940,N_6833);
xnor U7231 (N_7231,N_6855,N_6447);
nor U7232 (N_7232,N_6600,N_6978);
or U7233 (N_7233,N_7185,N_6897);
and U7234 (N_7234,N_6579,N_7042);
or U7235 (N_7235,N_6604,N_6844);
or U7236 (N_7236,N_6646,N_7048);
and U7237 (N_7237,N_6997,N_6641);
xor U7238 (N_7238,N_6862,N_6795);
nor U7239 (N_7239,N_6705,N_6427);
nand U7240 (N_7240,N_6704,N_6732);
xor U7241 (N_7241,N_6480,N_7057);
nor U7242 (N_7242,N_6537,N_6849);
nand U7243 (N_7243,N_6914,N_6644);
nand U7244 (N_7244,N_6466,N_6488);
xor U7245 (N_7245,N_6570,N_6626);
and U7246 (N_7246,N_6495,N_7179);
nor U7247 (N_7247,N_6610,N_7157);
nor U7248 (N_7248,N_6607,N_6818);
or U7249 (N_7249,N_7152,N_6931);
and U7250 (N_7250,N_7050,N_6758);
or U7251 (N_7251,N_6813,N_7079);
xnor U7252 (N_7252,N_7044,N_6785);
and U7253 (N_7253,N_6827,N_6460);
nand U7254 (N_7254,N_6798,N_6524);
and U7255 (N_7255,N_6472,N_6509);
nor U7256 (N_7256,N_6853,N_6635);
nand U7257 (N_7257,N_6558,N_7165);
xnor U7258 (N_7258,N_6918,N_6532);
nand U7259 (N_7259,N_6449,N_6531);
xor U7260 (N_7260,N_6973,N_6773);
and U7261 (N_7261,N_6576,N_6507);
nand U7262 (N_7262,N_6599,N_6834);
and U7263 (N_7263,N_6887,N_6432);
xnor U7264 (N_7264,N_7064,N_7020);
xor U7265 (N_7265,N_6678,N_6622);
xnor U7266 (N_7266,N_7025,N_6643);
nand U7267 (N_7267,N_6708,N_6968);
xor U7268 (N_7268,N_6400,N_7003);
and U7269 (N_7269,N_6774,N_7125);
nand U7270 (N_7270,N_7062,N_6976);
nor U7271 (N_7271,N_6805,N_7188);
or U7272 (N_7272,N_6982,N_6920);
nor U7273 (N_7273,N_7095,N_6696);
nor U7274 (N_7274,N_6766,N_6820);
nor U7275 (N_7275,N_7076,N_6603);
and U7276 (N_7276,N_7046,N_7136);
nor U7277 (N_7277,N_6498,N_6850);
nand U7278 (N_7278,N_7195,N_7001);
or U7279 (N_7279,N_6679,N_7181);
or U7280 (N_7280,N_7164,N_6601);
and U7281 (N_7281,N_6910,N_6979);
or U7282 (N_7282,N_6438,N_6631);
xnor U7283 (N_7283,N_6856,N_6896);
and U7284 (N_7284,N_6984,N_6542);
nand U7285 (N_7285,N_6926,N_6806);
nor U7286 (N_7286,N_6776,N_6444);
and U7287 (N_7287,N_7186,N_7105);
xor U7288 (N_7288,N_6523,N_6593);
xor U7289 (N_7289,N_6858,N_6456);
nor U7290 (N_7290,N_6753,N_6754);
nand U7291 (N_7291,N_6508,N_7128);
xnor U7292 (N_7292,N_7073,N_7060);
xnor U7293 (N_7293,N_6535,N_6494);
xor U7294 (N_7294,N_6487,N_7069);
and U7295 (N_7295,N_6411,N_6404);
nor U7296 (N_7296,N_7032,N_6421);
and U7297 (N_7297,N_6898,N_6836);
nor U7298 (N_7298,N_7016,N_7047);
or U7299 (N_7299,N_7187,N_6663);
or U7300 (N_7300,N_6602,N_6783);
or U7301 (N_7301,N_6950,N_7034);
xor U7302 (N_7302,N_7161,N_6623);
or U7303 (N_7303,N_6734,N_7040);
and U7304 (N_7304,N_7056,N_6782);
nor U7305 (N_7305,N_6762,N_6426);
or U7306 (N_7306,N_7124,N_6415);
or U7307 (N_7307,N_6406,N_6919);
nor U7308 (N_7308,N_7027,N_6983);
nor U7309 (N_7309,N_6408,N_6769);
or U7310 (N_7310,N_6668,N_6895);
xor U7311 (N_7311,N_6781,N_6865);
and U7312 (N_7312,N_6571,N_6788);
nor U7313 (N_7313,N_6716,N_7081);
and U7314 (N_7314,N_7013,N_6902);
nand U7315 (N_7315,N_6471,N_6761);
and U7316 (N_7316,N_7146,N_6760);
nand U7317 (N_7317,N_6666,N_6657);
nand U7318 (N_7318,N_6825,N_6845);
nor U7319 (N_7319,N_7119,N_6787);
xor U7320 (N_7320,N_6709,N_6917);
or U7321 (N_7321,N_6639,N_6402);
nand U7322 (N_7322,N_6733,N_6515);
nor U7323 (N_7323,N_6465,N_7134);
nand U7324 (N_7324,N_6980,N_6430);
and U7325 (N_7325,N_6727,N_6459);
and U7326 (N_7326,N_6803,N_6424);
and U7327 (N_7327,N_6491,N_7160);
xnor U7328 (N_7328,N_6837,N_6656);
nor U7329 (N_7329,N_6715,N_7054);
xnor U7330 (N_7330,N_7104,N_6549);
and U7331 (N_7331,N_6652,N_6520);
or U7332 (N_7332,N_6687,N_7170);
nor U7333 (N_7333,N_6930,N_6729);
and U7334 (N_7334,N_6777,N_6676);
xnor U7335 (N_7335,N_6752,N_7190);
and U7336 (N_7336,N_6768,N_6790);
nor U7337 (N_7337,N_6501,N_6786);
xor U7338 (N_7338,N_6497,N_6545);
nor U7339 (N_7339,N_6843,N_6922);
and U7340 (N_7340,N_7036,N_7051);
xnor U7341 (N_7341,N_7078,N_7087);
and U7342 (N_7342,N_6403,N_6975);
nor U7343 (N_7343,N_6838,N_7114);
or U7344 (N_7344,N_6992,N_6736);
and U7345 (N_7345,N_6547,N_6744);
nor U7346 (N_7346,N_7033,N_7116);
or U7347 (N_7347,N_6775,N_7140);
xor U7348 (N_7348,N_6701,N_6892);
or U7349 (N_7349,N_6530,N_7150);
xnor U7350 (N_7350,N_6550,N_6693);
nand U7351 (N_7351,N_6900,N_6672);
or U7352 (N_7352,N_7172,N_6913);
or U7353 (N_7353,N_6680,N_6953);
nor U7354 (N_7354,N_7012,N_6852);
or U7355 (N_7355,N_6698,N_7007);
xor U7356 (N_7356,N_7118,N_6492);
xor U7357 (N_7357,N_6453,N_6924);
and U7358 (N_7358,N_6546,N_6737);
and U7359 (N_7359,N_6413,N_7014);
and U7360 (N_7360,N_6442,N_6699);
xor U7361 (N_7361,N_7102,N_6955);
nand U7362 (N_7362,N_6987,N_7030);
or U7363 (N_7363,N_7077,N_6712);
xnor U7364 (N_7364,N_6630,N_6407);
nor U7365 (N_7365,N_6958,N_6743);
xor U7366 (N_7366,N_6948,N_6479);
nand U7367 (N_7367,N_6645,N_7002);
and U7368 (N_7368,N_6710,N_6934);
nand U7369 (N_7369,N_7167,N_6741);
nand U7370 (N_7370,N_6909,N_6586);
xor U7371 (N_7371,N_7065,N_7082);
or U7372 (N_7372,N_6510,N_7085);
nor U7373 (N_7373,N_7158,N_6792);
or U7374 (N_7374,N_6452,N_6677);
xor U7375 (N_7375,N_6594,N_6539);
nand U7376 (N_7376,N_7184,N_6969);
and U7377 (N_7377,N_7096,N_6817);
or U7378 (N_7378,N_6738,N_6685);
xor U7379 (N_7379,N_7139,N_6637);
nand U7380 (N_7380,N_6405,N_7121);
nand U7381 (N_7381,N_6560,N_7021);
xor U7382 (N_7382,N_6814,N_6629);
nand U7383 (N_7383,N_6885,N_6714);
xnor U7384 (N_7384,N_6526,N_7010);
and U7385 (N_7385,N_6740,N_7089);
nor U7386 (N_7386,N_6999,N_6533);
nor U7387 (N_7387,N_6966,N_6580);
nand U7388 (N_7388,N_7072,N_7059);
xnor U7389 (N_7389,N_6867,N_7198);
or U7390 (N_7390,N_6443,N_6927);
nand U7391 (N_7391,N_6911,N_6835);
nand U7392 (N_7392,N_7023,N_6730);
or U7393 (N_7393,N_7189,N_6717);
and U7394 (N_7394,N_6823,N_6832);
nand U7395 (N_7395,N_6901,N_7178);
nor U7396 (N_7396,N_6938,N_6974);
nor U7397 (N_7397,N_6642,N_6500);
and U7398 (N_7398,N_6731,N_7196);
xor U7399 (N_7399,N_6454,N_6554);
nor U7400 (N_7400,N_7145,N_6863);
or U7401 (N_7401,N_6534,N_7086);
nor U7402 (N_7402,N_6906,N_6611);
nor U7403 (N_7403,N_7074,N_6659);
nor U7404 (N_7404,N_6633,N_6912);
or U7405 (N_7405,N_6784,N_7008);
nor U7406 (N_7406,N_6990,N_6614);
xnor U7407 (N_7407,N_6527,N_6481);
nor U7408 (N_7408,N_6828,N_6561);
nor U7409 (N_7409,N_7005,N_7169);
and U7410 (N_7410,N_6821,N_7009);
or U7411 (N_7411,N_6949,N_7043);
nand U7412 (N_7412,N_7101,N_6871);
xnor U7413 (N_7413,N_6662,N_7045);
xnor U7414 (N_7414,N_6414,N_6860);
and U7415 (N_7415,N_6851,N_7006);
nand U7416 (N_7416,N_7156,N_7199);
or U7417 (N_7417,N_6625,N_6562);
xnor U7418 (N_7418,N_6578,N_7066);
and U7419 (N_7419,N_6985,N_6543);
nand U7420 (N_7420,N_7159,N_6707);
nand U7421 (N_7421,N_6961,N_6473);
nand U7422 (N_7422,N_6943,N_6634);
nand U7423 (N_7423,N_6582,N_6799);
and U7424 (N_7424,N_7163,N_7173);
and U7425 (N_7425,N_6723,N_6597);
or U7426 (N_7426,N_6700,N_6822);
or U7427 (N_7427,N_6640,N_6703);
nor U7428 (N_7428,N_6748,N_6932);
nand U7429 (N_7429,N_6915,N_6540);
nand U7430 (N_7430,N_6618,N_6812);
or U7431 (N_7431,N_6609,N_6410);
or U7432 (N_7432,N_6423,N_6875);
nor U7433 (N_7433,N_6962,N_6686);
xnor U7434 (N_7434,N_6746,N_6841);
and U7435 (N_7435,N_6559,N_6861);
nor U7436 (N_7436,N_6954,N_6496);
nor U7437 (N_7437,N_6991,N_6728);
nand U7438 (N_7438,N_6451,N_7084);
nor U7439 (N_7439,N_6477,N_6831);
nand U7440 (N_7440,N_7155,N_6907);
nand U7441 (N_7441,N_6998,N_6941);
xnor U7442 (N_7442,N_6857,N_6767);
xor U7443 (N_7443,N_6994,N_6638);
or U7444 (N_7444,N_7127,N_6942);
and U7445 (N_7445,N_7115,N_7123);
nand U7446 (N_7446,N_7068,N_6538);
or U7447 (N_7447,N_6409,N_7071);
nor U7448 (N_7448,N_6694,N_6811);
or U7449 (N_7449,N_6627,N_6720);
nor U7450 (N_7450,N_7100,N_6801);
nor U7451 (N_7451,N_6590,N_6725);
or U7452 (N_7452,N_6793,N_6870);
and U7453 (N_7453,N_6544,N_6702);
or U7454 (N_7454,N_6518,N_7004);
and U7455 (N_7455,N_6612,N_6484);
nand U7456 (N_7456,N_7183,N_6482);
xor U7457 (N_7457,N_6548,N_6879);
xor U7458 (N_7458,N_6598,N_6474);
nand U7459 (N_7459,N_6455,N_6890);
nor U7460 (N_7460,N_6566,N_6674);
xnor U7461 (N_7461,N_6905,N_6935);
nand U7462 (N_7462,N_6755,N_7049);
or U7463 (N_7463,N_7029,N_6493);
and U7464 (N_7464,N_7113,N_7018);
xor U7465 (N_7465,N_6660,N_6499);
nand U7466 (N_7466,N_7130,N_6574);
xor U7467 (N_7467,N_6996,N_6747);
nand U7468 (N_7468,N_7035,N_6970);
and U7469 (N_7469,N_6588,N_6947);
and U7470 (N_7470,N_7141,N_7015);
nor U7471 (N_7471,N_6742,N_6802);
or U7472 (N_7472,N_6468,N_6810);
or U7473 (N_7473,N_6711,N_7031);
and U7474 (N_7474,N_6563,N_6808);
xnor U7475 (N_7475,N_6461,N_7038);
xnor U7476 (N_7476,N_6536,N_6706);
and U7477 (N_7477,N_6756,N_6595);
or U7478 (N_7478,N_6891,N_6684);
xor U7479 (N_7479,N_6779,N_6908);
xor U7480 (N_7480,N_6431,N_6683);
nand U7481 (N_7481,N_6504,N_6511);
nand U7482 (N_7482,N_6995,N_6695);
or U7483 (N_7483,N_6726,N_7080);
nor U7484 (N_7484,N_7028,N_6416);
nor U7485 (N_7485,N_6819,N_6965);
and U7486 (N_7486,N_6529,N_6605);
or U7487 (N_7487,N_7166,N_6944);
or U7488 (N_7488,N_6718,N_6655);
and U7489 (N_7489,N_6401,N_6569);
or U7490 (N_7490,N_6555,N_7000);
nor U7491 (N_7491,N_6457,N_7149);
and U7492 (N_7492,N_6486,N_7168);
or U7493 (N_7493,N_6669,N_6959);
nand U7494 (N_7494,N_6688,N_6789);
and U7495 (N_7495,N_7019,N_6412);
xor U7496 (N_7496,N_6670,N_6809);
nand U7497 (N_7497,N_7192,N_7058);
nor U7498 (N_7498,N_6624,N_6521);
or U7499 (N_7499,N_6764,N_6616);
nor U7500 (N_7500,N_6878,N_6882);
or U7501 (N_7501,N_6437,N_7111);
nand U7502 (N_7502,N_7070,N_7148);
and U7503 (N_7503,N_7061,N_6724);
and U7504 (N_7504,N_6606,N_6689);
and U7505 (N_7505,N_6469,N_6757);
nor U7506 (N_7506,N_6770,N_7176);
nor U7507 (N_7507,N_6829,N_7171);
xor U7508 (N_7508,N_7129,N_6621);
or U7509 (N_7509,N_6815,N_7039);
or U7510 (N_7510,N_6750,N_6873);
or U7511 (N_7511,N_7180,N_6956);
nor U7512 (N_7512,N_6667,N_7098);
xor U7513 (N_7513,N_6957,N_6868);
and U7514 (N_7514,N_6854,N_7151);
or U7515 (N_7515,N_6681,N_6419);
xnor U7516 (N_7516,N_6682,N_7153);
nor U7517 (N_7517,N_6796,N_6771);
nand U7518 (N_7518,N_6876,N_6581);
and U7519 (N_7519,N_7138,N_6434);
nand U7520 (N_7520,N_6428,N_6651);
or U7521 (N_7521,N_6937,N_6847);
or U7522 (N_7522,N_6519,N_6433);
and U7523 (N_7523,N_6422,N_6977);
nand U7524 (N_7524,N_6636,N_7154);
or U7525 (N_7525,N_6505,N_6869);
nand U7526 (N_7526,N_6556,N_6928);
nor U7527 (N_7527,N_6513,N_6417);
and U7528 (N_7528,N_6525,N_6960);
or U7529 (N_7529,N_6440,N_6904);
nor U7530 (N_7530,N_6971,N_6516);
xor U7531 (N_7531,N_6441,N_6923);
and U7532 (N_7532,N_7037,N_6839);
xnor U7533 (N_7533,N_6502,N_6889);
or U7534 (N_7534,N_6528,N_7022);
nand U7535 (N_7535,N_7182,N_6583);
and U7536 (N_7536,N_6765,N_6506);
xor U7537 (N_7537,N_6745,N_6903);
xor U7538 (N_7538,N_7090,N_6661);
or U7539 (N_7539,N_7177,N_7106);
xor U7540 (N_7540,N_6617,N_6552);
xnor U7541 (N_7541,N_6425,N_7088);
nand U7542 (N_7542,N_6763,N_7122);
nor U7543 (N_7543,N_6650,N_6567);
xor U7544 (N_7544,N_6989,N_6591);
and U7545 (N_7545,N_6564,N_7174);
and U7546 (N_7546,N_6450,N_7108);
and U7547 (N_7547,N_7147,N_6436);
nand U7548 (N_7548,N_7197,N_7193);
and U7549 (N_7549,N_6791,N_6512);
xnor U7550 (N_7550,N_6816,N_6964);
nand U7551 (N_7551,N_6797,N_6489);
and U7552 (N_7552,N_6448,N_7162);
nand U7553 (N_7553,N_6963,N_6874);
nor U7554 (N_7554,N_6936,N_6587);
nand U7555 (N_7555,N_6772,N_6751);
nor U7556 (N_7556,N_6439,N_7142);
nor U7557 (N_7557,N_6503,N_7175);
nor U7558 (N_7558,N_6933,N_6899);
nor U7559 (N_7559,N_6490,N_6713);
nand U7560 (N_7560,N_6972,N_7143);
and U7561 (N_7561,N_6665,N_6551);
nand U7562 (N_7562,N_6848,N_7093);
and U7563 (N_7563,N_6420,N_6483);
and U7564 (N_7564,N_6719,N_6925);
nor U7565 (N_7565,N_6596,N_6804);
xnor U7566 (N_7566,N_6794,N_6648);
xnor U7567 (N_7567,N_6692,N_7017);
nand U7568 (N_7568,N_6671,N_6435);
nand U7569 (N_7569,N_7052,N_6780);
xor U7570 (N_7570,N_6826,N_7026);
nand U7571 (N_7571,N_6522,N_6585);
nand U7572 (N_7572,N_7099,N_7024);
nor U7573 (N_7573,N_6478,N_6514);
nor U7574 (N_7574,N_6986,N_6988);
or U7575 (N_7575,N_7126,N_6589);
and U7576 (N_7576,N_6981,N_6653);
nand U7577 (N_7577,N_6952,N_7041);
or U7578 (N_7578,N_6553,N_6945);
nand U7579 (N_7579,N_6673,N_6929);
nand U7580 (N_7580,N_6568,N_6575);
nand U7581 (N_7581,N_6664,N_6592);
nor U7582 (N_7582,N_7053,N_6429);
and U7583 (N_7583,N_6846,N_7137);
nor U7584 (N_7584,N_6735,N_6647);
and U7585 (N_7585,N_7055,N_6894);
nand U7586 (N_7586,N_6800,N_6697);
xnor U7587 (N_7587,N_6445,N_6446);
nor U7588 (N_7588,N_6759,N_6654);
nand U7589 (N_7589,N_6541,N_7011);
or U7590 (N_7590,N_6886,N_6577);
nand U7591 (N_7591,N_7117,N_6888);
xnor U7592 (N_7592,N_6476,N_6877);
nor U7593 (N_7593,N_7194,N_7091);
xor U7594 (N_7594,N_7135,N_7067);
nand U7595 (N_7595,N_6722,N_6675);
nand U7596 (N_7596,N_6658,N_7063);
xor U7597 (N_7597,N_6458,N_7120);
nor U7598 (N_7598,N_6749,N_6632);
nor U7599 (N_7599,N_6939,N_6778);
nor U7600 (N_7600,N_7109,N_6484);
nand U7601 (N_7601,N_6427,N_7188);
and U7602 (N_7602,N_7132,N_6636);
nor U7603 (N_7603,N_6601,N_6691);
and U7604 (N_7604,N_7113,N_6814);
nor U7605 (N_7605,N_7037,N_6675);
xor U7606 (N_7606,N_6819,N_7127);
and U7607 (N_7607,N_7048,N_7176);
and U7608 (N_7608,N_7079,N_7000);
xor U7609 (N_7609,N_6620,N_6642);
xor U7610 (N_7610,N_6475,N_6424);
nand U7611 (N_7611,N_6420,N_6904);
and U7612 (N_7612,N_7062,N_6635);
or U7613 (N_7613,N_6497,N_6849);
nor U7614 (N_7614,N_6693,N_6770);
nand U7615 (N_7615,N_6529,N_6714);
xor U7616 (N_7616,N_7139,N_6643);
and U7617 (N_7617,N_6972,N_6639);
nor U7618 (N_7618,N_7018,N_6751);
xor U7619 (N_7619,N_6856,N_6619);
and U7620 (N_7620,N_6810,N_7170);
and U7621 (N_7621,N_6847,N_6681);
or U7622 (N_7622,N_6904,N_6594);
nor U7623 (N_7623,N_6415,N_7185);
nand U7624 (N_7624,N_6983,N_6622);
or U7625 (N_7625,N_6459,N_6507);
or U7626 (N_7626,N_6532,N_6632);
and U7627 (N_7627,N_6922,N_6507);
xor U7628 (N_7628,N_6441,N_6717);
xnor U7629 (N_7629,N_7172,N_7043);
xor U7630 (N_7630,N_6754,N_7008);
nand U7631 (N_7631,N_6569,N_7058);
or U7632 (N_7632,N_7155,N_6781);
or U7633 (N_7633,N_6884,N_6901);
nand U7634 (N_7634,N_7154,N_6407);
nand U7635 (N_7635,N_6492,N_7085);
nor U7636 (N_7636,N_6963,N_7082);
nor U7637 (N_7637,N_6470,N_6720);
xor U7638 (N_7638,N_7184,N_6428);
nand U7639 (N_7639,N_6423,N_6438);
nor U7640 (N_7640,N_6957,N_6749);
or U7641 (N_7641,N_6443,N_6815);
nand U7642 (N_7642,N_6503,N_7100);
or U7643 (N_7643,N_7148,N_6642);
or U7644 (N_7644,N_7170,N_6516);
nand U7645 (N_7645,N_6571,N_6828);
and U7646 (N_7646,N_6484,N_6577);
nor U7647 (N_7647,N_6982,N_6984);
and U7648 (N_7648,N_6534,N_6719);
nor U7649 (N_7649,N_7068,N_7184);
or U7650 (N_7650,N_6938,N_6860);
and U7651 (N_7651,N_6705,N_7082);
and U7652 (N_7652,N_6684,N_7153);
nand U7653 (N_7653,N_6792,N_6695);
xnor U7654 (N_7654,N_6817,N_6813);
or U7655 (N_7655,N_6675,N_6685);
or U7656 (N_7656,N_6713,N_6907);
xnor U7657 (N_7657,N_7037,N_6666);
nand U7658 (N_7658,N_7028,N_6888);
or U7659 (N_7659,N_6416,N_6977);
nor U7660 (N_7660,N_6708,N_7116);
and U7661 (N_7661,N_6527,N_6648);
or U7662 (N_7662,N_6719,N_6667);
or U7663 (N_7663,N_6863,N_6496);
nand U7664 (N_7664,N_6656,N_7103);
and U7665 (N_7665,N_6542,N_6545);
or U7666 (N_7666,N_6486,N_6925);
nand U7667 (N_7667,N_7000,N_6574);
or U7668 (N_7668,N_6836,N_6654);
nor U7669 (N_7669,N_6403,N_6868);
xor U7670 (N_7670,N_6882,N_7160);
and U7671 (N_7671,N_6606,N_6440);
and U7672 (N_7672,N_7160,N_6893);
or U7673 (N_7673,N_6611,N_6984);
nand U7674 (N_7674,N_7008,N_7140);
nor U7675 (N_7675,N_6950,N_7075);
nand U7676 (N_7676,N_6652,N_6656);
nor U7677 (N_7677,N_6496,N_7161);
nor U7678 (N_7678,N_6568,N_6745);
or U7679 (N_7679,N_7023,N_6582);
or U7680 (N_7680,N_6824,N_6804);
and U7681 (N_7681,N_6913,N_6757);
nor U7682 (N_7682,N_6440,N_6599);
and U7683 (N_7683,N_7062,N_6480);
xnor U7684 (N_7684,N_6847,N_7089);
nand U7685 (N_7685,N_6862,N_6660);
and U7686 (N_7686,N_6820,N_6526);
nor U7687 (N_7687,N_7181,N_7172);
and U7688 (N_7688,N_6557,N_6534);
or U7689 (N_7689,N_6404,N_6655);
nor U7690 (N_7690,N_6566,N_6615);
xnor U7691 (N_7691,N_6955,N_6817);
and U7692 (N_7692,N_6865,N_6455);
nand U7693 (N_7693,N_6769,N_6960);
nor U7694 (N_7694,N_6691,N_7046);
and U7695 (N_7695,N_6932,N_6665);
nor U7696 (N_7696,N_7188,N_6405);
nand U7697 (N_7697,N_6612,N_6786);
nand U7698 (N_7698,N_6508,N_6883);
nand U7699 (N_7699,N_7072,N_6994);
or U7700 (N_7700,N_6503,N_6442);
nand U7701 (N_7701,N_6469,N_7002);
and U7702 (N_7702,N_6916,N_6549);
xnor U7703 (N_7703,N_6829,N_6592);
and U7704 (N_7704,N_7137,N_7184);
or U7705 (N_7705,N_6795,N_7126);
nand U7706 (N_7706,N_6821,N_6838);
nand U7707 (N_7707,N_6498,N_6409);
nor U7708 (N_7708,N_7009,N_6529);
xor U7709 (N_7709,N_6502,N_6424);
or U7710 (N_7710,N_6544,N_6931);
nor U7711 (N_7711,N_6968,N_7116);
nand U7712 (N_7712,N_7044,N_6870);
nor U7713 (N_7713,N_6797,N_6450);
nand U7714 (N_7714,N_7106,N_7154);
and U7715 (N_7715,N_6985,N_7075);
or U7716 (N_7716,N_6684,N_6922);
nor U7717 (N_7717,N_6571,N_7150);
nand U7718 (N_7718,N_6763,N_6406);
nand U7719 (N_7719,N_6961,N_6922);
xor U7720 (N_7720,N_7002,N_7133);
and U7721 (N_7721,N_6547,N_6475);
and U7722 (N_7722,N_6522,N_6747);
nor U7723 (N_7723,N_6798,N_6557);
nor U7724 (N_7724,N_6448,N_6511);
nand U7725 (N_7725,N_6815,N_6596);
nor U7726 (N_7726,N_6439,N_6459);
nor U7727 (N_7727,N_6471,N_6422);
xnor U7728 (N_7728,N_6491,N_6521);
nand U7729 (N_7729,N_7064,N_7172);
and U7730 (N_7730,N_6826,N_6738);
xnor U7731 (N_7731,N_6488,N_6944);
or U7732 (N_7732,N_6777,N_6786);
nor U7733 (N_7733,N_6877,N_6683);
xnor U7734 (N_7734,N_6519,N_6949);
and U7735 (N_7735,N_6616,N_6809);
and U7736 (N_7736,N_6875,N_6629);
nand U7737 (N_7737,N_6816,N_6576);
nor U7738 (N_7738,N_6418,N_6634);
and U7739 (N_7739,N_6769,N_6701);
and U7740 (N_7740,N_6875,N_6692);
nor U7741 (N_7741,N_6552,N_6607);
nand U7742 (N_7742,N_7098,N_6999);
nor U7743 (N_7743,N_7002,N_6818);
nor U7744 (N_7744,N_6760,N_7086);
xnor U7745 (N_7745,N_6780,N_6593);
or U7746 (N_7746,N_6719,N_6873);
and U7747 (N_7747,N_7157,N_6562);
or U7748 (N_7748,N_7129,N_6802);
xor U7749 (N_7749,N_6864,N_6661);
nand U7750 (N_7750,N_6619,N_6702);
xor U7751 (N_7751,N_6882,N_6448);
nand U7752 (N_7752,N_7079,N_6570);
nor U7753 (N_7753,N_6885,N_7175);
and U7754 (N_7754,N_6952,N_6460);
xor U7755 (N_7755,N_7141,N_6872);
and U7756 (N_7756,N_6499,N_6908);
or U7757 (N_7757,N_6705,N_6784);
and U7758 (N_7758,N_6716,N_7094);
nor U7759 (N_7759,N_6426,N_6407);
nor U7760 (N_7760,N_7125,N_7011);
or U7761 (N_7761,N_6695,N_6768);
and U7762 (N_7762,N_6948,N_6769);
nor U7763 (N_7763,N_6823,N_6485);
nor U7764 (N_7764,N_7195,N_7076);
and U7765 (N_7765,N_7168,N_6521);
xnor U7766 (N_7766,N_6730,N_7106);
xor U7767 (N_7767,N_6458,N_6936);
nor U7768 (N_7768,N_6757,N_6607);
nor U7769 (N_7769,N_6902,N_7040);
and U7770 (N_7770,N_6894,N_6535);
nor U7771 (N_7771,N_6530,N_6488);
xnor U7772 (N_7772,N_7018,N_6927);
xor U7773 (N_7773,N_6611,N_6681);
or U7774 (N_7774,N_6820,N_6706);
nand U7775 (N_7775,N_7103,N_6891);
nor U7776 (N_7776,N_6886,N_7035);
xor U7777 (N_7777,N_6745,N_6681);
or U7778 (N_7778,N_7129,N_7141);
nand U7779 (N_7779,N_7019,N_6935);
and U7780 (N_7780,N_6898,N_6576);
or U7781 (N_7781,N_7136,N_6694);
and U7782 (N_7782,N_6418,N_6813);
nand U7783 (N_7783,N_7070,N_6775);
nand U7784 (N_7784,N_6940,N_6737);
nand U7785 (N_7785,N_6906,N_7028);
nor U7786 (N_7786,N_7069,N_6965);
xnor U7787 (N_7787,N_6955,N_6628);
nor U7788 (N_7788,N_6436,N_6806);
nand U7789 (N_7789,N_6690,N_7195);
and U7790 (N_7790,N_7048,N_6622);
nand U7791 (N_7791,N_6561,N_7141);
xor U7792 (N_7792,N_6616,N_6846);
nand U7793 (N_7793,N_6790,N_6877);
and U7794 (N_7794,N_6765,N_6467);
nor U7795 (N_7795,N_6407,N_7146);
and U7796 (N_7796,N_7046,N_6633);
xnor U7797 (N_7797,N_6924,N_6776);
nor U7798 (N_7798,N_6554,N_6537);
or U7799 (N_7799,N_6532,N_6989);
or U7800 (N_7800,N_6944,N_7127);
nor U7801 (N_7801,N_6719,N_6454);
nor U7802 (N_7802,N_7123,N_7135);
nor U7803 (N_7803,N_6427,N_6779);
nand U7804 (N_7804,N_6906,N_6595);
or U7805 (N_7805,N_6811,N_7114);
nand U7806 (N_7806,N_6422,N_6650);
nor U7807 (N_7807,N_6773,N_6735);
and U7808 (N_7808,N_6852,N_6716);
and U7809 (N_7809,N_6806,N_6512);
and U7810 (N_7810,N_6835,N_6594);
nor U7811 (N_7811,N_6875,N_6776);
or U7812 (N_7812,N_6684,N_6633);
and U7813 (N_7813,N_6907,N_7144);
xor U7814 (N_7814,N_7119,N_6921);
or U7815 (N_7815,N_6984,N_7054);
nor U7816 (N_7816,N_6655,N_6763);
xor U7817 (N_7817,N_6909,N_6955);
nand U7818 (N_7818,N_7051,N_6409);
or U7819 (N_7819,N_6852,N_6459);
nand U7820 (N_7820,N_7140,N_6848);
nor U7821 (N_7821,N_7047,N_6551);
xor U7822 (N_7822,N_6964,N_6563);
nor U7823 (N_7823,N_6842,N_6910);
nand U7824 (N_7824,N_6673,N_6714);
nand U7825 (N_7825,N_6418,N_6526);
nor U7826 (N_7826,N_6658,N_7124);
xor U7827 (N_7827,N_7157,N_6802);
nor U7828 (N_7828,N_6876,N_6704);
nor U7829 (N_7829,N_6860,N_6842);
nand U7830 (N_7830,N_6581,N_7085);
and U7831 (N_7831,N_6567,N_6632);
and U7832 (N_7832,N_6772,N_6877);
nor U7833 (N_7833,N_7014,N_6690);
nand U7834 (N_7834,N_6719,N_6537);
nand U7835 (N_7835,N_6768,N_6834);
xnor U7836 (N_7836,N_7173,N_6998);
or U7837 (N_7837,N_6778,N_6710);
nand U7838 (N_7838,N_6978,N_6817);
nand U7839 (N_7839,N_6562,N_7163);
xor U7840 (N_7840,N_6772,N_6828);
and U7841 (N_7841,N_6746,N_7138);
and U7842 (N_7842,N_7090,N_6906);
xor U7843 (N_7843,N_7025,N_6823);
and U7844 (N_7844,N_6501,N_6486);
xor U7845 (N_7845,N_6633,N_7131);
or U7846 (N_7846,N_6975,N_6589);
nor U7847 (N_7847,N_6458,N_6559);
xnor U7848 (N_7848,N_7064,N_7132);
nor U7849 (N_7849,N_6536,N_6682);
nand U7850 (N_7850,N_6766,N_6797);
and U7851 (N_7851,N_6659,N_7156);
nand U7852 (N_7852,N_6975,N_6504);
nand U7853 (N_7853,N_6831,N_6819);
xnor U7854 (N_7854,N_6511,N_6865);
nand U7855 (N_7855,N_7117,N_6403);
xnor U7856 (N_7856,N_6947,N_6484);
nor U7857 (N_7857,N_7140,N_6452);
nand U7858 (N_7858,N_6922,N_6963);
nand U7859 (N_7859,N_7120,N_6960);
nand U7860 (N_7860,N_6419,N_6414);
nand U7861 (N_7861,N_6877,N_7039);
or U7862 (N_7862,N_6677,N_6919);
nand U7863 (N_7863,N_7081,N_7138);
nand U7864 (N_7864,N_6946,N_6975);
nand U7865 (N_7865,N_6602,N_6924);
nand U7866 (N_7866,N_6498,N_7154);
nor U7867 (N_7867,N_6552,N_6923);
nor U7868 (N_7868,N_6972,N_7106);
xnor U7869 (N_7869,N_7170,N_6413);
or U7870 (N_7870,N_6977,N_6710);
and U7871 (N_7871,N_6408,N_6773);
nor U7872 (N_7872,N_6411,N_6680);
nand U7873 (N_7873,N_6467,N_7080);
xnor U7874 (N_7874,N_7145,N_6823);
nor U7875 (N_7875,N_7191,N_6734);
nor U7876 (N_7876,N_6639,N_6664);
nand U7877 (N_7877,N_7000,N_6940);
nor U7878 (N_7878,N_7184,N_6856);
xnor U7879 (N_7879,N_6621,N_6561);
nand U7880 (N_7880,N_6467,N_6561);
and U7881 (N_7881,N_6751,N_6637);
and U7882 (N_7882,N_6707,N_6661);
xor U7883 (N_7883,N_6771,N_7126);
nand U7884 (N_7884,N_6680,N_6947);
nand U7885 (N_7885,N_7019,N_6637);
and U7886 (N_7886,N_6693,N_6494);
nor U7887 (N_7887,N_6615,N_6536);
or U7888 (N_7888,N_7194,N_6425);
xor U7889 (N_7889,N_6908,N_6937);
or U7890 (N_7890,N_7063,N_7130);
or U7891 (N_7891,N_6469,N_7037);
or U7892 (N_7892,N_6941,N_7017);
and U7893 (N_7893,N_6528,N_6564);
nor U7894 (N_7894,N_6846,N_7022);
xor U7895 (N_7895,N_7043,N_6749);
and U7896 (N_7896,N_6686,N_7041);
nor U7897 (N_7897,N_6614,N_6513);
or U7898 (N_7898,N_6538,N_7057);
xnor U7899 (N_7899,N_6552,N_7056);
xor U7900 (N_7900,N_7133,N_7081);
and U7901 (N_7901,N_7158,N_6722);
or U7902 (N_7902,N_6546,N_6749);
or U7903 (N_7903,N_6421,N_7099);
nand U7904 (N_7904,N_6618,N_6920);
and U7905 (N_7905,N_6422,N_6830);
xor U7906 (N_7906,N_6893,N_6793);
or U7907 (N_7907,N_6636,N_7112);
xor U7908 (N_7908,N_6475,N_7054);
or U7909 (N_7909,N_6807,N_6743);
nand U7910 (N_7910,N_6668,N_7076);
or U7911 (N_7911,N_6517,N_7117);
or U7912 (N_7912,N_6868,N_7079);
nand U7913 (N_7913,N_6726,N_6562);
or U7914 (N_7914,N_6906,N_6877);
xnor U7915 (N_7915,N_7073,N_6483);
or U7916 (N_7916,N_6537,N_6588);
or U7917 (N_7917,N_6734,N_6660);
nor U7918 (N_7918,N_6938,N_6613);
and U7919 (N_7919,N_6478,N_6423);
or U7920 (N_7920,N_6824,N_6740);
or U7921 (N_7921,N_6644,N_6734);
xor U7922 (N_7922,N_6486,N_6409);
xor U7923 (N_7923,N_6922,N_7018);
nand U7924 (N_7924,N_6714,N_6692);
nor U7925 (N_7925,N_6751,N_6588);
and U7926 (N_7926,N_7011,N_6480);
nor U7927 (N_7927,N_7121,N_6692);
or U7928 (N_7928,N_6539,N_6857);
nor U7929 (N_7929,N_6964,N_6439);
xnor U7930 (N_7930,N_7168,N_6786);
or U7931 (N_7931,N_6433,N_6817);
nand U7932 (N_7932,N_7113,N_6843);
and U7933 (N_7933,N_7157,N_6416);
nor U7934 (N_7934,N_7172,N_6894);
and U7935 (N_7935,N_6663,N_6708);
nand U7936 (N_7936,N_6805,N_6451);
or U7937 (N_7937,N_6939,N_7166);
nand U7938 (N_7938,N_6456,N_6673);
and U7939 (N_7939,N_7125,N_7064);
or U7940 (N_7940,N_7058,N_6774);
nor U7941 (N_7941,N_6689,N_6718);
nor U7942 (N_7942,N_7125,N_6735);
or U7943 (N_7943,N_6564,N_6427);
nor U7944 (N_7944,N_6562,N_7115);
nand U7945 (N_7945,N_6570,N_7170);
and U7946 (N_7946,N_6621,N_6632);
nand U7947 (N_7947,N_6999,N_6432);
and U7948 (N_7948,N_6575,N_7111);
nor U7949 (N_7949,N_6511,N_6748);
xor U7950 (N_7950,N_6806,N_7027);
nor U7951 (N_7951,N_7136,N_6819);
or U7952 (N_7952,N_6424,N_6809);
nor U7953 (N_7953,N_6635,N_6804);
xor U7954 (N_7954,N_6513,N_6865);
nand U7955 (N_7955,N_6919,N_7099);
or U7956 (N_7956,N_6899,N_7183);
nand U7957 (N_7957,N_6551,N_6480);
xor U7958 (N_7958,N_6776,N_7026);
or U7959 (N_7959,N_6582,N_6531);
xnor U7960 (N_7960,N_7118,N_6474);
nor U7961 (N_7961,N_6730,N_6758);
or U7962 (N_7962,N_6577,N_7166);
nand U7963 (N_7963,N_6787,N_7182);
and U7964 (N_7964,N_6804,N_6614);
nor U7965 (N_7965,N_6563,N_6540);
xor U7966 (N_7966,N_6620,N_6678);
xor U7967 (N_7967,N_6554,N_6808);
xor U7968 (N_7968,N_6704,N_7131);
nor U7969 (N_7969,N_6478,N_6422);
nand U7970 (N_7970,N_6910,N_6995);
xnor U7971 (N_7971,N_7156,N_6486);
nor U7972 (N_7972,N_6539,N_6702);
xor U7973 (N_7973,N_6839,N_6547);
nand U7974 (N_7974,N_6720,N_6485);
or U7975 (N_7975,N_6507,N_7120);
or U7976 (N_7976,N_6477,N_7185);
or U7977 (N_7977,N_6646,N_6572);
or U7978 (N_7978,N_6778,N_7001);
nand U7979 (N_7979,N_6995,N_6563);
or U7980 (N_7980,N_6802,N_6751);
xor U7981 (N_7981,N_7196,N_6984);
or U7982 (N_7982,N_7052,N_7089);
nand U7983 (N_7983,N_6972,N_6716);
or U7984 (N_7984,N_6731,N_7041);
nor U7985 (N_7985,N_6515,N_7145);
or U7986 (N_7986,N_6706,N_6726);
nand U7987 (N_7987,N_6857,N_6518);
xnor U7988 (N_7988,N_6872,N_6422);
or U7989 (N_7989,N_6547,N_6564);
xnor U7990 (N_7990,N_6630,N_6519);
and U7991 (N_7991,N_6969,N_6772);
nand U7992 (N_7992,N_6491,N_7199);
nand U7993 (N_7993,N_6877,N_7003);
xor U7994 (N_7994,N_7037,N_6587);
xor U7995 (N_7995,N_6995,N_7050);
xnor U7996 (N_7996,N_7017,N_6821);
xor U7997 (N_7997,N_6489,N_6859);
xnor U7998 (N_7998,N_7187,N_6878);
nand U7999 (N_7999,N_7197,N_6711);
or U8000 (N_8000,N_7794,N_7472);
nand U8001 (N_8001,N_7812,N_7240);
nand U8002 (N_8002,N_7647,N_7379);
nor U8003 (N_8003,N_7872,N_7238);
nor U8004 (N_8004,N_7578,N_7525);
and U8005 (N_8005,N_7893,N_7570);
and U8006 (N_8006,N_7418,N_7921);
xor U8007 (N_8007,N_7342,N_7832);
and U8008 (N_8008,N_7897,N_7603);
or U8009 (N_8009,N_7358,N_7308);
xor U8010 (N_8010,N_7512,N_7526);
and U8011 (N_8011,N_7749,N_7253);
xor U8012 (N_8012,N_7696,N_7429);
nor U8013 (N_8013,N_7902,N_7901);
or U8014 (N_8014,N_7631,N_7447);
or U8015 (N_8015,N_7702,N_7333);
nand U8016 (N_8016,N_7255,N_7881);
and U8017 (N_8017,N_7237,N_7280);
nor U8018 (N_8018,N_7935,N_7747);
or U8019 (N_8019,N_7368,N_7380);
xor U8020 (N_8020,N_7995,N_7576);
or U8021 (N_8021,N_7304,N_7653);
and U8022 (N_8022,N_7931,N_7299);
or U8023 (N_8023,N_7662,N_7937);
and U8024 (N_8024,N_7974,N_7353);
or U8025 (N_8025,N_7699,N_7571);
nor U8026 (N_8026,N_7998,N_7875);
xor U8027 (N_8027,N_7880,N_7431);
or U8028 (N_8028,N_7848,N_7396);
nand U8029 (N_8029,N_7797,N_7417);
nor U8030 (N_8030,N_7581,N_7329);
and U8031 (N_8031,N_7874,N_7854);
xor U8032 (N_8032,N_7544,N_7348);
xnor U8033 (N_8033,N_7265,N_7297);
nor U8034 (N_8034,N_7732,N_7674);
xor U8035 (N_8035,N_7269,N_7225);
xnor U8036 (N_8036,N_7487,N_7323);
nor U8037 (N_8037,N_7259,N_7252);
nor U8038 (N_8038,N_7464,N_7613);
xor U8039 (N_8039,N_7599,N_7973);
nand U8040 (N_8040,N_7783,N_7343);
nor U8041 (N_8041,N_7451,N_7499);
nand U8042 (N_8042,N_7898,N_7955);
xnor U8043 (N_8043,N_7870,N_7887);
nor U8044 (N_8044,N_7496,N_7750);
and U8045 (N_8045,N_7542,N_7740);
nand U8046 (N_8046,N_7231,N_7422);
nor U8047 (N_8047,N_7687,N_7939);
nor U8048 (N_8048,N_7878,N_7273);
nand U8049 (N_8049,N_7790,N_7501);
nor U8050 (N_8050,N_7957,N_7298);
nor U8051 (N_8051,N_7331,N_7286);
and U8052 (N_8052,N_7737,N_7940);
nor U8053 (N_8053,N_7816,N_7791);
and U8054 (N_8054,N_7554,N_7724);
nor U8055 (N_8055,N_7807,N_7932);
nand U8056 (N_8056,N_7612,N_7270);
nor U8057 (N_8057,N_7338,N_7624);
or U8058 (N_8058,N_7934,N_7315);
and U8059 (N_8059,N_7467,N_7719);
and U8060 (N_8060,N_7677,N_7637);
and U8061 (N_8061,N_7779,N_7520);
nand U8062 (N_8062,N_7210,N_7307);
and U8063 (N_8063,N_7885,N_7853);
nor U8064 (N_8064,N_7589,N_7636);
or U8065 (N_8065,N_7414,N_7793);
nor U8066 (N_8066,N_7310,N_7876);
and U8067 (N_8067,N_7558,N_7245);
and U8068 (N_8068,N_7466,N_7498);
nor U8069 (N_8069,N_7263,N_7650);
and U8070 (N_8070,N_7289,N_7508);
nand U8071 (N_8071,N_7376,N_7523);
xnor U8072 (N_8072,N_7679,N_7863);
nand U8073 (N_8073,N_7446,N_7585);
xnor U8074 (N_8074,N_7689,N_7775);
or U8075 (N_8075,N_7456,N_7519);
nand U8076 (N_8076,N_7730,N_7987);
or U8077 (N_8077,N_7611,N_7202);
and U8078 (N_8078,N_7648,N_7291);
xor U8079 (N_8079,N_7913,N_7820);
xnor U8080 (N_8080,N_7734,N_7758);
xnor U8081 (N_8081,N_7443,N_7610);
nand U8082 (N_8082,N_7882,N_7223);
or U8083 (N_8083,N_7781,N_7976);
or U8084 (N_8084,N_7547,N_7708);
or U8085 (N_8085,N_7627,N_7435);
xnor U8086 (N_8086,N_7938,N_7694);
or U8087 (N_8087,N_7577,N_7980);
or U8088 (N_8088,N_7306,N_7489);
xor U8089 (N_8089,N_7441,N_7565);
xnor U8090 (N_8090,N_7982,N_7201);
nor U8091 (N_8091,N_7909,N_7469);
nand U8092 (N_8092,N_7428,N_7262);
xnor U8093 (N_8093,N_7910,N_7860);
or U8094 (N_8094,N_7203,N_7841);
and U8095 (N_8095,N_7314,N_7411);
or U8096 (N_8096,N_7620,N_7671);
nor U8097 (N_8097,N_7596,N_7354);
nand U8098 (N_8098,N_7236,N_7274);
nor U8099 (N_8099,N_7319,N_7457);
nand U8100 (N_8100,N_7471,N_7945);
or U8101 (N_8101,N_7999,N_7246);
xnor U8102 (N_8102,N_7883,N_7320);
or U8103 (N_8103,N_7385,N_7318);
xnor U8104 (N_8104,N_7322,N_7328);
nor U8105 (N_8105,N_7264,N_7742);
nand U8106 (N_8106,N_7908,N_7470);
xor U8107 (N_8107,N_7409,N_7442);
and U8108 (N_8108,N_7907,N_7663);
nor U8109 (N_8109,N_7697,N_7805);
nor U8110 (N_8110,N_7335,N_7574);
xor U8111 (N_8111,N_7664,N_7356);
xor U8112 (N_8112,N_7561,N_7216);
nand U8113 (N_8113,N_7827,N_7215);
nor U8114 (N_8114,N_7529,N_7321);
and U8115 (N_8115,N_7929,N_7502);
nand U8116 (N_8116,N_7300,N_7959);
xor U8117 (N_8117,N_7733,N_7680);
or U8118 (N_8118,N_7421,N_7723);
or U8119 (N_8119,N_7248,N_7683);
xor U8120 (N_8120,N_7695,N_7224);
or U8121 (N_8121,N_7573,N_7731);
nand U8122 (N_8122,N_7864,N_7592);
or U8123 (N_8123,N_7716,N_7381);
and U8124 (N_8124,N_7922,N_7667);
nor U8125 (N_8125,N_7366,N_7281);
or U8126 (N_8126,N_7769,N_7293);
or U8127 (N_8127,N_7453,N_7904);
xor U8128 (N_8128,N_7420,N_7579);
nor U8129 (N_8129,N_7673,N_7383);
nor U8130 (N_8130,N_7767,N_7272);
or U8131 (N_8131,N_7958,N_7388);
and U8132 (N_8132,N_7686,N_7657);
and U8133 (N_8133,N_7389,N_7590);
or U8134 (N_8134,N_7205,N_7822);
or U8135 (N_8135,N_7211,N_7785);
xnor U8136 (N_8136,N_7652,N_7551);
nand U8137 (N_8137,N_7370,N_7642);
or U8138 (N_8138,N_7377,N_7969);
nor U8139 (N_8139,N_7247,N_7365);
and U8140 (N_8140,N_7254,N_7753);
or U8141 (N_8141,N_7847,N_7838);
or U8142 (N_8142,N_7886,N_7799);
xnor U8143 (N_8143,N_7659,N_7220);
and U8144 (N_8144,N_7609,N_7917);
xnor U8145 (N_8145,N_7433,N_7230);
and U8146 (N_8146,N_7474,N_7700);
and U8147 (N_8147,N_7595,N_7408);
or U8148 (N_8148,N_7317,N_7324);
or U8149 (N_8149,N_7560,N_7583);
nand U8150 (N_8150,N_7916,N_7510);
nand U8151 (N_8151,N_7926,N_7514);
nand U8152 (N_8152,N_7303,N_7622);
nand U8153 (N_8153,N_7994,N_7608);
nand U8154 (N_8154,N_7656,N_7960);
nor U8155 (N_8155,N_7754,N_7895);
nor U8156 (N_8156,N_7978,N_7538);
or U8157 (N_8157,N_7282,N_7972);
xnor U8158 (N_8158,N_7707,N_7729);
and U8159 (N_8159,N_7440,N_7840);
and U8160 (N_8160,N_7949,N_7533);
and U8161 (N_8161,N_7891,N_7384);
or U8162 (N_8162,N_7345,N_7339);
nor U8163 (N_8163,N_7531,N_7743);
nor U8164 (N_8164,N_7965,N_7504);
nor U8165 (N_8165,N_7855,N_7405);
or U8166 (N_8166,N_7406,N_7628);
or U8167 (N_8167,N_7575,N_7513);
xor U8168 (N_8168,N_7235,N_7851);
xnor U8169 (N_8169,N_7947,N_7705);
and U8170 (N_8170,N_7778,N_7550);
xor U8171 (N_8171,N_7903,N_7984);
nor U8172 (N_8172,N_7424,N_7744);
xor U8173 (N_8173,N_7675,N_7352);
nor U8174 (N_8174,N_7630,N_7941);
xnor U8175 (N_8175,N_7204,N_7761);
xnor U8176 (N_8176,N_7745,N_7437);
and U8177 (N_8177,N_7676,N_7334);
nand U8178 (N_8178,N_7398,N_7540);
or U8179 (N_8179,N_7803,N_7463);
nand U8180 (N_8180,N_7537,N_7445);
and U8181 (N_8181,N_7726,N_7226);
or U8182 (N_8182,N_7811,N_7332);
or U8183 (N_8183,N_7640,N_7587);
xor U8184 (N_8184,N_7927,N_7450);
and U8185 (N_8185,N_7682,N_7552);
nor U8186 (N_8186,N_7206,N_7771);
and U8187 (N_8187,N_7404,N_7266);
nor U8188 (N_8188,N_7942,N_7912);
nor U8189 (N_8189,N_7458,N_7290);
nor U8190 (N_8190,N_7983,N_7507);
or U8191 (N_8191,N_7244,N_7454);
or U8192 (N_8192,N_7207,N_7639);
nor U8193 (N_8193,N_7249,N_7536);
nor U8194 (N_8194,N_7776,N_7432);
or U8195 (N_8195,N_7490,N_7258);
nand U8196 (N_8196,N_7439,N_7839);
xnor U8197 (N_8197,N_7214,N_7371);
nand U8198 (N_8198,N_7241,N_7920);
nor U8199 (N_8199,N_7918,N_7643);
and U8200 (N_8200,N_7884,N_7626);
or U8201 (N_8201,N_7588,N_7294);
nor U8202 (N_8202,N_7473,N_7678);
xor U8203 (N_8203,N_7243,N_7752);
and U8204 (N_8204,N_7990,N_7954);
xnor U8205 (N_8205,N_7764,N_7715);
and U8206 (N_8206,N_7780,N_7867);
nand U8207 (N_8207,N_7364,N_7948);
and U8208 (N_8208,N_7486,N_7899);
nor U8209 (N_8209,N_7943,N_7234);
or U8210 (N_8210,N_7810,N_7232);
xor U8211 (N_8211,N_7539,N_7849);
nor U8212 (N_8212,N_7268,N_7792);
nor U8213 (N_8213,N_7415,N_7511);
or U8214 (N_8214,N_7509,N_7452);
nor U8215 (N_8215,N_7476,N_7591);
or U8216 (N_8216,N_7250,N_7722);
nor U8217 (N_8217,N_7692,N_7302);
nor U8218 (N_8218,N_7607,N_7548);
or U8219 (N_8219,N_7462,N_7900);
xnor U8220 (N_8220,N_7862,N_7936);
nor U8221 (N_8221,N_7685,N_7986);
nand U8222 (N_8222,N_7401,N_7660);
xor U8223 (N_8223,N_7967,N_7889);
or U8224 (N_8224,N_7768,N_7815);
and U8225 (N_8225,N_7992,N_7257);
and U8226 (N_8226,N_7833,N_7760);
nor U8227 (N_8227,N_7493,N_7218);
or U8228 (N_8228,N_7727,N_7861);
xor U8229 (N_8229,N_7506,N_7879);
nor U8230 (N_8230,N_7260,N_7615);
and U8231 (N_8231,N_7928,N_7925);
xnor U8232 (N_8232,N_7741,N_7981);
xnor U8233 (N_8233,N_7933,N_7228);
nand U8234 (N_8234,N_7826,N_7709);
and U8235 (N_8235,N_7373,N_7527);
nand U8236 (N_8236,N_7829,N_7459);
nand U8237 (N_8237,N_7713,N_7755);
nor U8238 (N_8238,N_7763,N_7301);
xor U8239 (N_8239,N_7997,N_7774);
and U8240 (N_8240,N_7394,N_7786);
xnor U8241 (N_8241,N_7968,N_7718);
and U8242 (N_8242,N_7888,N_7911);
nand U8243 (N_8243,N_7654,N_7277);
nor U8244 (N_8244,N_7563,N_7309);
and U8245 (N_8245,N_7766,N_7614);
or U8246 (N_8246,N_7979,N_7390);
or U8247 (N_8247,N_7905,N_7569);
and U8248 (N_8248,N_7746,N_7391);
nor U8249 (N_8249,N_7808,N_7950);
and U8250 (N_8250,N_7449,N_7546);
or U8251 (N_8251,N_7416,N_7661);
or U8252 (N_8252,N_7545,N_7691);
nand U8253 (N_8253,N_7562,N_7200);
nor U8254 (N_8254,N_7444,N_7222);
nand U8255 (N_8255,N_7535,N_7844);
or U8256 (N_8256,N_7946,N_7944);
xnor U8257 (N_8257,N_7890,N_7714);
nand U8258 (N_8258,N_7341,N_7495);
xor U8259 (N_8259,N_7284,N_7804);
and U8260 (N_8260,N_7465,N_7478);
nor U8261 (N_8261,N_7975,N_7633);
nand U8262 (N_8262,N_7584,N_7868);
xor U8263 (N_8263,N_7505,N_7710);
and U8264 (N_8264,N_7896,N_7279);
nor U8265 (N_8265,N_7412,N_7350);
or U8266 (N_8266,N_7485,N_7634);
xnor U8267 (N_8267,N_7488,N_7572);
and U8268 (N_8268,N_7582,N_7711);
nand U8269 (N_8269,N_7605,N_7209);
xor U8270 (N_8270,N_7430,N_7311);
nor U8271 (N_8271,N_7835,N_7261);
and U8272 (N_8272,N_7378,N_7287);
nor U8273 (N_8273,N_7991,N_7985);
xor U8274 (N_8274,N_7285,N_7555);
nor U8275 (N_8275,N_7482,N_7503);
or U8276 (N_8276,N_7316,N_7670);
or U8277 (N_8277,N_7859,N_7712);
xor U8278 (N_8278,N_7271,N_7357);
and U8279 (N_8279,N_7426,N_7480);
nand U8280 (N_8280,N_7953,N_7892);
xnor U8281 (N_8281,N_7728,N_7347);
xnor U8282 (N_8282,N_7483,N_7690);
xnor U8283 (N_8283,N_7625,N_7251);
nor U8284 (N_8284,N_7586,N_7326);
or U8285 (N_8285,N_7518,N_7491);
xnor U8286 (N_8286,N_7372,N_7641);
nand U8287 (N_8287,N_7276,N_7330);
and U8288 (N_8288,N_7966,N_7638);
xor U8289 (N_8289,N_7951,N_7602);
and U8290 (N_8290,N_7801,N_7484);
xor U8291 (N_8291,N_7403,N_7693);
nor U8292 (N_8292,N_7877,N_7387);
or U8293 (N_8293,N_7646,N_7813);
or U8294 (N_8294,N_7522,N_7468);
nor U8295 (N_8295,N_7566,N_7698);
and U8296 (N_8296,N_7382,N_7846);
xor U8297 (N_8297,N_7530,N_7632);
xnor U8298 (N_8298,N_7221,N_7930);
xor U8299 (N_8299,N_7756,N_7549);
or U8300 (N_8300,N_7564,N_7964);
nor U8301 (N_8301,N_7397,N_7425);
xnor U8302 (N_8302,N_7736,N_7725);
or U8303 (N_8303,N_7956,N_7337);
xnor U8304 (N_8304,N_7619,N_7601);
or U8305 (N_8305,N_7988,N_7762);
and U8306 (N_8306,N_7479,N_7971);
xor U8307 (N_8307,N_7809,N_7915);
and U8308 (N_8308,N_7344,N_7873);
nor U8309 (N_8309,N_7213,N_7393);
nand U8310 (N_8310,N_7806,N_7796);
and U8311 (N_8311,N_7295,N_7906);
nor U8312 (N_8312,N_7704,N_7386);
and U8313 (N_8313,N_7789,N_7651);
xor U8314 (N_8314,N_7233,N_7327);
nor U8315 (N_8315,N_7962,N_7534);
or U8316 (N_8316,N_7410,N_7720);
or U8317 (N_8317,N_7423,N_7823);
or U8318 (N_8318,N_7553,N_7703);
nor U8319 (N_8319,N_7278,N_7375);
and U8320 (N_8320,N_7748,N_7814);
xnor U8321 (N_8321,N_7834,N_7963);
xnor U8322 (N_8322,N_7645,N_7400);
and U8323 (N_8323,N_7606,N_7721);
or U8324 (N_8324,N_7821,N_7850);
xor U8325 (N_8325,N_7427,N_7593);
xor U8326 (N_8326,N_7757,N_7735);
or U8327 (N_8327,N_7494,N_7830);
nand U8328 (N_8328,N_7894,N_7770);
nor U8329 (N_8329,N_7312,N_7296);
xnor U8330 (N_8330,N_7856,N_7688);
and U8331 (N_8331,N_7831,N_7658);
nor U8332 (N_8332,N_7773,N_7784);
or U8333 (N_8333,N_7568,N_7340);
and U8334 (N_8334,N_7666,N_7701);
nor U8335 (N_8335,N_7865,N_7481);
or U8336 (N_8336,N_7461,N_7541);
xnor U8337 (N_8337,N_7436,N_7681);
nand U8338 (N_8338,N_7598,N_7288);
nand U8339 (N_8339,N_7395,N_7351);
nand U8340 (N_8340,N_7706,N_7597);
and U8341 (N_8341,N_7346,N_7788);
xor U8342 (N_8342,N_7914,N_7239);
and U8343 (N_8343,N_7919,N_7360);
nor U8344 (N_8344,N_7392,N_7374);
or U8345 (N_8345,N_7532,N_7361);
and U8346 (N_8346,N_7993,N_7208);
or U8347 (N_8347,N_7836,N_7623);
or U8348 (N_8348,N_7795,N_7739);
and U8349 (N_8349,N_7824,N_7594);
and U8350 (N_8350,N_7669,N_7212);
nor U8351 (N_8351,N_7516,N_7283);
and U8352 (N_8352,N_7543,N_7751);
xor U8353 (N_8353,N_7455,N_7672);
nor U8354 (N_8354,N_7313,N_7871);
xor U8355 (N_8355,N_7665,N_7492);
nand U8356 (N_8356,N_7819,N_7977);
and U8357 (N_8357,N_7524,N_7477);
or U8358 (N_8358,N_7655,N_7717);
and U8359 (N_8359,N_7837,N_7227);
or U8360 (N_8360,N_7616,N_7267);
and U8361 (N_8361,N_7399,N_7438);
nand U8362 (N_8362,N_7825,N_7852);
and U8363 (N_8363,N_7961,N_7604);
xnor U8364 (N_8364,N_7349,N_7800);
nand U8365 (N_8365,N_7242,N_7644);
and U8366 (N_8366,N_7559,N_7842);
or U8367 (N_8367,N_7460,N_7857);
nand U8368 (N_8368,N_7367,N_7500);
or U8369 (N_8369,N_7845,N_7325);
xnor U8370 (N_8370,N_7798,N_7363);
or U8371 (N_8371,N_7515,N_7434);
nor U8372 (N_8372,N_7362,N_7759);
nand U8373 (N_8373,N_7996,N_7818);
nor U8374 (N_8374,N_7475,N_7219);
or U8375 (N_8375,N_7292,N_7828);
or U8376 (N_8376,N_7924,N_7402);
nor U8377 (N_8377,N_7556,N_7497);
nor U8378 (N_8378,N_7738,N_7407);
xor U8379 (N_8379,N_7787,N_7600);
xnor U8380 (N_8380,N_7989,N_7448);
nor U8381 (N_8381,N_7413,N_7359);
and U8382 (N_8382,N_7635,N_7580);
xnor U8383 (N_8383,N_7869,N_7866);
and U8384 (N_8384,N_7649,N_7843);
xnor U8385 (N_8385,N_7952,N_7336);
or U8386 (N_8386,N_7668,N_7629);
nor U8387 (N_8387,N_7256,N_7305);
nand U8388 (N_8388,N_7617,N_7419);
xor U8389 (N_8389,N_7802,N_7229);
xnor U8390 (N_8390,N_7817,N_7528);
nand U8391 (N_8391,N_7772,N_7777);
or U8392 (N_8392,N_7858,N_7217);
or U8393 (N_8393,N_7765,N_7275);
or U8394 (N_8394,N_7782,N_7517);
or U8395 (N_8395,N_7923,N_7567);
or U8396 (N_8396,N_7618,N_7355);
nor U8397 (N_8397,N_7621,N_7684);
nor U8398 (N_8398,N_7970,N_7521);
nor U8399 (N_8399,N_7369,N_7557);
nand U8400 (N_8400,N_7844,N_7656);
nor U8401 (N_8401,N_7360,N_7643);
and U8402 (N_8402,N_7513,N_7275);
and U8403 (N_8403,N_7321,N_7607);
nand U8404 (N_8404,N_7260,N_7515);
and U8405 (N_8405,N_7462,N_7490);
xnor U8406 (N_8406,N_7354,N_7801);
xor U8407 (N_8407,N_7611,N_7807);
nand U8408 (N_8408,N_7558,N_7763);
or U8409 (N_8409,N_7398,N_7622);
nor U8410 (N_8410,N_7827,N_7365);
xor U8411 (N_8411,N_7216,N_7426);
xor U8412 (N_8412,N_7621,N_7884);
nor U8413 (N_8413,N_7345,N_7226);
nand U8414 (N_8414,N_7440,N_7276);
nand U8415 (N_8415,N_7875,N_7669);
or U8416 (N_8416,N_7641,N_7561);
xnor U8417 (N_8417,N_7223,N_7714);
nor U8418 (N_8418,N_7687,N_7338);
nand U8419 (N_8419,N_7779,N_7990);
nor U8420 (N_8420,N_7876,N_7205);
nand U8421 (N_8421,N_7356,N_7897);
or U8422 (N_8422,N_7404,N_7587);
or U8423 (N_8423,N_7256,N_7223);
and U8424 (N_8424,N_7595,N_7908);
nor U8425 (N_8425,N_7386,N_7444);
and U8426 (N_8426,N_7269,N_7239);
xnor U8427 (N_8427,N_7683,N_7852);
or U8428 (N_8428,N_7373,N_7800);
nor U8429 (N_8429,N_7262,N_7927);
or U8430 (N_8430,N_7870,N_7331);
and U8431 (N_8431,N_7285,N_7749);
nor U8432 (N_8432,N_7447,N_7954);
nor U8433 (N_8433,N_7214,N_7870);
or U8434 (N_8434,N_7559,N_7444);
nand U8435 (N_8435,N_7403,N_7746);
xor U8436 (N_8436,N_7338,N_7742);
and U8437 (N_8437,N_7896,N_7250);
and U8438 (N_8438,N_7881,N_7783);
nand U8439 (N_8439,N_7259,N_7258);
nand U8440 (N_8440,N_7425,N_7726);
nand U8441 (N_8441,N_7410,N_7657);
or U8442 (N_8442,N_7709,N_7441);
nor U8443 (N_8443,N_7738,N_7409);
nand U8444 (N_8444,N_7863,N_7356);
or U8445 (N_8445,N_7883,N_7955);
nor U8446 (N_8446,N_7758,N_7933);
nor U8447 (N_8447,N_7265,N_7374);
or U8448 (N_8448,N_7274,N_7390);
nor U8449 (N_8449,N_7804,N_7344);
xnor U8450 (N_8450,N_7280,N_7803);
nand U8451 (N_8451,N_7808,N_7207);
and U8452 (N_8452,N_7465,N_7534);
nor U8453 (N_8453,N_7706,N_7660);
nand U8454 (N_8454,N_7976,N_7857);
or U8455 (N_8455,N_7464,N_7962);
and U8456 (N_8456,N_7648,N_7376);
xor U8457 (N_8457,N_7290,N_7253);
nand U8458 (N_8458,N_7672,N_7761);
xnor U8459 (N_8459,N_7649,N_7303);
or U8460 (N_8460,N_7779,N_7962);
nand U8461 (N_8461,N_7443,N_7507);
nor U8462 (N_8462,N_7507,N_7790);
xnor U8463 (N_8463,N_7365,N_7764);
nand U8464 (N_8464,N_7227,N_7375);
or U8465 (N_8465,N_7331,N_7738);
and U8466 (N_8466,N_7711,N_7719);
or U8467 (N_8467,N_7691,N_7572);
nor U8468 (N_8468,N_7550,N_7616);
nand U8469 (N_8469,N_7331,N_7657);
or U8470 (N_8470,N_7915,N_7439);
or U8471 (N_8471,N_7347,N_7520);
nor U8472 (N_8472,N_7612,N_7455);
and U8473 (N_8473,N_7374,N_7730);
xor U8474 (N_8474,N_7824,N_7229);
or U8475 (N_8475,N_7607,N_7293);
xnor U8476 (N_8476,N_7769,N_7903);
nand U8477 (N_8477,N_7979,N_7766);
and U8478 (N_8478,N_7544,N_7465);
or U8479 (N_8479,N_7639,N_7283);
and U8480 (N_8480,N_7286,N_7975);
and U8481 (N_8481,N_7460,N_7314);
and U8482 (N_8482,N_7654,N_7995);
xnor U8483 (N_8483,N_7689,N_7878);
and U8484 (N_8484,N_7895,N_7739);
or U8485 (N_8485,N_7813,N_7709);
nand U8486 (N_8486,N_7218,N_7322);
nor U8487 (N_8487,N_7442,N_7959);
and U8488 (N_8488,N_7422,N_7920);
xor U8489 (N_8489,N_7241,N_7255);
nor U8490 (N_8490,N_7900,N_7667);
or U8491 (N_8491,N_7565,N_7830);
and U8492 (N_8492,N_7673,N_7730);
nor U8493 (N_8493,N_7916,N_7834);
nor U8494 (N_8494,N_7711,N_7311);
xnor U8495 (N_8495,N_7608,N_7233);
and U8496 (N_8496,N_7497,N_7360);
or U8497 (N_8497,N_7827,N_7812);
xor U8498 (N_8498,N_7973,N_7671);
and U8499 (N_8499,N_7952,N_7963);
xnor U8500 (N_8500,N_7390,N_7340);
or U8501 (N_8501,N_7382,N_7993);
xnor U8502 (N_8502,N_7909,N_7857);
nor U8503 (N_8503,N_7287,N_7253);
and U8504 (N_8504,N_7493,N_7394);
or U8505 (N_8505,N_7895,N_7555);
nand U8506 (N_8506,N_7893,N_7348);
or U8507 (N_8507,N_7628,N_7236);
or U8508 (N_8508,N_7942,N_7934);
nand U8509 (N_8509,N_7949,N_7225);
xor U8510 (N_8510,N_7794,N_7225);
xor U8511 (N_8511,N_7220,N_7977);
or U8512 (N_8512,N_7498,N_7205);
nor U8513 (N_8513,N_7369,N_7478);
nor U8514 (N_8514,N_7963,N_7685);
xnor U8515 (N_8515,N_7707,N_7868);
or U8516 (N_8516,N_7446,N_7352);
nand U8517 (N_8517,N_7747,N_7252);
xnor U8518 (N_8518,N_7947,N_7410);
nor U8519 (N_8519,N_7471,N_7344);
or U8520 (N_8520,N_7799,N_7446);
and U8521 (N_8521,N_7415,N_7321);
and U8522 (N_8522,N_7625,N_7769);
nand U8523 (N_8523,N_7566,N_7918);
or U8524 (N_8524,N_7565,N_7846);
nand U8525 (N_8525,N_7930,N_7691);
and U8526 (N_8526,N_7768,N_7621);
or U8527 (N_8527,N_7661,N_7272);
or U8528 (N_8528,N_7411,N_7828);
nor U8529 (N_8529,N_7698,N_7906);
or U8530 (N_8530,N_7530,N_7924);
nand U8531 (N_8531,N_7310,N_7861);
xnor U8532 (N_8532,N_7313,N_7459);
nor U8533 (N_8533,N_7260,N_7765);
or U8534 (N_8534,N_7737,N_7433);
or U8535 (N_8535,N_7691,N_7784);
or U8536 (N_8536,N_7438,N_7913);
nand U8537 (N_8537,N_7608,N_7638);
xor U8538 (N_8538,N_7567,N_7795);
and U8539 (N_8539,N_7755,N_7630);
and U8540 (N_8540,N_7656,N_7751);
or U8541 (N_8541,N_7866,N_7912);
xnor U8542 (N_8542,N_7757,N_7205);
or U8543 (N_8543,N_7504,N_7397);
nor U8544 (N_8544,N_7726,N_7875);
xnor U8545 (N_8545,N_7769,N_7855);
and U8546 (N_8546,N_7606,N_7781);
or U8547 (N_8547,N_7491,N_7935);
nand U8548 (N_8548,N_7681,N_7323);
and U8549 (N_8549,N_7276,N_7289);
nand U8550 (N_8550,N_7855,N_7694);
and U8551 (N_8551,N_7927,N_7571);
or U8552 (N_8552,N_7394,N_7487);
nand U8553 (N_8553,N_7984,N_7541);
or U8554 (N_8554,N_7852,N_7583);
nand U8555 (N_8555,N_7431,N_7281);
xnor U8556 (N_8556,N_7576,N_7204);
and U8557 (N_8557,N_7374,N_7947);
xnor U8558 (N_8558,N_7406,N_7703);
xnor U8559 (N_8559,N_7966,N_7666);
and U8560 (N_8560,N_7457,N_7497);
xor U8561 (N_8561,N_7983,N_7631);
xnor U8562 (N_8562,N_7437,N_7684);
nand U8563 (N_8563,N_7431,N_7558);
nor U8564 (N_8564,N_7447,N_7490);
xor U8565 (N_8565,N_7481,N_7600);
xor U8566 (N_8566,N_7991,N_7870);
nor U8567 (N_8567,N_7790,N_7723);
nand U8568 (N_8568,N_7360,N_7471);
nor U8569 (N_8569,N_7321,N_7205);
and U8570 (N_8570,N_7241,N_7969);
xor U8571 (N_8571,N_7518,N_7861);
nand U8572 (N_8572,N_7625,N_7994);
nand U8573 (N_8573,N_7562,N_7829);
and U8574 (N_8574,N_7626,N_7427);
xor U8575 (N_8575,N_7745,N_7725);
xnor U8576 (N_8576,N_7365,N_7941);
nor U8577 (N_8577,N_7908,N_7256);
nand U8578 (N_8578,N_7678,N_7959);
and U8579 (N_8579,N_7829,N_7758);
xor U8580 (N_8580,N_7246,N_7696);
nor U8581 (N_8581,N_7609,N_7703);
and U8582 (N_8582,N_7944,N_7505);
nor U8583 (N_8583,N_7820,N_7733);
nand U8584 (N_8584,N_7416,N_7738);
nand U8585 (N_8585,N_7684,N_7707);
xnor U8586 (N_8586,N_7791,N_7595);
nor U8587 (N_8587,N_7329,N_7870);
or U8588 (N_8588,N_7895,N_7972);
and U8589 (N_8589,N_7804,N_7233);
nand U8590 (N_8590,N_7378,N_7252);
xnor U8591 (N_8591,N_7723,N_7850);
nand U8592 (N_8592,N_7250,N_7371);
or U8593 (N_8593,N_7594,N_7939);
and U8594 (N_8594,N_7642,N_7632);
nor U8595 (N_8595,N_7413,N_7617);
or U8596 (N_8596,N_7867,N_7220);
xor U8597 (N_8597,N_7548,N_7611);
or U8598 (N_8598,N_7374,N_7367);
nor U8599 (N_8599,N_7802,N_7463);
nor U8600 (N_8600,N_7217,N_7609);
and U8601 (N_8601,N_7304,N_7929);
or U8602 (N_8602,N_7483,N_7325);
nand U8603 (N_8603,N_7682,N_7622);
nor U8604 (N_8604,N_7291,N_7421);
nor U8605 (N_8605,N_7842,N_7281);
nand U8606 (N_8606,N_7369,N_7724);
nand U8607 (N_8607,N_7444,N_7868);
and U8608 (N_8608,N_7913,N_7912);
nor U8609 (N_8609,N_7576,N_7312);
nor U8610 (N_8610,N_7419,N_7320);
nor U8611 (N_8611,N_7418,N_7868);
nand U8612 (N_8612,N_7826,N_7797);
nand U8613 (N_8613,N_7372,N_7371);
and U8614 (N_8614,N_7884,N_7529);
nor U8615 (N_8615,N_7803,N_7352);
xor U8616 (N_8616,N_7791,N_7852);
or U8617 (N_8617,N_7449,N_7923);
and U8618 (N_8618,N_7200,N_7323);
or U8619 (N_8619,N_7299,N_7773);
or U8620 (N_8620,N_7716,N_7736);
nand U8621 (N_8621,N_7859,N_7913);
nor U8622 (N_8622,N_7428,N_7356);
or U8623 (N_8623,N_7210,N_7658);
nor U8624 (N_8624,N_7837,N_7319);
xor U8625 (N_8625,N_7205,N_7273);
and U8626 (N_8626,N_7229,N_7879);
or U8627 (N_8627,N_7342,N_7213);
or U8628 (N_8628,N_7235,N_7423);
and U8629 (N_8629,N_7547,N_7387);
xor U8630 (N_8630,N_7787,N_7729);
nor U8631 (N_8631,N_7307,N_7745);
xnor U8632 (N_8632,N_7803,N_7694);
xnor U8633 (N_8633,N_7385,N_7679);
nor U8634 (N_8634,N_7211,N_7357);
nand U8635 (N_8635,N_7597,N_7356);
and U8636 (N_8636,N_7715,N_7245);
xor U8637 (N_8637,N_7889,N_7620);
and U8638 (N_8638,N_7237,N_7309);
and U8639 (N_8639,N_7784,N_7689);
or U8640 (N_8640,N_7776,N_7485);
or U8641 (N_8641,N_7219,N_7252);
xnor U8642 (N_8642,N_7605,N_7728);
xnor U8643 (N_8643,N_7219,N_7779);
and U8644 (N_8644,N_7769,N_7665);
nor U8645 (N_8645,N_7929,N_7845);
xor U8646 (N_8646,N_7743,N_7902);
and U8647 (N_8647,N_7790,N_7776);
xor U8648 (N_8648,N_7678,N_7232);
and U8649 (N_8649,N_7720,N_7849);
and U8650 (N_8650,N_7562,N_7906);
nor U8651 (N_8651,N_7293,N_7998);
nor U8652 (N_8652,N_7602,N_7576);
or U8653 (N_8653,N_7266,N_7511);
and U8654 (N_8654,N_7541,N_7511);
and U8655 (N_8655,N_7924,N_7520);
xor U8656 (N_8656,N_7615,N_7277);
or U8657 (N_8657,N_7315,N_7607);
or U8658 (N_8658,N_7598,N_7332);
nor U8659 (N_8659,N_7349,N_7480);
nor U8660 (N_8660,N_7389,N_7309);
or U8661 (N_8661,N_7515,N_7590);
nand U8662 (N_8662,N_7443,N_7939);
nor U8663 (N_8663,N_7627,N_7220);
nand U8664 (N_8664,N_7707,N_7361);
nor U8665 (N_8665,N_7542,N_7859);
nor U8666 (N_8666,N_7727,N_7487);
nand U8667 (N_8667,N_7866,N_7412);
or U8668 (N_8668,N_7211,N_7499);
or U8669 (N_8669,N_7815,N_7655);
nor U8670 (N_8670,N_7349,N_7880);
nor U8671 (N_8671,N_7473,N_7713);
xnor U8672 (N_8672,N_7668,N_7716);
and U8673 (N_8673,N_7848,N_7212);
nand U8674 (N_8674,N_7231,N_7661);
or U8675 (N_8675,N_7879,N_7346);
xor U8676 (N_8676,N_7532,N_7405);
and U8677 (N_8677,N_7761,N_7997);
nand U8678 (N_8678,N_7803,N_7842);
nand U8679 (N_8679,N_7852,N_7520);
nand U8680 (N_8680,N_7911,N_7994);
nand U8681 (N_8681,N_7900,N_7821);
nand U8682 (N_8682,N_7276,N_7566);
or U8683 (N_8683,N_7943,N_7706);
or U8684 (N_8684,N_7200,N_7864);
xor U8685 (N_8685,N_7517,N_7425);
and U8686 (N_8686,N_7647,N_7834);
nor U8687 (N_8687,N_7414,N_7871);
nor U8688 (N_8688,N_7842,N_7596);
xor U8689 (N_8689,N_7210,N_7398);
xnor U8690 (N_8690,N_7976,N_7462);
or U8691 (N_8691,N_7218,N_7740);
nor U8692 (N_8692,N_7442,N_7472);
and U8693 (N_8693,N_7667,N_7848);
and U8694 (N_8694,N_7815,N_7393);
and U8695 (N_8695,N_7295,N_7405);
nor U8696 (N_8696,N_7424,N_7907);
or U8697 (N_8697,N_7757,N_7628);
nor U8698 (N_8698,N_7332,N_7714);
nor U8699 (N_8699,N_7562,N_7300);
and U8700 (N_8700,N_7660,N_7698);
xnor U8701 (N_8701,N_7945,N_7931);
xnor U8702 (N_8702,N_7413,N_7382);
nor U8703 (N_8703,N_7526,N_7839);
xor U8704 (N_8704,N_7928,N_7637);
or U8705 (N_8705,N_7733,N_7301);
nor U8706 (N_8706,N_7618,N_7940);
and U8707 (N_8707,N_7344,N_7869);
nor U8708 (N_8708,N_7553,N_7349);
nand U8709 (N_8709,N_7880,N_7834);
xor U8710 (N_8710,N_7277,N_7384);
and U8711 (N_8711,N_7370,N_7922);
and U8712 (N_8712,N_7276,N_7748);
nor U8713 (N_8713,N_7735,N_7624);
nand U8714 (N_8714,N_7680,N_7606);
nand U8715 (N_8715,N_7366,N_7257);
nand U8716 (N_8716,N_7590,N_7488);
nor U8717 (N_8717,N_7877,N_7902);
nor U8718 (N_8718,N_7763,N_7408);
and U8719 (N_8719,N_7986,N_7255);
nor U8720 (N_8720,N_7314,N_7854);
or U8721 (N_8721,N_7506,N_7748);
xnor U8722 (N_8722,N_7945,N_7465);
or U8723 (N_8723,N_7807,N_7311);
nand U8724 (N_8724,N_7246,N_7385);
xor U8725 (N_8725,N_7508,N_7418);
xor U8726 (N_8726,N_7247,N_7938);
nor U8727 (N_8727,N_7685,N_7396);
or U8728 (N_8728,N_7761,N_7695);
and U8729 (N_8729,N_7802,N_7574);
or U8730 (N_8730,N_7321,N_7458);
and U8731 (N_8731,N_7314,N_7802);
nand U8732 (N_8732,N_7826,N_7742);
nor U8733 (N_8733,N_7822,N_7924);
nand U8734 (N_8734,N_7528,N_7438);
or U8735 (N_8735,N_7284,N_7823);
and U8736 (N_8736,N_7372,N_7236);
xnor U8737 (N_8737,N_7779,N_7418);
nand U8738 (N_8738,N_7429,N_7718);
and U8739 (N_8739,N_7925,N_7312);
or U8740 (N_8740,N_7415,N_7401);
nor U8741 (N_8741,N_7713,N_7535);
or U8742 (N_8742,N_7408,N_7346);
nand U8743 (N_8743,N_7532,N_7832);
nor U8744 (N_8744,N_7962,N_7254);
xnor U8745 (N_8745,N_7335,N_7268);
and U8746 (N_8746,N_7281,N_7854);
and U8747 (N_8747,N_7815,N_7895);
nor U8748 (N_8748,N_7384,N_7822);
nor U8749 (N_8749,N_7223,N_7618);
or U8750 (N_8750,N_7209,N_7277);
or U8751 (N_8751,N_7699,N_7761);
nor U8752 (N_8752,N_7686,N_7946);
nand U8753 (N_8753,N_7960,N_7258);
or U8754 (N_8754,N_7697,N_7250);
xnor U8755 (N_8755,N_7717,N_7528);
and U8756 (N_8756,N_7482,N_7878);
and U8757 (N_8757,N_7951,N_7815);
nand U8758 (N_8758,N_7722,N_7214);
and U8759 (N_8759,N_7387,N_7212);
nor U8760 (N_8760,N_7627,N_7510);
and U8761 (N_8761,N_7794,N_7620);
xor U8762 (N_8762,N_7735,N_7208);
nor U8763 (N_8763,N_7237,N_7764);
and U8764 (N_8764,N_7847,N_7774);
nor U8765 (N_8765,N_7517,N_7841);
xnor U8766 (N_8766,N_7379,N_7634);
nand U8767 (N_8767,N_7954,N_7786);
and U8768 (N_8768,N_7670,N_7790);
nand U8769 (N_8769,N_7362,N_7408);
nand U8770 (N_8770,N_7203,N_7891);
nor U8771 (N_8771,N_7847,N_7579);
nor U8772 (N_8772,N_7929,N_7445);
and U8773 (N_8773,N_7450,N_7441);
or U8774 (N_8774,N_7478,N_7953);
nor U8775 (N_8775,N_7341,N_7541);
nor U8776 (N_8776,N_7417,N_7701);
and U8777 (N_8777,N_7566,N_7807);
and U8778 (N_8778,N_7866,N_7559);
xnor U8779 (N_8779,N_7214,N_7343);
xnor U8780 (N_8780,N_7636,N_7585);
or U8781 (N_8781,N_7417,N_7621);
xnor U8782 (N_8782,N_7493,N_7644);
nand U8783 (N_8783,N_7317,N_7925);
nor U8784 (N_8784,N_7987,N_7581);
nor U8785 (N_8785,N_7690,N_7679);
or U8786 (N_8786,N_7411,N_7802);
or U8787 (N_8787,N_7916,N_7874);
nand U8788 (N_8788,N_7556,N_7521);
xor U8789 (N_8789,N_7351,N_7882);
nor U8790 (N_8790,N_7481,N_7422);
and U8791 (N_8791,N_7285,N_7675);
xor U8792 (N_8792,N_7206,N_7207);
and U8793 (N_8793,N_7727,N_7953);
or U8794 (N_8794,N_7383,N_7777);
nand U8795 (N_8795,N_7679,N_7362);
nand U8796 (N_8796,N_7525,N_7939);
xnor U8797 (N_8797,N_7269,N_7535);
nor U8798 (N_8798,N_7580,N_7954);
nand U8799 (N_8799,N_7847,N_7777);
xnor U8800 (N_8800,N_8259,N_8169);
and U8801 (N_8801,N_8280,N_8399);
nor U8802 (N_8802,N_8469,N_8562);
and U8803 (N_8803,N_8422,N_8224);
nor U8804 (N_8804,N_8671,N_8213);
or U8805 (N_8805,N_8576,N_8061);
and U8806 (N_8806,N_8225,N_8125);
nor U8807 (N_8807,N_8105,N_8048);
nand U8808 (N_8808,N_8240,N_8680);
xnor U8809 (N_8809,N_8111,N_8339);
or U8810 (N_8810,N_8792,N_8234);
nand U8811 (N_8811,N_8159,N_8349);
xor U8812 (N_8812,N_8538,N_8664);
or U8813 (N_8813,N_8455,N_8536);
and U8814 (N_8814,N_8679,N_8662);
xor U8815 (N_8815,N_8690,N_8047);
or U8816 (N_8816,N_8698,N_8618);
and U8817 (N_8817,N_8151,N_8470);
or U8818 (N_8818,N_8295,N_8477);
nand U8819 (N_8819,N_8539,N_8189);
nor U8820 (N_8820,N_8250,N_8075);
nor U8821 (N_8821,N_8244,N_8186);
xnor U8822 (N_8822,N_8092,N_8115);
xor U8823 (N_8823,N_8427,N_8214);
nand U8824 (N_8824,N_8388,N_8301);
or U8825 (N_8825,N_8443,N_8567);
or U8826 (N_8826,N_8086,N_8117);
nand U8827 (N_8827,N_8144,N_8438);
xnor U8828 (N_8828,N_8034,N_8681);
nand U8829 (N_8829,N_8683,N_8011);
and U8830 (N_8830,N_8030,N_8072);
nor U8831 (N_8831,N_8559,N_8794);
nand U8832 (N_8832,N_8327,N_8003);
xor U8833 (N_8833,N_8713,N_8708);
or U8834 (N_8834,N_8166,N_8094);
or U8835 (N_8835,N_8597,N_8445);
nor U8836 (N_8836,N_8797,N_8112);
and U8837 (N_8837,N_8419,N_8712);
nand U8838 (N_8838,N_8273,N_8572);
or U8839 (N_8839,N_8793,N_8300);
nand U8840 (N_8840,N_8025,N_8620);
or U8841 (N_8841,N_8089,N_8791);
xnor U8842 (N_8842,N_8376,N_8700);
nor U8843 (N_8843,N_8208,N_8465);
or U8844 (N_8844,N_8055,N_8499);
xor U8845 (N_8845,N_8175,N_8610);
and U8846 (N_8846,N_8473,N_8747);
nor U8847 (N_8847,N_8065,N_8303);
and U8848 (N_8848,N_8447,N_8436);
xor U8849 (N_8849,N_8717,N_8317);
or U8850 (N_8850,N_8164,N_8517);
or U8851 (N_8851,N_8340,N_8343);
xor U8852 (N_8852,N_8590,N_8570);
and U8853 (N_8853,N_8353,N_8421);
xnor U8854 (N_8854,N_8059,N_8685);
xor U8855 (N_8855,N_8533,N_8336);
and U8856 (N_8856,N_8254,N_8777);
xnor U8857 (N_8857,N_8724,N_8549);
or U8858 (N_8858,N_8631,N_8206);
and U8859 (N_8859,N_8192,N_8346);
or U8860 (N_8860,N_8589,N_8696);
nor U8861 (N_8861,N_8551,N_8401);
xor U8862 (N_8862,N_8150,N_8788);
and U8863 (N_8863,N_8644,N_8320);
nor U8864 (N_8864,N_8201,N_8594);
or U8865 (N_8865,N_8609,N_8433);
xnor U8866 (N_8866,N_8216,N_8351);
xnor U8867 (N_8867,N_8296,N_8358);
nor U8868 (N_8868,N_8449,N_8492);
or U8869 (N_8869,N_8135,N_8769);
or U8870 (N_8870,N_8534,N_8429);
nor U8871 (N_8871,N_8472,N_8402);
xnor U8872 (N_8872,N_8716,N_8621);
xnor U8873 (N_8873,N_8750,N_8658);
nand U8874 (N_8874,N_8742,N_8527);
and U8875 (N_8875,N_8302,N_8479);
nand U8876 (N_8876,N_8605,N_8196);
or U8877 (N_8877,N_8757,N_8434);
or U8878 (N_8878,N_8555,N_8475);
or U8879 (N_8879,N_8737,N_8264);
nand U8880 (N_8880,N_8446,N_8513);
xor U8881 (N_8881,N_8382,N_8318);
xnor U8882 (N_8882,N_8010,N_8299);
and U8883 (N_8883,N_8093,N_8348);
xnor U8884 (N_8884,N_8778,N_8341);
xnor U8885 (N_8885,N_8601,N_8198);
or U8886 (N_8886,N_8774,N_8078);
xor U8887 (N_8887,N_8420,N_8728);
and U8888 (N_8888,N_8227,N_8591);
xnor U8889 (N_8889,N_8640,N_8200);
xor U8890 (N_8890,N_8205,N_8754);
and U8891 (N_8891,N_8347,N_8223);
or U8892 (N_8892,N_8503,N_8408);
nor U8893 (N_8893,N_8123,N_8369);
xor U8894 (N_8894,N_8573,N_8678);
and U8895 (N_8895,N_8546,N_8004);
xor U8896 (N_8896,N_8370,N_8688);
or U8897 (N_8897,N_8697,N_8795);
and U8898 (N_8898,N_8173,N_8629);
nor U8899 (N_8899,N_8739,N_8614);
nand U8900 (N_8900,N_8691,N_8467);
or U8901 (N_8901,N_8087,N_8387);
nor U8902 (N_8902,N_8126,N_8523);
xnor U8903 (N_8903,N_8141,N_8246);
nand U8904 (N_8904,N_8577,N_8384);
xor U8905 (N_8905,N_8395,N_8765);
or U8906 (N_8906,N_8676,N_8294);
nand U8907 (N_8907,N_8560,N_8699);
and U8908 (N_8908,N_8583,N_8134);
and U8909 (N_8909,N_8319,N_8278);
and U8910 (N_8910,N_8608,N_8108);
nand U8911 (N_8911,N_8480,N_8406);
xnor U8912 (N_8912,N_8091,N_8185);
nand U8913 (N_8913,N_8623,N_8260);
and U8914 (N_8914,N_8116,N_8022);
nand U8915 (N_8915,N_8001,N_8038);
or U8916 (N_8916,N_8049,N_8487);
and U8917 (N_8917,N_8665,N_8068);
xor U8918 (N_8918,N_8693,N_8235);
xor U8919 (N_8919,N_8005,N_8316);
and U8920 (N_8920,N_8368,N_8329);
nand U8921 (N_8921,N_8053,N_8404);
or U8922 (N_8922,N_8062,N_8090);
xnor U8923 (N_8923,N_8652,N_8039);
or U8924 (N_8924,N_8071,N_8396);
or U8925 (N_8925,N_8361,N_8437);
xor U8926 (N_8926,N_8613,N_8174);
nor U8927 (N_8927,N_8079,N_8245);
nor U8928 (N_8928,N_8702,N_8645);
xnor U8929 (N_8929,N_8453,N_8454);
nand U8930 (N_8930,N_8036,N_8648);
nor U8931 (N_8931,N_8101,N_8617);
nor U8932 (N_8932,N_8498,N_8569);
xor U8933 (N_8933,N_8309,N_8655);
or U8934 (N_8934,N_8593,N_8097);
nand U8935 (N_8935,N_8770,N_8415);
xor U8936 (N_8936,N_8383,N_8506);
xor U8937 (N_8937,N_8096,N_8008);
nand U8938 (N_8938,N_8711,N_8416);
xnor U8939 (N_8939,N_8257,N_8323);
nor U8940 (N_8940,N_8760,N_8102);
nor U8941 (N_8941,N_8501,N_8464);
and U8942 (N_8942,N_8009,N_8554);
and U8943 (N_8943,N_8263,N_8571);
nor U8944 (N_8944,N_8315,N_8378);
and U8945 (N_8945,N_8720,N_8674);
and U8946 (N_8946,N_8553,N_8228);
nand U8947 (N_8947,N_8496,N_8675);
nand U8948 (N_8948,N_8391,N_8615);
nor U8949 (N_8949,N_8120,N_8740);
and U8950 (N_8950,N_8602,N_8290);
or U8951 (N_8951,N_8588,N_8050);
nor U8952 (N_8952,N_8110,N_8459);
nand U8953 (N_8953,N_8474,N_8535);
nand U8954 (N_8954,N_8154,N_8425);
nor U8955 (N_8955,N_8532,N_8771);
or U8956 (N_8956,N_8355,N_8289);
or U8957 (N_8957,N_8342,N_8160);
or U8958 (N_8958,N_8579,N_8667);
and U8959 (N_8959,N_8424,N_8218);
xor U8960 (N_8960,N_8460,N_8191);
xnor U8961 (N_8961,N_8485,N_8118);
and U8962 (N_8962,N_8650,N_8767);
nor U8963 (N_8963,N_8450,N_8360);
and U8964 (N_8964,N_8256,N_8431);
or U8965 (N_8965,N_8689,N_8148);
and U8966 (N_8966,N_8179,N_8133);
xnor U8967 (N_8967,N_8344,N_8721);
and U8968 (N_8968,N_8393,N_8452);
nand U8969 (N_8969,N_8345,N_8236);
nor U8970 (N_8970,N_8007,N_8633);
nand U8971 (N_8971,N_8237,N_8267);
xnor U8972 (N_8972,N_8018,N_8389);
nand U8973 (N_8973,N_8002,N_8611);
xor U8974 (N_8974,N_8232,N_8203);
xor U8975 (N_8975,N_8741,N_8321);
xnor U8976 (N_8976,N_8789,N_8563);
xor U8977 (N_8977,N_8514,N_8790);
nand U8978 (N_8978,N_8006,N_8574);
and U8979 (N_8979,N_8016,N_8687);
and U8980 (N_8980,N_8212,N_8332);
nand U8981 (N_8981,N_8181,N_8372);
nand U8982 (N_8982,N_8718,N_8627);
xor U8983 (N_8983,N_8584,N_8516);
nor U8984 (N_8984,N_8266,N_8283);
nand U8985 (N_8985,N_8511,N_8337);
or U8986 (N_8986,N_8156,N_8122);
nand U8987 (N_8987,N_8723,N_8619);
xor U8988 (N_8988,N_8275,N_8749);
xnor U8989 (N_8989,N_8738,N_8172);
and U8990 (N_8990,N_8411,N_8780);
or U8991 (N_8991,N_8064,N_8568);
nor U8992 (N_8992,N_8028,N_8195);
nor U8993 (N_8993,N_8409,N_8537);
nand U8994 (N_8994,N_8530,N_8385);
nor U8995 (N_8995,N_8162,N_8787);
nand U8996 (N_8996,N_8426,N_8442);
and U8997 (N_8997,N_8764,N_8131);
and U8998 (N_8998,N_8146,N_8586);
nand U8999 (N_8999,N_8145,N_8731);
or U9000 (N_9000,N_8701,N_8582);
nor U9001 (N_9001,N_8542,N_8132);
nor U9002 (N_9002,N_8103,N_8413);
or U9003 (N_9003,N_8277,N_8682);
and U9004 (N_9004,N_8157,N_8058);
nor U9005 (N_9005,N_8265,N_8291);
nand U9006 (N_9006,N_8733,N_8448);
and U9007 (N_9007,N_8081,N_8066);
xnor U9008 (N_9008,N_8276,N_8381);
nor U9009 (N_9009,N_8634,N_8715);
nand U9010 (N_9010,N_8736,N_8462);
and U9011 (N_9011,N_8782,N_8694);
nand U9012 (N_9012,N_8625,N_8488);
or U9013 (N_9013,N_8202,N_8364);
or U9014 (N_9014,N_8458,N_8070);
or U9015 (N_9015,N_8052,N_8779);
nand U9016 (N_9016,N_8466,N_8607);
or U9017 (N_9017,N_8761,N_8649);
or U9018 (N_9018,N_8439,N_8271);
nor U9019 (N_9019,N_8494,N_8167);
nand U9020 (N_9020,N_8684,N_8759);
nand U9021 (N_9021,N_8398,N_8063);
nand U9022 (N_9022,N_8270,N_8673);
xnor U9023 (N_9023,N_8666,N_8710);
or U9024 (N_9024,N_8281,N_8238);
and U9025 (N_9025,N_8178,N_8119);
nor U9026 (N_9026,N_8441,N_8635);
xnor U9027 (N_9027,N_8020,N_8215);
nor U9028 (N_9028,N_8706,N_8784);
and U9029 (N_9029,N_8067,N_8746);
xnor U9030 (N_9030,N_8657,N_8580);
xor U9031 (N_9031,N_8249,N_8219);
nor U9032 (N_9032,N_8188,N_8461);
nor U9033 (N_9033,N_8130,N_8558);
xnor U9034 (N_9034,N_8044,N_8233);
nor U9035 (N_9035,N_8753,N_8197);
xnor U9036 (N_9036,N_8489,N_8377);
nand U9037 (N_9037,N_8335,N_8177);
nand U9038 (N_9038,N_8239,N_8288);
or U9039 (N_9039,N_8221,N_8222);
nor U9040 (N_9040,N_8493,N_8362);
nand U9041 (N_9041,N_8149,N_8491);
nand U9042 (N_9042,N_8444,N_8194);
or U9043 (N_9043,N_8497,N_8677);
xor U9044 (N_9044,N_8379,N_8041);
or U9045 (N_9045,N_8155,N_8476);
xor U9046 (N_9046,N_8037,N_8138);
and U9047 (N_9047,N_8158,N_8056);
or U9048 (N_9048,N_8311,N_8029);
or U9049 (N_9049,N_8541,N_8531);
and U9050 (N_9050,N_8217,N_8756);
and U9051 (N_9051,N_8183,N_8253);
xnor U9052 (N_9052,N_8165,N_8104);
or U9053 (N_9053,N_8596,N_8478);
nand U9054 (N_9054,N_8705,N_8147);
nand U9055 (N_9055,N_8565,N_8204);
nor U9056 (N_9056,N_8528,N_8751);
xor U9057 (N_9057,N_8255,N_8483);
and U9058 (N_9058,N_8297,N_8084);
nor U9059 (N_9059,N_8663,N_8180);
xnor U9060 (N_9060,N_8729,N_8547);
and U9061 (N_9061,N_8324,N_8199);
xnor U9062 (N_9062,N_8734,N_8013);
nand U9063 (N_9063,N_8190,N_8307);
nor U9064 (N_9064,N_8502,N_8305);
xnor U9065 (N_9065,N_8153,N_8719);
xor U9066 (N_9066,N_8211,N_8354);
or U9067 (N_9067,N_8170,N_8540);
nand U9068 (N_9068,N_8672,N_8085);
and U9069 (N_9069,N_8763,N_8374);
xor U9070 (N_9070,N_8373,N_8703);
and U9071 (N_9071,N_8412,N_8550);
nand U9072 (N_9072,N_8414,N_8114);
and U9073 (N_9073,N_8587,N_8040);
xor U9074 (N_9074,N_8510,N_8262);
or U9075 (N_9075,N_8727,N_8077);
nor U9076 (N_9076,N_8035,N_8292);
nand U9077 (N_9077,N_8334,N_8268);
xor U9078 (N_9078,N_8636,N_8083);
xor U9079 (N_9079,N_8768,N_8637);
and U9080 (N_9080,N_8669,N_8392);
and U9081 (N_9081,N_8798,N_8612);
and U9082 (N_9082,N_8076,N_8367);
and U9083 (N_9083,N_8670,N_8099);
xor U9084 (N_9084,N_8333,N_8209);
nand U9085 (N_9085,N_8772,N_8410);
nand U9086 (N_9086,N_8661,N_8328);
nor U9087 (N_9087,N_8732,N_8557);
nand U9088 (N_9088,N_8785,N_8543);
nor U9089 (N_9089,N_8045,N_8088);
nand U9090 (N_9090,N_8113,N_8500);
nand U9091 (N_9091,N_8248,N_8730);
or U9092 (N_9092,N_8668,N_8024);
xor U9093 (N_9093,N_8752,N_8507);
nand U9094 (N_9094,N_8043,N_8735);
xor U9095 (N_9095,N_8285,N_8400);
xnor U9096 (N_9096,N_8241,N_8428);
nor U9097 (N_9097,N_8599,N_8137);
and U9098 (N_9098,N_8121,N_8272);
nor U9099 (N_9099,N_8632,N_8247);
and U9100 (N_9100,N_8628,N_8394);
xnor U9101 (N_9101,N_8060,N_8252);
or U9102 (N_9102,N_8312,N_8308);
nand U9103 (N_9103,N_8468,N_8293);
xor U9104 (N_9104,N_8495,N_8136);
or U9105 (N_9105,N_8592,N_8356);
and U9106 (N_9106,N_8026,N_8504);
xor U9107 (N_9107,N_8456,N_8220);
or U9108 (N_9108,N_8000,N_8585);
nand U9109 (N_9109,N_8545,N_8032);
nand U9110 (N_9110,N_8451,N_8624);
nand U9111 (N_9111,N_8725,N_8143);
or U9112 (N_9112,N_8529,N_8509);
nand U9113 (N_9113,N_8106,N_8080);
nand U9114 (N_9114,N_8418,N_8051);
nand U9115 (N_9115,N_8359,N_8519);
and U9116 (N_9116,N_8781,N_8371);
xor U9117 (N_9117,N_8298,N_8773);
nor U9118 (N_9118,N_8019,N_8352);
nor U9119 (N_9119,N_8098,N_8758);
nor U9120 (N_9120,N_8654,N_8326);
or U9121 (N_9121,N_8595,N_8692);
nand U9122 (N_9122,N_8552,N_8325);
xnor U9123 (N_9123,N_8630,N_8107);
nor U9124 (N_9124,N_8606,N_8653);
xnor U9125 (N_9125,N_8033,N_8745);
nor U9126 (N_9126,N_8365,N_8726);
and U9127 (N_9127,N_8338,N_8440);
or U9128 (N_9128,N_8193,N_8322);
nand U9129 (N_9129,N_8023,N_8603);
xnor U9130 (N_9130,N_8598,N_8482);
nand U9131 (N_9131,N_8100,N_8508);
and U9132 (N_9132,N_8457,N_8128);
or U9133 (N_9133,N_8082,N_8282);
or U9134 (N_9134,N_8207,N_8231);
or U9135 (N_9135,N_8380,N_8484);
and U9136 (N_9136,N_8168,N_8310);
and U9137 (N_9137,N_8704,N_8643);
or U9138 (N_9138,N_8521,N_8766);
nand U9139 (N_9139,N_8251,N_8184);
and U9140 (N_9140,N_8230,N_8659);
or U9141 (N_9141,N_8357,N_8313);
nor U9142 (N_9142,N_8622,N_8544);
nor U9143 (N_9143,N_8161,N_8171);
and U9144 (N_9144,N_8142,N_8287);
nor U9145 (N_9145,N_8176,N_8330);
nand U9146 (N_9146,N_8139,N_8490);
nand U9147 (N_9147,N_8522,N_8604);
xor U9148 (N_9148,N_8775,N_8258);
and U9149 (N_9149,N_8243,N_8027);
nor U9150 (N_9150,N_8274,N_8397);
and U9151 (N_9151,N_8363,N_8709);
nor U9152 (N_9152,N_8695,N_8269);
nor U9153 (N_9153,N_8639,N_8656);
xor U9154 (N_9154,N_8417,N_8042);
and U9155 (N_9155,N_8226,N_8375);
nand U9156 (N_9156,N_8074,N_8284);
or U9157 (N_9157,N_8481,N_8017);
xor U9158 (N_9158,N_8714,N_8279);
xnor U9159 (N_9159,N_8331,N_8129);
nand U9160 (N_9160,N_8486,N_8407);
nand U9161 (N_9161,N_8021,N_8647);
and U9162 (N_9162,N_8242,N_8520);
or U9163 (N_9163,N_8783,N_8564);
xnor U9164 (N_9164,N_8261,N_8304);
nand U9165 (N_9165,N_8046,N_8127);
and U9166 (N_9166,N_8432,N_8505);
xor U9167 (N_9167,N_8566,N_8799);
and U9168 (N_9168,N_8152,N_8423);
and U9169 (N_9169,N_8744,N_8163);
or U9170 (N_9170,N_8581,N_8642);
xor U9171 (N_9171,N_8762,N_8660);
nor U9172 (N_9172,N_8031,N_8600);
and U9173 (N_9173,N_8057,N_8786);
and U9174 (N_9174,N_8748,N_8286);
nor U9175 (N_9175,N_8403,N_8386);
nor U9176 (N_9176,N_8350,N_8575);
xor U9177 (N_9177,N_8638,N_8548);
nand U9178 (N_9178,N_8641,N_8686);
and U9179 (N_9179,N_8366,N_8755);
xnor U9180 (N_9180,N_8182,N_8390);
and U9181 (N_9181,N_8109,N_8140);
nand U9182 (N_9182,N_8722,N_8518);
nand U9183 (N_9183,N_8525,N_8616);
xor U9184 (N_9184,N_8012,N_8124);
nand U9185 (N_9185,N_8014,N_8015);
or U9186 (N_9186,N_8578,N_8776);
xor U9187 (N_9187,N_8561,N_8556);
nor U9188 (N_9188,N_8796,N_8651);
xnor U9189 (N_9189,N_8314,N_8526);
or U9190 (N_9190,N_8073,N_8512);
nor U9191 (N_9191,N_8524,N_8646);
nor U9192 (N_9192,N_8626,N_8515);
nand U9193 (N_9193,N_8707,N_8054);
nor U9194 (N_9194,N_8069,N_8210);
nand U9195 (N_9195,N_8095,N_8463);
nor U9196 (N_9196,N_8306,N_8405);
nand U9197 (N_9197,N_8430,N_8435);
nor U9198 (N_9198,N_8187,N_8471);
xor U9199 (N_9199,N_8229,N_8743);
xnor U9200 (N_9200,N_8641,N_8114);
and U9201 (N_9201,N_8750,N_8299);
xor U9202 (N_9202,N_8140,N_8507);
and U9203 (N_9203,N_8253,N_8319);
xnor U9204 (N_9204,N_8557,N_8701);
and U9205 (N_9205,N_8472,N_8059);
nand U9206 (N_9206,N_8721,N_8539);
nor U9207 (N_9207,N_8111,N_8474);
and U9208 (N_9208,N_8136,N_8655);
xor U9209 (N_9209,N_8560,N_8647);
nor U9210 (N_9210,N_8012,N_8163);
xnor U9211 (N_9211,N_8024,N_8312);
or U9212 (N_9212,N_8134,N_8618);
or U9213 (N_9213,N_8289,N_8032);
and U9214 (N_9214,N_8513,N_8226);
and U9215 (N_9215,N_8763,N_8465);
or U9216 (N_9216,N_8564,N_8101);
nor U9217 (N_9217,N_8648,N_8043);
nand U9218 (N_9218,N_8686,N_8428);
or U9219 (N_9219,N_8353,N_8515);
or U9220 (N_9220,N_8606,N_8660);
nand U9221 (N_9221,N_8284,N_8285);
or U9222 (N_9222,N_8013,N_8028);
and U9223 (N_9223,N_8532,N_8284);
nor U9224 (N_9224,N_8619,N_8334);
nand U9225 (N_9225,N_8732,N_8387);
xnor U9226 (N_9226,N_8240,N_8547);
nor U9227 (N_9227,N_8231,N_8079);
and U9228 (N_9228,N_8585,N_8713);
xor U9229 (N_9229,N_8411,N_8057);
nand U9230 (N_9230,N_8797,N_8389);
xnor U9231 (N_9231,N_8072,N_8714);
or U9232 (N_9232,N_8032,N_8231);
and U9233 (N_9233,N_8748,N_8329);
xor U9234 (N_9234,N_8131,N_8685);
nor U9235 (N_9235,N_8419,N_8482);
nor U9236 (N_9236,N_8779,N_8577);
nor U9237 (N_9237,N_8135,N_8415);
nand U9238 (N_9238,N_8403,N_8071);
nand U9239 (N_9239,N_8461,N_8146);
nor U9240 (N_9240,N_8648,N_8044);
and U9241 (N_9241,N_8070,N_8299);
xnor U9242 (N_9242,N_8718,N_8725);
xnor U9243 (N_9243,N_8156,N_8609);
and U9244 (N_9244,N_8317,N_8541);
nand U9245 (N_9245,N_8235,N_8681);
nand U9246 (N_9246,N_8087,N_8424);
xnor U9247 (N_9247,N_8031,N_8371);
xnor U9248 (N_9248,N_8425,N_8628);
or U9249 (N_9249,N_8658,N_8018);
nand U9250 (N_9250,N_8598,N_8241);
xor U9251 (N_9251,N_8680,N_8415);
or U9252 (N_9252,N_8619,N_8257);
or U9253 (N_9253,N_8432,N_8294);
and U9254 (N_9254,N_8017,N_8209);
xor U9255 (N_9255,N_8101,N_8702);
nor U9256 (N_9256,N_8495,N_8320);
nand U9257 (N_9257,N_8746,N_8101);
xor U9258 (N_9258,N_8273,N_8694);
and U9259 (N_9259,N_8138,N_8777);
xnor U9260 (N_9260,N_8424,N_8350);
or U9261 (N_9261,N_8748,N_8444);
or U9262 (N_9262,N_8361,N_8418);
or U9263 (N_9263,N_8393,N_8304);
and U9264 (N_9264,N_8765,N_8078);
or U9265 (N_9265,N_8224,N_8739);
nand U9266 (N_9266,N_8684,N_8308);
or U9267 (N_9267,N_8157,N_8764);
xnor U9268 (N_9268,N_8677,N_8010);
xnor U9269 (N_9269,N_8441,N_8083);
nor U9270 (N_9270,N_8173,N_8710);
and U9271 (N_9271,N_8228,N_8219);
nand U9272 (N_9272,N_8340,N_8743);
and U9273 (N_9273,N_8556,N_8345);
xnor U9274 (N_9274,N_8604,N_8658);
nor U9275 (N_9275,N_8091,N_8687);
and U9276 (N_9276,N_8595,N_8274);
nor U9277 (N_9277,N_8543,N_8635);
and U9278 (N_9278,N_8686,N_8206);
xnor U9279 (N_9279,N_8416,N_8223);
xnor U9280 (N_9280,N_8171,N_8638);
or U9281 (N_9281,N_8330,N_8642);
xnor U9282 (N_9282,N_8200,N_8411);
xnor U9283 (N_9283,N_8607,N_8703);
or U9284 (N_9284,N_8451,N_8732);
nor U9285 (N_9285,N_8171,N_8489);
and U9286 (N_9286,N_8322,N_8649);
xnor U9287 (N_9287,N_8068,N_8661);
nand U9288 (N_9288,N_8532,N_8370);
nand U9289 (N_9289,N_8605,N_8469);
nand U9290 (N_9290,N_8494,N_8304);
or U9291 (N_9291,N_8180,N_8355);
or U9292 (N_9292,N_8267,N_8609);
xnor U9293 (N_9293,N_8027,N_8441);
or U9294 (N_9294,N_8639,N_8604);
nand U9295 (N_9295,N_8637,N_8028);
and U9296 (N_9296,N_8086,N_8574);
xnor U9297 (N_9297,N_8424,N_8479);
and U9298 (N_9298,N_8425,N_8449);
xnor U9299 (N_9299,N_8395,N_8246);
or U9300 (N_9300,N_8638,N_8794);
nor U9301 (N_9301,N_8306,N_8145);
nor U9302 (N_9302,N_8347,N_8324);
nor U9303 (N_9303,N_8181,N_8696);
xor U9304 (N_9304,N_8311,N_8322);
or U9305 (N_9305,N_8100,N_8221);
nor U9306 (N_9306,N_8759,N_8428);
and U9307 (N_9307,N_8633,N_8180);
and U9308 (N_9308,N_8631,N_8379);
or U9309 (N_9309,N_8296,N_8560);
or U9310 (N_9310,N_8636,N_8344);
xnor U9311 (N_9311,N_8619,N_8188);
nand U9312 (N_9312,N_8714,N_8141);
nor U9313 (N_9313,N_8125,N_8044);
nand U9314 (N_9314,N_8722,N_8457);
xnor U9315 (N_9315,N_8596,N_8360);
or U9316 (N_9316,N_8091,N_8604);
nand U9317 (N_9317,N_8300,N_8164);
nor U9318 (N_9318,N_8233,N_8563);
xnor U9319 (N_9319,N_8341,N_8679);
and U9320 (N_9320,N_8488,N_8734);
xor U9321 (N_9321,N_8759,N_8584);
nor U9322 (N_9322,N_8046,N_8475);
nor U9323 (N_9323,N_8265,N_8581);
nor U9324 (N_9324,N_8786,N_8700);
or U9325 (N_9325,N_8649,N_8314);
nand U9326 (N_9326,N_8469,N_8411);
nand U9327 (N_9327,N_8560,N_8248);
nand U9328 (N_9328,N_8027,N_8224);
xnor U9329 (N_9329,N_8452,N_8127);
or U9330 (N_9330,N_8509,N_8204);
nor U9331 (N_9331,N_8354,N_8048);
or U9332 (N_9332,N_8730,N_8377);
nor U9333 (N_9333,N_8118,N_8528);
or U9334 (N_9334,N_8628,N_8096);
and U9335 (N_9335,N_8178,N_8785);
nand U9336 (N_9336,N_8741,N_8398);
nor U9337 (N_9337,N_8604,N_8227);
xnor U9338 (N_9338,N_8262,N_8318);
nor U9339 (N_9339,N_8238,N_8416);
nor U9340 (N_9340,N_8429,N_8786);
or U9341 (N_9341,N_8066,N_8266);
nand U9342 (N_9342,N_8071,N_8212);
nand U9343 (N_9343,N_8516,N_8284);
nand U9344 (N_9344,N_8355,N_8244);
nand U9345 (N_9345,N_8439,N_8032);
and U9346 (N_9346,N_8362,N_8517);
xor U9347 (N_9347,N_8718,N_8260);
nor U9348 (N_9348,N_8294,N_8125);
and U9349 (N_9349,N_8551,N_8394);
nand U9350 (N_9350,N_8649,N_8101);
nand U9351 (N_9351,N_8500,N_8793);
nor U9352 (N_9352,N_8052,N_8547);
nor U9353 (N_9353,N_8759,N_8794);
nor U9354 (N_9354,N_8237,N_8234);
and U9355 (N_9355,N_8248,N_8231);
and U9356 (N_9356,N_8113,N_8649);
nand U9357 (N_9357,N_8041,N_8118);
nor U9358 (N_9358,N_8249,N_8316);
nand U9359 (N_9359,N_8477,N_8062);
nand U9360 (N_9360,N_8475,N_8147);
nand U9361 (N_9361,N_8769,N_8092);
xnor U9362 (N_9362,N_8439,N_8713);
nor U9363 (N_9363,N_8086,N_8448);
nand U9364 (N_9364,N_8606,N_8748);
nand U9365 (N_9365,N_8626,N_8113);
and U9366 (N_9366,N_8749,N_8243);
or U9367 (N_9367,N_8755,N_8788);
or U9368 (N_9368,N_8748,N_8559);
xnor U9369 (N_9369,N_8321,N_8302);
nand U9370 (N_9370,N_8322,N_8782);
nand U9371 (N_9371,N_8384,N_8411);
nor U9372 (N_9372,N_8585,N_8006);
xnor U9373 (N_9373,N_8318,N_8731);
and U9374 (N_9374,N_8462,N_8121);
xor U9375 (N_9375,N_8195,N_8361);
or U9376 (N_9376,N_8103,N_8519);
xnor U9377 (N_9377,N_8538,N_8096);
nor U9378 (N_9378,N_8763,N_8326);
nand U9379 (N_9379,N_8479,N_8475);
nor U9380 (N_9380,N_8702,N_8110);
and U9381 (N_9381,N_8042,N_8238);
nor U9382 (N_9382,N_8466,N_8478);
and U9383 (N_9383,N_8567,N_8464);
nor U9384 (N_9384,N_8478,N_8319);
nand U9385 (N_9385,N_8466,N_8615);
or U9386 (N_9386,N_8649,N_8065);
nand U9387 (N_9387,N_8215,N_8218);
and U9388 (N_9388,N_8719,N_8154);
or U9389 (N_9389,N_8507,N_8519);
xor U9390 (N_9390,N_8457,N_8522);
xnor U9391 (N_9391,N_8074,N_8186);
and U9392 (N_9392,N_8324,N_8153);
and U9393 (N_9393,N_8201,N_8517);
or U9394 (N_9394,N_8668,N_8122);
or U9395 (N_9395,N_8487,N_8767);
nor U9396 (N_9396,N_8685,N_8391);
xnor U9397 (N_9397,N_8721,N_8009);
nand U9398 (N_9398,N_8449,N_8424);
xnor U9399 (N_9399,N_8297,N_8463);
or U9400 (N_9400,N_8036,N_8332);
or U9401 (N_9401,N_8462,N_8034);
nand U9402 (N_9402,N_8531,N_8078);
and U9403 (N_9403,N_8585,N_8623);
nand U9404 (N_9404,N_8045,N_8438);
xnor U9405 (N_9405,N_8728,N_8602);
and U9406 (N_9406,N_8141,N_8606);
nand U9407 (N_9407,N_8212,N_8746);
nor U9408 (N_9408,N_8103,N_8773);
and U9409 (N_9409,N_8660,N_8083);
nor U9410 (N_9410,N_8586,N_8256);
and U9411 (N_9411,N_8035,N_8257);
nand U9412 (N_9412,N_8075,N_8149);
or U9413 (N_9413,N_8281,N_8531);
nor U9414 (N_9414,N_8679,N_8466);
nand U9415 (N_9415,N_8181,N_8044);
xnor U9416 (N_9416,N_8305,N_8753);
nand U9417 (N_9417,N_8064,N_8096);
nor U9418 (N_9418,N_8166,N_8036);
xor U9419 (N_9419,N_8212,N_8272);
or U9420 (N_9420,N_8535,N_8251);
nand U9421 (N_9421,N_8639,N_8281);
nor U9422 (N_9422,N_8548,N_8658);
nor U9423 (N_9423,N_8233,N_8513);
nand U9424 (N_9424,N_8706,N_8655);
nor U9425 (N_9425,N_8218,N_8191);
nor U9426 (N_9426,N_8304,N_8569);
xnor U9427 (N_9427,N_8022,N_8632);
nor U9428 (N_9428,N_8644,N_8169);
xor U9429 (N_9429,N_8215,N_8666);
or U9430 (N_9430,N_8432,N_8309);
or U9431 (N_9431,N_8265,N_8122);
or U9432 (N_9432,N_8287,N_8653);
nand U9433 (N_9433,N_8236,N_8136);
or U9434 (N_9434,N_8663,N_8199);
xnor U9435 (N_9435,N_8299,N_8125);
nor U9436 (N_9436,N_8475,N_8027);
nor U9437 (N_9437,N_8373,N_8366);
or U9438 (N_9438,N_8419,N_8709);
and U9439 (N_9439,N_8143,N_8085);
and U9440 (N_9440,N_8595,N_8249);
or U9441 (N_9441,N_8510,N_8293);
and U9442 (N_9442,N_8254,N_8157);
and U9443 (N_9443,N_8772,N_8550);
xnor U9444 (N_9444,N_8717,N_8158);
nand U9445 (N_9445,N_8118,N_8065);
nand U9446 (N_9446,N_8251,N_8370);
or U9447 (N_9447,N_8424,N_8437);
nor U9448 (N_9448,N_8508,N_8620);
nand U9449 (N_9449,N_8210,N_8599);
xor U9450 (N_9450,N_8198,N_8300);
or U9451 (N_9451,N_8663,N_8059);
or U9452 (N_9452,N_8441,N_8294);
and U9453 (N_9453,N_8716,N_8002);
nand U9454 (N_9454,N_8553,N_8254);
nor U9455 (N_9455,N_8642,N_8533);
xor U9456 (N_9456,N_8714,N_8306);
xnor U9457 (N_9457,N_8645,N_8187);
xor U9458 (N_9458,N_8785,N_8774);
or U9459 (N_9459,N_8708,N_8382);
nor U9460 (N_9460,N_8288,N_8352);
xnor U9461 (N_9461,N_8395,N_8226);
nor U9462 (N_9462,N_8272,N_8131);
nor U9463 (N_9463,N_8622,N_8581);
nand U9464 (N_9464,N_8345,N_8532);
nor U9465 (N_9465,N_8280,N_8731);
and U9466 (N_9466,N_8678,N_8726);
nor U9467 (N_9467,N_8463,N_8791);
nand U9468 (N_9468,N_8672,N_8509);
xnor U9469 (N_9469,N_8536,N_8447);
and U9470 (N_9470,N_8196,N_8403);
and U9471 (N_9471,N_8139,N_8448);
nor U9472 (N_9472,N_8056,N_8162);
or U9473 (N_9473,N_8561,N_8025);
xor U9474 (N_9474,N_8067,N_8362);
or U9475 (N_9475,N_8323,N_8683);
nand U9476 (N_9476,N_8161,N_8533);
nor U9477 (N_9477,N_8299,N_8435);
and U9478 (N_9478,N_8769,N_8231);
and U9479 (N_9479,N_8503,N_8248);
and U9480 (N_9480,N_8158,N_8092);
or U9481 (N_9481,N_8757,N_8278);
nand U9482 (N_9482,N_8564,N_8352);
nand U9483 (N_9483,N_8046,N_8102);
nand U9484 (N_9484,N_8235,N_8388);
nand U9485 (N_9485,N_8785,N_8640);
nor U9486 (N_9486,N_8722,N_8176);
xor U9487 (N_9487,N_8433,N_8748);
xor U9488 (N_9488,N_8292,N_8235);
and U9489 (N_9489,N_8047,N_8580);
nand U9490 (N_9490,N_8503,N_8142);
nand U9491 (N_9491,N_8174,N_8254);
or U9492 (N_9492,N_8725,N_8198);
and U9493 (N_9493,N_8189,N_8518);
or U9494 (N_9494,N_8510,N_8097);
and U9495 (N_9495,N_8032,N_8278);
or U9496 (N_9496,N_8304,N_8593);
or U9497 (N_9497,N_8719,N_8780);
or U9498 (N_9498,N_8438,N_8053);
xnor U9499 (N_9499,N_8419,N_8034);
and U9500 (N_9500,N_8203,N_8128);
xor U9501 (N_9501,N_8278,N_8471);
xor U9502 (N_9502,N_8459,N_8798);
or U9503 (N_9503,N_8083,N_8727);
nand U9504 (N_9504,N_8357,N_8724);
or U9505 (N_9505,N_8648,N_8523);
and U9506 (N_9506,N_8301,N_8161);
and U9507 (N_9507,N_8169,N_8495);
or U9508 (N_9508,N_8040,N_8745);
xnor U9509 (N_9509,N_8308,N_8353);
or U9510 (N_9510,N_8356,N_8722);
and U9511 (N_9511,N_8243,N_8495);
nand U9512 (N_9512,N_8691,N_8576);
and U9513 (N_9513,N_8474,N_8052);
or U9514 (N_9514,N_8148,N_8270);
nand U9515 (N_9515,N_8276,N_8151);
nand U9516 (N_9516,N_8247,N_8654);
nand U9517 (N_9517,N_8013,N_8274);
nor U9518 (N_9518,N_8456,N_8352);
and U9519 (N_9519,N_8562,N_8128);
nand U9520 (N_9520,N_8601,N_8385);
and U9521 (N_9521,N_8763,N_8466);
and U9522 (N_9522,N_8783,N_8325);
and U9523 (N_9523,N_8668,N_8796);
nor U9524 (N_9524,N_8325,N_8227);
nor U9525 (N_9525,N_8456,N_8628);
nand U9526 (N_9526,N_8592,N_8249);
and U9527 (N_9527,N_8138,N_8209);
and U9528 (N_9528,N_8341,N_8054);
or U9529 (N_9529,N_8580,N_8277);
nor U9530 (N_9530,N_8423,N_8477);
nor U9531 (N_9531,N_8056,N_8088);
nand U9532 (N_9532,N_8675,N_8271);
xnor U9533 (N_9533,N_8592,N_8578);
and U9534 (N_9534,N_8080,N_8063);
and U9535 (N_9535,N_8181,N_8749);
or U9536 (N_9536,N_8295,N_8145);
xor U9537 (N_9537,N_8219,N_8444);
xnor U9538 (N_9538,N_8450,N_8017);
or U9539 (N_9539,N_8143,N_8372);
and U9540 (N_9540,N_8466,N_8087);
nand U9541 (N_9541,N_8406,N_8325);
and U9542 (N_9542,N_8672,N_8192);
or U9543 (N_9543,N_8476,N_8704);
and U9544 (N_9544,N_8432,N_8755);
or U9545 (N_9545,N_8116,N_8750);
nand U9546 (N_9546,N_8740,N_8781);
nand U9547 (N_9547,N_8356,N_8703);
xnor U9548 (N_9548,N_8133,N_8430);
xor U9549 (N_9549,N_8049,N_8555);
and U9550 (N_9550,N_8114,N_8608);
and U9551 (N_9551,N_8253,N_8179);
nand U9552 (N_9552,N_8509,N_8317);
or U9553 (N_9553,N_8587,N_8430);
nand U9554 (N_9554,N_8086,N_8303);
or U9555 (N_9555,N_8130,N_8250);
nand U9556 (N_9556,N_8264,N_8724);
nand U9557 (N_9557,N_8102,N_8754);
nor U9558 (N_9558,N_8317,N_8338);
nand U9559 (N_9559,N_8177,N_8146);
or U9560 (N_9560,N_8743,N_8626);
or U9561 (N_9561,N_8681,N_8364);
nand U9562 (N_9562,N_8345,N_8486);
xor U9563 (N_9563,N_8024,N_8122);
nand U9564 (N_9564,N_8348,N_8267);
or U9565 (N_9565,N_8728,N_8637);
nand U9566 (N_9566,N_8694,N_8642);
xor U9567 (N_9567,N_8273,N_8435);
nor U9568 (N_9568,N_8055,N_8185);
or U9569 (N_9569,N_8166,N_8319);
and U9570 (N_9570,N_8372,N_8496);
nand U9571 (N_9571,N_8544,N_8402);
nor U9572 (N_9572,N_8372,N_8121);
nand U9573 (N_9573,N_8200,N_8198);
and U9574 (N_9574,N_8786,N_8150);
xor U9575 (N_9575,N_8051,N_8480);
nand U9576 (N_9576,N_8773,N_8763);
nor U9577 (N_9577,N_8574,N_8290);
and U9578 (N_9578,N_8312,N_8125);
and U9579 (N_9579,N_8438,N_8690);
and U9580 (N_9580,N_8396,N_8505);
xor U9581 (N_9581,N_8123,N_8689);
nor U9582 (N_9582,N_8237,N_8735);
xor U9583 (N_9583,N_8731,N_8290);
and U9584 (N_9584,N_8443,N_8165);
nand U9585 (N_9585,N_8718,N_8201);
nor U9586 (N_9586,N_8261,N_8738);
or U9587 (N_9587,N_8011,N_8166);
nand U9588 (N_9588,N_8215,N_8480);
nand U9589 (N_9589,N_8489,N_8033);
nor U9590 (N_9590,N_8493,N_8284);
or U9591 (N_9591,N_8247,N_8073);
or U9592 (N_9592,N_8713,N_8651);
and U9593 (N_9593,N_8604,N_8190);
or U9594 (N_9594,N_8634,N_8606);
nor U9595 (N_9595,N_8678,N_8580);
nand U9596 (N_9596,N_8136,N_8491);
xnor U9597 (N_9597,N_8748,N_8491);
nor U9598 (N_9598,N_8071,N_8509);
nor U9599 (N_9599,N_8200,N_8576);
or U9600 (N_9600,N_8808,N_9333);
nand U9601 (N_9601,N_9045,N_9559);
nand U9602 (N_9602,N_8812,N_9195);
and U9603 (N_9603,N_9336,N_9399);
or U9604 (N_9604,N_9083,N_9299);
and U9605 (N_9605,N_9109,N_8986);
nand U9606 (N_9606,N_9519,N_9452);
or U9607 (N_9607,N_9079,N_9078);
or U9608 (N_9608,N_9408,N_9551);
and U9609 (N_9609,N_8824,N_8973);
nor U9610 (N_9610,N_9245,N_9449);
nor U9611 (N_9611,N_9517,N_9252);
and U9612 (N_9612,N_9190,N_9343);
or U9613 (N_9613,N_8977,N_8974);
and U9614 (N_9614,N_9272,N_8911);
or U9615 (N_9615,N_9447,N_8930);
and U9616 (N_9616,N_8840,N_9342);
nand U9617 (N_9617,N_9143,N_9367);
and U9618 (N_9618,N_8952,N_9063);
nor U9619 (N_9619,N_9315,N_9579);
xor U9620 (N_9620,N_9217,N_9129);
nand U9621 (N_9621,N_8941,N_9588);
nand U9622 (N_9622,N_9318,N_9265);
nor U9623 (N_9623,N_9193,N_9160);
nor U9624 (N_9624,N_9550,N_9199);
nand U9625 (N_9625,N_9073,N_9284);
nor U9626 (N_9626,N_9084,N_9498);
nor U9627 (N_9627,N_8886,N_9308);
or U9628 (N_9628,N_9472,N_9556);
nand U9629 (N_9629,N_8942,N_9263);
or U9630 (N_9630,N_8855,N_9506);
nor U9631 (N_9631,N_9025,N_9071);
or U9632 (N_9632,N_9441,N_9355);
nand U9633 (N_9633,N_9339,N_9224);
nand U9634 (N_9634,N_9474,N_9326);
xnor U9635 (N_9635,N_8932,N_9554);
nor U9636 (N_9636,N_9286,N_9391);
nor U9637 (N_9637,N_8921,N_9317);
nor U9638 (N_9638,N_8811,N_9323);
nor U9639 (N_9639,N_9487,N_8815);
nor U9640 (N_9640,N_8972,N_8806);
or U9641 (N_9641,N_9570,N_9510);
or U9642 (N_9642,N_9275,N_8926);
nor U9643 (N_9643,N_8990,N_8865);
or U9644 (N_9644,N_9163,N_9139);
and U9645 (N_9645,N_9029,N_9241);
and U9646 (N_9646,N_9102,N_8881);
xnor U9647 (N_9647,N_9370,N_9553);
nand U9648 (N_9648,N_8891,N_9536);
xnor U9649 (N_9649,N_9405,N_9234);
nand U9650 (N_9650,N_9122,N_9259);
nand U9651 (N_9651,N_9352,N_9169);
and U9652 (N_9652,N_9401,N_9386);
and U9653 (N_9653,N_9277,N_8982);
nor U9654 (N_9654,N_9431,N_9457);
nor U9655 (N_9655,N_9219,N_9243);
and U9656 (N_9656,N_9194,N_8895);
or U9657 (N_9657,N_8831,N_9146);
nand U9658 (N_9658,N_8861,N_9499);
xor U9659 (N_9659,N_9125,N_8801);
and U9660 (N_9660,N_9177,N_9189);
nor U9661 (N_9661,N_9521,N_9548);
xor U9662 (N_9662,N_9019,N_9211);
nor U9663 (N_9663,N_9206,N_9101);
or U9664 (N_9664,N_9053,N_9276);
nand U9665 (N_9665,N_9095,N_9170);
xor U9666 (N_9666,N_9520,N_9423);
nor U9667 (N_9667,N_9330,N_8864);
or U9668 (N_9668,N_9356,N_9113);
xnor U9669 (N_9669,N_9172,N_8838);
xor U9670 (N_9670,N_9329,N_9027);
xor U9671 (N_9671,N_9422,N_9372);
xor U9672 (N_9672,N_9127,N_8910);
nand U9673 (N_9673,N_9228,N_9567);
or U9674 (N_9674,N_9145,N_8892);
xnor U9675 (N_9675,N_9003,N_9017);
nand U9676 (N_9676,N_9018,N_8960);
nand U9677 (N_9677,N_9363,N_8913);
or U9678 (N_9678,N_9124,N_9512);
xnor U9679 (N_9679,N_9131,N_9229);
xor U9680 (N_9680,N_9320,N_9419);
and U9681 (N_9681,N_9142,N_9054);
and U9682 (N_9682,N_8834,N_8877);
xnor U9683 (N_9683,N_9393,N_9009);
nor U9684 (N_9684,N_9007,N_8897);
or U9685 (N_9685,N_9440,N_9255);
and U9686 (N_9686,N_9473,N_8890);
or U9687 (N_9687,N_9133,N_8968);
and U9688 (N_9688,N_9532,N_9198);
and U9689 (N_9689,N_9087,N_9149);
nand U9690 (N_9690,N_9258,N_9011);
xor U9691 (N_9691,N_9392,N_8872);
and U9692 (N_9692,N_8965,N_8916);
xor U9693 (N_9693,N_9060,N_9545);
and U9694 (N_9694,N_9591,N_9507);
nand U9695 (N_9695,N_9335,N_8918);
nand U9696 (N_9696,N_8951,N_8843);
nor U9697 (N_9697,N_9130,N_8820);
and U9698 (N_9698,N_9508,N_9213);
nor U9699 (N_9699,N_9572,N_9436);
xnor U9700 (N_9700,N_9119,N_9240);
and U9701 (N_9701,N_8888,N_8813);
nor U9702 (N_9702,N_8802,N_9106);
nand U9703 (N_9703,N_9411,N_9068);
or U9704 (N_9704,N_9048,N_8807);
nand U9705 (N_9705,N_9446,N_9467);
and U9706 (N_9706,N_8847,N_9218);
nor U9707 (N_9707,N_9069,N_9171);
nor U9708 (N_9708,N_9503,N_8809);
xnor U9709 (N_9709,N_9256,N_9385);
nor U9710 (N_9710,N_9033,N_8887);
and U9711 (N_9711,N_9103,N_9400);
nand U9712 (N_9712,N_9395,N_9024);
nand U9713 (N_9713,N_9042,N_9469);
or U9714 (N_9714,N_9088,N_9114);
or U9715 (N_9715,N_9464,N_9438);
xor U9716 (N_9716,N_9388,N_8849);
nor U9717 (N_9717,N_8954,N_9120);
or U9718 (N_9718,N_9273,N_9135);
xor U9719 (N_9719,N_8814,N_9126);
or U9720 (N_9720,N_9055,N_9344);
nand U9721 (N_9721,N_9562,N_9590);
or U9722 (N_9722,N_9274,N_9349);
nor U9723 (N_9723,N_9182,N_9346);
nand U9724 (N_9724,N_9176,N_9140);
nor U9725 (N_9725,N_9107,N_8837);
and U9726 (N_9726,N_9471,N_9597);
and U9727 (N_9727,N_9000,N_9051);
nand U9728 (N_9728,N_9123,N_9062);
or U9729 (N_9729,N_9537,N_9242);
xor U9730 (N_9730,N_9369,N_9093);
nor U9731 (N_9731,N_9075,N_8870);
and U9732 (N_9732,N_9233,N_9478);
nor U9733 (N_9733,N_8922,N_9066);
nand U9734 (N_9734,N_9207,N_9340);
nand U9735 (N_9735,N_9092,N_9465);
nand U9736 (N_9736,N_9566,N_9387);
and U9737 (N_9737,N_8854,N_9424);
nand U9738 (N_9738,N_8901,N_8874);
or U9739 (N_9739,N_9410,N_8860);
xnor U9740 (N_9740,N_9070,N_9137);
nand U9741 (N_9741,N_9046,N_9505);
or U9742 (N_9742,N_9351,N_8884);
nor U9743 (N_9743,N_8955,N_9525);
xnor U9744 (N_9744,N_9492,N_9489);
nand U9745 (N_9745,N_9496,N_9157);
or U9746 (N_9746,N_9244,N_9303);
or U9747 (N_9747,N_9064,N_9509);
xnor U9748 (N_9748,N_9577,N_9294);
nand U9749 (N_9749,N_9268,N_8876);
nand U9750 (N_9750,N_8915,N_9511);
xor U9751 (N_9751,N_9461,N_8894);
nor U9752 (N_9752,N_9350,N_8819);
or U9753 (N_9753,N_9292,N_9166);
xnor U9754 (N_9754,N_9576,N_8856);
or U9755 (N_9755,N_9573,N_8800);
and U9756 (N_9756,N_8833,N_9013);
or U9757 (N_9757,N_9281,N_9426);
nand U9758 (N_9758,N_8970,N_9050);
nor U9759 (N_9759,N_9183,N_9044);
nor U9760 (N_9760,N_9141,N_8904);
nand U9761 (N_9761,N_9155,N_9375);
xnor U9762 (N_9762,N_9210,N_8844);
nor U9763 (N_9763,N_9186,N_8853);
nor U9764 (N_9764,N_9285,N_9321);
and U9765 (N_9765,N_9491,N_9152);
nand U9766 (N_9766,N_9026,N_9100);
nor U9767 (N_9767,N_9112,N_9501);
nor U9768 (N_9768,N_9184,N_9288);
or U9769 (N_9769,N_9500,N_9082);
or U9770 (N_9770,N_8994,N_9444);
nor U9771 (N_9771,N_9547,N_9090);
nor U9772 (N_9772,N_9454,N_8832);
nor U9773 (N_9773,N_9202,N_9104);
nor U9774 (N_9774,N_8989,N_9533);
xor U9775 (N_9775,N_9428,N_8940);
or U9776 (N_9776,N_8944,N_9527);
xnor U9777 (N_9777,N_8917,N_9307);
or U9778 (N_9778,N_8927,N_9121);
nand U9779 (N_9779,N_9014,N_8842);
or U9780 (N_9780,N_9589,N_8803);
or U9781 (N_9781,N_9209,N_8938);
xnor U9782 (N_9782,N_9040,N_9514);
or U9783 (N_9783,N_9164,N_8804);
and U9784 (N_9784,N_9413,N_8988);
nor U9785 (N_9785,N_8909,N_9204);
or U9786 (N_9786,N_9089,N_9222);
nor U9787 (N_9787,N_9582,N_8950);
and U9788 (N_9788,N_8903,N_9175);
or U9789 (N_9789,N_9598,N_9065);
and U9790 (N_9790,N_9593,N_9168);
and U9791 (N_9791,N_9057,N_8871);
nand U9792 (N_9792,N_9552,N_9384);
nand U9793 (N_9793,N_8948,N_8983);
nor U9794 (N_9794,N_9358,N_8992);
xnor U9795 (N_9795,N_9235,N_8868);
and U9796 (N_9796,N_9008,N_9322);
and U9797 (N_9797,N_9522,N_9460);
nor U9798 (N_9798,N_9279,N_9015);
xor U9799 (N_9799,N_8829,N_9364);
xnor U9800 (N_9800,N_8996,N_8902);
and U9801 (N_9801,N_9156,N_9403);
nor U9802 (N_9802,N_8835,N_9434);
nand U9803 (N_9803,N_9291,N_9493);
and U9804 (N_9804,N_9254,N_8893);
and U9805 (N_9805,N_9477,N_9154);
or U9806 (N_9806,N_9542,N_8905);
xnor U9807 (N_9807,N_9382,N_9036);
and U9808 (N_9808,N_9442,N_8979);
nor U9809 (N_9809,N_9283,N_9415);
or U9810 (N_9810,N_9455,N_9325);
xnor U9811 (N_9811,N_9076,N_9420);
or U9812 (N_9812,N_8963,N_9594);
and U9813 (N_9813,N_9074,N_9586);
nand U9814 (N_9814,N_9389,N_8830);
nor U9815 (N_9815,N_8980,N_9353);
xnor U9816 (N_9816,N_8866,N_9041);
and U9817 (N_9817,N_9304,N_9497);
and U9818 (N_9818,N_9030,N_9324);
xor U9819 (N_9819,N_9249,N_8878);
or U9820 (N_9820,N_9429,N_9354);
or U9821 (N_9821,N_9257,N_8810);
nor U9822 (N_9822,N_9380,N_9584);
and U9823 (N_9823,N_9581,N_9407);
and U9824 (N_9824,N_9147,N_9148);
nand U9825 (N_9825,N_9309,N_9376);
nand U9826 (N_9826,N_9298,N_8969);
and U9827 (N_9827,N_9490,N_8880);
or U9828 (N_9828,N_9362,N_8859);
nor U9829 (N_9829,N_9230,N_8869);
or U9830 (N_9830,N_9031,N_9338);
nand U9831 (N_9831,N_8998,N_9223);
xor U9832 (N_9832,N_8867,N_9301);
nand U9833 (N_9833,N_9479,N_8934);
or U9834 (N_9834,N_9359,N_8959);
nor U9835 (N_9835,N_9115,N_9270);
nor U9836 (N_9836,N_9214,N_8999);
nor U9837 (N_9837,N_8825,N_9005);
nand U9838 (N_9838,N_9397,N_9248);
nor U9839 (N_9839,N_8845,N_8997);
nor U9840 (N_9840,N_9578,N_9374);
and U9841 (N_9841,N_9287,N_9534);
and U9842 (N_9842,N_9328,N_9221);
or U9843 (N_9843,N_8828,N_9049);
or U9844 (N_9844,N_9456,N_9494);
nand U9845 (N_9845,N_9406,N_9016);
nand U9846 (N_9846,N_9485,N_9312);
xor U9847 (N_9847,N_9531,N_9067);
and U9848 (N_9848,N_9368,N_9515);
or U9849 (N_9849,N_8981,N_8975);
xnor U9850 (N_9850,N_8826,N_9379);
nand U9851 (N_9851,N_8967,N_8857);
nand U9852 (N_9852,N_8827,N_8852);
xor U9853 (N_9853,N_8816,N_9282);
and U9854 (N_9854,N_9047,N_9111);
and U9855 (N_9855,N_9251,N_9231);
and U9856 (N_9856,N_9377,N_9458);
and U9857 (N_9857,N_8907,N_9022);
nor U9858 (N_9858,N_9038,N_9271);
and U9859 (N_9859,N_9425,N_9002);
and U9860 (N_9860,N_9185,N_9430);
xor U9861 (N_9861,N_9563,N_9037);
xnor U9862 (N_9862,N_9574,N_9568);
xnor U9863 (N_9863,N_8836,N_8889);
and U9864 (N_9864,N_9541,N_8933);
and U9865 (N_9865,N_8985,N_9437);
and U9866 (N_9866,N_8906,N_8945);
nand U9867 (N_9867,N_9390,N_9529);
nor U9868 (N_9868,N_9365,N_9159);
xnor U9869 (N_9869,N_9319,N_9094);
xor U9870 (N_9870,N_8898,N_9151);
xnor U9871 (N_9871,N_9345,N_9313);
nor U9872 (N_9872,N_9099,N_8912);
and U9873 (N_9873,N_9560,N_9488);
nor U9874 (N_9874,N_9311,N_9227);
nor U9875 (N_9875,N_9250,N_9052);
or U9876 (N_9876,N_9561,N_9264);
and U9877 (N_9877,N_9295,N_9158);
nor U9878 (N_9878,N_9238,N_9072);
nor U9879 (N_9879,N_8882,N_9450);
xnor U9880 (N_9880,N_9086,N_9153);
nand U9881 (N_9881,N_9435,N_9096);
nand U9882 (N_9882,N_9417,N_9571);
nand U9883 (N_9883,N_9475,N_9439);
nand U9884 (N_9884,N_8962,N_9549);
nor U9885 (N_9885,N_9144,N_9236);
nor U9886 (N_9886,N_9451,N_9381);
or U9887 (N_9887,N_9061,N_9305);
nand U9888 (N_9888,N_8935,N_9371);
nand U9889 (N_9889,N_9077,N_9278);
nor U9890 (N_9890,N_9530,N_9043);
nor U9891 (N_9891,N_9482,N_9513);
nor U9892 (N_9892,N_9179,N_9544);
nor U9893 (N_9893,N_9128,N_9575);
nand U9894 (N_9894,N_9416,N_9341);
or U9895 (N_9895,N_8931,N_9565);
xor U9896 (N_9896,N_9178,N_8956);
or U9897 (N_9897,N_9289,N_9136);
or U9898 (N_9898,N_9538,N_8851);
nor U9899 (N_9899,N_9188,N_9595);
nor U9900 (N_9900,N_9020,N_9010);
nand U9901 (N_9901,N_8805,N_9587);
nor U9902 (N_9902,N_8966,N_9483);
nand U9903 (N_9903,N_9059,N_9348);
and U9904 (N_9904,N_9476,N_9481);
xnor U9905 (N_9905,N_9528,N_9518);
xor U9906 (N_9906,N_9486,N_9132);
nor U9907 (N_9907,N_8929,N_8991);
nand U9908 (N_9908,N_9220,N_9334);
nand U9909 (N_9909,N_8961,N_8964);
and U9910 (N_9910,N_8925,N_9216);
or U9911 (N_9911,N_8818,N_9203);
and U9912 (N_9912,N_8993,N_9433);
or U9913 (N_9913,N_9269,N_9260);
nor U9914 (N_9914,N_8846,N_9585);
and U9915 (N_9915,N_9280,N_9332);
or U9916 (N_9916,N_9331,N_8937);
xor U9917 (N_9917,N_8896,N_8821);
nand U9918 (N_9918,N_9200,N_9357);
and U9919 (N_9919,N_8908,N_8875);
or U9920 (N_9920,N_9173,N_9596);
or U9921 (N_9921,N_9253,N_8971);
or U9922 (N_9922,N_9085,N_9028);
or U9923 (N_9923,N_9012,N_9310);
nor U9924 (N_9924,N_9197,N_9599);
xnor U9925 (N_9925,N_9466,N_8885);
and U9926 (N_9926,N_8883,N_9558);
nand U9927 (N_9927,N_8946,N_9502);
nor U9928 (N_9928,N_9162,N_9056);
and U9929 (N_9929,N_9316,N_9187);
or U9930 (N_9930,N_9138,N_9196);
or U9931 (N_9931,N_9246,N_9443);
xnor U9932 (N_9932,N_8848,N_9232);
or U9933 (N_9933,N_9418,N_9383);
and U9934 (N_9934,N_8899,N_8823);
nor U9935 (N_9935,N_9080,N_9373);
nor U9936 (N_9936,N_9004,N_9174);
xor U9937 (N_9937,N_8923,N_8939);
and U9938 (N_9938,N_9445,N_9237);
nor U9939 (N_9939,N_8943,N_9239);
nor U9940 (N_9940,N_9361,N_9448);
xnor U9941 (N_9941,N_9539,N_9409);
or U9942 (N_9942,N_9314,N_9524);
nor U9943 (N_9943,N_9215,N_9212);
or U9944 (N_9944,N_8817,N_9463);
nor U9945 (N_9945,N_9180,N_9366);
xor U9946 (N_9946,N_8862,N_8919);
xor U9947 (N_9947,N_9167,N_9580);
xor U9948 (N_9948,N_9404,N_8957);
nor U9949 (N_9949,N_9592,N_9226);
or U9950 (N_9950,N_9564,N_9347);
nand U9951 (N_9951,N_9150,N_9470);
nor U9952 (N_9952,N_8850,N_9297);
xor U9953 (N_9953,N_9327,N_9098);
xnor U9954 (N_9954,N_8976,N_9006);
xor U9955 (N_9955,N_8879,N_9504);
xnor U9956 (N_9956,N_9484,N_9421);
nor U9957 (N_9957,N_9396,N_9480);
nand U9958 (N_9958,N_9021,N_9118);
and U9959 (N_9959,N_9266,N_9290);
nor U9960 (N_9960,N_9453,N_8928);
nand U9961 (N_9961,N_8873,N_9191);
nand U9962 (N_9962,N_9495,N_9205);
nand U9963 (N_9963,N_9555,N_9097);
xnor U9964 (N_9964,N_9360,N_9540);
or U9965 (N_9965,N_9181,N_9557);
nor U9966 (N_9966,N_9569,N_8841);
nand U9967 (N_9967,N_9034,N_9058);
or U9968 (N_9968,N_8978,N_9394);
and U9969 (N_9969,N_8920,N_9001);
or U9970 (N_9970,N_8900,N_9108);
xor U9971 (N_9971,N_9402,N_8953);
xnor U9972 (N_9972,N_9300,N_9201);
xor U9973 (N_9973,N_8839,N_8987);
nand U9974 (N_9974,N_9546,N_9516);
nand U9975 (N_9975,N_9023,N_9117);
and U9976 (N_9976,N_9432,N_8924);
nor U9977 (N_9977,N_9105,N_9208);
xor U9978 (N_9978,N_9293,N_9091);
and U9979 (N_9979,N_9296,N_9414);
and U9980 (N_9980,N_8949,N_9523);
nand U9981 (N_9981,N_9459,N_9412);
and U9982 (N_9982,N_8958,N_9116);
xnor U9983 (N_9983,N_9306,N_9262);
or U9984 (N_9984,N_9427,N_8822);
nand U9985 (N_9985,N_8914,N_9134);
xnor U9986 (N_9986,N_9247,N_9225);
and U9987 (N_9987,N_9267,N_9302);
nor U9988 (N_9988,N_9110,N_9032);
and U9989 (N_9989,N_8936,N_9468);
nand U9990 (N_9990,N_9378,N_8858);
xor U9991 (N_9991,N_9081,N_9398);
or U9992 (N_9992,N_9165,N_8947);
nand U9993 (N_9993,N_9526,N_9337);
or U9994 (N_9994,N_9535,N_9161);
nand U9995 (N_9995,N_8984,N_9543);
xnor U9996 (N_9996,N_9192,N_9583);
xnor U9997 (N_9997,N_9039,N_9035);
xnor U9998 (N_9998,N_8863,N_9261);
xnor U9999 (N_9999,N_8995,N_9462);
xnor U10000 (N_10000,N_9097,N_9058);
nand U10001 (N_10001,N_9115,N_9030);
nand U10002 (N_10002,N_9113,N_9435);
nor U10003 (N_10003,N_9292,N_9293);
xor U10004 (N_10004,N_9052,N_9210);
or U10005 (N_10005,N_9341,N_9500);
nor U10006 (N_10006,N_9416,N_8813);
nor U10007 (N_10007,N_8966,N_8915);
and U10008 (N_10008,N_9348,N_9439);
xnor U10009 (N_10009,N_9375,N_8910);
nor U10010 (N_10010,N_9232,N_9184);
nor U10011 (N_10011,N_9217,N_9236);
nor U10012 (N_10012,N_9173,N_9177);
nand U10013 (N_10013,N_8848,N_9487);
xnor U10014 (N_10014,N_8870,N_9116);
nand U10015 (N_10015,N_9151,N_8929);
xnor U10016 (N_10016,N_9167,N_9176);
nor U10017 (N_10017,N_9330,N_9379);
nand U10018 (N_10018,N_9435,N_9141);
or U10019 (N_10019,N_8806,N_9253);
nand U10020 (N_10020,N_9359,N_9270);
nor U10021 (N_10021,N_9471,N_9526);
nor U10022 (N_10022,N_8896,N_9546);
nor U10023 (N_10023,N_9170,N_8803);
xor U10024 (N_10024,N_8955,N_9576);
nor U10025 (N_10025,N_9291,N_8969);
and U10026 (N_10026,N_8895,N_9148);
nand U10027 (N_10027,N_9194,N_9351);
nor U10028 (N_10028,N_9535,N_9065);
nand U10029 (N_10029,N_9123,N_9217);
or U10030 (N_10030,N_8975,N_9104);
or U10031 (N_10031,N_9100,N_9315);
xnor U10032 (N_10032,N_9321,N_8901);
xnor U10033 (N_10033,N_8998,N_9296);
xor U10034 (N_10034,N_9029,N_9501);
nor U10035 (N_10035,N_8882,N_8873);
xor U10036 (N_10036,N_9195,N_9332);
nor U10037 (N_10037,N_9039,N_9001);
nor U10038 (N_10038,N_9360,N_9347);
and U10039 (N_10039,N_9203,N_8916);
and U10040 (N_10040,N_8872,N_8898);
or U10041 (N_10041,N_9013,N_9150);
nor U10042 (N_10042,N_9358,N_9396);
nor U10043 (N_10043,N_9423,N_9586);
nand U10044 (N_10044,N_8937,N_9140);
nor U10045 (N_10045,N_9148,N_8809);
nor U10046 (N_10046,N_9117,N_9294);
nor U10047 (N_10047,N_9012,N_9536);
and U10048 (N_10048,N_9568,N_8862);
or U10049 (N_10049,N_9359,N_8859);
and U10050 (N_10050,N_9059,N_9227);
and U10051 (N_10051,N_9040,N_9143);
and U10052 (N_10052,N_9476,N_9193);
nor U10053 (N_10053,N_9286,N_9020);
nor U10054 (N_10054,N_9243,N_9589);
and U10055 (N_10055,N_9517,N_9120);
xnor U10056 (N_10056,N_9485,N_9507);
and U10057 (N_10057,N_9383,N_9405);
and U10058 (N_10058,N_9470,N_9596);
nand U10059 (N_10059,N_8881,N_9079);
or U10060 (N_10060,N_9296,N_9581);
and U10061 (N_10061,N_9428,N_8962);
and U10062 (N_10062,N_9166,N_8978);
xor U10063 (N_10063,N_9486,N_9344);
xor U10064 (N_10064,N_9576,N_9192);
or U10065 (N_10065,N_8861,N_9409);
nand U10066 (N_10066,N_9401,N_8910);
or U10067 (N_10067,N_9249,N_9576);
xor U10068 (N_10068,N_8826,N_8901);
xor U10069 (N_10069,N_9505,N_9497);
xnor U10070 (N_10070,N_9279,N_9359);
and U10071 (N_10071,N_9522,N_9570);
and U10072 (N_10072,N_9007,N_9255);
xnor U10073 (N_10073,N_9339,N_9284);
xor U10074 (N_10074,N_9578,N_9381);
xor U10075 (N_10075,N_8951,N_8967);
xor U10076 (N_10076,N_9509,N_8996);
nand U10077 (N_10077,N_9199,N_9007);
nand U10078 (N_10078,N_9299,N_8912);
nand U10079 (N_10079,N_8874,N_9374);
and U10080 (N_10080,N_8841,N_9362);
nor U10081 (N_10081,N_9593,N_9022);
xnor U10082 (N_10082,N_9583,N_8850);
and U10083 (N_10083,N_9188,N_9428);
xnor U10084 (N_10084,N_8809,N_8842);
xor U10085 (N_10085,N_9384,N_9126);
xnor U10086 (N_10086,N_8800,N_8964);
and U10087 (N_10087,N_9066,N_9074);
nand U10088 (N_10088,N_9475,N_9418);
nand U10089 (N_10089,N_9041,N_8907);
and U10090 (N_10090,N_9482,N_9083);
or U10091 (N_10091,N_9188,N_8818);
nor U10092 (N_10092,N_9202,N_9013);
and U10093 (N_10093,N_8895,N_9339);
or U10094 (N_10094,N_9488,N_9573);
or U10095 (N_10095,N_9591,N_8948);
xnor U10096 (N_10096,N_9107,N_9316);
and U10097 (N_10097,N_8845,N_9154);
nand U10098 (N_10098,N_9008,N_8956);
nor U10099 (N_10099,N_9523,N_8896);
xor U10100 (N_10100,N_9395,N_8991);
and U10101 (N_10101,N_9255,N_8912);
nand U10102 (N_10102,N_9317,N_9407);
or U10103 (N_10103,N_8980,N_9057);
nor U10104 (N_10104,N_9544,N_8804);
and U10105 (N_10105,N_8822,N_9573);
and U10106 (N_10106,N_9005,N_9035);
or U10107 (N_10107,N_8856,N_9155);
or U10108 (N_10108,N_8888,N_9279);
and U10109 (N_10109,N_9574,N_9512);
or U10110 (N_10110,N_9253,N_9116);
nor U10111 (N_10111,N_9044,N_9464);
or U10112 (N_10112,N_8819,N_9426);
nand U10113 (N_10113,N_8894,N_9384);
nand U10114 (N_10114,N_9154,N_9353);
or U10115 (N_10115,N_9546,N_8918);
or U10116 (N_10116,N_8934,N_9231);
or U10117 (N_10117,N_9162,N_9160);
nor U10118 (N_10118,N_9578,N_9330);
xor U10119 (N_10119,N_9147,N_8894);
or U10120 (N_10120,N_9181,N_9281);
nor U10121 (N_10121,N_9072,N_8804);
and U10122 (N_10122,N_9430,N_9572);
nand U10123 (N_10123,N_9050,N_8945);
nand U10124 (N_10124,N_9359,N_9418);
and U10125 (N_10125,N_9579,N_8949);
and U10126 (N_10126,N_9273,N_9426);
and U10127 (N_10127,N_8861,N_8911);
or U10128 (N_10128,N_9097,N_9255);
and U10129 (N_10129,N_9324,N_9015);
nand U10130 (N_10130,N_9335,N_9392);
nand U10131 (N_10131,N_9567,N_8927);
or U10132 (N_10132,N_8952,N_9246);
and U10133 (N_10133,N_8861,N_8807);
nor U10134 (N_10134,N_9353,N_9021);
and U10135 (N_10135,N_9001,N_9561);
xor U10136 (N_10136,N_9072,N_9433);
or U10137 (N_10137,N_8971,N_9281);
or U10138 (N_10138,N_8976,N_9222);
xnor U10139 (N_10139,N_9089,N_9422);
nor U10140 (N_10140,N_9027,N_9170);
xor U10141 (N_10141,N_9105,N_9134);
xor U10142 (N_10142,N_9085,N_9321);
xor U10143 (N_10143,N_8855,N_9168);
or U10144 (N_10144,N_9330,N_9444);
xnor U10145 (N_10145,N_9553,N_9330);
nand U10146 (N_10146,N_9144,N_8844);
or U10147 (N_10147,N_9283,N_9037);
xor U10148 (N_10148,N_9285,N_8898);
and U10149 (N_10149,N_9157,N_9143);
nand U10150 (N_10150,N_8949,N_9080);
nand U10151 (N_10151,N_9501,N_9291);
nor U10152 (N_10152,N_9100,N_8832);
xnor U10153 (N_10153,N_9122,N_8851);
xnor U10154 (N_10154,N_9444,N_8839);
or U10155 (N_10155,N_9067,N_9183);
xnor U10156 (N_10156,N_9187,N_8814);
nand U10157 (N_10157,N_9032,N_9515);
xor U10158 (N_10158,N_9326,N_8991);
or U10159 (N_10159,N_9022,N_9474);
or U10160 (N_10160,N_9430,N_9323);
nand U10161 (N_10161,N_9267,N_9453);
and U10162 (N_10162,N_9442,N_9545);
nand U10163 (N_10163,N_9482,N_9531);
or U10164 (N_10164,N_9591,N_8822);
xor U10165 (N_10165,N_8871,N_9273);
or U10166 (N_10166,N_9430,N_8919);
or U10167 (N_10167,N_9012,N_8974);
nor U10168 (N_10168,N_9260,N_9061);
xnor U10169 (N_10169,N_8907,N_9146);
nand U10170 (N_10170,N_9233,N_9430);
or U10171 (N_10171,N_8876,N_8850);
xor U10172 (N_10172,N_9289,N_8803);
or U10173 (N_10173,N_8902,N_8832);
xor U10174 (N_10174,N_9424,N_9246);
nor U10175 (N_10175,N_9175,N_8918);
and U10176 (N_10176,N_9270,N_9209);
and U10177 (N_10177,N_9327,N_8939);
nand U10178 (N_10178,N_9515,N_8965);
nand U10179 (N_10179,N_9588,N_8930);
and U10180 (N_10180,N_8852,N_8980);
nand U10181 (N_10181,N_8950,N_9278);
nand U10182 (N_10182,N_9518,N_8818);
and U10183 (N_10183,N_8975,N_9232);
or U10184 (N_10184,N_8883,N_8805);
and U10185 (N_10185,N_9134,N_9417);
or U10186 (N_10186,N_9152,N_8817);
nor U10187 (N_10187,N_8912,N_8860);
nand U10188 (N_10188,N_8845,N_9000);
nand U10189 (N_10189,N_8868,N_9332);
nand U10190 (N_10190,N_9283,N_9480);
or U10191 (N_10191,N_8845,N_8970);
nor U10192 (N_10192,N_9370,N_9061);
xor U10193 (N_10193,N_8951,N_9036);
nand U10194 (N_10194,N_8929,N_9409);
and U10195 (N_10195,N_9070,N_9175);
and U10196 (N_10196,N_8891,N_9008);
nor U10197 (N_10197,N_8801,N_9100);
nand U10198 (N_10198,N_8936,N_9067);
and U10199 (N_10199,N_9219,N_9203);
nor U10200 (N_10200,N_9489,N_8942);
nand U10201 (N_10201,N_9444,N_9052);
or U10202 (N_10202,N_9313,N_9218);
nor U10203 (N_10203,N_9509,N_8975);
or U10204 (N_10204,N_8850,N_9134);
xor U10205 (N_10205,N_9223,N_9105);
nand U10206 (N_10206,N_8852,N_8849);
xor U10207 (N_10207,N_9274,N_9404);
nor U10208 (N_10208,N_9380,N_9171);
and U10209 (N_10209,N_9355,N_9397);
nand U10210 (N_10210,N_8834,N_9207);
nand U10211 (N_10211,N_9116,N_8895);
or U10212 (N_10212,N_9229,N_9482);
nor U10213 (N_10213,N_8826,N_9334);
nand U10214 (N_10214,N_9462,N_9454);
nor U10215 (N_10215,N_8886,N_9484);
nand U10216 (N_10216,N_9461,N_9538);
nor U10217 (N_10217,N_9217,N_9580);
xnor U10218 (N_10218,N_9191,N_9413);
and U10219 (N_10219,N_9431,N_8841);
nor U10220 (N_10220,N_9486,N_9304);
or U10221 (N_10221,N_8952,N_9301);
or U10222 (N_10222,N_8832,N_8965);
and U10223 (N_10223,N_9104,N_9537);
or U10224 (N_10224,N_9564,N_9484);
or U10225 (N_10225,N_9398,N_9286);
or U10226 (N_10226,N_9064,N_9123);
and U10227 (N_10227,N_9308,N_9465);
and U10228 (N_10228,N_9077,N_9369);
and U10229 (N_10229,N_9571,N_9108);
or U10230 (N_10230,N_8915,N_9049);
nand U10231 (N_10231,N_9110,N_8827);
nor U10232 (N_10232,N_9166,N_9407);
xnor U10233 (N_10233,N_9553,N_8811);
nand U10234 (N_10234,N_9314,N_9406);
and U10235 (N_10235,N_9474,N_9476);
and U10236 (N_10236,N_9144,N_9537);
nor U10237 (N_10237,N_9225,N_9201);
and U10238 (N_10238,N_9197,N_9452);
xnor U10239 (N_10239,N_9413,N_9506);
and U10240 (N_10240,N_9405,N_8816);
or U10241 (N_10241,N_8971,N_9111);
nand U10242 (N_10242,N_9403,N_9368);
nor U10243 (N_10243,N_9137,N_9317);
or U10244 (N_10244,N_9058,N_9018);
or U10245 (N_10245,N_9471,N_8865);
nor U10246 (N_10246,N_9234,N_9337);
and U10247 (N_10247,N_9329,N_9046);
nor U10248 (N_10248,N_8907,N_9270);
or U10249 (N_10249,N_9377,N_9204);
nor U10250 (N_10250,N_8844,N_8930);
nor U10251 (N_10251,N_9033,N_9195);
nor U10252 (N_10252,N_9037,N_9233);
nand U10253 (N_10253,N_9292,N_9364);
or U10254 (N_10254,N_8853,N_8982);
or U10255 (N_10255,N_9277,N_9384);
and U10256 (N_10256,N_9187,N_8972);
nand U10257 (N_10257,N_9130,N_8940);
and U10258 (N_10258,N_9037,N_8808);
xor U10259 (N_10259,N_8874,N_8943);
or U10260 (N_10260,N_9068,N_9238);
nand U10261 (N_10261,N_8961,N_8815);
nor U10262 (N_10262,N_8809,N_9041);
xnor U10263 (N_10263,N_9560,N_9314);
and U10264 (N_10264,N_9198,N_9157);
nand U10265 (N_10265,N_9468,N_9538);
and U10266 (N_10266,N_8837,N_9464);
nor U10267 (N_10267,N_9025,N_9414);
xor U10268 (N_10268,N_8928,N_9208);
nand U10269 (N_10269,N_9369,N_9578);
xnor U10270 (N_10270,N_9584,N_9418);
or U10271 (N_10271,N_8992,N_9422);
and U10272 (N_10272,N_8837,N_9042);
and U10273 (N_10273,N_9314,N_9555);
or U10274 (N_10274,N_8804,N_9033);
nor U10275 (N_10275,N_9451,N_8861);
xnor U10276 (N_10276,N_8875,N_9578);
or U10277 (N_10277,N_8836,N_8874);
or U10278 (N_10278,N_9194,N_9091);
nor U10279 (N_10279,N_8847,N_9419);
or U10280 (N_10280,N_9028,N_8983);
xor U10281 (N_10281,N_8988,N_9503);
nand U10282 (N_10282,N_9098,N_8994);
xnor U10283 (N_10283,N_8882,N_8981);
nor U10284 (N_10284,N_9299,N_9555);
or U10285 (N_10285,N_9014,N_9352);
nor U10286 (N_10286,N_9285,N_9004);
or U10287 (N_10287,N_8810,N_9555);
and U10288 (N_10288,N_9390,N_8972);
or U10289 (N_10289,N_9392,N_9586);
and U10290 (N_10290,N_9344,N_9571);
nor U10291 (N_10291,N_8978,N_9409);
nor U10292 (N_10292,N_9534,N_8801);
xnor U10293 (N_10293,N_9057,N_9196);
nand U10294 (N_10294,N_8806,N_8830);
nor U10295 (N_10295,N_9503,N_9038);
or U10296 (N_10296,N_8883,N_8887);
nor U10297 (N_10297,N_8919,N_9310);
xor U10298 (N_10298,N_8875,N_8849);
and U10299 (N_10299,N_9134,N_8943);
and U10300 (N_10300,N_9220,N_8982);
or U10301 (N_10301,N_9375,N_9466);
and U10302 (N_10302,N_9267,N_8943);
or U10303 (N_10303,N_9538,N_9438);
nand U10304 (N_10304,N_8946,N_9396);
nor U10305 (N_10305,N_8885,N_9543);
nor U10306 (N_10306,N_9558,N_9150);
or U10307 (N_10307,N_9442,N_9312);
xor U10308 (N_10308,N_9515,N_9472);
nor U10309 (N_10309,N_9472,N_9398);
or U10310 (N_10310,N_9560,N_9543);
xor U10311 (N_10311,N_8949,N_9522);
or U10312 (N_10312,N_9297,N_8948);
or U10313 (N_10313,N_9577,N_9385);
and U10314 (N_10314,N_9296,N_9109);
and U10315 (N_10315,N_9540,N_8905);
xnor U10316 (N_10316,N_9187,N_8919);
nor U10317 (N_10317,N_9198,N_9229);
xnor U10318 (N_10318,N_8877,N_9521);
nor U10319 (N_10319,N_9589,N_9095);
or U10320 (N_10320,N_8838,N_9016);
nand U10321 (N_10321,N_9154,N_9568);
nand U10322 (N_10322,N_8936,N_8909);
nand U10323 (N_10323,N_9499,N_9081);
nor U10324 (N_10324,N_9229,N_9393);
or U10325 (N_10325,N_9334,N_9209);
nand U10326 (N_10326,N_9170,N_9365);
nor U10327 (N_10327,N_8889,N_9220);
or U10328 (N_10328,N_9108,N_9469);
nand U10329 (N_10329,N_9185,N_9488);
or U10330 (N_10330,N_9267,N_9266);
or U10331 (N_10331,N_9495,N_9537);
xor U10332 (N_10332,N_9218,N_9571);
and U10333 (N_10333,N_9302,N_9212);
nor U10334 (N_10334,N_8840,N_9237);
xnor U10335 (N_10335,N_9471,N_9448);
nor U10336 (N_10336,N_9160,N_9216);
or U10337 (N_10337,N_9170,N_9524);
nor U10338 (N_10338,N_9215,N_9408);
xor U10339 (N_10339,N_9544,N_9374);
nand U10340 (N_10340,N_8928,N_9441);
or U10341 (N_10341,N_9024,N_9303);
nor U10342 (N_10342,N_9151,N_9472);
and U10343 (N_10343,N_8872,N_9092);
nor U10344 (N_10344,N_9178,N_9549);
and U10345 (N_10345,N_8872,N_9373);
or U10346 (N_10346,N_9319,N_9133);
or U10347 (N_10347,N_9417,N_9364);
nand U10348 (N_10348,N_8913,N_9261);
and U10349 (N_10349,N_9386,N_9358);
nor U10350 (N_10350,N_9597,N_9059);
nor U10351 (N_10351,N_9355,N_9198);
xor U10352 (N_10352,N_9235,N_9538);
xor U10353 (N_10353,N_9562,N_9328);
nand U10354 (N_10354,N_9155,N_8933);
nand U10355 (N_10355,N_9541,N_9034);
or U10356 (N_10356,N_8912,N_9159);
or U10357 (N_10357,N_9100,N_9013);
nand U10358 (N_10358,N_9203,N_9180);
or U10359 (N_10359,N_8849,N_9166);
nor U10360 (N_10360,N_9072,N_8868);
xnor U10361 (N_10361,N_9185,N_9159);
and U10362 (N_10362,N_9003,N_9482);
nand U10363 (N_10363,N_9274,N_8891);
nand U10364 (N_10364,N_9224,N_9416);
nand U10365 (N_10365,N_9064,N_8874);
or U10366 (N_10366,N_9561,N_8954);
nor U10367 (N_10367,N_9128,N_8965);
nor U10368 (N_10368,N_9162,N_9566);
and U10369 (N_10369,N_9337,N_9101);
xor U10370 (N_10370,N_9509,N_9421);
nor U10371 (N_10371,N_9358,N_9145);
or U10372 (N_10372,N_8827,N_9423);
xnor U10373 (N_10373,N_9463,N_9206);
nand U10374 (N_10374,N_9250,N_9471);
and U10375 (N_10375,N_8982,N_9457);
nand U10376 (N_10376,N_8903,N_9400);
or U10377 (N_10377,N_9157,N_9021);
nor U10378 (N_10378,N_9066,N_9523);
and U10379 (N_10379,N_8987,N_9435);
nand U10380 (N_10380,N_9458,N_9008);
nand U10381 (N_10381,N_9235,N_9460);
nor U10382 (N_10382,N_9086,N_8850);
and U10383 (N_10383,N_8955,N_9084);
nand U10384 (N_10384,N_8843,N_9493);
xor U10385 (N_10385,N_9208,N_9138);
nor U10386 (N_10386,N_9527,N_9453);
xnor U10387 (N_10387,N_9044,N_9039);
and U10388 (N_10388,N_9279,N_9450);
nand U10389 (N_10389,N_9506,N_9246);
xnor U10390 (N_10390,N_8843,N_9429);
or U10391 (N_10391,N_9406,N_9089);
nor U10392 (N_10392,N_9120,N_8832);
xnor U10393 (N_10393,N_9004,N_8884);
or U10394 (N_10394,N_8900,N_9106);
nor U10395 (N_10395,N_9195,N_9273);
or U10396 (N_10396,N_8921,N_9529);
xnor U10397 (N_10397,N_9230,N_9305);
xor U10398 (N_10398,N_9497,N_9282);
nor U10399 (N_10399,N_8980,N_9444);
nand U10400 (N_10400,N_10005,N_10010);
nor U10401 (N_10401,N_10285,N_9793);
and U10402 (N_10402,N_10061,N_9717);
xor U10403 (N_10403,N_9718,N_9929);
and U10404 (N_10404,N_9787,N_9620);
or U10405 (N_10405,N_9915,N_9659);
or U10406 (N_10406,N_9873,N_9975);
nand U10407 (N_10407,N_10077,N_10128);
xnor U10408 (N_10408,N_10336,N_10323);
or U10409 (N_10409,N_10038,N_9698);
or U10410 (N_10410,N_9928,N_10385);
or U10411 (N_10411,N_9744,N_10017);
or U10412 (N_10412,N_9704,N_10083);
xnor U10413 (N_10413,N_9957,N_9752);
nor U10414 (N_10414,N_10252,N_9774);
and U10415 (N_10415,N_9769,N_10389);
nand U10416 (N_10416,N_9700,N_10256);
or U10417 (N_10417,N_10086,N_10383);
xnor U10418 (N_10418,N_10219,N_9932);
xnor U10419 (N_10419,N_9907,N_10136);
and U10420 (N_10420,N_10051,N_10041);
and U10421 (N_10421,N_10117,N_10014);
nand U10422 (N_10422,N_10342,N_9834);
or U10423 (N_10423,N_9759,N_9885);
nor U10424 (N_10424,N_9822,N_9808);
xnor U10425 (N_10425,N_9691,N_10200);
or U10426 (N_10426,N_9911,N_9823);
or U10427 (N_10427,N_10114,N_9825);
nand U10428 (N_10428,N_10045,N_10094);
xnor U10429 (N_10429,N_10042,N_10089);
nand U10430 (N_10430,N_9676,N_10222);
nor U10431 (N_10431,N_10076,N_10080);
and U10432 (N_10432,N_10217,N_9657);
and U10433 (N_10433,N_10243,N_10164);
nor U10434 (N_10434,N_9841,N_10177);
and U10435 (N_10435,N_9988,N_9810);
or U10436 (N_10436,N_10134,N_9962);
nor U10437 (N_10437,N_10269,N_10168);
or U10438 (N_10438,N_10171,N_9917);
nand U10439 (N_10439,N_10106,N_10102);
nor U10440 (N_10440,N_9938,N_9912);
or U10441 (N_10441,N_9770,N_10173);
nand U10442 (N_10442,N_10208,N_9900);
xnor U10443 (N_10443,N_10282,N_10143);
nor U10444 (N_10444,N_10221,N_9767);
xnor U10445 (N_10445,N_9966,N_9678);
nand U10446 (N_10446,N_10257,N_10211);
nand U10447 (N_10447,N_10375,N_10085);
or U10448 (N_10448,N_9943,N_9817);
or U10449 (N_10449,N_9609,N_9904);
nand U10450 (N_10450,N_9977,N_10107);
nand U10451 (N_10451,N_10268,N_10122);
nand U10452 (N_10452,N_9987,N_10155);
xor U10453 (N_10453,N_9629,N_9878);
or U10454 (N_10454,N_10392,N_9748);
or U10455 (N_10455,N_9790,N_10374);
nand U10456 (N_10456,N_9681,N_9833);
or U10457 (N_10457,N_9890,N_10115);
or U10458 (N_10458,N_10274,N_10071);
nand U10459 (N_10459,N_10299,N_9666);
nand U10460 (N_10460,N_9610,N_10334);
or U10461 (N_10461,N_9828,N_10396);
nor U10462 (N_10462,N_9933,N_9697);
nand U10463 (N_10463,N_10230,N_9997);
nand U10464 (N_10464,N_10063,N_9675);
and U10465 (N_10465,N_9974,N_10179);
nand U10466 (N_10466,N_10242,N_10146);
nand U10467 (N_10467,N_9632,N_10047);
nor U10468 (N_10468,N_9773,N_10391);
xnor U10469 (N_10469,N_9940,N_10174);
nor U10470 (N_10470,N_9923,N_9600);
xnor U10471 (N_10471,N_9756,N_9809);
and U10472 (N_10472,N_10281,N_10029);
xor U10473 (N_10473,N_9984,N_10103);
and U10474 (N_10474,N_9667,N_10328);
nor U10475 (N_10475,N_10119,N_10160);
or U10476 (N_10476,N_9916,N_10144);
nor U10477 (N_10477,N_10355,N_10125);
nand U10478 (N_10478,N_9648,N_10099);
nand U10479 (N_10479,N_9775,N_10040);
nor U10480 (N_10480,N_10367,N_9887);
and U10481 (N_10481,N_10170,N_9705);
xor U10482 (N_10482,N_10393,N_10277);
nor U10483 (N_10483,N_9639,N_9771);
and U10484 (N_10484,N_10187,N_10302);
nor U10485 (N_10485,N_10226,N_9628);
nand U10486 (N_10486,N_10255,N_9740);
nor U10487 (N_10487,N_9807,N_10152);
nor U10488 (N_10488,N_10167,N_9980);
nand U10489 (N_10489,N_10068,N_9763);
nand U10490 (N_10490,N_10388,N_9820);
or U10491 (N_10491,N_9982,N_9858);
xnor U10492 (N_10492,N_9983,N_10092);
or U10493 (N_10493,N_10009,N_10079);
and U10494 (N_10494,N_10223,N_10265);
nand U10495 (N_10495,N_10031,N_10198);
or U10496 (N_10496,N_9640,N_9970);
xnor U10497 (N_10497,N_10039,N_10258);
and U10498 (N_10498,N_9934,N_9779);
xnor U10499 (N_10499,N_9702,N_9680);
xnor U10500 (N_10500,N_9813,N_9614);
or U10501 (N_10501,N_10232,N_9690);
or U10502 (N_10502,N_10147,N_10327);
or U10503 (N_10503,N_10248,N_10306);
xor U10504 (N_10504,N_9796,N_9949);
nor U10505 (N_10505,N_10363,N_10091);
or U10506 (N_10506,N_10234,N_9944);
xor U10507 (N_10507,N_10348,N_9876);
xnor U10508 (N_10508,N_9647,N_10067);
and U10509 (N_10509,N_9608,N_9689);
and U10510 (N_10510,N_10227,N_10313);
xor U10511 (N_10511,N_10054,N_9630);
nor U10512 (N_10512,N_9784,N_10237);
nand U10513 (N_10513,N_10368,N_9935);
xor U10514 (N_10514,N_10350,N_10140);
or U10515 (N_10515,N_9894,N_10161);
xnor U10516 (N_10516,N_10332,N_9710);
or U10517 (N_10517,N_9905,N_9737);
nor U10518 (N_10518,N_9826,N_10390);
and U10519 (N_10519,N_9831,N_9844);
xor U10520 (N_10520,N_10113,N_9852);
nor U10521 (N_10521,N_10132,N_10296);
and U10522 (N_10522,N_9755,N_10149);
or U10523 (N_10523,N_10188,N_9643);
xor U10524 (N_10524,N_10397,N_9613);
or U10525 (N_10525,N_9783,N_10301);
nor U10526 (N_10526,N_9963,N_9816);
and U10527 (N_10527,N_9996,N_9764);
nand U10528 (N_10528,N_9967,N_9724);
and U10529 (N_10529,N_10059,N_9802);
or U10530 (N_10530,N_10037,N_9971);
nand U10531 (N_10531,N_9886,N_10084);
nor U10532 (N_10532,N_10294,N_9685);
or U10533 (N_10533,N_9703,N_9658);
nor U10534 (N_10534,N_9728,N_10073);
nor U10535 (N_10535,N_10111,N_10399);
and U10536 (N_10536,N_9747,N_10028);
xor U10537 (N_10537,N_10139,N_10153);
xor U10538 (N_10538,N_9662,N_10319);
nor U10539 (N_10539,N_10098,N_10126);
or U10540 (N_10540,N_9968,N_9664);
and U10541 (N_10541,N_9707,N_10004);
and U10542 (N_10542,N_9909,N_10166);
nand U10543 (N_10543,N_9645,N_9875);
nor U10544 (N_10544,N_10082,N_9794);
xnor U10545 (N_10545,N_10286,N_10271);
or U10546 (N_10546,N_10199,N_10052);
xnor U10547 (N_10547,N_9950,N_9765);
nand U10548 (N_10548,N_9897,N_10022);
and U10549 (N_10549,N_10100,N_10216);
xnor U10550 (N_10550,N_10361,N_9857);
nand U10551 (N_10551,N_10048,N_9776);
nor U10552 (N_10552,N_9835,N_10032);
or U10553 (N_10553,N_9877,N_10272);
or U10554 (N_10554,N_10185,N_10108);
or U10555 (N_10555,N_9832,N_9918);
and U10556 (N_10556,N_9979,N_10070);
nor U10557 (N_10557,N_10116,N_10305);
nor U10558 (N_10558,N_10395,N_9829);
and U10559 (N_10559,N_10324,N_9743);
and U10560 (N_10560,N_10293,N_10241);
or U10561 (N_10561,N_9761,N_9731);
nand U10562 (N_10562,N_10095,N_10338);
nand U10563 (N_10563,N_9670,N_9811);
xor U10564 (N_10564,N_10050,N_9624);
xnor U10565 (N_10565,N_9819,N_9625);
xnor U10566 (N_10566,N_10145,N_9661);
xor U10567 (N_10567,N_10353,N_9656);
or U10568 (N_10568,N_9735,N_9867);
nand U10569 (N_10569,N_9893,N_9960);
nand U10570 (N_10570,N_9649,N_10123);
nand U10571 (N_10571,N_10333,N_9799);
nor U10572 (N_10572,N_9855,N_9749);
nor U10573 (N_10573,N_10343,N_9840);
or U10574 (N_10574,N_10105,N_9981);
or U10575 (N_10575,N_10062,N_9880);
nand U10576 (N_10576,N_9604,N_9782);
and U10577 (N_10577,N_10142,N_9652);
and U10578 (N_10578,N_9695,N_9869);
or U10579 (N_10579,N_10024,N_9706);
nor U10580 (N_10580,N_9758,N_9851);
or U10581 (N_10581,N_10195,N_9633);
and U10582 (N_10582,N_10358,N_10056);
and U10583 (N_10583,N_10318,N_9827);
xnor U10584 (N_10584,N_10175,N_10228);
nand U10585 (N_10585,N_10259,N_9925);
nor U10586 (N_10586,N_9931,N_9872);
xor U10587 (N_10587,N_9946,N_10246);
nor U10588 (N_10588,N_9654,N_9908);
and U10589 (N_10589,N_10192,N_10315);
or U10590 (N_10590,N_10203,N_9621);
nand U10591 (N_10591,N_9688,N_10109);
and U10592 (N_10592,N_9843,N_10036);
nand U10593 (N_10593,N_9939,N_9617);
xnor U10594 (N_10594,N_9947,N_10326);
or U10595 (N_10595,N_9956,N_9976);
or U10596 (N_10596,N_9868,N_9607);
and U10597 (N_10597,N_9797,N_10018);
and U10598 (N_10598,N_10150,N_9815);
and U10599 (N_10599,N_9906,N_10197);
and U10600 (N_10600,N_10290,N_10307);
nor U10601 (N_10601,N_10381,N_9738);
nor U10602 (N_10602,N_10292,N_10210);
nor U10603 (N_10603,N_10349,N_9723);
nand U10604 (N_10604,N_9636,N_10156);
nor U10605 (N_10605,N_10060,N_9990);
xnor U10606 (N_10606,N_9682,N_9845);
xor U10607 (N_10607,N_10310,N_9641);
or U10608 (N_10608,N_9669,N_9745);
or U10609 (N_10609,N_9674,N_10157);
or U10610 (N_10610,N_9850,N_10371);
nor U10611 (N_10611,N_10093,N_10025);
nor U10612 (N_10612,N_10298,N_10159);
xnor U10613 (N_10613,N_10364,N_10283);
or U10614 (N_10614,N_9955,N_9945);
and U10615 (N_10615,N_9926,N_9660);
or U10616 (N_10616,N_10235,N_9646);
and U10617 (N_10617,N_9663,N_9969);
nand U10618 (N_10618,N_10003,N_9736);
xor U10619 (N_10619,N_10035,N_10339);
nor U10620 (N_10620,N_10069,N_9842);
or U10621 (N_10621,N_10129,N_9746);
xnor U10622 (N_10622,N_10345,N_9986);
nand U10623 (N_10623,N_9913,N_10141);
nor U10624 (N_10624,N_9921,N_10011);
xor U10625 (N_10625,N_9719,N_10236);
xnor U10626 (N_10626,N_10072,N_9615);
nand U10627 (N_10627,N_9623,N_9638);
nor U10628 (N_10628,N_10096,N_9619);
nand U10629 (N_10629,N_9994,N_10190);
and U10630 (N_10630,N_9612,N_10279);
xor U10631 (N_10631,N_10021,N_10378);
xnor U10632 (N_10632,N_10335,N_9611);
nand U10633 (N_10633,N_9824,N_9941);
and U10634 (N_10634,N_10206,N_10262);
and U10635 (N_10635,N_10341,N_9768);
and U10636 (N_10636,N_9711,N_10204);
and U10637 (N_10637,N_9952,N_9772);
or U10638 (N_10638,N_9884,N_9804);
nor U10639 (N_10639,N_9818,N_9665);
xor U10640 (N_10640,N_10066,N_10300);
and U10641 (N_10641,N_10314,N_9853);
and U10642 (N_10642,N_10225,N_10046);
nor U10643 (N_10643,N_10377,N_9701);
xnor U10644 (N_10644,N_10384,N_9668);
and U10645 (N_10645,N_10033,N_9896);
nand U10646 (N_10646,N_9863,N_10186);
nor U10647 (N_10647,N_9726,N_10194);
and U10648 (N_10648,N_9757,N_9992);
and U10649 (N_10649,N_9882,N_10231);
nor U10650 (N_10650,N_9800,N_10121);
and U10651 (N_10651,N_10133,N_9874);
nand U10652 (N_10652,N_10254,N_9965);
xor U10653 (N_10653,N_9734,N_9716);
xor U10654 (N_10654,N_9795,N_9898);
and U10655 (N_10655,N_9637,N_9777);
and U10656 (N_10656,N_9789,N_9605);
and U10657 (N_10657,N_9650,N_9751);
nand U10658 (N_10658,N_10250,N_10309);
xnor U10659 (N_10659,N_10370,N_9902);
nand U10660 (N_10660,N_10289,N_9948);
nand U10661 (N_10661,N_9914,N_9760);
or U10662 (N_10662,N_9753,N_9715);
xor U10663 (N_10663,N_10016,N_10316);
xnor U10664 (N_10664,N_9961,N_10382);
nand U10665 (N_10665,N_9786,N_10163);
nor U10666 (N_10666,N_10218,N_9714);
and U10667 (N_10667,N_9806,N_9847);
xnor U10668 (N_10668,N_10263,N_10304);
nor U10669 (N_10669,N_9644,N_10043);
xnor U10670 (N_10670,N_9778,N_10362);
nor U10671 (N_10671,N_9892,N_9603);
and U10672 (N_10672,N_9677,N_9683);
and U10673 (N_10673,N_10212,N_9830);
and U10674 (N_10674,N_10233,N_10130);
nand U10675 (N_10675,N_9972,N_10270);
nor U10676 (N_10676,N_10087,N_9791);
nor U10677 (N_10677,N_9616,N_10346);
nor U10678 (N_10678,N_9958,N_10201);
nand U10679 (N_10679,N_10118,N_9673);
nand U10680 (N_10680,N_9899,N_9634);
and U10681 (N_10681,N_10312,N_9995);
nor U10682 (N_10682,N_10297,N_10137);
nor U10683 (N_10683,N_9978,N_9848);
nand U10684 (N_10684,N_10064,N_9655);
xor U10685 (N_10685,N_10104,N_10273);
xor U10686 (N_10686,N_9739,N_10275);
xnor U10687 (N_10687,N_10280,N_9780);
xor U10688 (N_10688,N_10344,N_9901);
and U10689 (N_10689,N_9985,N_10207);
xnor U10690 (N_10690,N_9837,N_9895);
and U10691 (N_10691,N_10007,N_9762);
nand U10692 (N_10692,N_9708,N_10284);
nor U10693 (N_10693,N_9732,N_10261);
or U10694 (N_10694,N_10295,N_10347);
xor U10695 (N_10695,N_9821,N_9849);
and U10696 (N_10696,N_9722,N_9713);
nand U10697 (N_10697,N_9727,N_10006);
and U10698 (N_10698,N_10357,N_10205);
xnor U10699 (N_10699,N_10131,N_9999);
and U10700 (N_10700,N_9788,N_10182);
nor U10701 (N_10701,N_9888,N_10337);
xnor U10702 (N_10702,N_10249,N_9631);
nor U10703 (N_10703,N_10366,N_9712);
or U10704 (N_10704,N_9729,N_10331);
nand U10705 (N_10705,N_9964,N_9720);
nor U10706 (N_10706,N_10264,N_9672);
xor U10707 (N_10707,N_9951,N_10148);
xnor U10708 (N_10708,N_9864,N_10055);
and U10709 (N_10709,N_10379,N_9879);
nor U10710 (N_10710,N_9920,N_10320);
nor U10711 (N_10711,N_10245,N_10124);
or U10712 (N_10712,N_10239,N_9836);
or U10713 (N_10713,N_9910,N_10229);
nor U10714 (N_10714,N_9741,N_10090);
nor U10715 (N_10715,N_10325,N_10247);
xnor U10716 (N_10716,N_9725,N_10276);
or U10717 (N_10717,N_9626,N_9692);
nor U10718 (N_10718,N_10165,N_9602);
nand U10719 (N_10719,N_9927,N_9846);
nor U10720 (N_10720,N_9618,N_10376);
nor U10721 (N_10721,N_10238,N_10251);
and U10722 (N_10722,N_9959,N_9891);
xor U10723 (N_10723,N_10224,N_9973);
xnor U10724 (N_10724,N_10394,N_9805);
xor U10725 (N_10725,N_10373,N_10329);
or U10726 (N_10726,N_9919,N_10209);
xnor U10727 (N_10727,N_10074,N_10057);
or U10728 (N_10728,N_10311,N_9733);
xor U10729 (N_10729,N_10112,N_10330);
nor U10730 (N_10730,N_9687,N_9814);
and U10731 (N_10731,N_10213,N_10181);
and U10732 (N_10732,N_10278,N_10202);
and U10733 (N_10733,N_9865,N_9989);
or U10734 (N_10734,N_10183,N_9781);
or U10735 (N_10735,N_10097,N_10386);
nor U10736 (N_10736,N_10020,N_10027);
and U10737 (N_10737,N_9839,N_10044);
and U10738 (N_10738,N_9754,N_10291);
and U10739 (N_10739,N_9993,N_10380);
or U10740 (N_10740,N_9860,N_10012);
and U10741 (N_10741,N_10365,N_9785);
and U10742 (N_10742,N_10019,N_10008);
and U10743 (N_10743,N_9942,N_10002);
nand U10744 (N_10744,N_9953,N_10214);
or U10745 (N_10745,N_10078,N_10189);
xnor U10746 (N_10746,N_10321,N_10176);
nor U10747 (N_10747,N_9686,N_9696);
nand U10748 (N_10748,N_10354,N_9903);
and U10749 (N_10749,N_10088,N_9653);
xnor U10750 (N_10750,N_10191,N_10075);
nand U10751 (N_10751,N_9684,N_9601);
nor U10752 (N_10752,N_10110,N_10253);
xor U10753 (N_10753,N_10308,N_9991);
nor U10754 (N_10754,N_10359,N_9801);
and U10755 (N_10755,N_9679,N_10215);
xnor U10756 (N_10756,N_10081,N_10030);
or U10757 (N_10757,N_10184,N_10013);
or U10758 (N_10758,N_9866,N_10138);
xnor U10759 (N_10759,N_10023,N_10101);
nand U10760 (N_10760,N_10369,N_9998);
xor U10761 (N_10761,N_10220,N_9936);
or U10762 (N_10762,N_10172,N_10151);
or U10763 (N_10763,N_9924,N_9856);
nor U10764 (N_10764,N_10288,N_9930);
xnor U10765 (N_10765,N_9854,N_10244);
xor U10766 (N_10766,N_9742,N_9635);
and U10767 (N_10767,N_10317,N_10154);
nand U10768 (N_10768,N_9671,N_9651);
nand U10769 (N_10769,N_10360,N_9937);
nand U10770 (N_10770,N_10303,N_9861);
nand U10771 (N_10771,N_10352,N_10158);
nand U10772 (N_10772,N_10340,N_10120);
or U10773 (N_10773,N_10135,N_9803);
xnor U10774 (N_10774,N_10049,N_9798);
xor U10775 (N_10775,N_9792,N_9883);
nand U10776 (N_10776,N_10260,N_10356);
nand U10777 (N_10777,N_9922,N_9889);
xor U10778 (N_10778,N_10058,N_10266);
or U10779 (N_10779,N_9812,N_9627);
nor U10780 (N_10780,N_9859,N_9699);
nor U10781 (N_10781,N_10000,N_9693);
nand U10782 (N_10782,N_9750,N_10015);
nand U10783 (N_10783,N_10178,N_10127);
nor U10784 (N_10784,N_10034,N_10287);
and U10785 (N_10785,N_9622,N_10065);
nor U10786 (N_10786,N_10398,N_10351);
or U10787 (N_10787,N_9721,N_10387);
xor U10788 (N_10788,N_10026,N_10162);
and U10789 (N_10789,N_10193,N_10372);
nand U10790 (N_10790,N_9694,N_10180);
nand U10791 (N_10791,N_9766,N_9730);
xnor U10792 (N_10792,N_9881,N_10240);
xor U10793 (N_10793,N_10001,N_10053);
nand U10794 (N_10794,N_9954,N_9838);
nand U10795 (N_10795,N_9870,N_10322);
or U10796 (N_10796,N_9862,N_10169);
nand U10797 (N_10797,N_9642,N_9871);
nand U10798 (N_10798,N_10196,N_9606);
and U10799 (N_10799,N_10267,N_9709);
nor U10800 (N_10800,N_10298,N_9945);
or U10801 (N_10801,N_10386,N_10104);
and U10802 (N_10802,N_9688,N_9821);
xor U10803 (N_10803,N_10340,N_10127);
and U10804 (N_10804,N_10116,N_10270);
nor U10805 (N_10805,N_9600,N_10164);
and U10806 (N_10806,N_10336,N_10180);
xnor U10807 (N_10807,N_10022,N_10273);
nand U10808 (N_10808,N_10045,N_10246);
xor U10809 (N_10809,N_10225,N_10025);
xnor U10810 (N_10810,N_10260,N_10267);
and U10811 (N_10811,N_9694,N_9998);
and U10812 (N_10812,N_9815,N_9925);
nand U10813 (N_10813,N_9849,N_10337);
nor U10814 (N_10814,N_10177,N_9925);
and U10815 (N_10815,N_9691,N_10288);
xnor U10816 (N_10816,N_9910,N_10167);
and U10817 (N_10817,N_9750,N_9896);
xnor U10818 (N_10818,N_10010,N_9898);
nor U10819 (N_10819,N_9829,N_10229);
xor U10820 (N_10820,N_9912,N_9923);
or U10821 (N_10821,N_10170,N_10259);
or U10822 (N_10822,N_9657,N_10060);
or U10823 (N_10823,N_10058,N_9855);
xor U10824 (N_10824,N_9823,N_10019);
or U10825 (N_10825,N_9712,N_10172);
and U10826 (N_10826,N_10398,N_9745);
or U10827 (N_10827,N_9893,N_9852);
or U10828 (N_10828,N_9794,N_9605);
xor U10829 (N_10829,N_10369,N_9921);
or U10830 (N_10830,N_9933,N_10135);
or U10831 (N_10831,N_10380,N_10042);
nor U10832 (N_10832,N_9977,N_10256);
or U10833 (N_10833,N_9852,N_10373);
xnor U10834 (N_10834,N_10058,N_10333);
nand U10835 (N_10835,N_10079,N_9972);
nor U10836 (N_10836,N_9911,N_10217);
xnor U10837 (N_10837,N_9670,N_10136);
nor U10838 (N_10838,N_10201,N_10307);
or U10839 (N_10839,N_10253,N_9994);
nor U10840 (N_10840,N_9970,N_9705);
nor U10841 (N_10841,N_9765,N_9826);
and U10842 (N_10842,N_10178,N_10128);
nor U10843 (N_10843,N_9820,N_10051);
and U10844 (N_10844,N_10285,N_9777);
nor U10845 (N_10845,N_10031,N_9916);
or U10846 (N_10846,N_9930,N_9703);
nor U10847 (N_10847,N_10377,N_9611);
and U10848 (N_10848,N_9737,N_9814);
nor U10849 (N_10849,N_10353,N_9622);
nor U10850 (N_10850,N_10029,N_10209);
and U10851 (N_10851,N_10303,N_10056);
or U10852 (N_10852,N_10216,N_10054);
nand U10853 (N_10853,N_9999,N_9824);
nand U10854 (N_10854,N_10238,N_10209);
xor U10855 (N_10855,N_10302,N_10375);
and U10856 (N_10856,N_10331,N_9617);
and U10857 (N_10857,N_10315,N_10053);
and U10858 (N_10858,N_10066,N_10107);
nand U10859 (N_10859,N_9733,N_10267);
nor U10860 (N_10860,N_10139,N_9876);
and U10861 (N_10861,N_9841,N_10075);
nor U10862 (N_10862,N_9905,N_10079);
xor U10863 (N_10863,N_9890,N_9879);
and U10864 (N_10864,N_10209,N_9636);
nor U10865 (N_10865,N_10289,N_10309);
xnor U10866 (N_10866,N_10131,N_10082);
and U10867 (N_10867,N_10016,N_10192);
and U10868 (N_10868,N_9616,N_9690);
and U10869 (N_10869,N_9776,N_9725);
nor U10870 (N_10870,N_9661,N_10225);
and U10871 (N_10871,N_9647,N_9639);
or U10872 (N_10872,N_10043,N_10099);
or U10873 (N_10873,N_10092,N_9973);
and U10874 (N_10874,N_9838,N_9895);
xor U10875 (N_10875,N_10090,N_9878);
nand U10876 (N_10876,N_9907,N_9999);
or U10877 (N_10877,N_10377,N_9667);
or U10878 (N_10878,N_9886,N_9607);
nor U10879 (N_10879,N_10001,N_9674);
and U10880 (N_10880,N_10346,N_10090);
nor U10881 (N_10881,N_9646,N_9614);
xor U10882 (N_10882,N_10013,N_10312);
and U10883 (N_10883,N_9979,N_9604);
or U10884 (N_10884,N_10390,N_10183);
or U10885 (N_10885,N_9977,N_10158);
nand U10886 (N_10886,N_9699,N_10181);
and U10887 (N_10887,N_9892,N_10299);
or U10888 (N_10888,N_9982,N_10354);
xnor U10889 (N_10889,N_10243,N_9707);
or U10890 (N_10890,N_10008,N_10023);
or U10891 (N_10891,N_9887,N_10359);
and U10892 (N_10892,N_10154,N_10061);
nor U10893 (N_10893,N_9890,N_9690);
xor U10894 (N_10894,N_10062,N_10381);
xnor U10895 (N_10895,N_9621,N_9781);
nor U10896 (N_10896,N_10070,N_9656);
nand U10897 (N_10897,N_9602,N_10399);
nor U10898 (N_10898,N_9645,N_9806);
or U10899 (N_10899,N_9805,N_9715);
and U10900 (N_10900,N_10054,N_9872);
xnor U10901 (N_10901,N_9885,N_10192);
nor U10902 (N_10902,N_9725,N_10007);
or U10903 (N_10903,N_9897,N_10373);
nand U10904 (N_10904,N_9780,N_10076);
nand U10905 (N_10905,N_9807,N_9608);
nand U10906 (N_10906,N_9869,N_9850);
nor U10907 (N_10907,N_10189,N_9836);
or U10908 (N_10908,N_10064,N_10393);
nor U10909 (N_10909,N_10124,N_10226);
nand U10910 (N_10910,N_10340,N_9793);
nand U10911 (N_10911,N_10293,N_9977);
xnor U10912 (N_10912,N_10070,N_9917);
nor U10913 (N_10913,N_9874,N_10314);
and U10914 (N_10914,N_10092,N_10137);
nand U10915 (N_10915,N_10041,N_9681);
xnor U10916 (N_10916,N_9658,N_10119);
or U10917 (N_10917,N_9793,N_9764);
nand U10918 (N_10918,N_9966,N_9925);
or U10919 (N_10919,N_10222,N_10049);
xnor U10920 (N_10920,N_10039,N_9988);
or U10921 (N_10921,N_9854,N_9950);
and U10922 (N_10922,N_9778,N_9681);
nand U10923 (N_10923,N_10210,N_10134);
or U10924 (N_10924,N_10322,N_10009);
nand U10925 (N_10925,N_10066,N_9644);
xnor U10926 (N_10926,N_9736,N_9899);
xor U10927 (N_10927,N_10286,N_10282);
or U10928 (N_10928,N_10049,N_9972);
xor U10929 (N_10929,N_9610,N_10304);
nand U10930 (N_10930,N_9874,N_10130);
nor U10931 (N_10931,N_10043,N_9885);
and U10932 (N_10932,N_10275,N_9966);
xor U10933 (N_10933,N_10029,N_10071);
and U10934 (N_10934,N_10003,N_9849);
nor U10935 (N_10935,N_10012,N_9980);
nand U10936 (N_10936,N_9965,N_10301);
xor U10937 (N_10937,N_10179,N_9883);
and U10938 (N_10938,N_10003,N_9891);
and U10939 (N_10939,N_10246,N_9775);
or U10940 (N_10940,N_10222,N_10333);
or U10941 (N_10941,N_9834,N_9719);
xnor U10942 (N_10942,N_9886,N_9840);
and U10943 (N_10943,N_10113,N_10344);
xor U10944 (N_10944,N_9978,N_9831);
nand U10945 (N_10945,N_9939,N_9950);
nand U10946 (N_10946,N_10081,N_10239);
and U10947 (N_10947,N_10219,N_9852);
nor U10948 (N_10948,N_9660,N_9621);
xnor U10949 (N_10949,N_9976,N_9662);
or U10950 (N_10950,N_9761,N_9900);
xnor U10951 (N_10951,N_10062,N_10335);
nor U10952 (N_10952,N_9761,N_10066);
nor U10953 (N_10953,N_10217,N_10241);
or U10954 (N_10954,N_10174,N_9990);
nand U10955 (N_10955,N_9607,N_10125);
xor U10956 (N_10956,N_10096,N_9882);
nor U10957 (N_10957,N_9803,N_9604);
nor U10958 (N_10958,N_9807,N_10363);
nor U10959 (N_10959,N_10328,N_10354);
xnor U10960 (N_10960,N_10182,N_9886);
xor U10961 (N_10961,N_10050,N_10180);
nor U10962 (N_10962,N_10126,N_9897);
nand U10963 (N_10963,N_9657,N_10186);
xnor U10964 (N_10964,N_10129,N_9649);
xor U10965 (N_10965,N_10124,N_9974);
nand U10966 (N_10966,N_10260,N_9869);
and U10967 (N_10967,N_9871,N_9927);
nand U10968 (N_10968,N_9809,N_9941);
nand U10969 (N_10969,N_10140,N_10332);
xnor U10970 (N_10970,N_10332,N_9989);
xor U10971 (N_10971,N_10149,N_10161);
nand U10972 (N_10972,N_9838,N_9627);
or U10973 (N_10973,N_10388,N_10315);
xor U10974 (N_10974,N_10212,N_10270);
xnor U10975 (N_10975,N_10277,N_9785);
xnor U10976 (N_10976,N_10135,N_10273);
or U10977 (N_10977,N_10377,N_10182);
xor U10978 (N_10978,N_10302,N_10290);
nand U10979 (N_10979,N_9957,N_10252);
nand U10980 (N_10980,N_9884,N_10058);
xor U10981 (N_10981,N_10103,N_10388);
nand U10982 (N_10982,N_10228,N_10312);
xnor U10983 (N_10983,N_10258,N_10125);
and U10984 (N_10984,N_10244,N_9611);
nand U10985 (N_10985,N_9746,N_9633);
or U10986 (N_10986,N_9665,N_10065);
nor U10987 (N_10987,N_10303,N_10097);
nand U10988 (N_10988,N_10328,N_9815);
xor U10989 (N_10989,N_10178,N_9822);
nand U10990 (N_10990,N_10287,N_9844);
nor U10991 (N_10991,N_9905,N_10159);
nor U10992 (N_10992,N_9908,N_10293);
nor U10993 (N_10993,N_9944,N_10369);
xnor U10994 (N_10994,N_10368,N_10271);
xor U10995 (N_10995,N_9999,N_9648);
nand U10996 (N_10996,N_10275,N_9698);
nor U10997 (N_10997,N_9818,N_9772);
nand U10998 (N_10998,N_9710,N_10010);
xor U10999 (N_10999,N_9780,N_9852);
and U11000 (N_11000,N_9916,N_9666);
nand U11001 (N_11001,N_9653,N_10133);
xor U11002 (N_11002,N_9824,N_10395);
nor U11003 (N_11003,N_9859,N_10351);
or U11004 (N_11004,N_10280,N_9959);
and U11005 (N_11005,N_9965,N_9796);
nand U11006 (N_11006,N_9952,N_9984);
xnor U11007 (N_11007,N_10366,N_9613);
or U11008 (N_11008,N_10112,N_9928);
nand U11009 (N_11009,N_10026,N_10085);
xor U11010 (N_11010,N_9668,N_10280);
nand U11011 (N_11011,N_9906,N_9748);
or U11012 (N_11012,N_9731,N_10267);
nor U11013 (N_11013,N_10313,N_10008);
nand U11014 (N_11014,N_9652,N_10329);
or U11015 (N_11015,N_10064,N_10332);
or U11016 (N_11016,N_9816,N_9925);
xnor U11017 (N_11017,N_10152,N_10321);
nor U11018 (N_11018,N_10127,N_9843);
nand U11019 (N_11019,N_9810,N_10275);
and U11020 (N_11020,N_10315,N_10160);
or U11021 (N_11021,N_10304,N_10375);
nand U11022 (N_11022,N_9921,N_10047);
and U11023 (N_11023,N_9626,N_9710);
nor U11024 (N_11024,N_10327,N_9722);
xor U11025 (N_11025,N_9808,N_9627);
or U11026 (N_11026,N_10257,N_10233);
nor U11027 (N_11027,N_10260,N_9896);
and U11028 (N_11028,N_9984,N_9724);
nand U11029 (N_11029,N_9642,N_9695);
nor U11030 (N_11030,N_9968,N_10238);
or U11031 (N_11031,N_9751,N_9931);
xnor U11032 (N_11032,N_10047,N_10225);
xnor U11033 (N_11033,N_9891,N_10147);
or U11034 (N_11034,N_9997,N_10080);
nand U11035 (N_11035,N_10225,N_9856);
xnor U11036 (N_11036,N_10313,N_10223);
nand U11037 (N_11037,N_9671,N_9924);
or U11038 (N_11038,N_10139,N_9711);
or U11039 (N_11039,N_10097,N_10379);
nand U11040 (N_11040,N_9880,N_10341);
or U11041 (N_11041,N_10157,N_10317);
nand U11042 (N_11042,N_10150,N_10011);
nand U11043 (N_11043,N_9936,N_9995);
and U11044 (N_11044,N_10209,N_9975);
nor U11045 (N_11045,N_9799,N_10213);
and U11046 (N_11046,N_9796,N_10293);
xnor U11047 (N_11047,N_10361,N_10231);
or U11048 (N_11048,N_10327,N_9788);
and U11049 (N_11049,N_10347,N_9984);
nand U11050 (N_11050,N_10071,N_10381);
nor U11051 (N_11051,N_10225,N_9625);
and U11052 (N_11052,N_9630,N_9914);
or U11053 (N_11053,N_9983,N_10088);
xnor U11054 (N_11054,N_10057,N_10374);
and U11055 (N_11055,N_10218,N_9666);
nand U11056 (N_11056,N_9643,N_9736);
and U11057 (N_11057,N_9735,N_10006);
or U11058 (N_11058,N_9935,N_9976);
and U11059 (N_11059,N_10148,N_10126);
xnor U11060 (N_11060,N_10155,N_10225);
nand U11061 (N_11061,N_10023,N_10327);
nor U11062 (N_11062,N_9845,N_9786);
xor U11063 (N_11063,N_9603,N_9811);
nor U11064 (N_11064,N_9999,N_10073);
and U11065 (N_11065,N_9759,N_9999);
xor U11066 (N_11066,N_9852,N_10269);
nor U11067 (N_11067,N_10111,N_10185);
or U11068 (N_11068,N_10155,N_10295);
and U11069 (N_11069,N_9611,N_10156);
and U11070 (N_11070,N_10165,N_10289);
and U11071 (N_11071,N_9880,N_9955);
or U11072 (N_11072,N_9777,N_9668);
and U11073 (N_11073,N_10042,N_10311);
and U11074 (N_11074,N_10137,N_10000);
or U11075 (N_11075,N_10164,N_9795);
or U11076 (N_11076,N_10371,N_10099);
nand U11077 (N_11077,N_9675,N_9608);
nand U11078 (N_11078,N_9755,N_9707);
and U11079 (N_11079,N_9817,N_10351);
or U11080 (N_11080,N_10015,N_9733);
or U11081 (N_11081,N_9724,N_10331);
xor U11082 (N_11082,N_9787,N_10169);
and U11083 (N_11083,N_9921,N_10165);
and U11084 (N_11084,N_9881,N_9842);
or U11085 (N_11085,N_9641,N_9715);
xor U11086 (N_11086,N_9754,N_10021);
nor U11087 (N_11087,N_9991,N_9926);
nor U11088 (N_11088,N_9841,N_9941);
nor U11089 (N_11089,N_10284,N_9870);
nor U11090 (N_11090,N_10339,N_9948);
xor U11091 (N_11091,N_10224,N_10296);
nor U11092 (N_11092,N_10018,N_9668);
xnor U11093 (N_11093,N_9681,N_9657);
and U11094 (N_11094,N_9939,N_10264);
and U11095 (N_11095,N_9605,N_10080);
and U11096 (N_11096,N_9678,N_9849);
nor U11097 (N_11097,N_9615,N_9768);
nor U11098 (N_11098,N_9801,N_10139);
nand U11099 (N_11099,N_9863,N_9706);
nand U11100 (N_11100,N_10116,N_9701);
and U11101 (N_11101,N_9728,N_9919);
nor U11102 (N_11102,N_9739,N_9797);
xnor U11103 (N_11103,N_10144,N_9864);
nand U11104 (N_11104,N_10018,N_9612);
or U11105 (N_11105,N_9612,N_10127);
or U11106 (N_11106,N_9694,N_10388);
nand U11107 (N_11107,N_10167,N_10381);
or U11108 (N_11108,N_9977,N_10260);
or U11109 (N_11109,N_9900,N_9699);
nor U11110 (N_11110,N_10083,N_10054);
xnor U11111 (N_11111,N_9779,N_9878);
nor U11112 (N_11112,N_9790,N_10090);
or U11113 (N_11113,N_9694,N_9613);
nand U11114 (N_11114,N_9819,N_10155);
or U11115 (N_11115,N_9860,N_10049);
nand U11116 (N_11116,N_9835,N_9776);
nor U11117 (N_11117,N_10151,N_9974);
and U11118 (N_11118,N_10222,N_10066);
nor U11119 (N_11119,N_9911,N_9664);
xor U11120 (N_11120,N_9993,N_10275);
nand U11121 (N_11121,N_9615,N_9650);
or U11122 (N_11122,N_9783,N_9873);
and U11123 (N_11123,N_10374,N_9978);
or U11124 (N_11124,N_9892,N_10145);
nor U11125 (N_11125,N_9631,N_10354);
or U11126 (N_11126,N_9991,N_9776);
and U11127 (N_11127,N_9768,N_10267);
and U11128 (N_11128,N_10386,N_9812);
xor U11129 (N_11129,N_9989,N_9709);
nor U11130 (N_11130,N_10129,N_9700);
and U11131 (N_11131,N_10234,N_9914);
and U11132 (N_11132,N_10112,N_9601);
and U11133 (N_11133,N_9924,N_9871);
or U11134 (N_11134,N_9778,N_9755);
nor U11135 (N_11135,N_10164,N_10237);
xor U11136 (N_11136,N_9804,N_9973);
or U11137 (N_11137,N_10033,N_9974);
or U11138 (N_11138,N_9643,N_9719);
or U11139 (N_11139,N_10175,N_9927);
and U11140 (N_11140,N_9861,N_10182);
nand U11141 (N_11141,N_10284,N_10390);
or U11142 (N_11142,N_10348,N_9890);
or U11143 (N_11143,N_9916,N_10112);
nor U11144 (N_11144,N_9935,N_9986);
nand U11145 (N_11145,N_10297,N_10219);
or U11146 (N_11146,N_10033,N_10338);
and U11147 (N_11147,N_10350,N_9872);
nand U11148 (N_11148,N_10101,N_10325);
nor U11149 (N_11149,N_10042,N_10151);
xnor U11150 (N_11150,N_10275,N_9996);
nand U11151 (N_11151,N_9764,N_9635);
or U11152 (N_11152,N_9720,N_10223);
or U11153 (N_11153,N_10341,N_9670);
xnor U11154 (N_11154,N_9779,N_9860);
xor U11155 (N_11155,N_9909,N_9960);
or U11156 (N_11156,N_9702,N_9906);
nand U11157 (N_11157,N_10258,N_9808);
and U11158 (N_11158,N_10148,N_9740);
and U11159 (N_11159,N_9805,N_9773);
xnor U11160 (N_11160,N_9844,N_10137);
nor U11161 (N_11161,N_9957,N_10318);
xnor U11162 (N_11162,N_10292,N_9697);
nand U11163 (N_11163,N_10268,N_9947);
or U11164 (N_11164,N_9756,N_9708);
and U11165 (N_11165,N_9737,N_9745);
nand U11166 (N_11166,N_9749,N_10056);
xnor U11167 (N_11167,N_9622,N_10326);
nor U11168 (N_11168,N_10188,N_9629);
nor U11169 (N_11169,N_9737,N_9709);
xnor U11170 (N_11170,N_9882,N_10265);
nor U11171 (N_11171,N_9615,N_9904);
and U11172 (N_11172,N_9739,N_10051);
or U11173 (N_11173,N_10094,N_10012);
nor U11174 (N_11174,N_9729,N_9741);
nor U11175 (N_11175,N_9846,N_9828);
xor U11176 (N_11176,N_9905,N_10337);
or U11177 (N_11177,N_10071,N_10121);
and U11178 (N_11178,N_9619,N_9755);
or U11179 (N_11179,N_10055,N_9612);
nand U11180 (N_11180,N_9601,N_9600);
and U11181 (N_11181,N_9650,N_10236);
and U11182 (N_11182,N_10045,N_10155);
xor U11183 (N_11183,N_9651,N_10359);
nor U11184 (N_11184,N_9661,N_9861);
xnor U11185 (N_11185,N_10213,N_10097);
or U11186 (N_11186,N_10284,N_10354);
nor U11187 (N_11187,N_9847,N_9771);
xor U11188 (N_11188,N_10240,N_10304);
xor U11189 (N_11189,N_10062,N_9753);
or U11190 (N_11190,N_10149,N_9664);
nor U11191 (N_11191,N_9892,N_10314);
xor U11192 (N_11192,N_10096,N_10391);
and U11193 (N_11193,N_10141,N_10347);
nor U11194 (N_11194,N_10286,N_9753);
nor U11195 (N_11195,N_10305,N_9673);
and U11196 (N_11196,N_10232,N_9914);
and U11197 (N_11197,N_10167,N_9937);
xnor U11198 (N_11198,N_9735,N_10033);
xnor U11199 (N_11199,N_10126,N_9812);
nand U11200 (N_11200,N_10686,N_10988);
and U11201 (N_11201,N_10808,N_10641);
xor U11202 (N_11202,N_11060,N_11162);
nand U11203 (N_11203,N_11171,N_10456);
and U11204 (N_11204,N_10601,N_10602);
nor U11205 (N_11205,N_10718,N_10961);
and U11206 (N_11206,N_11124,N_11091);
or U11207 (N_11207,N_11042,N_11054);
nand U11208 (N_11208,N_10584,N_11051);
xor U11209 (N_11209,N_10532,N_10692);
xnor U11210 (N_11210,N_11057,N_10603);
nand U11211 (N_11211,N_10680,N_11035);
nor U11212 (N_11212,N_10870,N_10559);
nor U11213 (N_11213,N_10535,N_10514);
or U11214 (N_11214,N_10931,N_10442);
or U11215 (N_11215,N_11021,N_11183);
or U11216 (N_11216,N_10834,N_10461);
nor U11217 (N_11217,N_10430,N_10866);
nor U11218 (N_11218,N_10951,N_11081);
nand U11219 (N_11219,N_10582,N_10463);
and U11220 (N_11220,N_10417,N_10520);
nand U11221 (N_11221,N_11096,N_11003);
or U11222 (N_11222,N_10590,N_10581);
or U11223 (N_11223,N_11000,N_10803);
or U11224 (N_11224,N_10760,N_10571);
and U11225 (N_11225,N_10861,N_11182);
or U11226 (N_11226,N_10560,N_10886);
nor U11227 (N_11227,N_10794,N_10972);
nor U11228 (N_11228,N_10495,N_10966);
and U11229 (N_11229,N_10554,N_10478);
nand U11230 (N_11230,N_10848,N_10657);
nand U11231 (N_11231,N_11150,N_10466);
nor U11232 (N_11232,N_11020,N_11193);
xnor U11233 (N_11233,N_10492,N_11058);
xor U11234 (N_11234,N_10565,N_10955);
and U11235 (N_11235,N_10599,N_11041);
nor U11236 (N_11236,N_10432,N_10898);
nand U11237 (N_11237,N_10837,N_11009);
and U11238 (N_11238,N_10850,N_10756);
nand U11239 (N_11239,N_10428,N_11194);
or U11240 (N_11240,N_10563,N_11053);
nor U11241 (N_11241,N_11069,N_10690);
nor U11242 (N_11242,N_10637,N_10426);
nand U11243 (N_11243,N_10856,N_10684);
or U11244 (N_11244,N_10632,N_10780);
and U11245 (N_11245,N_11098,N_11139);
and U11246 (N_11246,N_11191,N_10618);
xnor U11247 (N_11247,N_11110,N_10800);
and U11248 (N_11248,N_10784,N_10516);
xnor U11249 (N_11249,N_10405,N_10630);
nor U11250 (N_11250,N_10928,N_10607);
nor U11251 (N_11251,N_10593,N_10896);
xor U11252 (N_11252,N_10673,N_10990);
and U11253 (N_11253,N_10653,N_10859);
and U11254 (N_11254,N_10422,N_10869);
and U11255 (N_11255,N_10787,N_11169);
nor U11256 (N_11256,N_11026,N_10893);
xor U11257 (N_11257,N_11146,N_10579);
and U11258 (N_11258,N_10408,N_10687);
xnor U11259 (N_11259,N_10773,N_10615);
nor U11260 (N_11260,N_10711,N_10853);
xor U11261 (N_11261,N_11100,N_11056);
xnor U11262 (N_11262,N_10746,N_10851);
and U11263 (N_11263,N_10830,N_11032);
nor U11264 (N_11264,N_10811,N_10863);
and U11265 (N_11265,N_11031,N_11185);
and U11266 (N_11266,N_10805,N_10598);
xor U11267 (N_11267,N_10524,N_10675);
nand U11268 (N_11268,N_10788,N_11155);
nor U11269 (N_11269,N_11163,N_10839);
and U11270 (N_11270,N_10676,N_10564);
xnor U11271 (N_11271,N_10908,N_10454);
or U11272 (N_11272,N_10505,N_10846);
or U11273 (N_11273,N_10439,N_11095);
xnor U11274 (N_11274,N_10977,N_10715);
nand U11275 (N_11275,N_10433,N_10576);
and U11276 (N_11276,N_11006,N_10752);
nor U11277 (N_11277,N_10651,N_11038);
nor U11278 (N_11278,N_10731,N_10726);
and U11279 (N_11279,N_10522,N_11055);
nand U11280 (N_11280,N_10538,N_10915);
or U11281 (N_11281,N_11074,N_10695);
or U11282 (N_11282,N_10566,N_11092);
nor U11283 (N_11283,N_11174,N_10874);
xnor U11284 (N_11284,N_10665,N_10710);
xor U11285 (N_11285,N_11187,N_10663);
and U11286 (N_11286,N_10763,N_10660);
xnor U11287 (N_11287,N_10424,N_10625);
and U11288 (N_11288,N_10713,N_10844);
xor U11289 (N_11289,N_10646,N_10407);
nand U11290 (N_11290,N_11131,N_10926);
and U11291 (N_11291,N_10555,N_11173);
nor U11292 (N_11292,N_10714,N_10472);
xor U11293 (N_11293,N_10515,N_10790);
xnor U11294 (N_11294,N_11080,N_10556);
nand U11295 (N_11295,N_10943,N_11125);
nand U11296 (N_11296,N_10677,N_10785);
nand U11297 (N_11297,N_11177,N_10883);
nor U11298 (N_11298,N_10523,N_10789);
or U11299 (N_11299,N_10455,N_10936);
nor U11300 (N_11300,N_11152,N_10628);
or U11301 (N_11301,N_10580,N_10412);
xor U11302 (N_11302,N_10828,N_10669);
and U11303 (N_11303,N_11186,N_10768);
or U11304 (N_11304,N_11168,N_10735);
xnor U11305 (N_11305,N_11180,N_10402);
and U11306 (N_11306,N_10403,N_10659);
or U11307 (N_11307,N_11199,N_11130);
xnor U11308 (N_11308,N_10567,N_10799);
nand U11309 (N_11309,N_10624,N_11044);
nor U11310 (N_11310,N_10414,N_10613);
nor U11311 (N_11311,N_10815,N_10434);
and U11312 (N_11312,N_11024,N_10871);
or U11313 (N_11313,N_11103,N_10450);
and U11314 (N_11314,N_10410,N_10553);
or U11315 (N_11315,N_11153,N_10994);
nand U11316 (N_11316,N_11076,N_10526);
or U11317 (N_11317,N_11105,N_10777);
and U11318 (N_11318,N_10849,N_10451);
nand U11319 (N_11319,N_10840,N_10502);
or U11320 (N_11320,N_10948,N_11065);
nor U11321 (N_11321,N_10823,N_10476);
and U11322 (N_11322,N_10724,N_10647);
nor U11323 (N_11323,N_10652,N_10758);
or U11324 (N_11324,N_10499,N_10699);
xor U11325 (N_11325,N_10448,N_11166);
xor U11326 (N_11326,N_10479,N_10864);
and U11327 (N_11327,N_10689,N_10767);
and U11328 (N_11328,N_11114,N_11008);
xor U11329 (N_11329,N_11197,N_10674);
xnor U11330 (N_11330,N_10987,N_10529);
xor U11331 (N_11331,N_10513,N_11039);
xnor U11332 (N_11332,N_10645,N_10757);
or U11333 (N_11333,N_10818,N_10501);
nand U11334 (N_11334,N_10542,N_11101);
or U11335 (N_11335,N_10667,N_11178);
nor U11336 (N_11336,N_10539,N_10435);
or U11337 (N_11337,N_11135,N_11147);
and U11338 (N_11338,N_10493,N_11160);
nor U11339 (N_11339,N_10879,N_11047);
xnor U11340 (N_11340,N_10950,N_10901);
and U11341 (N_11341,N_10895,N_10927);
xor U11342 (N_11342,N_10894,N_10678);
nand U11343 (N_11343,N_10500,N_11002);
or U11344 (N_11344,N_10740,N_10816);
and U11345 (N_11345,N_10610,N_11090);
nand U11346 (N_11346,N_10427,N_11107);
nor U11347 (N_11347,N_10983,N_11070);
xnor U11348 (N_11348,N_11083,N_10989);
or U11349 (N_11349,N_10916,N_10964);
nand U11350 (N_11350,N_10981,N_11001);
nand U11351 (N_11351,N_10445,N_10709);
and U11352 (N_11352,N_11075,N_11025);
nor U11353 (N_11353,N_10764,N_10875);
or U11354 (N_11354,N_10570,N_10540);
or U11355 (N_11355,N_11145,N_10852);
nand U11356 (N_11356,N_10716,N_10934);
xor U11357 (N_11357,N_10587,N_10804);
and U11358 (N_11358,N_10619,N_10732);
and U11359 (N_11359,N_10993,N_10545);
or U11360 (N_11360,N_10881,N_10719);
nand U11361 (N_11361,N_11007,N_10820);
nand U11362 (N_11362,N_10795,N_10945);
nor U11363 (N_11363,N_10420,N_10986);
nor U11364 (N_11364,N_10832,N_10939);
xor U11365 (N_11365,N_10829,N_10616);
nor U11366 (N_11366,N_10855,N_10666);
or U11367 (N_11367,N_11141,N_10594);
nor U11368 (N_11368,N_10998,N_10958);
nor U11369 (N_11369,N_10888,N_11167);
or U11370 (N_11370,N_10507,N_11013);
xor U11371 (N_11371,N_10544,N_10679);
or U11372 (N_11372,N_10457,N_10462);
nor U11373 (N_11373,N_11102,N_10867);
xor U11374 (N_11374,N_11028,N_10668);
nor U11375 (N_11375,N_11071,N_10723);
and U11376 (N_11376,N_10779,N_11018);
xor U11377 (N_11377,N_10798,N_10868);
xnor U11378 (N_11378,N_10793,N_10586);
nand U11379 (N_11379,N_10985,N_10890);
xnor U11380 (N_11380,N_11108,N_10683);
nor U11381 (N_11381,N_10591,N_10952);
nand U11382 (N_11382,N_11159,N_10940);
nand U11383 (N_11383,N_11190,N_10494);
or U11384 (N_11384,N_11086,N_10585);
or U11385 (N_11385,N_10425,N_10980);
or U11386 (N_11386,N_10503,N_10892);
xnor U11387 (N_11387,N_10569,N_11078);
xnor U11388 (N_11388,N_10459,N_10708);
and U11389 (N_11389,N_10473,N_10534);
or U11390 (N_11390,N_10743,N_10845);
xor U11391 (N_11391,N_11136,N_11094);
xor U11392 (N_11392,N_10842,N_11115);
nand U11393 (N_11393,N_10865,N_10992);
and U11394 (N_11394,N_11085,N_10596);
nand U11395 (N_11395,N_10877,N_10400);
xnor U11396 (N_11396,N_10819,N_10949);
nand U11397 (N_11397,N_10791,N_10860);
nand U11398 (N_11398,N_11132,N_10761);
and U11399 (N_11399,N_10588,N_10976);
and U11400 (N_11400,N_10919,N_10991);
nor U11401 (N_11401,N_11104,N_11109);
xor U11402 (N_11402,N_10750,N_10612);
nor U11403 (N_11403,N_10648,N_10906);
and U11404 (N_11404,N_10662,N_10491);
or U11405 (N_11405,N_10480,N_11005);
xor U11406 (N_11406,N_10626,N_10826);
and U11407 (N_11407,N_10975,N_10464);
xor U11408 (N_11408,N_11034,N_10490);
xnor U11409 (N_11409,N_11120,N_10749);
and U11410 (N_11410,N_10720,N_10418);
xnor U11411 (N_11411,N_11142,N_10882);
nor U11412 (N_11412,N_11176,N_10910);
nor U11413 (N_11413,N_10772,N_10727);
nand U11414 (N_11414,N_10781,N_10485);
xor U11415 (N_11415,N_10912,N_10629);
or U11416 (N_11416,N_10775,N_11154);
nand U11417 (N_11417,N_10688,N_10941);
and U11418 (N_11418,N_10621,N_11046);
or U11419 (N_11419,N_10960,N_11122);
xnor U11420 (N_11420,N_10944,N_11172);
or U11421 (N_11421,N_11134,N_10982);
nand U11422 (N_11422,N_10835,N_11052);
or U11423 (N_11423,N_10914,N_10631);
xor U11424 (N_11424,N_10909,N_10738);
or U11425 (N_11425,N_10600,N_10452);
xor U11426 (N_11426,N_10627,N_10814);
and U11427 (N_11427,N_11099,N_10801);
nor U11428 (N_11428,N_11027,N_10918);
nand U11429 (N_11429,N_11037,N_10970);
nor U11430 (N_11430,N_10670,N_10510);
xor U11431 (N_11431,N_10401,N_10921);
and U11432 (N_11432,N_10880,N_10622);
nand U11433 (N_11433,N_10444,N_10460);
or U11434 (N_11434,N_10971,N_10953);
and U11435 (N_11435,N_11010,N_10744);
and U11436 (N_11436,N_10857,N_10900);
nand U11437 (N_11437,N_10736,N_10449);
and U11438 (N_11438,N_10568,N_10447);
nor U11439 (N_11439,N_11188,N_10691);
xor U11440 (N_11440,N_10656,N_10946);
xor U11441 (N_11441,N_10620,N_10833);
xor U11442 (N_11442,N_10640,N_10962);
nor U11443 (N_11443,N_11004,N_10717);
or U11444 (N_11444,N_10937,N_10932);
or U11445 (N_11445,N_10617,N_10644);
xor U11446 (N_11446,N_10712,N_10745);
nand U11447 (N_11447,N_10705,N_10753);
nand U11448 (N_11448,N_11040,N_10595);
or U11449 (N_11449,N_10742,N_10959);
nand U11450 (N_11450,N_11111,N_10899);
nand U11451 (N_11451,N_11161,N_10655);
and U11452 (N_11452,N_10809,N_10694);
nand U11453 (N_11453,N_11014,N_10506);
xor U11454 (N_11454,N_11068,N_10623);
nor U11455 (N_11455,N_10889,N_11093);
nand U11456 (N_11456,N_10557,N_10443);
nor U11457 (N_11457,N_10702,N_10649);
nand U11458 (N_11458,N_10671,N_10697);
nand U11459 (N_11459,N_10891,N_11088);
xnor U11460 (N_11460,N_10920,N_10481);
xnor U11461 (N_11461,N_10550,N_10562);
and U11462 (N_11462,N_10606,N_10583);
or U11463 (N_11463,N_10887,N_10498);
and U11464 (N_11464,N_10872,N_11116);
nor U11465 (N_11465,N_11048,N_10947);
xor U11466 (N_11466,N_10415,N_10905);
nor U11467 (N_11467,N_11113,N_10527);
xor U11468 (N_11468,N_10437,N_11181);
and U11469 (N_11469,N_11126,N_10796);
xor U11470 (N_11470,N_10807,N_10774);
xnor U11471 (N_11471,N_10822,N_10973);
or U11472 (N_11472,N_10817,N_10517);
xor U11473 (N_11473,N_11045,N_10551);
xnor U11474 (N_11474,N_10634,N_10821);
and U11475 (N_11475,N_10547,N_11022);
xor U11476 (N_11476,N_10733,N_10897);
or U11477 (N_11477,N_10813,N_10797);
and U11478 (N_11478,N_10783,N_10923);
nor U11479 (N_11479,N_10664,N_10831);
nor U11480 (N_11480,N_10843,N_10995);
xnor U11481 (N_11481,N_11119,N_11165);
or U11482 (N_11482,N_11192,N_11140);
or U11483 (N_11483,N_10924,N_10786);
and U11484 (N_11484,N_10838,N_10737);
or U11485 (N_11485,N_10770,N_10812);
or U11486 (N_11486,N_11143,N_10543);
xor U11487 (N_11487,N_11158,N_10605);
and U11488 (N_11488,N_10636,N_10537);
nand U11489 (N_11489,N_11059,N_10438);
and U11490 (N_11490,N_10486,N_11087);
and U11491 (N_11491,N_10754,N_10474);
or U11492 (N_11492,N_10873,N_10913);
nand U11493 (N_11493,N_10672,N_11164);
nand U11494 (N_11494,N_10984,N_11189);
nand U11495 (N_11495,N_10825,N_10876);
xnor U11496 (N_11496,N_10802,N_11149);
and U11497 (N_11497,N_10458,N_10903);
and U11498 (N_11498,N_11029,N_10531);
xor U11499 (N_11499,N_11066,N_10766);
xor U11500 (N_11500,N_10696,N_10858);
nor U11501 (N_11501,N_10416,N_10609);
nor U11502 (N_11502,N_10525,N_10701);
xnor U11503 (N_11503,N_11106,N_11063);
xnor U11504 (N_11504,N_10465,N_10475);
and U11505 (N_11505,N_10483,N_11097);
xor U11506 (N_11506,N_10650,N_10762);
nor U11507 (N_11507,N_10963,N_10854);
or U11508 (N_11508,N_11133,N_11129);
nor U11509 (N_11509,N_11156,N_10935);
and U11510 (N_11510,N_10824,N_11016);
and U11511 (N_11511,N_11067,N_10488);
or U11512 (N_11512,N_11019,N_10759);
xor U11513 (N_11513,N_10413,N_10658);
or U11514 (N_11514,N_10453,N_10643);
xnor U11515 (N_11515,N_10572,N_10721);
xnor U11516 (N_11516,N_10611,N_10575);
or U11517 (N_11517,N_10885,N_10771);
or U11518 (N_11518,N_11036,N_11138);
nand U11519 (N_11519,N_10925,N_10954);
nand U11520 (N_11520,N_10968,N_10755);
or U11521 (N_11521,N_11157,N_10608);
nor U11522 (N_11522,N_10902,N_10552);
xnor U11523 (N_11523,N_10969,N_10996);
nor U11524 (N_11524,N_10827,N_10654);
and U11525 (N_11525,N_10446,N_11084);
and U11526 (N_11526,N_10633,N_10508);
or U11527 (N_11527,N_10978,N_10884);
and U11528 (N_11528,N_10421,N_10518);
nand U11529 (N_11529,N_10778,N_10782);
or U11530 (N_11530,N_10578,N_10470);
xnor U11531 (N_11531,N_11184,N_10748);
or U11532 (N_11532,N_10706,N_11079);
nor U11533 (N_11533,N_10878,N_10792);
xor U11534 (N_11534,N_10776,N_10703);
and U11535 (N_11535,N_10406,N_11073);
nor U11536 (N_11536,N_10979,N_10635);
xnor U11537 (N_11537,N_10577,N_11015);
nor U11538 (N_11538,N_10836,N_10734);
or U11539 (N_11539,N_11077,N_10521);
nand U11540 (N_11540,N_10722,N_10419);
or U11541 (N_11541,N_10751,N_10546);
nor U11542 (N_11542,N_10489,N_10471);
nor U11543 (N_11543,N_10862,N_11137);
xor U11544 (N_11544,N_10440,N_11030);
or U11545 (N_11545,N_10693,N_10592);
xnor U11546 (N_11546,N_10469,N_10504);
nor U11547 (N_11547,N_10642,N_11082);
or U11548 (N_11548,N_11023,N_10614);
and U11549 (N_11549,N_11012,N_11144);
and U11550 (N_11550,N_11198,N_11064);
nand U11551 (N_11551,N_10511,N_10841);
nand U11552 (N_11552,N_10436,N_10965);
and U11553 (N_11553,N_10541,N_10638);
nor U11554 (N_11554,N_11112,N_10431);
nor U11555 (N_11555,N_11061,N_11043);
nor U11556 (N_11556,N_10904,N_11196);
xor U11557 (N_11557,N_10967,N_11050);
nor U11558 (N_11558,N_10661,N_10974);
or U11559 (N_11559,N_10639,N_10938);
or U11560 (N_11560,N_10681,N_10685);
xor U11561 (N_11561,N_10729,N_10533);
nand U11562 (N_11562,N_10997,N_11117);
or U11563 (N_11563,N_10956,N_10739);
and U11564 (N_11564,N_10911,N_10573);
and U11565 (N_11565,N_11151,N_10704);
nand U11566 (N_11566,N_10741,N_10536);
and U11567 (N_11567,N_11123,N_11062);
or U11568 (N_11568,N_10574,N_10847);
and U11569 (N_11569,N_11118,N_10806);
and U11570 (N_11570,N_10549,N_10528);
xor U11571 (N_11571,N_10423,N_11033);
or U11572 (N_11572,N_10730,N_10597);
or U11573 (N_11573,N_10769,N_10441);
or U11574 (N_11574,N_10409,N_10477);
and U11575 (N_11575,N_10682,N_11089);
xor U11576 (N_11576,N_10930,N_10707);
or U11577 (N_11577,N_11072,N_11179);
xor U11578 (N_11578,N_11017,N_10411);
or U11579 (N_11579,N_11170,N_10484);
nor U11580 (N_11580,N_11121,N_10530);
or U11581 (N_11581,N_10512,N_10700);
nand U11582 (N_11582,N_10999,N_10482);
nand U11583 (N_11583,N_10942,N_10957);
and U11584 (N_11584,N_10487,N_11049);
nor U11585 (N_11585,N_11128,N_10933);
or U11586 (N_11586,N_11195,N_10497);
xnor U11587 (N_11587,N_10907,N_10558);
nand U11588 (N_11588,N_10725,N_10728);
xnor U11589 (N_11589,N_11175,N_10509);
or U11590 (N_11590,N_10467,N_10404);
or U11591 (N_11591,N_10561,N_10810);
or U11592 (N_11592,N_10519,N_10468);
xnor U11593 (N_11593,N_10589,N_10429);
and U11594 (N_11594,N_10548,N_10604);
or U11595 (N_11595,N_10698,N_10765);
and U11596 (N_11596,N_10747,N_10922);
and U11597 (N_11597,N_10929,N_10496);
nor U11598 (N_11598,N_11127,N_11011);
and U11599 (N_11599,N_11148,N_10917);
nand U11600 (N_11600,N_10463,N_10417);
or U11601 (N_11601,N_10681,N_10406);
xnor U11602 (N_11602,N_10485,N_10648);
nand U11603 (N_11603,N_10731,N_10762);
or U11604 (N_11604,N_10472,N_10663);
xor U11605 (N_11605,N_11051,N_11155);
xnor U11606 (N_11606,N_10597,N_10485);
nor U11607 (N_11607,N_10519,N_10753);
nor U11608 (N_11608,N_10607,N_10927);
or U11609 (N_11609,N_11154,N_10648);
or U11610 (N_11610,N_11165,N_10565);
nor U11611 (N_11611,N_10943,N_10931);
and U11612 (N_11612,N_10403,N_10835);
xor U11613 (N_11613,N_11000,N_11146);
and U11614 (N_11614,N_10888,N_10605);
and U11615 (N_11615,N_10562,N_10728);
nand U11616 (N_11616,N_10971,N_10985);
nor U11617 (N_11617,N_10957,N_10923);
nand U11618 (N_11618,N_10472,N_10785);
nor U11619 (N_11619,N_11080,N_10632);
xnor U11620 (N_11620,N_10659,N_10513);
nand U11621 (N_11621,N_11016,N_10447);
nor U11622 (N_11622,N_10703,N_10566);
nor U11623 (N_11623,N_10677,N_10683);
nand U11624 (N_11624,N_10815,N_10419);
and U11625 (N_11625,N_11110,N_10651);
xor U11626 (N_11626,N_10763,N_10817);
nand U11627 (N_11627,N_11072,N_11019);
or U11628 (N_11628,N_11125,N_10876);
nand U11629 (N_11629,N_10959,N_11102);
nand U11630 (N_11630,N_11002,N_10609);
xnor U11631 (N_11631,N_10549,N_10458);
and U11632 (N_11632,N_10650,N_10608);
and U11633 (N_11633,N_10981,N_10749);
nor U11634 (N_11634,N_10479,N_10417);
or U11635 (N_11635,N_10577,N_11153);
or U11636 (N_11636,N_10453,N_11091);
or U11637 (N_11637,N_10876,N_10647);
nand U11638 (N_11638,N_10475,N_10738);
or U11639 (N_11639,N_11133,N_11172);
nor U11640 (N_11640,N_10823,N_10846);
nand U11641 (N_11641,N_10685,N_10944);
nand U11642 (N_11642,N_10756,N_11181);
and U11643 (N_11643,N_10574,N_10773);
or U11644 (N_11644,N_10838,N_10401);
or U11645 (N_11645,N_10851,N_11092);
nand U11646 (N_11646,N_10785,N_10974);
nand U11647 (N_11647,N_10541,N_10903);
xor U11648 (N_11648,N_10982,N_10552);
or U11649 (N_11649,N_10678,N_10793);
xnor U11650 (N_11650,N_10759,N_10621);
nand U11651 (N_11651,N_10443,N_10688);
and U11652 (N_11652,N_10710,N_10818);
xnor U11653 (N_11653,N_10918,N_11037);
and U11654 (N_11654,N_10735,N_10519);
and U11655 (N_11655,N_10638,N_10628);
nor U11656 (N_11656,N_10966,N_10756);
or U11657 (N_11657,N_10984,N_10444);
or U11658 (N_11658,N_10949,N_10780);
xnor U11659 (N_11659,N_10571,N_10716);
or U11660 (N_11660,N_10886,N_10638);
xnor U11661 (N_11661,N_11071,N_10957);
or U11662 (N_11662,N_10647,N_10568);
xnor U11663 (N_11663,N_10435,N_10635);
xor U11664 (N_11664,N_10580,N_10823);
nor U11665 (N_11665,N_10544,N_11095);
nand U11666 (N_11666,N_10426,N_10794);
and U11667 (N_11667,N_11017,N_11098);
nand U11668 (N_11668,N_10419,N_11022);
nand U11669 (N_11669,N_11145,N_10613);
xnor U11670 (N_11670,N_11131,N_10584);
xor U11671 (N_11671,N_10419,N_10477);
or U11672 (N_11672,N_10987,N_10788);
xnor U11673 (N_11673,N_10749,N_10934);
nor U11674 (N_11674,N_11094,N_10890);
xnor U11675 (N_11675,N_10740,N_11028);
or U11676 (N_11676,N_10900,N_10501);
nand U11677 (N_11677,N_10852,N_10770);
and U11678 (N_11678,N_11110,N_10428);
and U11679 (N_11679,N_10706,N_10537);
or U11680 (N_11680,N_10908,N_10497);
or U11681 (N_11681,N_11006,N_10792);
xnor U11682 (N_11682,N_10944,N_10727);
and U11683 (N_11683,N_11195,N_10871);
xnor U11684 (N_11684,N_10615,N_10447);
nor U11685 (N_11685,N_10768,N_11015);
xor U11686 (N_11686,N_10521,N_10767);
or U11687 (N_11687,N_10704,N_10476);
nand U11688 (N_11688,N_10837,N_10852);
or U11689 (N_11689,N_11099,N_10715);
xor U11690 (N_11690,N_10945,N_10769);
or U11691 (N_11691,N_10726,N_10478);
nand U11692 (N_11692,N_10783,N_11190);
xnor U11693 (N_11693,N_10748,N_10514);
nor U11694 (N_11694,N_11170,N_10730);
and U11695 (N_11695,N_10676,N_10846);
and U11696 (N_11696,N_10951,N_11144);
or U11697 (N_11697,N_10720,N_11016);
nand U11698 (N_11698,N_10559,N_10861);
xnor U11699 (N_11699,N_11171,N_11051);
or U11700 (N_11700,N_10669,N_10763);
nand U11701 (N_11701,N_10689,N_10933);
or U11702 (N_11702,N_10465,N_11086);
or U11703 (N_11703,N_10514,N_10789);
nand U11704 (N_11704,N_10455,N_11197);
or U11705 (N_11705,N_11049,N_10425);
nor U11706 (N_11706,N_10691,N_11113);
and U11707 (N_11707,N_10688,N_10540);
xnor U11708 (N_11708,N_10948,N_10769);
nand U11709 (N_11709,N_10744,N_10500);
and U11710 (N_11710,N_11167,N_10835);
nand U11711 (N_11711,N_10476,N_10940);
nor U11712 (N_11712,N_10471,N_11080);
xnor U11713 (N_11713,N_10446,N_10577);
nand U11714 (N_11714,N_10637,N_10924);
nand U11715 (N_11715,N_10451,N_10864);
or U11716 (N_11716,N_11029,N_10998);
nand U11717 (N_11717,N_10506,N_10919);
nor U11718 (N_11718,N_10474,N_10654);
xor U11719 (N_11719,N_10745,N_11049);
nand U11720 (N_11720,N_10453,N_10553);
or U11721 (N_11721,N_10855,N_10567);
nor U11722 (N_11722,N_11193,N_11171);
xor U11723 (N_11723,N_10547,N_11011);
nand U11724 (N_11724,N_10721,N_10743);
nor U11725 (N_11725,N_10765,N_10840);
nor U11726 (N_11726,N_10959,N_11021);
or U11727 (N_11727,N_11146,N_10813);
and U11728 (N_11728,N_10682,N_10775);
and U11729 (N_11729,N_10509,N_10939);
or U11730 (N_11730,N_10716,N_10497);
or U11731 (N_11731,N_10569,N_10545);
nor U11732 (N_11732,N_11172,N_10784);
and U11733 (N_11733,N_10997,N_10765);
nor U11734 (N_11734,N_10838,N_10547);
nor U11735 (N_11735,N_10540,N_10433);
and U11736 (N_11736,N_11171,N_10531);
nor U11737 (N_11737,N_10864,N_10589);
nor U11738 (N_11738,N_10723,N_10661);
nand U11739 (N_11739,N_10838,N_10616);
or U11740 (N_11740,N_10588,N_10494);
and U11741 (N_11741,N_10945,N_10854);
or U11742 (N_11742,N_10721,N_10731);
nand U11743 (N_11743,N_10989,N_10732);
nor U11744 (N_11744,N_11039,N_10658);
xnor U11745 (N_11745,N_11038,N_10514);
xor U11746 (N_11746,N_10857,N_10824);
xnor U11747 (N_11747,N_10955,N_10555);
xnor U11748 (N_11748,N_10572,N_10675);
nand U11749 (N_11749,N_10621,N_10401);
nand U11750 (N_11750,N_10785,N_10614);
nand U11751 (N_11751,N_11120,N_10461);
nor U11752 (N_11752,N_10514,N_11026);
and U11753 (N_11753,N_10512,N_10570);
nand U11754 (N_11754,N_10436,N_10579);
nor U11755 (N_11755,N_11156,N_10690);
xnor U11756 (N_11756,N_11120,N_10901);
xor U11757 (N_11757,N_10770,N_10881);
xor U11758 (N_11758,N_10625,N_11046);
and U11759 (N_11759,N_10461,N_11170);
and U11760 (N_11760,N_10955,N_10688);
or U11761 (N_11761,N_11000,N_11120);
nand U11762 (N_11762,N_10904,N_10847);
xnor U11763 (N_11763,N_11105,N_11127);
nor U11764 (N_11764,N_11102,N_10484);
nand U11765 (N_11765,N_10896,N_10891);
or U11766 (N_11766,N_10977,N_10610);
xor U11767 (N_11767,N_11038,N_10952);
nand U11768 (N_11768,N_11063,N_10898);
xor U11769 (N_11769,N_10513,N_11085);
nor U11770 (N_11770,N_11027,N_10947);
nor U11771 (N_11771,N_10513,N_11104);
nand U11772 (N_11772,N_10546,N_11174);
nand U11773 (N_11773,N_10620,N_10692);
xor U11774 (N_11774,N_10527,N_10691);
xor U11775 (N_11775,N_10476,N_10843);
nor U11776 (N_11776,N_10624,N_11042);
or U11777 (N_11777,N_10449,N_11145);
nor U11778 (N_11778,N_11079,N_11037);
or U11779 (N_11779,N_10983,N_10560);
and U11780 (N_11780,N_10969,N_10431);
xor U11781 (N_11781,N_11015,N_10702);
nor U11782 (N_11782,N_10763,N_10473);
nor U11783 (N_11783,N_10571,N_10868);
xnor U11784 (N_11784,N_10975,N_10604);
nand U11785 (N_11785,N_10720,N_10834);
or U11786 (N_11786,N_10466,N_10691);
nor U11787 (N_11787,N_10485,N_10685);
xnor U11788 (N_11788,N_10468,N_10530);
or U11789 (N_11789,N_11135,N_10985);
nand U11790 (N_11790,N_11018,N_10615);
xnor U11791 (N_11791,N_11092,N_11132);
and U11792 (N_11792,N_10527,N_10600);
and U11793 (N_11793,N_11051,N_10856);
xnor U11794 (N_11794,N_11048,N_11099);
xnor U11795 (N_11795,N_10568,N_11016);
nand U11796 (N_11796,N_10532,N_10978);
nand U11797 (N_11797,N_10764,N_10952);
nand U11798 (N_11798,N_10734,N_11132);
or U11799 (N_11799,N_10816,N_10712);
or U11800 (N_11800,N_11049,N_10686);
nand U11801 (N_11801,N_10926,N_10832);
and U11802 (N_11802,N_10565,N_11013);
xor U11803 (N_11803,N_10944,N_10416);
nand U11804 (N_11804,N_10426,N_11029);
nand U11805 (N_11805,N_11028,N_11180);
nor U11806 (N_11806,N_11075,N_10897);
or U11807 (N_11807,N_10921,N_10520);
xor U11808 (N_11808,N_10581,N_11005);
nand U11809 (N_11809,N_10523,N_11094);
nor U11810 (N_11810,N_10421,N_10718);
or U11811 (N_11811,N_11104,N_11111);
and U11812 (N_11812,N_11042,N_11013);
xor U11813 (N_11813,N_11043,N_10632);
or U11814 (N_11814,N_11045,N_10696);
xor U11815 (N_11815,N_10612,N_10742);
and U11816 (N_11816,N_11133,N_10551);
nand U11817 (N_11817,N_10556,N_10646);
nor U11818 (N_11818,N_11024,N_10419);
nand U11819 (N_11819,N_11082,N_11098);
nor U11820 (N_11820,N_10599,N_10891);
nand U11821 (N_11821,N_10619,N_10538);
nor U11822 (N_11822,N_11097,N_11081);
and U11823 (N_11823,N_11197,N_10968);
nand U11824 (N_11824,N_10449,N_10580);
nor U11825 (N_11825,N_10980,N_11146);
nand U11826 (N_11826,N_10592,N_10640);
nor U11827 (N_11827,N_11090,N_10832);
nor U11828 (N_11828,N_10431,N_10798);
xor U11829 (N_11829,N_11029,N_10852);
and U11830 (N_11830,N_11063,N_10670);
and U11831 (N_11831,N_11123,N_10872);
xor U11832 (N_11832,N_10898,N_10412);
nand U11833 (N_11833,N_11017,N_10824);
or U11834 (N_11834,N_10743,N_10875);
and U11835 (N_11835,N_10648,N_11081);
and U11836 (N_11836,N_10630,N_10684);
nor U11837 (N_11837,N_11124,N_11021);
nand U11838 (N_11838,N_10554,N_10605);
and U11839 (N_11839,N_10704,N_10885);
and U11840 (N_11840,N_10569,N_10911);
or U11841 (N_11841,N_10804,N_10706);
and U11842 (N_11842,N_10437,N_10742);
nand U11843 (N_11843,N_10609,N_10658);
nor U11844 (N_11844,N_10408,N_11077);
nor U11845 (N_11845,N_10534,N_10935);
nor U11846 (N_11846,N_10949,N_10454);
nor U11847 (N_11847,N_10912,N_11158);
nor U11848 (N_11848,N_11193,N_11122);
xnor U11849 (N_11849,N_10572,N_11161);
nor U11850 (N_11850,N_11085,N_11072);
xnor U11851 (N_11851,N_10679,N_10904);
xor U11852 (N_11852,N_11139,N_11055);
and U11853 (N_11853,N_10625,N_10523);
xnor U11854 (N_11854,N_10934,N_10875);
nor U11855 (N_11855,N_10660,N_10893);
nand U11856 (N_11856,N_10586,N_11176);
nand U11857 (N_11857,N_10489,N_10607);
and U11858 (N_11858,N_10566,N_10880);
nand U11859 (N_11859,N_10721,N_11184);
or U11860 (N_11860,N_11120,N_10713);
nand U11861 (N_11861,N_11142,N_10813);
or U11862 (N_11862,N_10738,N_10943);
and U11863 (N_11863,N_11105,N_10867);
or U11864 (N_11864,N_11084,N_10516);
or U11865 (N_11865,N_10453,N_10917);
xnor U11866 (N_11866,N_10617,N_10418);
nand U11867 (N_11867,N_10504,N_10763);
nand U11868 (N_11868,N_10981,N_10656);
nand U11869 (N_11869,N_10520,N_11104);
nand U11870 (N_11870,N_10656,N_10686);
nand U11871 (N_11871,N_10942,N_11026);
xor U11872 (N_11872,N_11176,N_10577);
xnor U11873 (N_11873,N_10682,N_10824);
nor U11874 (N_11874,N_10816,N_10795);
nor U11875 (N_11875,N_10780,N_10938);
nand U11876 (N_11876,N_10677,N_11008);
nor U11877 (N_11877,N_10946,N_10697);
nor U11878 (N_11878,N_11147,N_10571);
or U11879 (N_11879,N_10882,N_10606);
xor U11880 (N_11880,N_11159,N_11086);
xor U11881 (N_11881,N_10852,N_10463);
nor U11882 (N_11882,N_10772,N_10519);
xnor U11883 (N_11883,N_10497,N_11041);
nor U11884 (N_11884,N_10447,N_10792);
xnor U11885 (N_11885,N_10806,N_11128);
or U11886 (N_11886,N_10421,N_11097);
nor U11887 (N_11887,N_11156,N_11161);
nand U11888 (N_11888,N_10727,N_10543);
and U11889 (N_11889,N_10897,N_10832);
nor U11890 (N_11890,N_11104,N_10760);
and U11891 (N_11891,N_11087,N_10782);
xnor U11892 (N_11892,N_10585,N_11078);
nand U11893 (N_11893,N_10699,N_11115);
nand U11894 (N_11894,N_11012,N_10716);
xor U11895 (N_11895,N_10533,N_10621);
nor U11896 (N_11896,N_10783,N_11173);
nor U11897 (N_11897,N_10698,N_10588);
nand U11898 (N_11898,N_11048,N_11013);
xnor U11899 (N_11899,N_11002,N_11101);
and U11900 (N_11900,N_10750,N_10608);
and U11901 (N_11901,N_10715,N_11170);
nand U11902 (N_11902,N_10409,N_10426);
nand U11903 (N_11903,N_10660,N_10545);
nand U11904 (N_11904,N_10737,N_10882);
xnor U11905 (N_11905,N_10885,N_10741);
nor U11906 (N_11906,N_10512,N_10810);
nor U11907 (N_11907,N_10695,N_10848);
xnor U11908 (N_11908,N_10859,N_10877);
and U11909 (N_11909,N_11174,N_11074);
and U11910 (N_11910,N_10472,N_10698);
xor U11911 (N_11911,N_11196,N_11014);
xor U11912 (N_11912,N_10718,N_11077);
nor U11913 (N_11913,N_11195,N_11164);
nor U11914 (N_11914,N_11166,N_10425);
and U11915 (N_11915,N_10965,N_10807);
or U11916 (N_11916,N_10886,N_11144);
xor U11917 (N_11917,N_10749,N_11032);
and U11918 (N_11918,N_10569,N_11058);
nand U11919 (N_11919,N_11022,N_11065);
nor U11920 (N_11920,N_10446,N_10459);
nor U11921 (N_11921,N_10603,N_10746);
and U11922 (N_11922,N_10448,N_10965);
nor U11923 (N_11923,N_10773,N_10777);
xnor U11924 (N_11924,N_10986,N_10405);
nand U11925 (N_11925,N_10452,N_11060);
or U11926 (N_11926,N_10764,N_10557);
or U11927 (N_11927,N_11122,N_10552);
nor U11928 (N_11928,N_11133,N_11025);
xor U11929 (N_11929,N_10765,N_10770);
nand U11930 (N_11930,N_10657,N_11196);
nor U11931 (N_11931,N_10464,N_10531);
nand U11932 (N_11932,N_11122,N_10662);
and U11933 (N_11933,N_10543,N_10520);
xnor U11934 (N_11934,N_10958,N_10411);
or U11935 (N_11935,N_11117,N_11156);
nor U11936 (N_11936,N_10596,N_11190);
and U11937 (N_11937,N_10961,N_10782);
and U11938 (N_11938,N_10739,N_10899);
xnor U11939 (N_11939,N_11163,N_10592);
or U11940 (N_11940,N_10537,N_10783);
xor U11941 (N_11941,N_10985,N_10547);
nand U11942 (N_11942,N_11069,N_11023);
nand U11943 (N_11943,N_10402,N_10845);
xnor U11944 (N_11944,N_10570,N_11027);
or U11945 (N_11945,N_10965,N_10750);
or U11946 (N_11946,N_10913,N_10968);
and U11947 (N_11947,N_10893,N_10433);
nor U11948 (N_11948,N_11193,N_10935);
or U11949 (N_11949,N_10465,N_11096);
and U11950 (N_11950,N_10761,N_10690);
or U11951 (N_11951,N_11146,N_11171);
nor U11952 (N_11952,N_10776,N_11064);
and U11953 (N_11953,N_11177,N_11075);
nor U11954 (N_11954,N_10602,N_10580);
nand U11955 (N_11955,N_11092,N_10690);
and U11956 (N_11956,N_10782,N_11069);
nand U11957 (N_11957,N_10712,N_10561);
xor U11958 (N_11958,N_10712,N_10493);
and U11959 (N_11959,N_10450,N_10757);
and U11960 (N_11960,N_10850,N_10452);
xor U11961 (N_11961,N_10554,N_10994);
nand U11962 (N_11962,N_10467,N_10592);
or U11963 (N_11963,N_10512,N_11194);
or U11964 (N_11964,N_10898,N_10872);
or U11965 (N_11965,N_10515,N_10973);
nand U11966 (N_11966,N_10835,N_11153);
or U11967 (N_11967,N_10557,N_10969);
and U11968 (N_11968,N_10777,N_10883);
or U11969 (N_11969,N_10533,N_11001);
nor U11970 (N_11970,N_10776,N_10606);
nand U11971 (N_11971,N_10584,N_11007);
nand U11972 (N_11972,N_11094,N_10796);
nor U11973 (N_11973,N_10815,N_10852);
xor U11974 (N_11974,N_10847,N_11100);
and U11975 (N_11975,N_10592,N_10490);
or U11976 (N_11976,N_10998,N_10417);
or U11977 (N_11977,N_10714,N_10798);
or U11978 (N_11978,N_10872,N_10972);
nor U11979 (N_11979,N_10762,N_10794);
nand U11980 (N_11980,N_11027,N_10945);
or U11981 (N_11981,N_11116,N_10873);
and U11982 (N_11982,N_10470,N_10670);
and U11983 (N_11983,N_10976,N_10651);
nor U11984 (N_11984,N_10935,N_11180);
or U11985 (N_11985,N_10998,N_11065);
nand U11986 (N_11986,N_10738,N_10986);
nand U11987 (N_11987,N_10881,N_10487);
xor U11988 (N_11988,N_10760,N_10978);
xnor U11989 (N_11989,N_10718,N_10929);
or U11990 (N_11990,N_10431,N_10855);
or U11991 (N_11991,N_11057,N_10527);
and U11992 (N_11992,N_10754,N_11145);
and U11993 (N_11993,N_11027,N_10499);
nand U11994 (N_11994,N_10459,N_10406);
nor U11995 (N_11995,N_10442,N_11021);
and U11996 (N_11996,N_11198,N_10868);
nor U11997 (N_11997,N_10646,N_10657);
nor U11998 (N_11998,N_11068,N_11179);
xnor U11999 (N_11999,N_11194,N_10651);
nor U12000 (N_12000,N_11308,N_11563);
nand U12001 (N_12001,N_11301,N_11987);
and U12002 (N_12002,N_11786,N_11835);
nand U12003 (N_12003,N_11392,N_11274);
nand U12004 (N_12004,N_11819,N_11204);
nor U12005 (N_12005,N_11750,N_11899);
or U12006 (N_12006,N_11494,N_11638);
and U12007 (N_12007,N_11711,N_11415);
and U12008 (N_12008,N_11995,N_11649);
or U12009 (N_12009,N_11503,N_11782);
nor U12010 (N_12010,N_11557,N_11895);
and U12011 (N_12011,N_11860,N_11481);
nor U12012 (N_12012,N_11227,N_11810);
and U12013 (N_12013,N_11996,N_11844);
xnor U12014 (N_12014,N_11695,N_11861);
nor U12015 (N_12015,N_11656,N_11634);
nor U12016 (N_12016,N_11215,N_11236);
xnor U12017 (N_12017,N_11344,N_11476);
and U12018 (N_12018,N_11769,N_11959);
and U12019 (N_12019,N_11334,N_11555);
nand U12020 (N_12020,N_11228,N_11752);
nand U12021 (N_12021,N_11836,N_11238);
or U12022 (N_12022,N_11556,N_11382);
or U12023 (N_12023,N_11672,N_11580);
nand U12024 (N_12024,N_11551,N_11424);
nand U12025 (N_12025,N_11902,N_11277);
or U12026 (N_12026,N_11840,N_11407);
and U12027 (N_12027,N_11571,N_11375);
nand U12028 (N_12028,N_11327,N_11218);
nand U12029 (N_12029,N_11621,N_11882);
and U12030 (N_12030,N_11522,N_11982);
and U12031 (N_12031,N_11604,N_11578);
and U12032 (N_12032,N_11312,N_11340);
nand U12033 (N_12033,N_11395,N_11814);
nand U12034 (N_12034,N_11406,N_11332);
xor U12035 (N_12035,N_11449,N_11792);
and U12036 (N_12036,N_11279,N_11720);
nand U12037 (N_12037,N_11520,N_11355);
nor U12038 (N_12038,N_11842,N_11582);
and U12039 (N_12039,N_11213,N_11953);
nand U12040 (N_12040,N_11714,N_11525);
nor U12041 (N_12041,N_11960,N_11774);
xor U12042 (N_12042,N_11343,N_11856);
and U12043 (N_12043,N_11313,N_11824);
nor U12044 (N_12044,N_11947,N_11806);
and U12045 (N_12045,N_11888,N_11922);
nand U12046 (N_12046,N_11230,N_11793);
nand U12047 (N_12047,N_11261,N_11956);
nand U12048 (N_12048,N_11402,N_11874);
nand U12049 (N_12049,N_11877,N_11225);
or U12050 (N_12050,N_11660,N_11643);
nand U12051 (N_12051,N_11504,N_11541);
nor U12052 (N_12052,N_11862,N_11791);
and U12053 (N_12053,N_11853,N_11387);
xnor U12054 (N_12054,N_11579,N_11433);
nor U12055 (N_12055,N_11299,N_11916);
nor U12056 (N_12056,N_11281,N_11409);
or U12057 (N_12057,N_11278,N_11463);
xnor U12058 (N_12058,N_11794,N_11413);
xnor U12059 (N_12059,N_11813,N_11434);
nand U12060 (N_12060,N_11822,N_11348);
nand U12061 (N_12061,N_11891,N_11529);
nand U12062 (N_12062,N_11289,N_11918);
or U12063 (N_12063,N_11833,N_11359);
nand U12064 (N_12064,N_11200,N_11843);
or U12065 (N_12065,N_11364,N_11753);
nand U12066 (N_12066,N_11287,N_11746);
xor U12067 (N_12067,N_11469,N_11455);
xnor U12068 (N_12068,N_11785,N_11724);
or U12069 (N_12069,N_11485,N_11229);
or U12070 (N_12070,N_11589,N_11298);
nor U12071 (N_12071,N_11478,N_11954);
xnor U12072 (N_12072,N_11905,N_11770);
and U12073 (N_12073,N_11762,N_11544);
xnor U12074 (N_12074,N_11797,N_11626);
xor U12075 (N_12075,N_11821,N_11901);
nor U12076 (N_12076,N_11913,N_11764);
nand U12077 (N_12077,N_11264,N_11548);
xnor U12078 (N_12078,N_11667,N_11633);
or U12079 (N_12079,N_11351,N_11925);
nand U12080 (N_12080,N_11690,N_11595);
and U12081 (N_12081,N_11659,N_11430);
or U12082 (N_12082,N_11788,N_11222);
or U12083 (N_12083,N_11631,N_11868);
nand U12084 (N_12084,N_11800,N_11262);
or U12085 (N_12085,N_11491,N_11795);
xnor U12086 (N_12086,N_11374,N_11965);
xor U12087 (N_12087,N_11350,N_11319);
nor U12088 (N_12088,N_11999,N_11592);
nor U12089 (N_12089,N_11698,N_11475);
or U12090 (N_12090,N_11484,N_11779);
nand U12091 (N_12091,N_11207,N_11851);
nand U12092 (N_12092,N_11725,N_11524);
nand U12093 (N_12093,N_11887,N_11684);
or U12094 (N_12094,N_11256,N_11624);
and U12095 (N_12095,N_11271,N_11776);
and U12096 (N_12096,N_11285,N_11342);
and U12097 (N_12097,N_11546,N_11910);
and U12098 (N_12098,N_11609,N_11325);
xor U12099 (N_12099,N_11818,N_11234);
xor U12100 (N_12100,N_11966,N_11629);
or U12101 (N_12101,N_11586,N_11329);
nand U12102 (N_12102,N_11828,N_11907);
and U12103 (N_12103,N_11331,N_11553);
nand U12104 (N_12104,N_11976,N_11534);
or U12105 (N_12105,N_11937,N_11687);
xnor U12106 (N_12106,N_11993,N_11400);
nand U12107 (N_12107,N_11948,N_11863);
nand U12108 (N_12108,N_11991,N_11318);
and U12109 (N_12109,N_11543,N_11326);
nor U12110 (N_12110,N_11671,N_11642);
xor U12111 (N_12111,N_11908,N_11854);
and U12112 (N_12112,N_11946,N_11566);
xor U12113 (N_12113,N_11981,N_11865);
and U12114 (N_12114,N_11816,N_11619);
xnor U12115 (N_12115,N_11284,N_11871);
or U12116 (N_12116,N_11425,N_11789);
xor U12117 (N_12117,N_11527,N_11533);
and U12118 (N_12118,N_11630,N_11602);
nor U12119 (N_12119,N_11386,N_11783);
nand U12120 (N_12120,N_11558,N_11657);
nor U12121 (N_12121,N_11886,N_11303);
nor U12122 (N_12122,N_11474,N_11502);
nand U12123 (N_12123,N_11323,N_11712);
nor U12124 (N_12124,N_11896,N_11738);
nor U12125 (N_12125,N_11992,N_11510);
xor U12126 (N_12126,N_11740,N_11385);
nand U12127 (N_12127,N_11670,N_11858);
and U12128 (N_12128,N_11569,N_11461);
and U12129 (N_12129,N_11678,N_11757);
and U12130 (N_12130,N_11482,N_11646);
or U12131 (N_12131,N_11676,N_11466);
and U12132 (N_12132,N_11926,N_11243);
nor U12133 (N_12133,N_11934,N_11496);
nand U12134 (N_12134,N_11390,N_11611);
nor U12135 (N_12135,N_11654,N_11499);
xnor U12136 (N_12136,N_11439,N_11700);
or U12137 (N_12137,N_11202,N_11932);
nand U12138 (N_12138,N_11384,N_11517);
nand U12139 (N_12139,N_11250,N_11453);
xor U12140 (N_12140,N_11610,N_11539);
nor U12141 (N_12141,N_11322,N_11706);
nand U12142 (N_12142,N_11435,N_11226);
nor U12143 (N_12143,N_11574,N_11962);
nand U12144 (N_12144,N_11246,N_11214);
nor U12145 (N_12145,N_11928,N_11912);
nor U12146 (N_12146,N_11980,N_11817);
and U12147 (N_12147,N_11870,N_11295);
xnor U12148 (N_12148,N_11235,N_11837);
xor U12149 (N_12149,N_11457,N_11975);
and U12150 (N_12150,N_11664,N_11761);
nor U12151 (N_12151,N_11587,N_11935);
nand U12152 (N_12152,N_11944,N_11538);
nand U12153 (N_12153,N_11767,N_11661);
nand U12154 (N_12154,N_11969,N_11411);
nor U12155 (N_12155,N_11603,N_11315);
or U12156 (N_12156,N_11362,N_11458);
or U12157 (N_12157,N_11943,N_11560);
xnor U12158 (N_12158,N_11696,N_11669);
nand U12159 (N_12159,N_11704,N_11617);
xor U12160 (N_12160,N_11366,N_11903);
and U12161 (N_12161,N_11988,N_11428);
or U12162 (N_12162,N_11713,N_11967);
xor U12163 (N_12163,N_11697,N_11490);
nand U12164 (N_12164,N_11426,N_11663);
nand U12165 (N_12165,N_11998,N_11924);
nand U12166 (N_12166,N_11211,N_11722);
or U12167 (N_12167,N_11662,N_11984);
and U12168 (N_12168,N_11939,N_11347);
and U12169 (N_12169,N_11547,N_11247);
or U12170 (N_12170,N_11938,N_11952);
and U12171 (N_12171,N_11884,N_11258);
nor U12172 (N_12172,N_11760,N_11607);
xor U12173 (N_12173,N_11321,N_11694);
nand U12174 (N_12174,N_11268,N_11869);
or U12175 (N_12175,N_11275,N_11872);
xnor U12176 (N_12176,N_11518,N_11705);
or U12177 (N_12177,N_11577,N_11773);
nand U12178 (N_12178,N_11388,N_11812);
and U12179 (N_12179,N_11983,N_11508);
nand U12180 (N_12180,N_11930,N_11365);
nor U12181 (N_12181,N_11997,N_11823);
and U12182 (N_12182,N_11894,N_11873);
or U12183 (N_12183,N_11808,N_11622);
or U12184 (N_12184,N_11216,N_11221);
xnor U12185 (N_12185,N_11208,N_11727);
and U12186 (N_12186,N_11237,N_11639);
xnor U12187 (N_12187,N_11825,N_11650);
or U12188 (N_12188,N_11304,N_11625);
and U12189 (N_12189,N_11371,N_11742);
and U12190 (N_12190,N_11989,N_11807);
nand U12191 (N_12191,N_11272,N_11632);
or U12192 (N_12192,N_11479,N_11708);
nor U12193 (N_12193,N_11772,N_11446);
or U12194 (N_12194,N_11809,N_11205);
nor U12195 (N_12195,N_11283,N_11790);
or U12196 (N_12196,N_11487,N_11964);
nor U12197 (N_12197,N_11605,N_11691);
nor U12198 (N_12198,N_11233,N_11701);
nand U12199 (N_12199,N_11735,N_11920);
xnor U12200 (N_12200,N_11263,N_11591);
and U12201 (N_12201,N_11741,N_11929);
nor U12202 (N_12202,N_11505,N_11909);
xnor U12203 (N_12203,N_11743,N_11521);
nand U12204 (N_12204,N_11796,N_11550);
or U12205 (N_12205,N_11500,N_11468);
or U12206 (N_12206,N_11758,N_11565);
and U12207 (N_12207,N_11804,N_11889);
nand U12208 (N_12208,N_11472,N_11368);
and U12209 (N_12209,N_11291,N_11432);
nand U12210 (N_12210,N_11867,N_11376);
nor U12211 (N_12211,N_11972,N_11542);
and U12212 (N_12212,N_11979,N_11330);
or U12213 (N_12213,N_11341,N_11847);
and U12214 (N_12214,N_11568,N_11217);
nand U12215 (N_12215,N_11459,N_11644);
or U12216 (N_12216,N_11801,N_11751);
or U12217 (N_12217,N_11438,N_11512);
xor U12218 (N_12218,N_11201,N_11219);
nand U12219 (N_12219,N_11253,N_11974);
nand U12220 (N_12220,N_11464,N_11251);
xnor U12221 (N_12221,N_11931,N_11399);
nor U12222 (N_12222,N_11549,N_11561);
and U12223 (N_12223,N_11683,N_11336);
or U12224 (N_12224,N_11356,N_11585);
or U12225 (N_12225,N_11766,N_11440);
nand U12226 (N_12226,N_11370,N_11486);
xor U12227 (N_12227,N_11483,N_11443);
and U12228 (N_12228,N_11682,N_11637);
nor U12229 (N_12229,N_11452,N_11802);
and U12230 (N_12230,N_11248,N_11456);
xor U12231 (N_12231,N_11688,N_11827);
or U12232 (N_12232,N_11497,N_11745);
or U12233 (N_12233,N_11501,N_11460);
nand U12234 (N_12234,N_11570,N_11620);
xnor U12235 (N_12235,N_11404,N_11875);
nand U12236 (N_12236,N_11396,N_11748);
and U12237 (N_12237,N_11436,N_11380);
xor U12238 (N_12238,N_11519,N_11919);
nand U12239 (N_12239,N_11509,N_11883);
or U12240 (N_12240,N_11480,N_11955);
or U12241 (N_12241,N_11950,N_11848);
or U12242 (N_12242,N_11220,N_11707);
and U12243 (N_12243,N_11307,N_11613);
nand U12244 (N_12244,N_11677,N_11737);
nand U12245 (N_12245,N_11957,N_11257);
nand U12246 (N_12246,N_11328,N_11703);
or U12247 (N_12247,N_11680,N_11598);
nor U12248 (N_12248,N_11333,N_11266);
or U12249 (N_12249,N_11635,N_11876);
or U12250 (N_12250,N_11345,N_11850);
or U12251 (N_12251,N_11986,N_11838);
or U12252 (N_12252,N_11968,N_11276);
xnor U12253 (N_12253,N_11805,N_11798);
and U12254 (N_12254,N_11379,N_11921);
and U12255 (N_12255,N_11803,N_11405);
xnor U12256 (N_12256,N_11885,N_11606);
nand U12257 (N_12257,N_11906,N_11628);
or U12258 (N_12258,N_11584,N_11576);
xnor U12259 (N_12259,N_11590,N_11410);
or U12260 (N_12260,N_11515,N_11488);
nand U12261 (N_12261,N_11447,N_11210);
xnor U12262 (N_12262,N_11337,N_11958);
nor U12263 (N_12263,N_11841,N_11293);
nand U12264 (N_12264,N_11780,N_11363);
and U12265 (N_12265,N_11422,N_11242);
and U12266 (N_12266,N_11652,N_11721);
xor U12267 (N_12267,N_11573,N_11693);
nor U12268 (N_12268,N_11575,N_11254);
or U12269 (N_12269,N_11911,N_11777);
nand U12270 (N_12270,N_11310,N_11961);
and U12271 (N_12271,N_11239,N_11734);
nand U12272 (N_12272,N_11526,N_11597);
nor U12273 (N_12273,N_11224,N_11730);
nand U12274 (N_12274,N_11465,N_11942);
or U12275 (N_12275,N_11477,N_11267);
nor U12276 (N_12276,N_11349,N_11338);
nand U12277 (N_12277,N_11346,N_11489);
and U12278 (N_12278,N_11645,N_11702);
xor U12279 (N_12279,N_11615,N_11747);
or U12280 (N_12280,N_11493,N_11692);
xnor U12281 (N_12281,N_11799,N_11361);
or U12282 (N_12282,N_11623,N_11401);
or U12283 (N_12283,N_11397,N_11674);
nand U12284 (N_12284,N_11973,N_11897);
nand U12285 (N_12285,N_11270,N_11431);
xor U12286 (N_12286,N_11528,N_11269);
nor U12287 (N_12287,N_11616,N_11296);
nor U12288 (N_12288,N_11900,N_11545);
xor U12289 (N_12289,N_11710,N_11904);
nand U12290 (N_12290,N_11427,N_11594);
and U12291 (N_12291,N_11437,N_11826);
nand U12292 (N_12292,N_11249,N_11709);
xor U12293 (N_12293,N_11588,N_11492);
nand U12294 (N_12294,N_11451,N_11360);
and U12295 (N_12295,N_11936,N_11655);
and U12296 (N_12296,N_11245,N_11914);
and U12297 (N_12297,N_11300,N_11627);
nand U12298 (N_12298,N_11839,N_11846);
xor U12299 (N_12299,N_11414,N_11951);
nor U12300 (N_12300,N_11880,N_11255);
or U12301 (N_12301,N_11732,N_11286);
nor U12302 (N_12302,N_11915,N_11442);
and U12303 (N_12303,N_11971,N_11755);
or U12304 (N_12304,N_11716,N_11845);
nor U12305 (N_12305,N_11679,N_11423);
nand U12306 (N_12306,N_11288,N_11666);
or U12307 (N_12307,N_11990,N_11892);
xnor U12308 (N_12308,N_11394,N_11316);
or U12309 (N_12309,N_11731,N_11581);
nor U12310 (N_12310,N_11290,N_11879);
nor U12311 (N_12311,N_11324,N_11530);
or U12312 (N_12312,N_11759,N_11358);
nand U12313 (N_12313,N_11335,N_11567);
xor U12314 (N_12314,N_11294,N_11665);
xor U12315 (N_12315,N_11945,N_11749);
or U12316 (N_12316,N_11830,N_11686);
nor U12317 (N_12317,N_11717,N_11306);
xor U12318 (N_12318,N_11618,N_11554);
nor U12319 (N_12319,N_11855,N_11421);
nand U12320 (N_12320,N_11282,N_11507);
or U12321 (N_12321,N_11206,N_11377);
or U12322 (N_12322,N_11600,N_11240);
nand U12323 (N_12323,N_11612,N_11923);
xnor U12324 (N_12324,N_11829,N_11864);
nor U12325 (N_12325,N_11369,N_11495);
xor U12326 (N_12326,N_11537,N_11754);
nor U12327 (N_12327,N_11259,N_11866);
nor U12328 (N_12328,N_11244,N_11601);
and U12329 (N_12329,N_11815,N_11699);
nor U12330 (N_12330,N_11552,N_11647);
nand U12331 (N_12331,N_11391,N_11689);
nand U12332 (N_12332,N_11881,N_11531);
and U12333 (N_12333,N_11949,N_11297);
or U12334 (N_12334,N_11393,N_11352);
and U12335 (N_12335,N_11583,N_11292);
nand U12336 (N_12336,N_11260,N_11473);
and U12337 (N_12337,N_11784,N_11719);
nand U12338 (N_12338,N_11765,N_11941);
or U12339 (N_12339,N_11540,N_11454);
and U12340 (N_12340,N_11450,N_11614);
or U12341 (N_12341,N_11978,N_11763);
and U12342 (N_12342,N_11498,N_11559);
or U12343 (N_12343,N_11317,N_11859);
xnor U12344 (N_12344,N_11771,N_11513);
nand U12345 (N_12345,N_11744,N_11985);
or U12346 (N_12346,N_11636,N_11232);
xor U12347 (N_12347,N_11523,N_11265);
nand U12348 (N_12348,N_11564,N_11212);
nor U12349 (N_12349,N_11940,N_11408);
and U12350 (N_12350,N_11852,N_11878);
xnor U12351 (N_12351,N_11445,N_11917);
or U12352 (N_12352,N_11715,N_11203);
nor U12353 (N_12353,N_11471,N_11963);
nand U12354 (N_12354,N_11653,N_11311);
or U12355 (N_12355,N_11516,N_11536);
nor U12356 (N_12356,N_11448,N_11231);
nor U12357 (N_12357,N_11733,N_11280);
or U12358 (N_12358,N_11718,N_11994);
and U12359 (N_12359,N_11357,N_11470);
nand U12360 (N_12360,N_11412,N_11898);
nand U12361 (N_12361,N_11681,N_11223);
nand U12362 (N_12362,N_11302,N_11608);
nor U12363 (N_12363,N_11927,N_11648);
nor U12364 (N_12364,N_11933,N_11511);
nor U12365 (N_12365,N_11768,N_11685);
xnor U12366 (N_12366,N_11756,N_11441);
xor U12367 (N_12367,N_11389,N_11977);
nand U12368 (N_12368,N_11353,N_11572);
xnor U12369 (N_12369,N_11252,N_11314);
nand U12370 (N_12370,N_11673,N_11831);
nor U12371 (N_12371,N_11420,N_11398);
nand U12372 (N_12372,N_11890,N_11354);
and U12373 (N_12373,N_11811,N_11593);
and U12374 (N_12374,N_11429,N_11419);
xnor U12375 (N_12375,N_11367,N_11383);
xor U12376 (N_12376,N_11739,N_11736);
and U12377 (N_12377,N_11599,N_11775);
nor U12378 (N_12378,N_11462,N_11658);
nor U12379 (N_12379,N_11467,N_11535);
and U12380 (N_12380,N_11834,N_11832);
nor U12381 (N_12381,N_11820,N_11444);
and U12382 (N_12382,N_11640,N_11506);
nand U12383 (N_12383,N_11320,N_11416);
nand U12384 (N_12384,N_11723,N_11778);
xnor U12385 (N_12385,N_11372,N_11668);
and U12386 (N_12386,N_11849,N_11596);
xor U12387 (N_12387,N_11728,N_11675);
xnor U12388 (N_12388,N_11273,N_11339);
nor U12389 (N_12389,N_11417,N_11726);
or U12390 (N_12390,N_11857,N_11241);
and U12391 (N_12391,N_11209,N_11729);
xnor U12392 (N_12392,N_11309,N_11781);
nor U12393 (N_12393,N_11514,N_11651);
nor U12394 (N_12394,N_11378,N_11403);
xor U12395 (N_12395,N_11787,N_11418);
and U12396 (N_12396,N_11373,N_11305);
xnor U12397 (N_12397,N_11893,N_11641);
nor U12398 (N_12398,N_11970,N_11562);
nor U12399 (N_12399,N_11381,N_11532);
xor U12400 (N_12400,N_11574,N_11992);
and U12401 (N_12401,N_11749,N_11708);
xnor U12402 (N_12402,N_11918,N_11361);
and U12403 (N_12403,N_11300,N_11383);
or U12404 (N_12404,N_11665,N_11530);
or U12405 (N_12405,N_11487,N_11745);
xor U12406 (N_12406,N_11242,N_11445);
and U12407 (N_12407,N_11251,N_11871);
or U12408 (N_12408,N_11576,N_11402);
nand U12409 (N_12409,N_11573,N_11928);
and U12410 (N_12410,N_11524,N_11257);
xnor U12411 (N_12411,N_11605,N_11810);
xor U12412 (N_12412,N_11595,N_11373);
or U12413 (N_12413,N_11741,N_11849);
xor U12414 (N_12414,N_11954,N_11494);
and U12415 (N_12415,N_11278,N_11957);
and U12416 (N_12416,N_11505,N_11478);
nor U12417 (N_12417,N_11503,N_11824);
and U12418 (N_12418,N_11778,N_11833);
xor U12419 (N_12419,N_11381,N_11446);
nand U12420 (N_12420,N_11495,N_11819);
nand U12421 (N_12421,N_11865,N_11994);
nor U12422 (N_12422,N_11359,N_11985);
and U12423 (N_12423,N_11814,N_11654);
xor U12424 (N_12424,N_11726,N_11551);
or U12425 (N_12425,N_11243,N_11549);
nand U12426 (N_12426,N_11630,N_11939);
xnor U12427 (N_12427,N_11939,N_11291);
and U12428 (N_12428,N_11652,N_11283);
nor U12429 (N_12429,N_11518,N_11429);
and U12430 (N_12430,N_11595,N_11483);
or U12431 (N_12431,N_11481,N_11850);
nor U12432 (N_12432,N_11568,N_11812);
nand U12433 (N_12433,N_11260,N_11805);
nand U12434 (N_12434,N_11875,N_11509);
or U12435 (N_12435,N_11390,N_11730);
nor U12436 (N_12436,N_11332,N_11903);
xor U12437 (N_12437,N_11437,N_11404);
and U12438 (N_12438,N_11298,N_11318);
nor U12439 (N_12439,N_11825,N_11894);
and U12440 (N_12440,N_11281,N_11373);
xor U12441 (N_12441,N_11936,N_11622);
or U12442 (N_12442,N_11909,N_11627);
and U12443 (N_12443,N_11857,N_11928);
nand U12444 (N_12444,N_11303,N_11908);
nand U12445 (N_12445,N_11669,N_11377);
nand U12446 (N_12446,N_11706,N_11386);
xor U12447 (N_12447,N_11207,N_11831);
and U12448 (N_12448,N_11473,N_11677);
and U12449 (N_12449,N_11547,N_11644);
and U12450 (N_12450,N_11428,N_11764);
or U12451 (N_12451,N_11206,N_11572);
and U12452 (N_12452,N_11808,N_11897);
and U12453 (N_12453,N_11329,N_11822);
nand U12454 (N_12454,N_11679,N_11233);
nand U12455 (N_12455,N_11357,N_11992);
or U12456 (N_12456,N_11762,N_11769);
and U12457 (N_12457,N_11315,N_11235);
and U12458 (N_12458,N_11550,N_11854);
or U12459 (N_12459,N_11567,N_11472);
or U12460 (N_12460,N_11662,N_11947);
and U12461 (N_12461,N_11707,N_11473);
and U12462 (N_12462,N_11529,N_11911);
nand U12463 (N_12463,N_11856,N_11860);
and U12464 (N_12464,N_11378,N_11469);
nand U12465 (N_12465,N_11711,N_11805);
nor U12466 (N_12466,N_11705,N_11503);
nor U12467 (N_12467,N_11363,N_11345);
xor U12468 (N_12468,N_11335,N_11858);
nand U12469 (N_12469,N_11524,N_11465);
nand U12470 (N_12470,N_11860,N_11333);
and U12471 (N_12471,N_11635,N_11294);
xor U12472 (N_12472,N_11497,N_11556);
xor U12473 (N_12473,N_11881,N_11518);
and U12474 (N_12474,N_11559,N_11406);
and U12475 (N_12475,N_11610,N_11967);
xor U12476 (N_12476,N_11777,N_11695);
and U12477 (N_12477,N_11366,N_11777);
and U12478 (N_12478,N_11798,N_11231);
and U12479 (N_12479,N_11905,N_11516);
nor U12480 (N_12480,N_11288,N_11952);
nor U12481 (N_12481,N_11936,N_11495);
nor U12482 (N_12482,N_11887,N_11768);
or U12483 (N_12483,N_11461,N_11206);
nand U12484 (N_12484,N_11833,N_11904);
xnor U12485 (N_12485,N_11556,N_11491);
or U12486 (N_12486,N_11933,N_11367);
nor U12487 (N_12487,N_11483,N_11958);
xnor U12488 (N_12488,N_11527,N_11768);
xor U12489 (N_12489,N_11791,N_11937);
nand U12490 (N_12490,N_11756,N_11641);
nand U12491 (N_12491,N_11380,N_11705);
xnor U12492 (N_12492,N_11309,N_11507);
xnor U12493 (N_12493,N_11676,N_11888);
xor U12494 (N_12494,N_11232,N_11573);
nor U12495 (N_12495,N_11814,N_11486);
nor U12496 (N_12496,N_11261,N_11685);
and U12497 (N_12497,N_11780,N_11830);
nand U12498 (N_12498,N_11431,N_11522);
xor U12499 (N_12499,N_11834,N_11652);
and U12500 (N_12500,N_11995,N_11998);
and U12501 (N_12501,N_11244,N_11801);
and U12502 (N_12502,N_11479,N_11295);
nand U12503 (N_12503,N_11918,N_11230);
or U12504 (N_12504,N_11787,N_11470);
and U12505 (N_12505,N_11361,N_11521);
nor U12506 (N_12506,N_11535,N_11338);
or U12507 (N_12507,N_11255,N_11260);
and U12508 (N_12508,N_11287,N_11843);
and U12509 (N_12509,N_11291,N_11628);
xor U12510 (N_12510,N_11554,N_11267);
nand U12511 (N_12511,N_11205,N_11669);
xnor U12512 (N_12512,N_11337,N_11296);
nand U12513 (N_12513,N_11702,N_11928);
and U12514 (N_12514,N_11917,N_11744);
or U12515 (N_12515,N_11814,N_11729);
or U12516 (N_12516,N_11231,N_11879);
and U12517 (N_12517,N_11824,N_11361);
and U12518 (N_12518,N_11428,N_11978);
nor U12519 (N_12519,N_11966,N_11790);
and U12520 (N_12520,N_11256,N_11815);
and U12521 (N_12521,N_11710,N_11464);
xnor U12522 (N_12522,N_11830,N_11201);
or U12523 (N_12523,N_11687,N_11524);
nand U12524 (N_12524,N_11709,N_11226);
or U12525 (N_12525,N_11691,N_11588);
nor U12526 (N_12526,N_11283,N_11660);
or U12527 (N_12527,N_11500,N_11473);
nand U12528 (N_12528,N_11287,N_11517);
and U12529 (N_12529,N_11235,N_11899);
or U12530 (N_12530,N_11524,N_11771);
and U12531 (N_12531,N_11829,N_11531);
nand U12532 (N_12532,N_11846,N_11919);
nor U12533 (N_12533,N_11304,N_11880);
nor U12534 (N_12534,N_11595,N_11963);
and U12535 (N_12535,N_11498,N_11810);
nor U12536 (N_12536,N_11812,N_11370);
nor U12537 (N_12537,N_11359,N_11802);
nor U12538 (N_12538,N_11262,N_11934);
nor U12539 (N_12539,N_11246,N_11430);
or U12540 (N_12540,N_11834,N_11461);
or U12541 (N_12541,N_11484,N_11826);
nor U12542 (N_12542,N_11954,N_11501);
nand U12543 (N_12543,N_11618,N_11792);
or U12544 (N_12544,N_11399,N_11917);
nor U12545 (N_12545,N_11366,N_11681);
or U12546 (N_12546,N_11952,N_11704);
or U12547 (N_12547,N_11254,N_11256);
nor U12548 (N_12548,N_11676,N_11863);
or U12549 (N_12549,N_11697,N_11618);
and U12550 (N_12550,N_11805,N_11958);
nand U12551 (N_12551,N_11803,N_11399);
xor U12552 (N_12552,N_11204,N_11288);
xor U12553 (N_12553,N_11676,N_11501);
nor U12554 (N_12554,N_11275,N_11508);
and U12555 (N_12555,N_11530,N_11202);
and U12556 (N_12556,N_11412,N_11978);
xor U12557 (N_12557,N_11340,N_11678);
nand U12558 (N_12558,N_11891,N_11480);
and U12559 (N_12559,N_11654,N_11360);
nor U12560 (N_12560,N_11877,N_11924);
and U12561 (N_12561,N_11488,N_11544);
and U12562 (N_12562,N_11977,N_11412);
xnor U12563 (N_12563,N_11653,N_11930);
nor U12564 (N_12564,N_11335,N_11298);
xnor U12565 (N_12565,N_11302,N_11224);
or U12566 (N_12566,N_11308,N_11303);
and U12567 (N_12567,N_11848,N_11558);
nor U12568 (N_12568,N_11432,N_11961);
nor U12569 (N_12569,N_11283,N_11479);
nor U12570 (N_12570,N_11675,N_11381);
nor U12571 (N_12571,N_11349,N_11708);
nor U12572 (N_12572,N_11675,N_11523);
xnor U12573 (N_12573,N_11207,N_11917);
nand U12574 (N_12574,N_11941,N_11851);
and U12575 (N_12575,N_11531,N_11265);
xor U12576 (N_12576,N_11582,N_11488);
nor U12577 (N_12577,N_11976,N_11871);
or U12578 (N_12578,N_11246,N_11350);
or U12579 (N_12579,N_11388,N_11604);
and U12580 (N_12580,N_11834,N_11668);
or U12581 (N_12581,N_11996,N_11372);
nand U12582 (N_12582,N_11634,N_11642);
nand U12583 (N_12583,N_11836,N_11283);
nor U12584 (N_12584,N_11720,N_11966);
nand U12585 (N_12585,N_11285,N_11210);
or U12586 (N_12586,N_11601,N_11228);
xor U12587 (N_12587,N_11265,N_11732);
and U12588 (N_12588,N_11601,N_11388);
xor U12589 (N_12589,N_11287,N_11473);
or U12590 (N_12590,N_11295,N_11377);
nand U12591 (N_12591,N_11720,N_11960);
nor U12592 (N_12592,N_11599,N_11959);
or U12593 (N_12593,N_11540,N_11532);
and U12594 (N_12594,N_11348,N_11307);
nand U12595 (N_12595,N_11203,N_11332);
or U12596 (N_12596,N_11600,N_11301);
nor U12597 (N_12597,N_11324,N_11521);
xor U12598 (N_12598,N_11430,N_11844);
nor U12599 (N_12599,N_11481,N_11567);
nand U12600 (N_12600,N_11496,N_11544);
nand U12601 (N_12601,N_11414,N_11459);
xnor U12602 (N_12602,N_11396,N_11496);
nor U12603 (N_12603,N_11371,N_11313);
or U12604 (N_12604,N_11397,N_11894);
nand U12605 (N_12605,N_11411,N_11857);
and U12606 (N_12606,N_11644,N_11613);
xnor U12607 (N_12607,N_11325,N_11508);
and U12608 (N_12608,N_11345,N_11842);
nor U12609 (N_12609,N_11802,N_11467);
or U12610 (N_12610,N_11649,N_11484);
nand U12611 (N_12611,N_11490,N_11694);
xor U12612 (N_12612,N_11927,N_11679);
nand U12613 (N_12613,N_11634,N_11888);
nor U12614 (N_12614,N_11789,N_11844);
xnor U12615 (N_12615,N_11761,N_11505);
xor U12616 (N_12616,N_11207,N_11304);
xnor U12617 (N_12617,N_11438,N_11963);
nand U12618 (N_12618,N_11612,N_11958);
or U12619 (N_12619,N_11269,N_11275);
nand U12620 (N_12620,N_11955,N_11950);
nand U12621 (N_12621,N_11527,N_11950);
xor U12622 (N_12622,N_11816,N_11908);
or U12623 (N_12623,N_11375,N_11801);
nand U12624 (N_12624,N_11304,N_11680);
nor U12625 (N_12625,N_11641,N_11299);
nor U12626 (N_12626,N_11641,N_11940);
and U12627 (N_12627,N_11456,N_11724);
xor U12628 (N_12628,N_11321,N_11414);
and U12629 (N_12629,N_11914,N_11671);
nor U12630 (N_12630,N_11807,N_11749);
nand U12631 (N_12631,N_11839,N_11553);
and U12632 (N_12632,N_11836,N_11447);
or U12633 (N_12633,N_11981,N_11368);
or U12634 (N_12634,N_11999,N_11831);
nand U12635 (N_12635,N_11830,N_11687);
nand U12636 (N_12636,N_11403,N_11687);
or U12637 (N_12637,N_11307,N_11825);
nor U12638 (N_12638,N_11768,N_11980);
and U12639 (N_12639,N_11468,N_11872);
nand U12640 (N_12640,N_11420,N_11319);
nand U12641 (N_12641,N_11768,N_11886);
xor U12642 (N_12642,N_11871,N_11985);
and U12643 (N_12643,N_11398,N_11278);
xnor U12644 (N_12644,N_11896,N_11353);
and U12645 (N_12645,N_11520,N_11719);
xnor U12646 (N_12646,N_11853,N_11818);
xnor U12647 (N_12647,N_11567,N_11362);
nor U12648 (N_12648,N_11707,N_11891);
xor U12649 (N_12649,N_11986,N_11417);
nor U12650 (N_12650,N_11673,N_11468);
xor U12651 (N_12651,N_11298,N_11901);
xor U12652 (N_12652,N_11835,N_11951);
nand U12653 (N_12653,N_11273,N_11316);
nand U12654 (N_12654,N_11255,N_11757);
and U12655 (N_12655,N_11435,N_11912);
xor U12656 (N_12656,N_11680,N_11766);
xnor U12657 (N_12657,N_11581,N_11989);
nand U12658 (N_12658,N_11434,N_11937);
xor U12659 (N_12659,N_11890,N_11987);
xor U12660 (N_12660,N_11882,N_11449);
nand U12661 (N_12661,N_11999,N_11236);
and U12662 (N_12662,N_11734,N_11750);
nor U12663 (N_12663,N_11251,N_11795);
nor U12664 (N_12664,N_11540,N_11836);
or U12665 (N_12665,N_11295,N_11437);
or U12666 (N_12666,N_11605,N_11971);
nor U12667 (N_12667,N_11339,N_11357);
nand U12668 (N_12668,N_11565,N_11290);
nand U12669 (N_12669,N_11985,N_11573);
xnor U12670 (N_12670,N_11507,N_11925);
nor U12671 (N_12671,N_11821,N_11764);
nand U12672 (N_12672,N_11772,N_11950);
nand U12673 (N_12673,N_11312,N_11968);
and U12674 (N_12674,N_11576,N_11776);
nor U12675 (N_12675,N_11489,N_11341);
and U12676 (N_12676,N_11552,N_11343);
nor U12677 (N_12677,N_11259,N_11411);
nor U12678 (N_12678,N_11916,N_11868);
xor U12679 (N_12679,N_11444,N_11216);
nand U12680 (N_12680,N_11572,N_11747);
or U12681 (N_12681,N_11379,N_11284);
or U12682 (N_12682,N_11545,N_11940);
or U12683 (N_12683,N_11840,N_11945);
xnor U12684 (N_12684,N_11787,N_11926);
nand U12685 (N_12685,N_11353,N_11311);
nand U12686 (N_12686,N_11603,N_11361);
or U12687 (N_12687,N_11467,N_11566);
nand U12688 (N_12688,N_11295,N_11595);
xnor U12689 (N_12689,N_11420,N_11853);
nand U12690 (N_12690,N_11967,N_11939);
nand U12691 (N_12691,N_11934,N_11914);
and U12692 (N_12692,N_11318,N_11384);
nor U12693 (N_12693,N_11885,N_11824);
or U12694 (N_12694,N_11879,N_11599);
xor U12695 (N_12695,N_11868,N_11978);
and U12696 (N_12696,N_11843,N_11822);
nand U12697 (N_12697,N_11969,N_11679);
xnor U12698 (N_12698,N_11806,N_11638);
xor U12699 (N_12699,N_11711,N_11311);
xor U12700 (N_12700,N_11869,N_11583);
or U12701 (N_12701,N_11489,N_11829);
xor U12702 (N_12702,N_11417,N_11250);
nand U12703 (N_12703,N_11693,N_11333);
nand U12704 (N_12704,N_11810,N_11410);
or U12705 (N_12705,N_11627,N_11500);
or U12706 (N_12706,N_11294,N_11451);
nor U12707 (N_12707,N_11436,N_11485);
nand U12708 (N_12708,N_11348,N_11977);
or U12709 (N_12709,N_11249,N_11986);
and U12710 (N_12710,N_11990,N_11921);
xor U12711 (N_12711,N_11228,N_11749);
or U12712 (N_12712,N_11915,N_11879);
xnor U12713 (N_12713,N_11764,N_11709);
and U12714 (N_12714,N_11830,N_11892);
or U12715 (N_12715,N_11545,N_11340);
xnor U12716 (N_12716,N_11523,N_11955);
xor U12717 (N_12717,N_11790,N_11479);
and U12718 (N_12718,N_11375,N_11878);
and U12719 (N_12719,N_11928,N_11395);
nand U12720 (N_12720,N_11297,N_11358);
and U12721 (N_12721,N_11490,N_11688);
or U12722 (N_12722,N_11428,N_11914);
or U12723 (N_12723,N_11677,N_11266);
nor U12724 (N_12724,N_11320,N_11398);
xnor U12725 (N_12725,N_11413,N_11434);
and U12726 (N_12726,N_11301,N_11646);
or U12727 (N_12727,N_11324,N_11457);
nor U12728 (N_12728,N_11289,N_11329);
nand U12729 (N_12729,N_11549,N_11408);
or U12730 (N_12730,N_11501,N_11778);
and U12731 (N_12731,N_11984,N_11604);
or U12732 (N_12732,N_11354,N_11390);
xnor U12733 (N_12733,N_11835,N_11557);
or U12734 (N_12734,N_11986,N_11916);
or U12735 (N_12735,N_11477,N_11748);
and U12736 (N_12736,N_11418,N_11776);
and U12737 (N_12737,N_11853,N_11815);
nand U12738 (N_12738,N_11435,N_11598);
and U12739 (N_12739,N_11513,N_11746);
xor U12740 (N_12740,N_11760,N_11931);
nor U12741 (N_12741,N_11795,N_11361);
xor U12742 (N_12742,N_11416,N_11598);
nor U12743 (N_12743,N_11647,N_11384);
and U12744 (N_12744,N_11900,N_11402);
and U12745 (N_12745,N_11353,N_11665);
or U12746 (N_12746,N_11426,N_11251);
xnor U12747 (N_12747,N_11949,N_11463);
and U12748 (N_12748,N_11750,N_11575);
or U12749 (N_12749,N_11518,N_11456);
xor U12750 (N_12750,N_11232,N_11946);
xor U12751 (N_12751,N_11648,N_11911);
xor U12752 (N_12752,N_11757,N_11236);
or U12753 (N_12753,N_11266,N_11451);
and U12754 (N_12754,N_11273,N_11923);
and U12755 (N_12755,N_11319,N_11560);
or U12756 (N_12756,N_11280,N_11884);
or U12757 (N_12757,N_11707,N_11329);
xnor U12758 (N_12758,N_11596,N_11700);
and U12759 (N_12759,N_11997,N_11972);
or U12760 (N_12760,N_11968,N_11277);
and U12761 (N_12761,N_11613,N_11290);
nand U12762 (N_12762,N_11860,N_11727);
nor U12763 (N_12763,N_11539,N_11274);
or U12764 (N_12764,N_11589,N_11226);
nor U12765 (N_12765,N_11716,N_11697);
or U12766 (N_12766,N_11502,N_11791);
xor U12767 (N_12767,N_11598,N_11928);
or U12768 (N_12768,N_11387,N_11677);
xnor U12769 (N_12769,N_11902,N_11599);
nand U12770 (N_12770,N_11458,N_11228);
xor U12771 (N_12771,N_11385,N_11688);
or U12772 (N_12772,N_11431,N_11647);
nand U12773 (N_12773,N_11959,N_11408);
nand U12774 (N_12774,N_11247,N_11225);
nor U12775 (N_12775,N_11658,N_11517);
nand U12776 (N_12776,N_11924,N_11838);
nand U12777 (N_12777,N_11520,N_11428);
nand U12778 (N_12778,N_11478,N_11247);
xnor U12779 (N_12779,N_11482,N_11614);
or U12780 (N_12780,N_11760,N_11582);
nor U12781 (N_12781,N_11807,N_11860);
nor U12782 (N_12782,N_11996,N_11353);
and U12783 (N_12783,N_11717,N_11792);
xor U12784 (N_12784,N_11775,N_11343);
nor U12785 (N_12785,N_11742,N_11596);
and U12786 (N_12786,N_11652,N_11408);
or U12787 (N_12787,N_11297,N_11265);
nand U12788 (N_12788,N_11222,N_11302);
nor U12789 (N_12789,N_11308,N_11313);
xor U12790 (N_12790,N_11728,N_11257);
and U12791 (N_12791,N_11612,N_11622);
xor U12792 (N_12792,N_11648,N_11635);
and U12793 (N_12793,N_11746,N_11621);
nor U12794 (N_12794,N_11221,N_11238);
or U12795 (N_12795,N_11941,N_11954);
nor U12796 (N_12796,N_11864,N_11495);
nand U12797 (N_12797,N_11691,N_11378);
nor U12798 (N_12798,N_11932,N_11563);
or U12799 (N_12799,N_11892,N_11457);
and U12800 (N_12800,N_12073,N_12490);
nand U12801 (N_12801,N_12045,N_12398);
and U12802 (N_12802,N_12611,N_12781);
nand U12803 (N_12803,N_12279,N_12081);
nand U12804 (N_12804,N_12711,N_12480);
or U12805 (N_12805,N_12746,N_12732);
or U12806 (N_12806,N_12177,N_12683);
xor U12807 (N_12807,N_12248,N_12071);
and U12808 (N_12808,N_12531,N_12054);
xnor U12809 (N_12809,N_12691,N_12134);
nand U12810 (N_12810,N_12438,N_12430);
nor U12811 (N_12811,N_12464,N_12470);
or U12812 (N_12812,N_12640,N_12622);
xor U12813 (N_12813,N_12239,N_12420);
and U12814 (N_12814,N_12339,N_12079);
and U12815 (N_12815,N_12665,N_12387);
nor U12816 (N_12816,N_12779,N_12338);
nand U12817 (N_12817,N_12199,N_12331);
xnor U12818 (N_12818,N_12039,N_12208);
nand U12819 (N_12819,N_12591,N_12244);
and U12820 (N_12820,N_12778,N_12380);
xnor U12821 (N_12821,N_12587,N_12201);
or U12822 (N_12822,N_12427,N_12566);
or U12823 (N_12823,N_12588,N_12447);
nor U12824 (N_12824,N_12213,N_12151);
and U12825 (N_12825,N_12685,N_12247);
nor U12826 (N_12826,N_12735,N_12602);
nor U12827 (N_12827,N_12756,N_12075);
nand U12828 (N_12828,N_12590,N_12273);
nor U12829 (N_12829,N_12596,N_12312);
nor U12830 (N_12830,N_12658,N_12743);
xnor U12831 (N_12831,N_12061,N_12226);
xor U12832 (N_12832,N_12488,N_12451);
nor U12833 (N_12833,N_12599,N_12368);
xor U12834 (N_12834,N_12124,N_12722);
nand U12835 (N_12835,N_12540,N_12193);
or U12836 (N_12836,N_12576,N_12684);
xnor U12837 (N_12837,N_12332,N_12388);
and U12838 (N_12838,N_12625,N_12059);
nand U12839 (N_12839,N_12313,N_12027);
xor U12840 (N_12840,N_12284,N_12639);
and U12841 (N_12841,N_12409,N_12173);
nor U12842 (N_12842,N_12594,N_12696);
nand U12843 (N_12843,N_12532,N_12498);
or U12844 (N_12844,N_12355,N_12334);
xor U12845 (N_12845,N_12162,N_12125);
xor U12846 (N_12846,N_12314,N_12769);
nor U12847 (N_12847,N_12783,N_12495);
xor U12848 (N_12848,N_12363,N_12772);
nand U12849 (N_12849,N_12616,N_12174);
nor U12850 (N_12850,N_12318,N_12621);
nor U12851 (N_12851,N_12615,N_12237);
or U12852 (N_12852,N_12787,N_12433);
xor U12853 (N_12853,N_12015,N_12270);
or U12854 (N_12854,N_12041,N_12670);
nor U12855 (N_12855,N_12004,N_12219);
or U12856 (N_12856,N_12589,N_12399);
and U12857 (N_12857,N_12094,N_12389);
nand U12858 (N_12858,N_12579,N_12148);
or U12859 (N_12859,N_12565,N_12036);
nor U12860 (N_12860,N_12697,N_12262);
or U12861 (N_12861,N_12227,N_12757);
or U12862 (N_12862,N_12462,N_12394);
nor U12863 (N_12863,N_12517,N_12373);
and U12864 (N_12864,N_12644,N_12428);
nor U12865 (N_12865,N_12090,N_12062);
or U12866 (N_12866,N_12630,N_12144);
or U12867 (N_12867,N_12283,N_12725);
and U12868 (N_12868,N_12403,N_12136);
nor U12869 (N_12869,N_12421,N_12216);
and U12870 (N_12870,N_12286,N_12108);
or U12871 (N_12871,N_12224,N_12407);
nor U12872 (N_12872,N_12305,N_12269);
or U12873 (N_12873,N_12505,N_12768);
nand U12874 (N_12874,N_12546,N_12606);
and U12875 (N_12875,N_12731,N_12051);
xnor U12876 (N_12876,N_12196,N_12763);
or U12877 (N_12877,N_12664,N_12537);
xnor U12878 (N_12878,N_12063,N_12249);
or U12879 (N_12879,N_12453,N_12548);
nor U12880 (N_12880,N_12165,N_12310);
or U12881 (N_12881,N_12150,N_12281);
nand U12882 (N_12882,N_12533,N_12709);
nor U12883 (N_12883,N_12088,N_12350);
and U12884 (N_12884,N_12138,N_12450);
and U12885 (N_12885,N_12098,N_12460);
nor U12886 (N_12886,N_12483,N_12232);
xor U12887 (N_12887,N_12489,N_12544);
nand U12888 (N_12888,N_12432,N_12740);
nor U12889 (N_12889,N_12189,N_12021);
or U12890 (N_12890,N_12386,N_12390);
xnor U12891 (N_12891,N_12157,N_12065);
nor U12892 (N_12892,N_12475,N_12619);
nand U12893 (N_12893,N_12478,N_12677);
nand U12894 (N_12894,N_12229,N_12082);
xnor U12895 (N_12895,N_12295,N_12518);
xnor U12896 (N_12896,N_12033,N_12245);
or U12897 (N_12897,N_12751,N_12121);
or U12898 (N_12898,N_12184,N_12205);
xnor U12899 (N_12899,N_12440,N_12688);
xor U12900 (N_12900,N_12256,N_12442);
or U12901 (N_12901,N_12741,N_12477);
or U12902 (N_12902,N_12492,N_12123);
or U12903 (N_12903,N_12734,N_12646);
nand U12904 (N_12904,N_12209,N_12534);
and U12905 (N_12905,N_12127,N_12365);
nor U12906 (N_12906,N_12142,N_12200);
nand U12907 (N_12907,N_12005,N_12713);
nand U12908 (N_12908,N_12666,N_12364);
and U12909 (N_12909,N_12119,N_12745);
and U12910 (N_12910,N_12494,N_12328);
and U12911 (N_12911,N_12042,N_12261);
or U12912 (N_12912,N_12449,N_12774);
xor U12913 (N_12913,N_12406,N_12726);
or U12914 (N_12914,N_12794,N_12673);
or U12915 (N_12915,N_12309,N_12647);
or U12916 (N_12916,N_12105,N_12155);
xor U12917 (N_12917,N_12603,N_12107);
xor U12918 (N_12918,N_12096,N_12435);
and U12919 (N_12919,N_12454,N_12303);
or U12920 (N_12920,N_12613,N_12182);
nor U12921 (N_12921,N_12559,N_12292);
xor U12922 (N_12922,N_12300,N_12211);
nor U12923 (N_12923,N_12308,N_12325);
nor U12924 (N_12924,N_12265,N_12167);
nor U12925 (N_12925,N_12641,N_12567);
nand U12926 (N_12926,N_12422,N_12680);
nor U12927 (N_12927,N_12057,N_12360);
xor U12928 (N_12928,N_12795,N_12649);
xnor U12929 (N_12929,N_12058,N_12321);
nor U12930 (N_12930,N_12040,N_12744);
nor U12931 (N_12931,N_12500,N_12584);
nand U12932 (N_12932,N_12676,N_12299);
and U12933 (N_12933,N_12396,N_12733);
xor U12934 (N_12934,N_12258,N_12612);
or U12935 (N_12935,N_12048,N_12401);
or U12936 (N_12936,N_12788,N_12149);
or U12937 (N_12937,N_12719,N_12180);
or U12938 (N_12938,N_12761,N_12474);
and U12939 (N_12939,N_12547,N_12271);
nand U12940 (N_12940,N_12571,N_12444);
or U12941 (N_12941,N_12549,N_12607);
and U12942 (N_12942,N_12264,N_12780);
xnor U12943 (N_12943,N_12514,N_12439);
nand U12944 (N_12944,N_12163,N_12341);
xor U12945 (N_12945,N_12706,N_12070);
and U12946 (N_12946,N_12304,N_12476);
nand U12947 (N_12947,N_12714,N_12293);
or U12948 (N_12948,N_12158,N_12595);
nand U12949 (N_12949,N_12146,N_12662);
nand U12950 (N_12950,N_12347,N_12323);
nor U12951 (N_12951,N_12797,N_12570);
or U12952 (N_12952,N_12792,N_12551);
and U12953 (N_12953,N_12424,N_12789);
nor U12954 (N_12954,N_12154,N_12472);
nand U12955 (N_12955,N_12516,N_12623);
nor U12956 (N_12956,N_12049,N_12637);
or U12957 (N_12957,N_12352,N_12679);
nand U12958 (N_12958,N_12538,N_12749);
or U12959 (N_12959,N_12132,N_12324);
or U12960 (N_12960,N_12234,N_12605);
xnor U12961 (N_12961,N_12333,N_12416);
and U12962 (N_12962,N_12723,N_12340);
and U12963 (N_12963,N_12561,N_12100);
nor U12964 (N_12964,N_12361,N_12122);
nand U12965 (N_12965,N_12717,N_12598);
and U12966 (N_12966,N_12160,N_12291);
and U12967 (N_12967,N_12747,N_12259);
or U12968 (N_12968,N_12484,N_12228);
and U12969 (N_12969,N_12114,N_12542);
or U12970 (N_12970,N_12393,N_12446);
nand U12971 (N_12971,N_12097,N_12786);
or U12972 (N_12972,N_12089,N_12569);
or U12973 (N_12973,N_12025,N_12190);
nand U12974 (N_12974,N_12301,N_12586);
nor U12975 (N_12975,N_12520,N_12738);
xor U12976 (N_12976,N_12465,N_12212);
and U12977 (N_12977,N_12263,N_12012);
and U12978 (N_12978,N_12507,N_12554);
nor U12979 (N_12979,N_12539,N_12766);
nor U12980 (N_12980,N_12034,N_12001);
xnor U12981 (N_12981,N_12186,N_12230);
and U12982 (N_12982,N_12242,N_12408);
nand U12983 (N_12983,N_12557,N_12486);
xnor U12984 (N_12984,N_12515,N_12115);
nor U12985 (N_12985,N_12203,N_12471);
nand U12986 (N_12986,N_12139,N_12656);
xor U12987 (N_12987,N_12585,N_12626);
nand U12988 (N_12988,N_12701,N_12102);
nand U12989 (N_12989,N_12614,N_12103);
nor U12990 (N_12990,N_12636,N_12461);
nand U12991 (N_12991,N_12702,N_12175);
or U12992 (N_12992,N_12275,N_12770);
nand U12993 (N_12993,N_12133,N_12068);
nand U12994 (N_12994,N_12050,N_12671);
nor U12995 (N_12995,N_12060,N_12316);
xnor U12996 (N_12996,N_12536,N_12580);
nand U12997 (N_12997,N_12511,N_12760);
nand U12998 (N_12998,N_12366,N_12790);
xnor U12999 (N_12999,N_12276,N_12093);
or U13000 (N_13000,N_12415,N_12522);
xor U13001 (N_13001,N_12431,N_12633);
nor U13002 (N_13002,N_12043,N_12377);
nor U13003 (N_13003,N_12319,N_12631);
nand U13004 (N_13004,N_12535,N_12254);
nand U13005 (N_13005,N_12240,N_12499);
nor U13006 (N_13006,N_12066,N_12581);
and U13007 (N_13007,N_12251,N_12443);
and U13008 (N_13008,N_12436,N_12220);
xnor U13009 (N_13009,N_12217,N_12192);
nor U13010 (N_13010,N_12412,N_12330);
nor U13011 (N_13011,N_12092,N_12573);
nand U13012 (N_13012,N_12653,N_12690);
nand U13013 (N_13013,N_12512,N_12349);
nand U13014 (N_13014,N_12397,N_12693);
nor U13015 (N_13015,N_12502,N_12392);
and U13016 (N_13016,N_12624,N_12290);
xor U13017 (N_13017,N_12335,N_12469);
xor U13018 (N_13018,N_12140,N_12267);
nor U13019 (N_13019,N_12404,N_12455);
and U13020 (N_13020,N_12600,N_12378);
and U13021 (N_13021,N_12253,N_12326);
nand U13022 (N_13022,N_12562,N_12171);
nor U13023 (N_13023,N_12592,N_12638);
and U13024 (N_13024,N_12705,N_12503);
and U13025 (N_13025,N_12715,N_12410);
or U13026 (N_13026,N_12374,N_12423);
and U13027 (N_13027,N_12750,N_12654);
nand U13028 (N_13028,N_12381,N_12185);
nand U13029 (N_13029,N_12764,N_12692);
nand U13030 (N_13030,N_12748,N_12370);
nand U13031 (N_13031,N_12222,N_12306);
nor U13032 (N_13032,N_12675,N_12117);
xnor U13033 (N_13033,N_12445,N_12737);
xnor U13034 (N_13034,N_12037,N_12775);
nor U13035 (N_13035,N_12456,N_12014);
and U13036 (N_13036,N_12101,N_12651);
and U13037 (N_13037,N_12007,N_12266);
or U13038 (N_13038,N_12545,N_12672);
nor U13039 (N_13039,N_12129,N_12504);
nor U13040 (N_13040,N_12597,N_12032);
nand U13041 (N_13041,N_12329,N_12011);
and U13042 (N_13042,N_12112,N_12215);
or U13043 (N_13043,N_12437,N_12187);
nor U13044 (N_13044,N_12345,N_12609);
and U13045 (N_13045,N_12391,N_12031);
and U13046 (N_13046,N_12116,N_12371);
and U13047 (N_13047,N_12047,N_12218);
and U13048 (N_13048,N_12231,N_12348);
nand U13049 (N_13049,N_12730,N_12161);
or U13050 (N_13050,N_12635,N_12022);
or U13051 (N_13051,N_12235,N_12686);
xnor U13052 (N_13052,N_12003,N_12320);
nor U13053 (N_13053,N_12556,N_12009);
xnor U13054 (N_13054,N_12257,N_12225);
xnor U13055 (N_13055,N_12179,N_12091);
or U13056 (N_13056,N_12362,N_12289);
and U13057 (N_13057,N_12601,N_12233);
nor U13058 (N_13058,N_12016,N_12659);
xor U13059 (N_13059,N_12356,N_12467);
nand U13060 (N_13060,N_12152,N_12052);
nand U13061 (N_13061,N_12297,N_12118);
nor U13062 (N_13062,N_12564,N_12210);
or U13063 (N_13063,N_12418,N_12681);
xnor U13064 (N_13064,N_12188,N_12642);
nor U13065 (N_13065,N_12742,N_12541);
nor U13066 (N_13066,N_12669,N_12652);
nand U13067 (N_13067,N_12298,N_12035);
nor U13068 (N_13068,N_12491,N_12194);
or U13069 (N_13069,N_12078,N_12523);
nand U13070 (N_13070,N_12689,N_12385);
nor U13071 (N_13071,N_12181,N_12776);
nor U13072 (N_13072,N_12459,N_12250);
nand U13073 (N_13073,N_12657,N_12074);
xnor U13074 (N_13074,N_12682,N_12583);
nor U13075 (N_13075,N_12575,N_12720);
or U13076 (N_13076,N_12120,N_12246);
and U13077 (N_13077,N_12145,N_12558);
and U13078 (N_13078,N_12076,N_12353);
nor U13079 (N_13079,N_12086,N_12315);
xnor U13080 (N_13080,N_12466,N_12243);
nand U13081 (N_13081,N_12288,N_12238);
nand U13082 (N_13082,N_12147,N_12425);
nor U13083 (N_13083,N_12191,N_12650);
nor U13084 (N_13084,N_12317,N_12170);
and U13085 (N_13085,N_12487,N_12496);
nor U13086 (N_13086,N_12553,N_12026);
or U13087 (N_13087,N_12367,N_12067);
and U13088 (N_13088,N_12668,N_12582);
xor U13089 (N_13089,N_12777,N_12277);
nor U13090 (N_13090,N_12574,N_12204);
nand U13091 (N_13091,N_12207,N_12080);
nand U13092 (N_13092,N_12645,N_12020);
nand U13093 (N_13093,N_12023,N_12527);
or U13094 (N_13094,N_12010,N_12434);
nor U13095 (N_13095,N_12593,N_12643);
and U13096 (N_13096,N_12452,N_12056);
nor U13097 (N_13097,N_12767,N_12354);
and U13098 (N_13098,N_12166,N_12628);
xnor U13099 (N_13099,N_12799,N_12302);
and U13100 (N_13100,N_12064,N_12024);
xnor U13101 (N_13101,N_12798,N_12441);
and U13102 (N_13102,N_12106,N_12383);
or U13103 (N_13103,N_12513,N_12728);
xnor U13104 (N_13104,N_12784,N_12530);
nor U13105 (N_13105,N_12721,N_12759);
and U13106 (N_13106,N_12716,N_12274);
nor U13107 (N_13107,N_12796,N_12578);
xnor U13108 (N_13108,N_12159,N_12137);
xnor U13109 (N_13109,N_12130,N_12202);
nor U13110 (N_13110,N_12627,N_12358);
or U13111 (N_13111,N_12634,N_12791);
and U13112 (N_13112,N_12084,N_12169);
and U13113 (N_13113,N_12506,N_12176);
xnor U13114 (N_13114,N_12285,N_12294);
xor U13115 (N_13115,N_12085,N_12044);
nor U13116 (N_13116,N_12272,N_12473);
nor U13117 (N_13117,N_12069,N_12164);
xnor U13118 (N_13118,N_12699,N_12346);
and U13119 (N_13119,N_12754,N_12405);
or U13120 (N_13120,N_12482,N_12694);
nor U13121 (N_13121,N_12156,N_12729);
xnor U13122 (N_13122,N_12758,N_12402);
nor U13123 (N_13123,N_12663,N_12083);
xnor U13124 (N_13124,N_12604,N_12710);
nor U13125 (N_13125,N_12241,N_12655);
nor U13126 (N_13126,N_12153,N_12030);
nor U13127 (N_13127,N_12135,N_12762);
xnor U13128 (N_13128,N_12379,N_12343);
nand U13129 (N_13129,N_12501,N_12429);
nor U13130 (N_13130,N_12006,N_12753);
nor U13131 (N_13131,N_12287,N_12525);
nand U13132 (N_13132,N_12519,N_12206);
nor U13133 (N_13133,N_12555,N_12577);
xnor U13134 (N_13134,N_12311,N_12687);
nand U13135 (N_13135,N_12695,N_12375);
or U13136 (N_13136,N_12785,N_12183);
xnor U13137 (N_13137,N_12620,N_12413);
and U13138 (N_13138,N_12793,N_12327);
xor U13139 (N_13139,N_12357,N_12718);
and U13140 (N_13140,N_12463,N_12131);
xnor U13141 (N_13141,N_12736,N_12278);
or U13142 (N_13142,N_12497,N_12674);
and U13143 (N_13143,N_12017,N_12707);
xnor U13144 (N_13144,N_12128,N_12002);
nand U13145 (N_13145,N_12568,N_12493);
nor U13146 (N_13146,N_12110,N_12104);
and U13147 (N_13147,N_12481,N_12724);
and U13148 (N_13148,N_12099,N_12143);
xnor U13149 (N_13149,N_12700,N_12055);
or U13150 (N_13150,N_12029,N_12126);
and U13151 (N_13151,N_12280,N_12018);
nor U13152 (N_13152,N_12667,N_12426);
and U13153 (N_13153,N_12755,N_12528);
nor U13154 (N_13154,N_12529,N_12252);
and U13155 (N_13155,N_12485,N_12168);
or U13156 (N_13156,N_12550,N_12648);
and U13157 (N_13157,N_12369,N_12342);
xnor U13158 (N_13158,N_12197,N_12282);
nor U13159 (N_13159,N_12457,N_12198);
nor U13160 (N_13160,N_12337,N_12268);
or U13161 (N_13161,N_12221,N_12296);
nand U13162 (N_13162,N_12141,N_12382);
nor U13163 (N_13163,N_12629,N_12563);
nand U13164 (N_13164,N_12307,N_12414);
and U13165 (N_13165,N_12053,N_12077);
xnor U13166 (N_13166,N_12113,N_12526);
nor U13167 (N_13167,N_12552,N_12727);
and U13168 (N_13168,N_12411,N_12524);
xor U13169 (N_13169,N_12468,N_12038);
xnor U13170 (N_13170,N_12255,N_12395);
nand U13171 (N_13171,N_12417,N_12178);
and U13172 (N_13172,N_12771,N_12752);
and U13173 (N_13173,N_12660,N_12479);
xnor U13174 (N_13174,N_12000,N_12322);
xor U13175 (N_13175,N_12678,N_12223);
nor U13176 (N_13176,N_12195,N_12509);
nand U13177 (N_13177,N_12712,N_12704);
or U13178 (N_13178,N_12632,N_12608);
and U13179 (N_13179,N_12572,N_12236);
nor U13180 (N_13180,N_12765,N_12400);
nor U13181 (N_13181,N_12510,N_12448);
xnor U13182 (N_13182,N_12111,N_12344);
xor U13183 (N_13183,N_12610,N_12508);
nand U13184 (N_13184,N_12384,N_12372);
xnor U13185 (N_13185,N_12661,N_12019);
xor U13186 (N_13186,N_12618,N_12109);
xnor U13187 (N_13187,N_12351,N_12376);
and U13188 (N_13188,N_12560,N_12013);
or U13189 (N_13189,N_12214,N_12739);
or U13190 (N_13190,N_12419,N_12072);
and U13191 (N_13191,N_12708,N_12336);
or U13192 (N_13192,N_12172,N_12458);
and U13193 (N_13193,N_12260,N_12703);
nand U13194 (N_13194,N_12543,N_12028);
nand U13195 (N_13195,N_12782,N_12095);
nand U13196 (N_13196,N_12046,N_12617);
nor U13197 (N_13197,N_12521,N_12087);
xnor U13198 (N_13198,N_12008,N_12773);
nand U13199 (N_13199,N_12698,N_12359);
and U13200 (N_13200,N_12246,N_12295);
or U13201 (N_13201,N_12796,N_12029);
or U13202 (N_13202,N_12717,N_12602);
xor U13203 (N_13203,N_12225,N_12682);
nor U13204 (N_13204,N_12744,N_12159);
nand U13205 (N_13205,N_12297,N_12448);
and U13206 (N_13206,N_12258,N_12321);
and U13207 (N_13207,N_12084,N_12154);
and U13208 (N_13208,N_12174,N_12631);
xor U13209 (N_13209,N_12441,N_12677);
xnor U13210 (N_13210,N_12351,N_12435);
and U13211 (N_13211,N_12076,N_12572);
or U13212 (N_13212,N_12522,N_12232);
nand U13213 (N_13213,N_12427,N_12739);
and U13214 (N_13214,N_12454,N_12366);
and U13215 (N_13215,N_12298,N_12129);
or U13216 (N_13216,N_12488,N_12596);
nand U13217 (N_13217,N_12034,N_12229);
nand U13218 (N_13218,N_12660,N_12472);
nand U13219 (N_13219,N_12039,N_12151);
nor U13220 (N_13220,N_12417,N_12485);
nor U13221 (N_13221,N_12644,N_12049);
nor U13222 (N_13222,N_12430,N_12626);
nor U13223 (N_13223,N_12323,N_12481);
or U13224 (N_13224,N_12031,N_12397);
nor U13225 (N_13225,N_12797,N_12538);
and U13226 (N_13226,N_12723,N_12611);
xor U13227 (N_13227,N_12557,N_12279);
nor U13228 (N_13228,N_12647,N_12268);
nand U13229 (N_13229,N_12729,N_12544);
nand U13230 (N_13230,N_12387,N_12101);
nand U13231 (N_13231,N_12571,N_12727);
or U13232 (N_13232,N_12120,N_12162);
nor U13233 (N_13233,N_12461,N_12414);
nor U13234 (N_13234,N_12183,N_12527);
and U13235 (N_13235,N_12395,N_12605);
nand U13236 (N_13236,N_12312,N_12447);
xnor U13237 (N_13237,N_12293,N_12199);
and U13238 (N_13238,N_12586,N_12328);
xnor U13239 (N_13239,N_12564,N_12471);
xor U13240 (N_13240,N_12490,N_12482);
nand U13241 (N_13241,N_12191,N_12702);
and U13242 (N_13242,N_12249,N_12036);
xnor U13243 (N_13243,N_12653,N_12479);
nor U13244 (N_13244,N_12716,N_12224);
nor U13245 (N_13245,N_12565,N_12015);
nor U13246 (N_13246,N_12565,N_12220);
and U13247 (N_13247,N_12346,N_12338);
nor U13248 (N_13248,N_12797,N_12734);
or U13249 (N_13249,N_12540,N_12754);
nor U13250 (N_13250,N_12120,N_12044);
xnor U13251 (N_13251,N_12006,N_12661);
nand U13252 (N_13252,N_12491,N_12388);
nor U13253 (N_13253,N_12061,N_12346);
nand U13254 (N_13254,N_12048,N_12010);
nor U13255 (N_13255,N_12465,N_12270);
nand U13256 (N_13256,N_12094,N_12166);
or U13257 (N_13257,N_12568,N_12516);
nor U13258 (N_13258,N_12043,N_12761);
nand U13259 (N_13259,N_12674,N_12444);
xor U13260 (N_13260,N_12248,N_12573);
and U13261 (N_13261,N_12220,N_12242);
or U13262 (N_13262,N_12711,N_12062);
xor U13263 (N_13263,N_12252,N_12110);
xor U13264 (N_13264,N_12718,N_12131);
xnor U13265 (N_13265,N_12166,N_12794);
and U13266 (N_13266,N_12432,N_12530);
nor U13267 (N_13267,N_12497,N_12711);
xor U13268 (N_13268,N_12248,N_12273);
nand U13269 (N_13269,N_12073,N_12449);
nor U13270 (N_13270,N_12626,N_12458);
nor U13271 (N_13271,N_12232,N_12506);
or U13272 (N_13272,N_12602,N_12090);
and U13273 (N_13273,N_12511,N_12224);
nand U13274 (N_13274,N_12524,N_12448);
nand U13275 (N_13275,N_12233,N_12521);
and U13276 (N_13276,N_12076,N_12228);
xnor U13277 (N_13277,N_12023,N_12215);
nand U13278 (N_13278,N_12382,N_12209);
nor U13279 (N_13279,N_12102,N_12598);
nand U13280 (N_13280,N_12060,N_12157);
or U13281 (N_13281,N_12611,N_12260);
xnor U13282 (N_13282,N_12471,N_12217);
xor U13283 (N_13283,N_12599,N_12033);
nor U13284 (N_13284,N_12119,N_12360);
nand U13285 (N_13285,N_12320,N_12701);
and U13286 (N_13286,N_12200,N_12084);
nor U13287 (N_13287,N_12153,N_12463);
xor U13288 (N_13288,N_12300,N_12719);
nand U13289 (N_13289,N_12330,N_12158);
nor U13290 (N_13290,N_12446,N_12035);
nor U13291 (N_13291,N_12687,N_12014);
xor U13292 (N_13292,N_12617,N_12096);
xor U13293 (N_13293,N_12124,N_12739);
or U13294 (N_13294,N_12444,N_12373);
nor U13295 (N_13295,N_12500,N_12111);
and U13296 (N_13296,N_12348,N_12092);
or U13297 (N_13297,N_12208,N_12094);
xor U13298 (N_13298,N_12391,N_12468);
nor U13299 (N_13299,N_12164,N_12175);
and U13300 (N_13300,N_12463,N_12662);
xor U13301 (N_13301,N_12429,N_12202);
and U13302 (N_13302,N_12076,N_12364);
xor U13303 (N_13303,N_12355,N_12408);
nor U13304 (N_13304,N_12048,N_12694);
and U13305 (N_13305,N_12120,N_12025);
or U13306 (N_13306,N_12526,N_12261);
nand U13307 (N_13307,N_12661,N_12727);
xor U13308 (N_13308,N_12788,N_12580);
xor U13309 (N_13309,N_12111,N_12270);
and U13310 (N_13310,N_12612,N_12330);
or U13311 (N_13311,N_12342,N_12333);
and U13312 (N_13312,N_12568,N_12741);
xor U13313 (N_13313,N_12322,N_12217);
nand U13314 (N_13314,N_12308,N_12773);
nand U13315 (N_13315,N_12415,N_12409);
nor U13316 (N_13316,N_12497,N_12054);
or U13317 (N_13317,N_12170,N_12684);
or U13318 (N_13318,N_12094,N_12771);
or U13319 (N_13319,N_12308,N_12190);
xor U13320 (N_13320,N_12257,N_12235);
nand U13321 (N_13321,N_12757,N_12040);
nand U13322 (N_13322,N_12267,N_12519);
xnor U13323 (N_13323,N_12077,N_12167);
xnor U13324 (N_13324,N_12543,N_12529);
xor U13325 (N_13325,N_12188,N_12598);
or U13326 (N_13326,N_12673,N_12278);
and U13327 (N_13327,N_12420,N_12007);
and U13328 (N_13328,N_12156,N_12291);
or U13329 (N_13329,N_12338,N_12582);
and U13330 (N_13330,N_12421,N_12646);
and U13331 (N_13331,N_12466,N_12366);
and U13332 (N_13332,N_12237,N_12372);
xor U13333 (N_13333,N_12047,N_12447);
nand U13334 (N_13334,N_12188,N_12741);
or U13335 (N_13335,N_12066,N_12095);
xnor U13336 (N_13336,N_12794,N_12681);
nand U13337 (N_13337,N_12637,N_12232);
xnor U13338 (N_13338,N_12575,N_12127);
nand U13339 (N_13339,N_12251,N_12658);
xor U13340 (N_13340,N_12617,N_12742);
or U13341 (N_13341,N_12582,N_12298);
nand U13342 (N_13342,N_12527,N_12634);
or U13343 (N_13343,N_12772,N_12554);
and U13344 (N_13344,N_12303,N_12527);
and U13345 (N_13345,N_12572,N_12681);
nor U13346 (N_13346,N_12565,N_12671);
nor U13347 (N_13347,N_12519,N_12384);
xor U13348 (N_13348,N_12475,N_12322);
nor U13349 (N_13349,N_12136,N_12545);
nor U13350 (N_13350,N_12165,N_12630);
or U13351 (N_13351,N_12250,N_12451);
xor U13352 (N_13352,N_12764,N_12796);
xor U13353 (N_13353,N_12378,N_12755);
and U13354 (N_13354,N_12220,N_12082);
nand U13355 (N_13355,N_12263,N_12644);
or U13356 (N_13356,N_12392,N_12533);
and U13357 (N_13357,N_12617,N_12302);
xor U13358 (N_13358,N_12786,N_12647);
xnor U13359 (N_13359,N_12095,N_12349);
and U13360 (N_13360,N_12251,N_12797);
or U13361 (N_13361,N_12752,N_12167);
nand U13362 (N_13362,N_12730,N_12382);
or U13363 (N_13363,N_12337,N_12519);
xnor U13364 (N_13364,N_12107,N_12333);
xor U13365 (N_13365,N_12425,N_12170);
or U13366 (N_13366,N_12609,N_12319);
nor U13367 (N_13367,N_12490,N_12729);
and U13368 (N_13368,N_12049,N_12115);
nor U13369 (N_13369,N_12637,N_12645);
and U13370 (N_13370,N_12327,N_12348);
and U13371 (N_13371,N_12174,N_12219);
nand U13372 (N_13372,N_12307,N_12500);
and U13373 (N_13373,N_12368,N_12392);
nor U13374 (N_13374,N_12380,N_12029);
nor U13375 (N_13375,N_12729,N_12026);
nor U13376 (N_13376,N_12417,N_12235);
nand U13377 (N_13377,N_12410,N_12582);
nor U13378 (N_13378,N_12520,N_12390);
or U13379 (N_13379,N_12382,N_12115);
and U13380 (N_13380,N_12501,N_12366);
xnor U13381 (N_13381,N_12221,N_12622);
xnor U13382 (N_13382,N_12553,N_12550);
or U13383 (N_13383,N_12670,N_12428);
and U13384 (N_13384,N_12084,N_12337);
nor U13385 (N_13385,N_12131,N_12321);
nand U13386 (N_13386,N_12759,N_12743);
or U13387 (N_13387,N_12186,N_12698);
nor U13388 (N_13388,N_12645,N_12440);
xnor U13389 (N_13389,N_12275,N_12135);
xnor U13390 (N_13390,N_12521,N_12333);
or U13391 (N_13391,N_12171,N_12708);
nor U13392 (N_13392,N_12387,N_12617);
or U13393 (N_13393,N_12174,N_12095);
and U13394 (N_13394,N_12517,N_12741);
nand U13395 (N_13395,N_12378,N_12047);
or U13396 (N_13396,N_12785,N_12779);
and U13397 (N_13397,N_12556,N_12555);
nor U13398 (N_13398,N_12655,N_12357);
nor U13399 (N_13399,N_12546,N_12207);
nor U13400 (N_13400,N_12207,N_12497);
or U13401 (N_13401,N_12555,N_12370);
or U13402 (N_13402,N_12593,N_12506);
nand U13403 (N_13403,N_12771,N_12499);
or U13404 (N_13404,N_12279,N_12198);
and U13405 (N_13405,N_12513,N_12245);
and U13406 (N_13406,N_12413,N_12253);
or U13407 (N_13407,N_12777,N_12640);
xor U13408 (N_13408,N_12275,N_12317);
xor U13409 (N_13409,N_12009,N_12552);
xnor U13410 (N_13410,N_12007,N_12741);
and U13411 (N_13411,N_12753,N_12138);
nand U13412 (N_13412,N_12422,N_12395);
or U13413 (N_13413,N_12265,N_12326);
nor U13414 (N_13414,N_12380,N_12538);
and U13415 (N_13415,N_12160,N_12511);
or U13416 (N_13416,N_12318,N_12258);
nor U13417 (N_13417,N_12365,N_12595);
or U13418 (N_13418,N_12446,N_12477);
nor U13419 (N_13419,N_12307,N_12514);
or U13420 (N_13420,N_12422,N_12420);
and U13421 (N_13421,N_12167,N_12232);
nor U13422 (N_13422,N_12320,N_12363);
xor U13423 (N_13423,N_12541,N_12456);
xnor U13424 (N_13424,N_12123,N_12124);
nand U13425 (N_13425,N_12651,N_12782);
and U13426 (N_13426,N_12331,N_12373);
nor U13427 (N_13427,N_12601,N_12729);
and U13428 (N_13428,N_12018,N_12473);
and U13429 (N_13429,N_12446,N_12454);
or U13430 (N_13430,N_12721,N_12142);
and U13431 (N_13431,N_12494,N_12642);
nor U13432 (N_13432,N_12483,N_12340);
or U13433 (N_13433,N_12325,N_12518);
nand U13434 (N_13434,N_12551,N_12325);
xor U13435 (N_13435,N_12475,N_12171);
or U13436 (N_13436,N_12551,N_12230);
xor U13437 (N_13437,N_12338,N_12039);
or U13438 (N_13438,N_12453,N_12387);
nand U13439 (N_13439,N_12697,N_12722);
and U13440 (N_13440,N_12609,N_12058);
xor U13441 (N_13441,N_12732,N_12132);
xor U13442 (N_13442,N_12003,N_12467);
and U13443 (N_13443,N_12474,N_12539);
xor U13444 (N_13444,N_12132,N_12261);
xor U13445 (N_13445,N_12718,N_12198);
or U13446 (N_13446,N_12777,N_12437);
nor U13447 (N_13447,N_12652,N_12326);
xnor U13448 (N_13448,N_12695,N_12439);
nand U13449 (N_13449,N_12502,N_12029);
nand U13450 (N_13450,N_12441,N_12240);
nand U13451 (N_13451,N_12644,N_12248);
nor U13452 (N_13452,N_12729,N_12476);
nand U13453 (N_13453,N_12406,N_12711);
xor U13454 (N_13454,N_12792,N_12711);
or U13455 (N_13455,N_12639,N_12548);
nand U13456 (N_13456,N_12528,N_12089);
nor U13457 (N_13457,N_12289,N_12678);
nand U13458 (N_13458,N_12088,N_12455);
nor U13459 (N_13459,N_12594,N_12740);
xor U13460 (N_13460,N_12487,N_12705);
nand U13461 (N_13461,N_12749,N_12134);
and U13462 (N_13462,N_12585,N_12706);
or U13463 (N_13463,N_12572,N_12710);
xor U13464 (N_13464,N_12475,N_12507);
nor U13465 (N_13465,N_12196,N_12513);
nor U13466 (N_13466,N_12085,N_12532);
nand U13467 (N_13467,N_12355,N_12135);
nor U13468 (N_13468,N_12342,N_12672);
nor U13469 (N_13469,N_12574,N_12304);
or U13470 (N_13470,N_12541,N_12540);
xnor U13471 (N_13471,N_12230,N_12233);
nand U13472 (N_13472,N_12790,N_12578);
nor U13473 (N_13473,N_12757,N_12709);
nand U13474 (N_13474,N_12676,N_12264);
and U13475 (N_13475,N_12224,N_12590);
nor U13476 (N_13476,N_12051,N_12151);
or U13477 (N_13477,N_12486,N_12148);
nor U13478 (N_13478,N_12197,N_12264);
nor U13479 (N_13479,N_12530,N_12093);
nor U13480 (N_13480,N_12210,N_12637);
nand U13481 (N_13481,N_12688,N_12557);
nand U13482 (N_13482,N_12658,N_12469);
nand U13483 (N_13483,N_12774,N_12648);
nand U13484 (N_13484,N_12749,N_12573);
xor U13485 (N_13485,N_12456,N_12216);
xnor U13486 (N_13486,N_12684,N_12237);
or U13487 (N_13487,N_12481,N_12110);
and U13488 (N_13488,N_12590,N_12085);
nand U13489 (N_13489,N_12772,N_12029);
nor U13490 (N_13490,N_12361,N_12435);
nand U13491 (N_13491,N_12137,N_12041);
or U13492 (N_13492,N_12632,N_12643);
or U13493 (N_13493,N_12144,N_12056);
xnor U13494 (N_13494,N_12363,N_12120);
nor U13495 (N_13495,N_12464,N_12741);
nor U13496 (N_13496,N_12429,N_12132);
nor U13497 (N_13497,N_12697,N_12159);
xnor U13498 (N_13498,N_12701,N_12652);
nand U13499 (N_13499,N_12342,N_12127);
and U13500 (N_13500,N_12649,N_12557);
xnor U13501 (N_13501,N_12384,N_12470);
nor U13502 (N_13502,N_12679,N_12242);
nand U13503 (N_13503,N_12005,N_12159);
nor U13504 (N_13504,N_12000,N_12694);
nand U13505 (N_13505,N_12010,N_12268);
xnor U13506 (N_13506,N_12107,N_12708);
and U13507 (N_13507,N_12201,N_12395);
xnor U13508 (N_13508,N_12219,N_12370);
xor U13509 (N_13509,N_12704,N_12782);
and U13510 (N_13510,N_12568,N_12754);
and U13511 (N_13511,N_12755,N_12533);
nor U13512 (N_13512,N_12389,N_12742);
xnor U13513 (N_13513,N_12371,N_12219);
nand U13514 (N_13514,N_12619,N_12646);
nor U13515 (N_13515,N_12505,N_12480);
or U13516 (N_13516,N_12248,N_12233);
xnor U13517 (N_13517,N_12006,N_12371);
and U13518 (N_13518,N_12320,N_12150);
nand U13519 (N_13519,N_12391,N_12317);
nor U13520 (N_13520,N_12214,N_12116);
and U13521 (N_13521,N_12155,N_12000);
nor U13522 (N_13522,N_12188,N_12468);
nor U13523 (N_13523,N_12522,N_12266);
or U13524 (N_13524,N_12761,N_12662);
and U13525 (N_13525,N_12632,N_12711);
or U13526 (N_13526,N_12153,N_12404);
nor U13527 (N_13527,N_12647,N_12083);
or U13528 (N_13528,N_12791,N_12780);
nand U13529 (N_13529,N_12438,N_12343);
nand U13530 (N_13530,N_12093,N_12714);
and U13531 (N_13531,N_12681,N_12030);
or U13532 (N_13532,N_12290,N_12176);
nand U13533 (N_13533,N_12606,N_12482);
and U13534 (N_13534,N_12299,N_12309);
nand U13535 (N_13535,N_12093,N_12743);
nand U13536 (N_13536,N_12677,N_12061);
nor U13537 (N_13537,N_12276,N_12419);
xnor U13538 (N_13538,N_12373,N_12301);
nor U13539 (N_13539,N_12314,N_12533);
nor U13540 (N_13540,N_12705,N_12615);
or U13541 (N_13541,N_12204,N_12695);
nor U13542 (N_13542,N_12129,N_12679);
xnor U13543 (N_13543,N_12241,N_12768);
nand U13544 (N_13544,N_12611,N_12682);
or U13545 (N_13545,N_12016,N_12400);
xor U13546 (N_13546,N_12725,N_12710);
or U13547 (N_13547,N_12430,N_12597);
and U13548 (N_13548,N_12716,N_12071);
and U13549 (N_13549,N_12337,N_12497);
nand U13550 (N_13550,N_12719,N_12516);
xor U13551 (N_13551,N_12438,N_12284);
or U13552 (N_13552,N_12604,N_12145);
xor U13553 (N_13553,N_12298,N_12138);
and U13554 (N_13554,N_12783,N_12215);
nor U13555 (N_13555,N_12409,N_12425);
and U13556 (N_13556,N_12512,N_12153);
or U13557 (N_13557,N_12773,N_12742);
nand U13558 (N_13558,N_12211,N_12163);
xnor U13559 (N_13559,N_12767,N_12693);
or U13560 (N_13560,N_12381,N_12023);
nand U13561 (N_13561,N_12480,N_12552);
nand U13562 (N_13562,N_12190,N_12606);
and U13563 (N_13563,N_12048,N_12172);
and U13564 (N_13564,N_12197,N_12644);
xor U13565 (N_13565,N_12358,N_12199);
nor U13566 (N_13566,N_12020,N_12705);
or U13567 (N_13567,N_12789,N_12177);
nand U13568 (N_13568,N_12383,N_12665);
nand U13569 (N_13569,N_12477,N_12591);
nand U13570 (N_13570,N_12567,N_12157);
xnor U13571 (N_13571,N_12128,N_12308);
nor U13572 (N_13572,N_12072,N_12509);
nor U13573 (N_13573,N_12651,N_12532);
or U13574 (N_13574,N_12747,N_12642);
nand U13575 (N_13575,N_12380,N_12098);
xor U13576 (N_13576,N_12163,N_12309);
nor U13577 (N_13577,N_12410,N_12250);
or U13578 (N_13578,N_12011,N_12440);
nand U13579 (N_13579,N_12674,N_12495);
nor U13580 (N_13580,N_12115,N_12224);
nand U13581 (N_13581,N_12172,N_12147);
nand U13582 (N_13582,N_12517,N_12284);
xnor U13583 (N_13583,N_12570,N_12086);
nand U13584 (N_13584,N_12139,N_12431);
or U13585 (N_13585,N_12038,N_12352);
xor U13586 (N_13586,N_12305,N_12024);
and U13587 (N_13587,N_12128,N_12357);
nor U13588 (N_13588,N_12525,N_12607);
nor U13589 (N_13589,N_12337,N_12400);
nor U13590 (N_13590,N_12547,N_12649);
nor U13591 (N_13591,N_12362,N_12504);
nand U13592 (N_13592,N_12509,N_12653);
or U13593 (N_13593,N_12079,N_12547);
xnor U13594 (N_13594,N_12528,N_12768);
nor U13595 (N_13595,N_12027,N_12716);
nor U13596 (N_13596,N_12197,N_12291);
xnor U13597 (N_13597,N_12190,N_12205);
nor U13598 (N_13598,N_12197,N_12371);
nor U13599 (N_13599,N_12337,N_12192);
or U13600 (N_13600,N_12902,N_13229);
xor U13601 (N_13601,N_13515,N_13011);
nand U13602 (N_13602,N_12836,N_12866);
nor U13603 (N_13603,N_13311,N_13263);
nor U13604 (N_13604,N_13210,N_13201);
and U13605 (N_13605,N_13153,N_13059);
and U13606 (N_13606,N_12935,N_13048);
or U13607 (N_13607,N_13445,N_13232);
xnor U13608 (N_13608,N_12811,N_13408);
xnor U13609 (N_13609,N_13248,N_13168);
or U13610 (N_13610,N_13301,N_13243);
nand U13611 (N_13611,N_13100,N_13335);
or U13612 (N_13612,N_13547,N_13390);
and U13613 (N_13613,N_13298,N_12861);
xor U13614 (N_13614,N_12807,N_13411);
xor U13615 (N_13615,N_13249,N_13043);
and U13616 (N_13616,N_12883,N_12851);
xor U13617 (N_13617,N_13065,N_12808);
nor U13618 (N_13618,N_12986,N_13215);
nor U13619 (N_13619,N_13258,N_13129);
nand U13620 (N_13620,N_12812,N_13045);
or U13621 (N_13621,N_13133,N_13510);
nor U13622 (N_13622,N_13016,N_13125);
or U13623 (N_13623,N_12805,N_13091);
nor U13624 (N_13624,N_13211,N_13173);
and U13625 (N_13625,N_12910,N_12835);
or U13626 (N_13626,N_13368,N_13039);
or U13627 (N_13627,N_13521,N_13351);
xor U13628 (N_13628,N_13049,N_12936);
and U13629 (N_13629,N_13018,N_13165);
or U13630 (N_13630,N_12955,N_13349);
xor U13631 (N_13631,N_12884,N_12945);
and U13632 (N_13632,N_12991,N_12845);
xnor U13633 (N_13633,N_13115,N_13325);
xnor U13634 (N_13634,N_13545,N_13527);
nor U13635 (N_13635,N_12973,N_13227);
or U13636 (N_13636,N_12939,N_13312);
xor U13637 (N_13637,N_13599,N_13481);
nor U13638 (N_13638,N_13340,N_13145);
or U13639 (N_13639,N_13446,N_13402);
or U13640 (N_13640,N_12843,N_13486);
and U13641 (N_13641,N_13314,N_12891);
nor U13642 (N_13642,N_12852,N_13162);
xnor U13643 (N_13643,N_13093,N_13352);
or U13644 (N_13644,N_13562,N_12961);
xnor U13645 (N_13645,N_13254,N_12922);
nand U13646 (N_13646,N_13507,N_13102);
xnor U13647 (N_13647,N_13084,N_13556);
xor U13648 (N_13648,N_13242,N_12975);
xor U13649 (N_13649,N_13364,N_12987);
nor U13650 (N_13650,N_13041,N_13096);
nand U13651 (N_13651,N_13321,N_13158);
nor U13652 (N_13652,N_13310,N_13555);
xor U13653 (N_13653,N_13070,N_13002);
or U13654 (N_13654,N_12875,N_13013);
nor U13655 (N_13655,N_12850,N_12924);
nand U13656 (N_13656,N_13577,N_13206);
xor U13657 (N_13657,N_13323,N_12989);
nand U13658 (N_13658,N_13347,N_13166);
nand U13659 (N_13659,N_13470,N_13116);
or U13660 (N_13660,N_13338,N_13451);
nand U13661 (N_13661,N_12854,N_13092);
and U13662 (N_13662,N_13006,N_13108);
nand U13663 (N_13663,N_13294,N_13267);
nand U13664 (N_13664,N_12860,N_13044);
nand U13665 (N_13665,N_13038,N_13150);
xnor U13666 (N_13666,N_13588,N_12899);
xor U13667 (N_13667,N_13063,N_13530);
or U13668 (N_13668,N_13421,N_13057);
or U13669 (N_13669,N_13117,N_13224);
or U13670 (N_13670,N_13480,N_13066);
or U13671 (N_13671,N_13028,N_13259);
xor U13672 (N_13672,N_12901,N_13400);
and U13673 (N_13673,N_13078,N_13441);
or U13674 (N_13674,N_13275,N_12879);
or U13675 (N_13675,N_13439,N_13274);
or U13676 (N_13676,N_13053,N_12914);
or U13677 (N_13677,N_13429,N_13292);
xor U13678 (N_13678,N_13186,N_13075);
and U13679 (N_13679,N_13250,N_13533);
or U13680 (N_13680,N_13273,N_13171);
and U13681 (N_13681,N_13074,N_12909);
or U13682 (N_13682,N_13388,N_13436);
and U13683 (N_13683,N_12847,N_13058);
nor U13684 (N_13684,N_12948,N_13401);
nor U13685 (N_13685,N_13404,N_12809);
or U13686 (N_13686,N_12967,N_13218);
or U13687 (N_13687,N_13184,N_13185);
nor U13688 (N_13688,N_13373,N_13362);
nand U13689 (N_13689,N_13094,N_13103);
and U13690 (N_13690,N_13328,N_12857);
and U13691 (N_13691,N_13268,N_13147);
nand U13692 (N_13692,N_12890,N_13559);
nor U13693 (N_13693,N_12983,N_12828);
and U13694 (N_13694,N_13146,N_13122);
xnor U13695 (N_13695,N_13357,N_13080);
nand U13696 (N_13696,N_13426,N_13468);
xor U13697 (N_13697,N_12876,N_13576);
nor U13698 (N_13698,N_13437,N_12824);
nand U13699 (N_13699,N_13138,N_13331);
nor U13700 (N_13700,N_13255,N_13004);
nand U13701 (N_13701,N_13285,N_13568);
and U13702 (N_13702,N_13288,N_12965);
nand U13703 (N_13703,N_13289,N_13159);
or U13704 (N_13704,N_13386,N_13354);
and U13705 (N_13705,N_13477,N_13350);
nand U13706 (N_13706,N_12974,N_13219);
xor U13707 (N_13707,N_13130,N_13544);
nand U13708 (N_13708,N_12814,N_13461);
nand U13709 (N_13709,N_13187,N_13047);
nand U13710 (N_13710,N_13356,N_12923);
or U13711 (N_13711,N_13235,N_12840);
nor U13712 (N_13712,N_12963,N_12918);
xor U13713 (N_13713,N_13179,N_13501);
nand U13714 (N_13714,N_13203,N_13052);
nor U13715 (N_13715,N_13113,N_13198);
xnor U13716 (N_13716,N_13346,N_13464);
or U13717 (N_13717,N_13230,N_13019);
nand U13718 (N_13718,N_13431,N_13241);
or U13719 (N_13719,N_13316,N_12900);
nand U13720 (N_13720,N_13180,N_13355);
nor U13721 (N_13721,N_12893,N_12816);
nand U13722 (N_13722,N_13286,N_12804);
or U13723 (N_13723,N_13353,N_13370);
nor U13724 (N_13724,N_13300,N_13278);
and U13725 (N_13725,N_13157,N_12855);
xor U13726 (N_13726,N_13478,N_12964);
and U13727 (N_13727,N_13160,N_12877);
and U13728 (N_13728,N_13391,N_12817);
or U13729 (N_13729,N_13418,N_13376);
or U13730 (N_13730,N_12881,N_13560);
nor U13731 (N_13731,N_12865,N_12966);
nand U13732 (N_13732,N_12815,N_12976);
xnor U13733 (N_13733,N_13022,N_13106);
nand U13734 (N_13734,N_13430,N_13597);
nand U13735 (N_13735,N_13265,N_12917);
or U13736 (N_13736,N_12906,N_12959);
nor U13737 (N_13737,N_13309,N_13008);
nor U13738 (N_13738,N_13483,N_12903);
and U13739 (N_13739,N_12954,N_13367);
and U13740 (N_13740,N_13296,N_13514);
or U13741 (N_13741,N_13155,N_13226);
and U13742 (N_13742,N_13405,N_13504);
xnor U13743 (N_13743,N_12980,N_13037);
nand U13744 (N_13744,N_13508,N_13010);
and U13745 (N_13745,N_13466,N_13459);
or U13746 (N_13746,N_13029,N_12921);
xnor U13747 (N_13747,N_13281,N_12950);
xnor U13748 (N_13748,N_12862,N_12997);
nor U13749 (N_13749,N_13064,N_13270);
or U13750 (N_13750,N_13543,N_13499);
and U13751 (N_13751,N_13313,N_13432);
nand U13752 (N_13752,N_13438,N_13287);
xnor U13753 (N_13753,N_13536,N_13455);
or U13754 (N_13754,N_13399,N_13120);
nor U13755 (N_13755,N_12984,N_13453);
and U13756 (N_13756,N_13060,N_12803);
xor U13757 (N_13757,N_13498,N_13083);
nor U13758 (N_13758,N_13377,N_13295);
nor U13759 (N_13759,N_13419,N_13079);
nand U13760 (N_13760,N_12888,N_13322);
xnor U13761 (N_13761,N_13382,N_13552);
nor U13762 (N_13762,N_13553,N_13088);
and U13763 (N_13763,N_13591,N_13191);
nor U13764 (N_13764,N_13345,N_13398);
nor U13765 (N_13765,N_12905,N_13087);
and U13766 (N_13766,N_13542,N_13111);
nor U13767 (N_13767,N_13546,N_13297);
nor U13768 (N_13768,N_12969,N_13566);
nand U13769 (N_13769,N_13086,N_12826);
or U13770 (N_13770,N_13360,N_13154);
or U13771 (N_13771,N_13372,N_13344);
xnor U13772 (N_13772,N_12833,N_12993);
nand U13773 (N_13773,N_13442,N_13590);
nand U13774 (N_13774,N_12821,N_13014);
or U13775 (N_13775,N_13409,N_12818);
xor U13776 (N_13776,N_12943,N_13460);
and U13777 (N_13777,N_13077,N_12834);
xor U13778 (N_13778,N_13465,N_13395);
nor U13779 (N_13779,N_13329,N_13516);
nor U13780 (N_13780,N_13374,N_12896);
and U13781 (N_13781,N_13489,N_13105);
nand U13782 (N_13782,N_13234,N_13476);
or U13783 (N_13783,N_12977,N_12856);
nor U13784 (N_13784,N_13522,N_12806);
or U13785 (N_13785,N_12869,N_13375);
and U13786 (N_13786,N_12904,N_13387);
nor U13787 (N_13787,N_13269,N_13448);
nand U13788 (N_13788,N_12907,N_13161);
nand U13789 (N_13789,N_13511,N_13450);
nor U13790 (N_13790,N_13023,N_13118);
xnor U13791 (N_13791,N_13126,N_13239);
or U13792 (N_13792,N_13482,N_13366);
nor U13793 (N_13793,N_12819,N_13561);
nor U13794 (N_13794,N_13535,N_12813);
nor U13795 (N_13795,N_13214,N_13512);
xnor U13796 (N_13796,N_12827,N_13558);
nor U13797 (N_13797,N_13121,N_12885);
nor U13798 (N_13798,N_12931,N_13557);
and U13799 (N_13799,N_13358,N_13193);
or U13800 (N_13800,N_13012,N_12928);
xnor U13801 (N_13801,N_12978,N_13564);
or U13802 (N_13802,N_13341,N_12942);
and U13803 (N_13803,N_13003,N_13035);
and U13804 (N_13804,N_13209,N_13379);
nand U13805 (N_13805,N_13484,N_13256);
nor U13806 (N_13806,N_13406,N_13582);
xnor U13807 (N_13807,N_13090,N_13061);
and U13808 (N_13808,N_13085,N_12820);
and U13809 (N_13809,N_12968,N_13479);
or U13810 (N_13810,N_13149,N_12990);
nand U13811 (N_13811,N_12933,N_13383);
xor U13812 (N_13812,N_13359,N_13237);
and U13813 (N_13813,N_13593,N_12971);
or U13814 (N_13814,N_13233,N_12870);
nand U13815 (N_13815,N_13332,N_13107);
nand U13816 (N_13816,N_13271,N_13208);
nand U13817 (N_13817,N_13524,N_13572);
xnor U13818 (N_13818,N_13139,N_13592);
or U13819 (N_13819,N_13005,N_13134);
or U13820 (N_13820,N_13320,N_12837);
nand U13821 (N_13821,N_13307,N_13110);
xnor U13822 (N_13822,N_13565,N_12823);
or U13823 (N_13823,N_13491,N_13410);
and U13824 (N_13824,N_12982,N_12864);
or U13825 (N_13825,N_13069,N_13142);
nand U13826 (N_13826,N_13051,N_12842);
nor U13827 (N_13827,N_13495,N_12958);
xor U13828 (N_13828,N_13452,N_12995);
nand U13829 (N_13829,N_12882,N_12892);
or U13830 (N_13830,N_13303,N_13033);
and U13831 (N_13831,N_13497,N_13097);
xnor U13832 (N_13832,N_12846,N_13407);
xor U13833 (N_13833,N_13277,N_12831);
and U13834 (N_13834,N_13579,N_13257);
and U13835 (N_13835,N_13318,N_13163);
nand U13836 (N_13836,N_13571,N_12853);
xor U13837 (N_13837,N_13236,N_13493);
and U13838 (N_13838,N_13587,N_13425);
or U13839 (N_13839,N_13081,N_13526);
nor U13840 (N_13840,N_13422,N_12940);
and U13841 (N_13841,N_13570,N_13128);
nand U13842 (N_13842,N_13473,N_13595);
and U13843 (N_13843,N_13127,N_13394);
nand U13844 (N_13844,N_13024,N_13260);
nand U13845 (N_13845,N_13585,N_13393);
or U13846 (N_13846,N_13471,N_13414);
nor U13847 (N_13847,N_12880,N_13469);
or U13848 (N_13848,N_13549,N_13299);
nor U13849 (N_13849,N_12895,N_13290);
xor U13850 (N_13850,N_13334,N_13055);
and U13851 (N_13851,N_13076,N_13433);
xor U13852 (N_13852,N_12946,N_12839);
xnor U13853 (N_13853,N_13098,N_13026);
nand U13854 (N_13854,N_13537,N_13056);
and U13855 (N_13855,N_13027,N_13046);
nor U13856 (N_13856,N_12897,N_13413);
nor U13857 (N_13857,N_13458,N_13594);
xor U13858 (N_13858,N_13474,N_13279);
and U13859 (N_13859,N_13040,N_13140);
and U13860 (N_13860,N_13443,N_13104);
or U13861 (N_13861,N_13365,N_13326);
and U13862 (N_13862,N_12911,N_13073);
nand U13863 (N_13863,N_13222,N_12867);
nor U13864 (N_13864,N_13183,N_12979);
nand U13865 (N_13865,N_13415,N_13444);
xor U13866 (N_13866,N_13178,N_12872);
xnor U13867 (N_13867,N_13282,N_13156);
xnor U13868 (N_13868,N_13449,N_13220);
or U13869 (N_13869,N_13135,N_12801);
and U13870 (N_13870,N_13584,N_12919);
nand U13871 (N_13871,N_13095,N_13308);
nor U13872 (N_13872,N_13252,N_13554);
nor U13873 (N_13873,N_13505,N_13071);
and U13874 (N_13874,N_13540,N_13563);
xnor U13875 (N_13875,N_13324,N_13330);
and U13876 (N_13876,N_13475,N_13050);
nor U13877 (N_13877,N_13315,N_13124);
or U13878 (N_13878,N_13333,N_13099);
and U13879 (N_13879,N_12962,N_13175);
and U13880 (N_13880,N_12830,N_13200);
and U13881 (N_13881,N_13068,N_12999);
and U13882 (N_13882,N_13337,N_12871);
and U13883 (N_13883,N_12972,N_13196);
xor U13884 (N_13884,N_13141,N_13131);
and U13885 (N_13885,N_13247,N_12912);
xnor U13886 (N_13886,N_12941,N_13136);
xor U13887 (N_13887,N_13447,N_13251);
or U13888 (N_13888,N_13575,N_13223);
and U13889 (N_13889,N_13336,N_13389);
and U13890 (N_13890,N_13164,N_13463);
nand U13891 (N_13891,N_12998,N_13291);
and U13892 (N_13892,N_13380,N_12947);
or U13893 (N_13893,N_13031,N_12938);
nand U13894 (N_13894,N_13132,N_13221);
or U13895 (N_13895,N_13598,N_12848);
and U13896 (N_13896,N_13195,N_13101);
nand U13897 (N_13897,N_12810,N_13551);
and U13898 (N_13898,N_13488,N_13392);
xor U13899 (N_13899,N_13262,N_12985);
or U13900 (N_13900,N_13240,N_12858);
and U13901 (N_13901,N_13494,N_13548);
xnor U13902 (N_13902,N_13174,N_13015);
xnor U13903 (N_13903,N_13462,N_13204);
and U13904 (N_13904,N_13062,N_13397);
nor U13905 (N_13905,N_13054,N_13518);
nor U13906 (N_13906,N_12925,N_12800);
nand U13907 (N_13907,N_13534,N_13412);
or U13908 (N_13908,N_13246,N_12929);
xor U13909 (N_13909,N_13148,N_13532);
xor U13910 (N_13910,N_13109,N_13283);
nand U13911 (N_13911,N_13496,N_13212);
nor U13912 (N_13912,N_13190,N_13596);
nor U13913 (N_13913,N_13245,N_13513);
nand U13914 (N_13914,N_12878,N_13306);
xor U13915 (N_13915,N_12932,N_12934);
and U13916 (N_13916,N_13114,N_13021);
nor U13917 (N_13917,N_12916,N_13181);
or U13918 (N_13918,N_13567,N_12956);
nand U13919 (N_13919,N_12949,N_13030);
or U13920 (N_13920,N_13228,N_12953);
and U13921 (N_13921,N_12859,N_13385);
nand U13922 (N_13922,N_13020,N_12944);
or U13923 (N_13923,N_13317,N_13172);
nor U13924 (N_13924,N_13467,N_13042);
nand U13925 (N_13925,N_12915,N_13363);
xor U13926 (N_13926,N_13416,N_13384);
and U13927 (N_13927,N_13280,N_13517);
xnor U13928 (N_13928,N_13169,N_13520);
or U13929 (N_13929,N_12894,N_12957);
and U13930 (N_13930,N_13569,N_13428);
and U13931 (N_13931,N_13202,N_13361);
nand U13932 (N_13932,N_12981,N_13266);
and U13933 (N_13933,N_13082,N_13529);
nand U13934 (N_13934,N_13225,N_12825);
nand U13935 (N_13935,N_12832,N_13472);
nor U13936 (N_13936,N_13025,N_12951);
nor U13937 (N_13937,N_12822,N_12908);
or U13938 (N_13938,N_13550,N_13381);
nor U13939 (N_13939,N_13177,N_13586);
and U13940 (N_13940,N_13509,N_13238);
and U13941 (N_13941,N_13589,N_13339);
or U13942 (N_13942,N_13152,N_13189);
nor U13943 (N_13943,N_13284,N_13417);
nor U13944 (N_13944,N_13199,N_13342);
xor U13945 (N_13945,N_13580,N_13538);
nand U13946 (N_13946,N_13205,N_13423);
nor U13947 (N_13947,N_13371,N_13119);
nand U13948 (N_13948,N_12952,N_13369);
xnor U13949 (N_13949,N_13072,N_13144);
nor U13950 (N_13950,N_13487,N_13378);
nand U13951 (N_13951,N_13457,N_12996);
nor U13952 (N_13952,N_13523,N_13305);
nor U13953 (N_13953,N_13216,N_12988);
nand U13954 (N_13954,N_13192,N_12829);
nand U13955 (N_13955,N_13574,N_13454);
and U13956 (N_13956,N_13424,N_13420);
nor U13957 (N_13957,N_13583,N_13261);
xor U13958 (N_13958,N_12960,N_12920);
nand U13959 (N_13959,N_13231,N_13519);
nor U13960 (N_13960,N_12887,N_13170);
or U13961 (N_13961,N_13067,N_13343);
xnor U13962 (N_13962,N_12927,N_13143);
nor U13963 (N_13963,N_13541,N_12841);
xor U13964 (N_13964,N_13017,N_13276);
nor U13965 (N_13965,N_13167,N_13293);
and U13966 (N_13966,N_13502,N_13253);
or U13967 (N_13967,N_13500,N_12849);
and U13968 (N_13968,N_13207,N_12930);
xnor U13969 (N_13969,N_13435,N_13327);
nor U13970 (N_13970,N_12863,N_12873);
nand U13971 (N_13971,N_13528,N_13434);
and U13972 (N_13972,N_12889,N_12886);
nand U13973 (N_13973,N_13000,N_12802);
nand U13974 (N_13974,N_12926,N_13302);
nor U13975 (N_13975,N_13001,N_12913);
nor U13976 (N_13976,N_13213,N_13490);
xor U13977 (N_13977,N_13506,N_13581);
and U13978 (N_13978,N_13182,N_13188);
xnor U13979 (N_13979,N_13112,N_12992);
xor U13980 (N_13980,N_13007,N_13573);
and U13981 (N_13981,N_13319,N_13194);
nand U13982 (N_13982,N_12868,N_13403);
and U13983 (N_13983,N_12937,N_13396);
nand U13984 (N_13984,N_13123,N_13503);
nand U13985 (N_13985,N_13272,N_13244);
or U13986 (N_13986,N_13151,N_13427);
or U13987 (N_13987,N_12874,N_12838);
nor U13988 (N_13988,N_13456,N_12994);
nor U13989 (N_13989,N_13264,N_13009);
or U13990 (N_13990,N_13032,N_13089);
nor U13991 (N_13991,N_13137,N_13539);
nand U13992 (N_13992,N_13578,N_13034);
xnor U13993 (N_13993,N_13197,N_12898);
nor U13994 (N_13994,N_13176,N_13440);
nor U13995 (N_13995,N_13525,N_13531);
and U13996 (N_13996,N_13304,N_13485);
nor U13997 (N_13997,N_13348,N_12970);
nor U13998 (N_13998,N_13217,N_12844);
nor U13999 (N_13999,N_13036,N_13492);
nand U14000 (N_14000,N_13226,N_13132);
and U14001 (N_14001,N_12905,N_12913);
xnor U14002 (N_14002,N_13217,N_13380);
and U14003 (N_14003,N_13031,N_12921);
and U14004 (N_14004,N_13238,N_13438);
nor U14005 (N_14005,N_13134,N_13193);
xor U14006 (N_14006,N_13463,N_13491);
nand U14007 (N_14007,N_13197,N_12941);
or U14008 (N_14008,N_13075,N_13164);
nand U14009 (N_14009,N_13567,N_12947);
xor U14010 (N_14010,N_13070,N_12937);
nor U14011 (N_14011,N_12882,N_13365);
or U14012 (N_14012,N_12942,N_13385);
or U14013 (N_14013,N_13304,N_13542);
and U14014 (N_14014,N_13168,N_13468);
nand U14015 (N_14015,N_13396,N_12907);
nor U14016 (N_14016,N_13299,N_13355);
nand U14017 (N_14017,N_13089,N_13579);
or U14018 (N_14018,N_13533,N_13045);
nand U14019 (N_14019,N_12820,N_13497);
or U14020 (N_14020,N_13325,N_13064);
and U14021 (N_14021,N_13065,N_13036);
nand U14022 (N_14022,N_12812,N_13220);
and U14023 (N_14023,N_13366,N_13569);
nor U14024 (N_14024,N_13297,N_12818);
xor U14025 (N_14025,N_13179,N_13478);
and U14026 (N_14026,N_13033,N_13421);
and U14027 (N_14027,N_13107,N_12840);
xnor U14028 (N_14028,N_12900,N_13001);
and U14029 (N_14029,N_13560,N_13116);
nand U14030 (N_14030,N_13006,N_13450);
nor U14031 (N_14031,N_13265,N_13558);
or U14032 (N_14032,N_13480,N_13343);
xor U14033 (N_14033,N_13144,N_13522);
or U14034 (N_14034,N_13506,N_13507);
xor U14035 (N_14035,N_12834,N_13031);
or U14036 (N_14036,N_13027,N_13262);
nor U14037 (N_14037,N_13366,N_12817);
nor U14038 (N_14038,N_12964,N_12801);
xnor U14039 (N_14039,N_13016,N_13377);
nor U14040 (N_14040,N_13259,N_13376);
and U14041 (N_14041,N_13088,N_12808);
nor U14042 (N_14042,N_13336,N_13016);
nor U14043 (N_14043,N_13124,N_13370);
nor U14044 (N_14044,N_12953,N_13529);
xnor U14045 (N_14045,N_13028,N_13555);
or U14046 (N_14046,N_13398,N_13287);
xnor U14047 (N_14047,N_13279,N_13136);
xor U14048 (N_14048,N_13490,N_12986);
nor U14049 (N_14049,N_12803,N_13087);
or U14050 (N_14050,N_13422,N_13494);
nand U14051 (N_14051,N_13295,N_13417);
nand U14052 (N_14052,N_13555,N_12905);
nor U14053 (N_14053,N_13283,N_13002);
and U14054 (N_14054,N_13086,N_13031);
nor U14055 (N_14055,N_13146,N_12846);
xor U14056 (N_14056,N_13155,N_12861);
nor U14057 (N_14057,N_12891,N_13489);
xnor U14058 (N_14058,N_12818,N_13312);
nor U14059 (N_14059,N_13366,N_13530);
nand U14060 (N_14060,N_13250,N_12885);
and U14061 (N_14061,N_13534,N_13361);
xor U14062 (N_14062,N_13069,N_13285);
nor U14063 (N_14063,N_13244,N_13315);
nand U14064 (N_14064,N_13525,N_13463);
nor U14065 (N_14065,N_13310,N_13001);
or U14066 (N_14066,N_12886,N_13454);
nor U14067 (N_14067,N_13197,N_13154);
or U14068 (N_14068,N_13086,N_12952);
nand U14069 (N_14069,N_13147,N_12837);
nor U14070 (N_14070,N_13085,N_12969);
and U14071 (N_14071,N_12901,N_13288);
or U14072 (N_14072,N_13079,N_13517);
or U14073 (N_14073,N_13063,N_13136);
and U14074 (N_14074,N_13597,N_12982);
or U14075 (N_14075,N_12978,N_13591);
nor U14076 (N_14076,N_13456,N_13247);
and U14077 (N_14077,N_13301,N_13222);
nor U14078 (N_14078,N_13026,N_12996);
nand U14079 (N_14079,N_13206,N_12814);
and U14080 (N_14080,N_13051,N_12913);
xnor U14081 (N_14081,N_12865,N_13357);
nand U14082 (N_14082,N_13077,N_13355);
and U14083 (N_14083,N_13007,N_13580);
nand U14084 (N_14084,N_13590,N_13513);
or U14085 (N_14085,N_12811,N_13097);
xor U14086 (N_14086,N_12912,N_12961);
nor U14087 (N_14087,N_12882,N_13271);
nor U14088 (N_14088,N_13420,N_12922);
nor U14089 (N_14089,N_13072,N_13126);
nor U14090 (N_14090,N_13588,N_12867);
nor U14091 (N_14091,N_13274,N_12984);
nor U14092 (N_14092,N_13322,N_13053);
or U14093 (N_14093,N_12847,N_13527);
or U14094 (N_14094,N_12997,N_13096);
and U14095 (N_14095,N_12920,N_13289);
nand U14096 (N_14096,N_13066,N_13504);
or U14097 (N_14097,N_13460,N_12966);
xnor U14098 (N_14098,N_13303,N_13525);
nor U14099 (N_14099,N_13443,N_13033);
nor U14100 (N_14100,N_13373,N_13493);
xnor U14101 (N_14101,N_13505,N_13221);
xnor U14102 (N_14102,N_12810,N_12836);
xor U14103 (N_14103,N_13374,N_12910);
or U14104 (N_14104,N_12838,N_13106);
nor U14105 (N_14105,N_13464,N_13569);
nor U14106 (N_14106,N_13381,N_12814);
xor U14107 (N_14107,N_13405,N_12854);
and U14108 (N_14108,N_13554,N_13491);
nor U14109 (N_14109,N_12814,N_13428);
or U14110 (N_14110,N_12903,N_12915);
and U14111 (N_14111,N_13032,N_13409);
xor U14112 (N_14112,N_13047,N_13372);
xor U14113 (N_14113,N_13379,N_13114);
xor U14114 (N_14114,N_13406,N_12981);
and U14115 (N_14115,N_13177,N_12974);
nand U14116 (N_14116,N_13468,N_13507);
nand U14117 (N_14117,N_13571,N_13193);
and U14118 (N_14118,N_12833,N_13356);
or U14119 (N_14119,N_13052,N_12938);
xor U14120 (N_14120,N_13141,N_12818);
and U14121 (N_14121,N_13243,N_13133);
or U14122 (N_14122,N_12830,N_13530);
nor U14123 (N_14123,N_13249,N_13331);
nor U14124 (N_14124,N_13474,N_12858);
nand U14125 (N_14125,N_13147,N_12843);
and U14126 (N_14126,N_13546,N_13034);
nand U14127 (N_14127,N_13090,N_13396);
and U14128 (N_14128,N_13342,N_13030);
xor U14129 (N_14129,N_13368,N_12999);
and U14130 (N_14130,N_12810,N_13190);
and U14131 (N_14131,N_13349,N_13142);
nor U14132 (N_14132,N_13405,N_13283);
nand U14133 (N_14133,N_13533,N_13453);
nor U14134 (N_14134,N_13247,N_12996);
nand U14135 (N_14135,N_12841,N_13491);
and U14136 (N_14136,N_12995,N_13494);
or U14137 (N_14137,N_12862,N_13524);
nand U14138 (N_14138,N_13329,N_12948);
and U14139 (N_14139,N_12878,N_13286);
and U14140 (N_14140,N_13060,N_13145);
and U14141 (N_14141,N_13153,N_12890);
xnor U14142 (N_14142,N_13550,N_13545);
xnor U14143 (N_14143,N_12916,N_13528);
nor U14144 (N_14144,N_13262,N_13471);
or U14145 (N_14145,N_13259,N_13065);
nor U14146 (N_14146,N_13451,N_13041);
and U14147 (N_14147,N_13297,N_13430);
nand U14148 (N_14148,N_13119,N_13053);
nor U14149 (N_14149,N_13123,N_13358);
xor U14150 (N_14150,N_13518,N_13447);
xnor U14151 (N_14151,N_13061,N_13402);
nor U14152 (N_14152,N_13177,N_13479);
nand U14153 (N_14153,N_13401,N_13361);
xnor U14154 (N_14154,N_13596,N_13008);
nor U14155 (N_14155,N_13389,N_13415);
nand U14156 (N_14156,N_13572,N_13320);
or U14157 (N_14157,N_13335,N_12810);
nand U14158 (N_14158,N_13594,N_13246);
or U14159 (N_14159,N_12986,N_13316);
nand U14160 (N_14160,N_12821,N_12895);
or U14161 (N_14161,N_12861,N_13021);
and U14162 (N_14162,N_13085,N_13424);
xnor U14163 (N_14163,N_13447,N_13088);
or U14164 (N_14164,N_12875,N_13043);
nor U14165 (N_14165,N_12849,N_13373);
nand U14166 (N_14166,N_13251,N_13422);
and U14167 (N_14167,N_13378,N_13043);
nand U14168 (N_14168,N_13563,N_13198);
or U14169 (N_14169,N_12830,N_12911);
nor U14170 (N_14170,N_13055,N_13423);
and U14171 (N_14171,N_13568,N_13458);
xnor U14172 (N_14172,N_13520,N_12905);
nor U14173 (N_14173,N_13135,N_13386);
nand U14174 (N_14174,N_13389,N_13458);
or U14175 (N_14175,N_12991,N_13102);
xnor U14176 (N_14176,N_13422,N_12972);
nand U14177 (N_14177,N_13063,N_13004);
and U14178 (N_14178,N_13385,N_13125);
or U14179 (N_14179,N_13300,N_13260);
or U14180 (N_14180,N_13325,N_12880);
xnor U14181 (N_14181,N_13373,N_12978);
and U14182 (N_14182,N_12836,N_12913);
or U14183 (N_14183,N_13134,N_12861);
nor U14184 (N_14184,N_13349,N_12867);
xor U14185 (N_14185,N_13440,N_13478);
nor U14186 (N_14186,N_13521,N_13418);
nand U14187 (N_14187,N_13393,N_12906);
xor U14188 (N_14188,N_13082,N_12896);
and U14189 (N_14189,N_13179,N_13152);
nor U14190 (N_14190,N_13242,N_13397);
and U14191 (N_14191,N_13012,N_12978);
or U14192 (N_14192,N_13536,N_13208);
and U14193 (N_14193,N_13123,N_13162);
nor U14194 (N_14194,N_12868,N_13390);
or U14195 (N_14195,N_13547,N_13218);
nor U14196 (N_14196,N_13181,N_13117);
and U14197 (N_14197,N_13307,N_12871);
nand U14198 (N_14198,N_12840,N_12918);
nor U14199 (N_14199,N_13389,N_12975);
and U14200 (N_14200,N_13224,N_13006);
and U14201 (N_14201,N_13153,N_13425);
nor U14202 (N_14202,N_13160,N_13123);
xnor U14203 (N_14203,N_13075,N_13163);
or U14204 (N_14204,N_12887,N_13408);
or U14205 (N_14205,N_13218,N_13462);
and U14206 (N_14206,N_13466,N_12932);
or U14207 (N_14207,N_13087,N_13231);
or U14208 (N_14208,N_13548,N_13041);
and U14209 (N_14209,N_12953,N_12997);
nand U14210 (N_14210,N_12883,N_13523);
nor U14211 (N_14211,N_13140,N_12836);
nor U14212 (N_14212,N_13348,N_13192);
nand U14213 (N_14213,N_12998,N_12931);
nand U14214 (N_14214,N_13441,N_13083);
xnor U14215 (N_14215,N_13019,N_13114);
or U14216 (N_14216,N_13053,N_12993);
or U14217 (N_14217,N_13052,N_13231);
xor U14218 (N_14218,N_12841,N_13363);
nor U14219 (N_14219,N_13398,N_13532);
nand U14220 (N_14220,N_13422,N_13536);
or U14221 (N_14221,N_12941,N_13429);
and U14222 (N_14222,N_12845,N_12956);
or U14223 (N_14223,N_12935,N_13197);
or U14224 (N_14224,N_13568,N_13263);
and U14225 (N_14225,N_13476,N_13490);
or U14226 (N_14226,N_13519,N_13359);
and U14227 (N_14227,N_12981,N_13017);
xnor U14228 (N_14228,N_13439,N_13089);
nor U14229 (N_14229,N_12901,N_13478);
or U14230 (N_14230,N_13554,N_13207);
nand U14231 (N_14231,N_13137,N_13192);
nand U14232 (N_14232,N_13130,N_13381);
and U14233 (N_14233,N_13256,N_13521);
and U14234 (N_14234,N_13124,N_12940);
and U14235 (N_14235,N_13206,N_13193);
xnor U14236 (N_14236,N_13484,N_13118);
or U14237 (N_14237,N_12996,N_13523);
or U14238 (N_14238,N_12846,N_13079);
nand U14239 (N_14239,N_12933,N_13212);
and U14240 (N_14240,N_13207,N_13386);
nor U14241 (N_14241,N_13377,N_12968);
and U14242 (N_14242,N_13371,N_13049);
xor U14243 (N_14243,N_12807,N_13409);
nand U14244 (N_14244,N_13281,N_13524);
and U14245 (N_14245,N_13524,N_13287);
xnor U14246 (N_14246,N_13409,N_12828);
and U14247 (N_14247,N_12814,N_13488);
and U14248 (N_14248,N_12912,N_13571);
nor U14249 (N_14249,N_13381,N_13271);
nor U14250 (N_14250,N_13389,N_13285);
and U14251 (N_14251,N_13140,N_13117);
and U14252 (N_14252,N_13276,N_13231);
xnor U14253 (N_14253,N_13385,N_13398);
xor U14254 (N_14254,N_13392,N_13053);
xnor U14255 (N_14255,N_13281,N_12892);
nor U14256 (N_14256,N_13374,N_12992);
or U14257 (N_14257,N_13567,N_13520);
xor U14258 (N_14258,N_12939,N_13158);
xor U14259 (N_14259,N_13214,N_12854);
nor U14260 (N_14260,N_13155,N_13515);
nand U14261 (N_14261,N_13013,N_12982);
or U14262 (N_14262,N_13554,N_13524);
xnor U14263 (N_14263,N_13426,N_13533);
nand U14264 (N_14264,N_13125,N_13384);
nor U14265 (N_14265,N_13097,N_13460);
xor U14266 (N_14266,N_12851,N_13069);
nand U14267 (N_14267,N_13068,N_12994);
and U14268 (N_14268,N_12849,N_12831);
xnor U14269 (N_14269,N_13592,N_13330);
nand U14270 (N_14270,N_13404,N_13279);
nor U14271 (N_14271,N_12811,N_13548);
nand U14272 (N_14272,N_13357,N_13217);
xor U14273 (N_14273,N_13433,N_12945);
xor U14274 (N_14274,N_13209,N_12897);
nand U14275 (N_14275,N_12964,N_13011);
xnor U14276 (N_14276,N_13375,N_13176);
and U14277 (N_14277,N_13130,N_13328);
or U14278 (N_14278,N_12857,N_13282);
nor U14279 (N_14279,N_13264,N_13212);
nand U14280 (N_14280,N_13024,N_13577);
xor U14281 (N_14281,N_13343,N_12866);
or U14282 (N_14282,N_13372,N_12997);
and U14283 (N_14283,N_13552,N_13016);
xnor U14284 (N_14284,N_12931,N_13005);
nor U14285 (N_14285,N_13332,N_13528);
or U14286 (N_14286,N_12928,N_13207);
nand U14287 (N_14287,N_13436,N_12985);
or U14288 (N_14288,N_13445,N_13366);
or U14289 (N_14289,N_12952,N_13145);
or U14290 (N_14290,N_13065,N_12895);
nand U14291 (N_14291,N_13221,N_12840);
xnor U14292 (N_14292,N_13501,N_13332);
nand U14293 (N_14293,N_12881,N_13010);
nor U14294 (N_14294,N_13125,N_12887);
xnor U14295 (N_14295,N_12846,N_13060);
and U14296 (N_14296,N_13567,N_13144);
or U14297 (N_14297,N_13400,N_12885);
and U14298 (N_14298,N_13442,N_13200);
nor U14299 (N_14299,N_12827,N_12971);
and U14300 (N_14300,N_12888,N_13370);
xnor U14301 (N_14301,N_12958,N_13086);
xor U14302 (N_14302,N_13308,N_13350);
or U14303 (N_14303,N_13242,N_13529);
and U14304 (N_14304,N_13453,N_13296);
xor U14305 (N_14305,N_13033,N_13202);
xnor U14306 (N_14306,N_13231,N_12910);
and U14307 (N_14307,N_13395,N_12995);
or U14308 (N_14308,N_13415,N_13115);
nor U14309 (N_14309,N_13506,N_13144);
or U14310 (N_14310,N_13116,N_13361);
nor U14311 (N_14311,N_13382,N_13365);
nor U14312 (N_14312,N_12910,N_13068);
and U14313 (N_14313,N_13119,N_13527);
or U14314 (N_14314,N_13442,N_12886);
xnor U14315 (N_14315,N_13161,N_13542);
and U14316 (N_14316,N_12858,N_13304);
or U14317 (N_14317,N_13037,N_13129);
or U14318 (N_14318,N_13260,N_12929);
and U14319 (N_14319,N_13219,N_13205);
and U14320 (N_14320,N_13211,N_13104);
or U14321 (N_14321,N_13179,N_12969);
nand U14322 (N_14322,N_13526,N_13104);
nor U14323 (N_14323,N_13115,N_12942);
and U14324 (N_14324,N_13213,N_12846);
nand U14325 (N_14325,N_13121,N_13536);
or U14326 (N_14326,N_13272,N_13329);
and U14327 (N_14327,N_13444,N_13321);
xor U14328 (N_14328,N_13199,N_13422);
or U14329 (N_14329,N_13140,N_13192);
or U14330 (N_14330,N_13570,N_12806);
nor U14331 (N_14331,N_12891,N_13004);
and U14332 (N_14332,N_13545,N_13568);
nor U14333 (N_14333,N_13010,N_12808);
or U14334 (N_14334,N_12834,N_13297);
and U14335 (N_14335,N_13314,N_13590);
nand U14336 (N_14336,N_13590,N_12936);
xnor U14337 (N_14337,N_13582,N_13283);
nor U14338 (N_14338,N_13372,N_13159);
and U14339 (N_14339,N_13058,N_13083);
nand U14340 (N_14340,N_13034,N_13403);
and U14341 (N_14341,N_13424,N_13145);
nand U14342 (N_14342,N_12801,N_13485);
nand U14343 (N_14343,N_13443,N_13204);
nand U14344 (N_14344,N_13514,N_13055);
nor U14345 (N_14345,N_13486,N_13190);
xnor U14346 (N_14346,N_13183,N_12825);
xor U14347 (N_14347,N_13194,N_13367);
and U14348 (N_14348,N_13457,N_13176);
nand U14349 (N_14349,N_13073,N_13028);
and U14350 (N_14350,N_13352,N_13486);
and U14351 (N_14351,N_13293,N_13365);
xor U14352 (N_14352,N_13532,N_13392);
or U14353 (N_14353,N_13094,N_13156);
nor U14354 (N_14354,N_13176,N_13307);
nand U14355 (N_14355,N_12825,N_13522);
or U14356 (N_14356,N_13340,N_13042);
nand U14357 (N_14357,N_13292,N_13052);
and U14358 (N_14358,N_13481,N_12815);
nor U14359 (N_14359,N_13024,N_13459);
nand U14360 (N_14360,N_13091,N_13385);
or U14361 (N_14361,N_13565,N_13183);
nor U14362 (N_14362,N_12966,N_12941);
nand U14363 (N_14363,N_13030,N_13173);
nor U14364 (N_14364,N_12822,N_13564);
xnor U14365 (N_14365,N_12890,N_12998);
nor U14366 (N_14366,N_12879,N_12959);
xor U14367 (N_14367,N_13086,N_13313);
or U14368 (N_14368,N_12855,N_13386);
xor U14369 (N_14369,N_13445,N_12951);
or U14370 (N_14370,N_13509,N_13252);
or U14371 (N_14371,N_13018,N_13347);
nor U14372 (N_14372,N_13079,N_13130);
nor U14373 (N_14373,N_13470,N_13325);
nor U14374 (N_14374,N_13418,N_13146);
and U14375 (N_14375,N_13245,N_13407);
xnor U14376 (N_14376,N_13251,N_12890);
xor U14377 (N_14377,N_13374,N_13320);
nand U14378 (N_14378,N_13442,N_13282);
or U14379 (N_14379,N_13223,N_13453);
and U14380 (N_14380,N_13579,N_12851);
and U14381 (N_14381,N_12902,N_13221);
nor U14382 (N_14382,N_13472,N_13456);
xor U14383 (N_14383,N_13135,N_13138);
and U14384 (N_14384,N_13067,N_13174);
nand U14385 (N_14385,N_12881,N_13381);
nor U14386 (N_14386,N_13214,N_13398);
and U14387 (N_14387,N_13209,N_13169);
or U14388 (N_14388,N_13569,N_13057);
and U14389 (N_14389,N_13541,N_13164);
nand U14390 (N_14390,N_13152,N_12830);
or U14391 (N_14391,N_13520,N_12997);
nand U14392 (N_14392,N_13223,N_12826);
or U14393 (N_14393,N_13585,N_13419);
nor U14394 (N_14394,N_13368,N_13553);
nor U14395 (N_14395,N_12835,N_13392);
and U14396 (N_14396,N_13173,N_12851);
nor U14397 (N_14397,N_13586,N_13316);
nand U14398 (N_14398,N_13430,N_13177);
xor U14399 (N_14399,N_13503,N_12930);
and U14400 (N_14400,N_14348,N_13662);
nor U14401 (N_14401,N_14105,N_14259);
or U14402 (N_14402,N_13800,N_14099);
nand U14403 (N_14403,N_14014,N_13888);
nand U14404 (N_14404,N_14016,N_13901);
or U14405 (N_14405,N_13826,N_13953);
and U14406 (N_14406,N_13728,N_14243);
nand U14407 (N_14407,N_14296,N_14080);
xnor U14408 (N_14408,N_14366,N_14053);
nor U14409 (N_14409,N_14361,N_13945);
nor U14410 (N_14410,N_13988,N_13760);
and U14411 (N_14411,N_14026,N_13978);
or U14412 (N_14412,N_14077,N_14272);
nand U14413 (N_14413,N_14204,N_13845);
xnor U14414 (N_14414,N_13610,N_14322);
and U14415 (N_14415,N_14205,N_14142);
and U14416 (N_14416,N_13828,N_13984);
and U14417 (N_14417,N_13714,N_13718);
xnor U14418 (N_14418,N_13770,N_13995);
and U14419 (N_14419,N_13708,N_14254);
or U14420 (N_14420,N_13773,N_13885);
xor U14421 (N_14421,N_14223,N_14236);
and U14422 (N_14422,N_14240,N_13739);
nand U14423 (N_14423,N_13791,N_13874);
nand U14424 (N_14424,N_13702,N_13906);
and U14425 (N_14425,N_13759,N_14028);
xnor U14426 (N_14426,N_14210,N_13858);
nor U14427 (N_14427,N_13848,N_14244);
or U14428 (N_14428,N_14226,N_13705);
or U14429 (N_14429,N_14275,N_13694);
or U14430 (N_14430,N_14224,N_14112);
and U14431 (N_14431,N_14397,N_13623);
nor U14432 (N_14432,N_13713,N_14158);
and U14433 (N_14433,N_13833,N_13651);
nor U14434 (N_14434,N_13832,N_14034);
or U14435 (N_14435,N_13980,N_14008);
and U14436 (N_14436,N_14374,N_13789);
and U14437 (N_14437,N_14277,N_13947);
nand U14438 (N_14438,N_14357,N_14081);
nand U14439 (N_14439,N_13682,N_13799);
or U14440 (N_14440,N_14285,N_13747);
xnor U14441 (N_14441,N_14358,N_13745);
nor U14442 (N_14442,N_13639,N_14246);
nor U14443 (N_14443,N_14027,N_13740);
xnor U14444 (N_14444,N_13814,N_14315);
and U14445 (N_14445,N_13626,N_13923);
xor U14446 (N_14446,N_14117,N_14318);
xor U14447 (N_14447,N_13765,N_13805);
xor U14448 (N_14448,N_14006,N_13824);
and U14449 (N_14449,N_14376,N_14161);
and U14450 (N_14450,N_14326,N_14089);
or U14451 (N_14451,N_14106,N_14237);
nor U14452 (N_14452,N_14169,N_13783);
nand U14453 (N_14453,N_13924,N_14068);
and U14454 (N_14454,N_14183,N_14368);
or U14455 (N_14455,N_13998,N_13720);
nand U14456 (N_14456,N_14151,N_14005);
or U14457 (N_14457,N_14062,N_13693);
nand U14458 (N_14458,N_13683,N_14010);
xnor U14459 (N_14459,N_14302,N_14152);
and U14460 (N_14460,N_14353,N_14156);
xnor U14461 (N_14461,N_13959,N_14058);
and U14462 (N_14462,N_13719,N_14121);
and U14463 (N_14463,N_14104,N_13798);
and U14464 (N_14464,N_14371,N_13827);
xnor U14465 (N_14465,N_14095,N_14346);
nor U14466 (N_14466,N_13685,N_14188);
nor U14467 (N_14467,N_13853,N_14388);
or U14468 (N_14468,N_14198,N_13608);
or U14469 (N_14469,N_13734,N_13815);
xor U14470 (N_14470,N_14050,N_13601);
nor U14471 (N_14471,N_13878,N_13629);
or U14472 (N_14472,N_13939,N_14291);
xnor U14473 (N_14473,N_14163,N_13768);
nor U14474 (N_14474,N_13616,N_13876);
nor U14475 (N_14475,N_14092,N_14234);
and U14476 (N_14476,N_14219,N_14263);
and U14477 (N_14477,N_14343,N_14056);
nand U14478 (N_14478,N_13696,N_14057);
nor U14479 (N_14479,N_14147,N_13905);
nand U14480 (N_14480,N_14093,N_14300);
xor U14481 (N_14481,N_14290,N_14137);
nand U14482 (N_14482,N_14076,N_13919);
xor U14483 (N_14483,N_14308,N_13709);
nor U14484 (N_14484,N_14084,N_13836);
and U14485 (N_14485,N_14177,N_14394);
xnor U14486 (N_14486,N_14009,N_14019);
or U14487 (N_14487,N_14088,N_14136);
nor U14488 (N_14488,N_13717,N_13668);
or U14489 (N_14489,N_14323,N_14030);
and U14490 (N_14490,N_13781,N_14230);
nor U14491 (N_14491,N_13870,N_14091);
nor U14492 (N_14492,N_14222,N_14273);
nor U14493 (N_14493,N_13687,N_14004);
and U14494 (N_14494,N_14317,N_14135);
xnor U14495 (N_14495,N_14072,N_13964);
nor U14496 (N_14496,N_13890,N_13809);
xnor U14497 (N_14497,N_13692,N_14020);
xnor U14498 (N_14498,N_13674,N_13772);
nand U14499 (N_14499,N_14002,N_14231);
xnor U14500 (N_14500,N_14003,N_14113);
xnor U14501 (N_14501,N_13859,N_14297);
or U14502 (N_14502,N_14261,N_14286);
xnor U14503 (N_14503,N_14209,N_14118);
and U14504 (N_14504,N_13787,N_14383);
or U14505 (N_14505,N_13647,N_14214);
or U14506 (N_14506,N_13981,N_13999);
and U14507 (N_14507,N_13819,N_13864);
or U14508 (N_14508,N_13688,N_14036);
or U14509 (N_14509,N_14220,N_14375);
or U14510 (N_14510,N_13695,N_14110);
nand U14511 (N_14511,N_13985,N_14289);
nand U14512 (N_14512,N_14173,N_13806);
or U14513 (N_14513,N_14085,N_13899);
nand U14514 (N_14514,N_13605,N_14190);
nand U14515 (N_14515,N_14398,N_14011);
and U14516 (N_14516,N_13612,N_14039);
or U14517 (N_14517,N_13837,N_13942);
and U14518 (N_14518,N_14241,N_13821);
xor U14519 (N_14519,N_13676,N_14215);
nor U14520 (N_14520,N_13993,N_14201);
or U14521 (N_14521,N_14377,N_14100);
or U14522 (N_14522,N_13755,N_13842);
nor U14523 (N_14523,N_13996,N_14166);
and U14524 (N_14524,N_14330,N_13897);
nor U14525 (N_14525,N_14359,N_13810);
and U14526 (N_14526,N_14124,N_13710);
nand U14527 (N_14527,N_13977,N_14086);
or U14528 (N_14528,N_13929,N_14387);
and U14529 (N_14529,N_14310,N_13927);
or U14530 (N_14530,N_13743,N_13788);
or U14531 (N_14531,N_13991,N_13746);
or U14532 (N_14532,N_14336,N_13920);
nor U14533 (N_14533,N_14252,N_14208);
and U14534 (N_14534,N_13603,N_13944);
nand U14535 (N_14535,N_14265,N_14054);
nor U14536 (N_14536,N_13829,N_14172);
nor U14537 (N_14537,N_14340,N_13952);
nand U14538 (N_14538,N_13872,N_13856);
and U14539 (N_14539,N_13949,N_14024);
or U14540 (N_14540,N_13830,N_13635);
and U14541 (N_14541,N_13754,N_14157);
nand U14542 (N_14542,N_13753,N_13887);
or U14543 (N_14543,N_13970,N_14070);
nor U14544 (N_14544,N_13611,N_14127);
and U14545 (N_14545,N_13666,N_14335);
nand U14546 (N_14546,N_13792,N_13802);
xnor U14547 (N_14547,N_13844,N_13911);
and U14548 (N_14548,N_13721,N_14149);
nor U14549 (N_14549,N_14128,N_14354);
xor U14550 (N_14550,N_14074,N_14351);
nand U14551 (N_14551,N_13646,N_14046);
and U14552 (N_14552,N_14212,N_13909);
xnor U14553 (N_14553,N_13699,N_14203);
xnor U14554 (N_14554,N_13777,N_13780);
and U14555 (N_14555,N_14350,N_14242);
xnor U14556 (N_14556,N_14094,N_14271);
nor U14557 (N_14557,N_14262,N_14369);
and U14558 (N_14558,N_14274,N_13868);
nor U14559 (N_14559,N_14170,N_13922);
xor U14560 (N_14560,N_13618,N_14162);
nand U14561 (N_14561,N_13613,N_14258);
xor U14562 (N_14562,N_13757,N_13994);
and U14563 (N_14563,N_14281,N_14116);
xnor U14564 (N_14564,N_14111,N_14207);
and U14565 (N_14565,N_14373,N_13982);
xnor U14566 (N_14566,N_13643,N_14276);
nand U14567 (N_14567,N_13684,N_13895);
nand U14568 (N_14568,N_13931,N_13748);
nor U14569 (N_14569,N_14256,N_13936);
nand U14570 (N_14570,N_14144,N_14123);
or U14571 (N_14571,N_13751,N_14356);
nor U14572 (N_14572,N_13937,N_14052);
nor U14573 (N_14573,N_13658,N_13889);
or U14574 (N_14574,N_13741,N_13659);
nor U14575 (N_14575,N_13989,N_14381);
xor U14576 (N_14576,N_13934,N_14245);
nor U14577 (N_14577,N_13904,N_14060);
nor U14578 (N_14578,N_13678,N_14066);
nand U14579 (N_14579,N_14329,N_14097);
or U14580 (N_14580,N_13722,N_14159);
nand U14581 (N_14581,N_13804,N_13776);
or U14582 (N_14582,N_13943,N_13892);
nand U14583 (N_14583,N_13869,N_14293);
xnor U14584 (N_14584,N_14269,N_13910);
and U14585 (N_14585,N_13915,N_13912);
and U14586 (N_14586,N_13928,N_14248);
nor U14587 (N_14587,N_14197,N_13862);
or U14588 (N_14588,N_13778,N_13767);
or U14589 (N_14589,N_14143,N_14055);
or U14590 (N_14590,N_13818,N_13762);
nor U14591 (N_14591,N_13958,N_13846);
or U14592 (N_14592,N_14328,N_14184);
xnor U14593 (N_14593,N_13997,N_14031);
nand U14594 (N_14594,N_14264,N_13961);
and U14595 (N_14595,N_14185,N_14141);
nand U14596 (N_14596,N_14392,N_14041);
and U14597 (N_14597,N_13983,N_13744);
nand U14598 (N_14598,N_13973,N_14165);
and U14599 (N_14599,N_13992,N_13786);
xor U14600 (N_14600,N_13893,N_13725);
xnor U14601 (N_14601,N_14306,N_13811);
nand U14602 (N_14602,N_14362,N_13664);
and U14603 (N_14603,N_13737,N_13667);
or U14604 (N_14604,N_14253,N_13896);
nor U14605 (N_14605,N_13921,N_13794);
nand U14606 (N_14606,N_14313,N_14364);
nand U14607 (N_14607,N_13817,N_13816);
or U14608 (N_14608,N_14206,N_13614);
or U14609 (N_14609,N_14319,N_14217);
xor U14610 (N_14610,N_14191,N_13857);
nor U14611 (N_14611,N_13948,N_13752);
nand U14612 (N_14612,N_14193,N_14033);
and U14613 (N_14613,N_13609,N_13913);
nand U14614 (N_14614,N_13839,N_14139);
nor U14615 (N_14615,N_13962,N_13677);
xnor U14616 (N_14616,N_14301,N_13966);
nor U14617 (N_14617,N_13951,N_13680);
xor U14618 (N_14618,N_14181,N_13715);
xnor U14619 (N_14619,N_13628,N_14071);
and U14620 (N_14620,N_13831,N_13903);
xor U14621 (N_14621,N_13935,N_14187);
or U14622 (N_14622,N_13974,N_14042);
nor U14623 (N_14623,N_14233,N_13823);
nor U14624 (N_14624,N_14132,N_14096);
and U14625 (N_14625,N_14090,N_13665);
nor U14626 (N_14626,N_13622,N_14101);
and U14627 (N_14627,N_13813,N_13729);
or U14628 (N_14628,N_14114,N_13712);
nand U14629 (N_14629,N_13670,N_14321);
or U14630 (N_14630,N_13672,N_14180);
xor U14631 (N_14631,N_13812,N_13960);
nand U14632 (N_14632,N_13671,N_14316);
nor U14633 (N_14633,N_14038,N_13979);
nor U14634 (N_14634,N_13891,N_14001);
and U14635 (N_14635,N_14171,N_14379);
nand U14636 (N_14636,N_14320,N_13652);
and U14637 (N_14637,N_14102,N_13916);
and U14638 (N_14638,N_13607,N_13645);
or U14639 (N_14639,N_13766,N_14078);
and U14640 (N_14640,N_13758,N_14138);
or U14641 (N_14641,N_13775,N_13849);
xor U14642 (N_14642,N_13669,N_14238);
and U14643 (N_14643,N_13843,N_14047);
nor U14644 (N_14644,N_13782,N_14098);
nor U14645 (N_14645,N_14126,N_13764);
or U14646 (N_14646,N_13852,N_13884);
xnor U14647 (N_14647,N_14225,N_14294);
nand U14648 (N_14648,N_14017,N_14334);
and U14649 (N_14649,N_14349,N_13797);
nand U14650 (N_14650,N_14043,N_14247);
xor U14651 (N_14651,N_14389,N_14202);
nor U14652 (N_14652,N_14342,N_14292);
and U14653 (N_14653,N_13617,N_14109);
xor U14654 (N_14654,N_14048,N_14153);
nand U14655 (N_14655,N_13624,N_13908);
nand U14656 (N_14656,N_14175,N_14295);
nand U14657 (N_14657,N_14051,N_14179);
or U14658 (N_14658,N_13679,N_13855);
and U14659 (N_14659,N_14073,N_14199);
nand U14660 (N_14660,N_14399,N_13971);
and U14661 (N_14661,N_13986,N_14160);
xor U14662 (N_14662,N_13825,N_13793);
or U14663 (N_14663,N_13946,N_13838);
xor U14664 (N_14664,N_14324,N_14069);
and U14665 (N_14665,N_14395,N_14391);
nand U14666 (N_14666,N_13606,N_14176);
and U14667 (N_14667,N_14327,N_14079);
nand U14668 (N_14668,N_13653,N_14385);
xor U14669 (N_14669,N_14154,N_14363);
or U14670 (N_14670,N_13881,N_14115);
and U14671 (N_14671,N_13726,N_13871);
and U14672 (N_14672,N_14287,N_13763);
or U14673 (N_14673,N_13630,N_14186);
nand U14674 (N_14674,N_13681,N_14122);
and U14675 (N_14675,N_14390,N_13663);
nand U14676 (N_14676,N_14174,N_14284);
xor U14677 (N_14677,N_14338,N_14229);
and U14678 (N_14678,N_13987,N_13956);
and U14679 (N_14679,N_13615,N_13650);
and U14680 (N_14680,N_13940,N_14333);
and U14681 (N_14681,N_13769,N_13861);
xnor U14682 (N_14682,N_13865,N_14299);
xor U14683 (N_14683,N_14396,N_13867);
or U14684 (N_14684,N_13941,N_14372);
nand U14685 (N_14685,N_13882,N_13883);
nor U14686 (N_14686,N_14148,N_14133);
or U14687 (N_14687,N_14305,N_14270);
xor U14688 (N_14688,N_14213,N_13847);
nand U14689 (N_14689,N_13689,N_14064);
nor U14690 (N_14690,N_13627,N_13634);
and U14691 (N_14691,N_14192,N_14182);
nand U14692 (N_14692,N_13785,N_14119);
and U14693 (N_14693,N_13727,N_14007);
and U14694 (N_14694,N_13700,N_14083);
xor U14695 (N_14695,N_14022,N_14125);
nand U14696 (N_14696,N_14018,N_13620);
nand U14697 (N_14697,N_14380,N_14279);
xor U14698 (N_14698,N_14013,N_13841);
and U14699 (N_14699,N_14061,N_13854);
nor U14700 (N_14700,N_13736,N_13673);
or U14701 (N_14701,N_13796,N_13733);
nand U14702 (N_14702,N_14168,N_14251);
xor U14703 (N_14703,N_14065,N_14370);
xnor U14704 (N_14704,N_14035,N_14129);
and U14705 (N_14705,N_13863,N_14140);
xnor U14706 (N_14706,N_13600,N_14393);
nor U14707 (N_14707,N_14345,N_14307);
and U14708 (N_14708,N_13918,N_13976);
or U14709 (N_14709,N_13771,N_13732);
nand U14710 (N_14710,N_13724,N_14260);
nor U14711 (N_14711,N_13808,N_13648);
and U14712 (N_14712,N_14312,N_13950);
nand U14713 (N_14713,N_13990,N_13749);
nand U14714 (N_14714,N_14355,N_13917);
nor U14715 (N_14715,N_13698,N_13660);
nor U14716 (N_14716,N_13784,N_13822);
nand U14717 (N_14717,N_14282,N_14195);
and U14718 (N_14718,N_14032,N_14025);
xor U14719 (N_14719,N_13902,N_13914);
nand U14720 (N_14720,N_13779,N_14365);
nor U14721 (N_14721,N_13691,N_14146);
nand U14722 (N_14722,N_13965,N_13835);
xnor U14723 (N_14723,N_14044,N_13619);
nand U14724 (N_14724,N_14200,N_14029);
nor U14725 (N_14725,N_14167,N_14131);
xnor U14726 (N_14726,N_14255,N_14309);
nor U14727 (N_14727,N_14063,N_13774);
nor U14728 (N_14728,N_13790,N_14332);
or U14729 (N_14729,N_13969,N_14367);
nor U14730 (N_14730,N_13640,N_14164);
and U14731 (N_14731,N_13750,N_13731);
nand U14732 (N_14732,N_13641,N_13898);
and U14733 (N_14733,N_13735,N_13850);
or U14734 (N_14734,N_14107,N_13707);
nor U14735 (N_14735,N_14347,N_13900);
xor U14736 (N_14736,N_14303,N_14023);
and U14737 (N_14737,N_14045,N_13654);
nand U14738 (N_14738,N_13873,N_13834);
nand U14739 (N_14739,N_13840,N_14268);
and U14740 (N_14740,N_14232,N_14049);
and U14741 (N_14741,N_13742,N_14216);
and U14742 (N_14742,N_13851,N_14103);
or U14743 (N_14743,N_14134,N_14304);
or U14744 (N_14744,N_13636,N_14130);
xnor U14745 (N_14745,N_14194,N_14314);
nand U14746 (N_14746,N_13756,N_14384);
and U14747 (N_14747,N_13690,N_13801);
xor U14748 (N_14748,N_13730,N_14283);
or U14749 (N_14749,N_14278,N_13886);
xor U14750 (N_14750,N_13738,N_14189);
nand U14751 (N_14751,N_14120,N_13632);
and U14752 (N_14752,N_14311,N_14059);
and U14753 (N_14753,N_13723,N_13697);
xnor U14754 (N_14754,N_13963,N_14360);
and U14755 (N_14755,N_13875,N_13656);
and U14756 (N_14756,N_14021,N_14067);
and U14757 (N_14757,N_13761,N_14075);
or U14758 (N_14758,N_13820,N_14298);
and U14759 (N_14759,N_14218,N_13706);
nor U14760 (N_14760,N_13938,N_14280);
and U14761 (N_14761,N_13957,N_13866);
nor U14762 (N_14762,N_14000,N_14211);
or U14763 (N_14763,N_14386,N_14040);
and U14764 (N_14764,N_13716,N_13955);
and U14765 (N_14765,N_13930,N_13894);
xnor U14766 (N_14766,N_13633,N_14331);
nand U14767 (N_14767,N_13625,N_13637);
and U14768 (N_14768,N_13631,N_14352);
nand U14769 (N_14769,N_13703,N_14178);
nor U14770 (N_14770,N_14325,N_13803);
or U14771 (N_14771,N_13649,N_13657);
nor U14772 (N_14772,N_13954,N_14378);
and U14773 (N_14773,N_13711,N_14266);
nand U14774 (N_14774,N_13675,N_13602);
or U14775 (N_14775,N_13972,N_14235);
and U14776 (N_14776,N_13933,N_14382);
or U14777 (N_14777,N_14239,N_14087);
xnor U14778 (N_14778,N_14221,N_13926);
and U14779 (N_14779,N_14037,N_14267);
nand U14780 (N_14780,N_13968,N_14015);
and U14781 (N_14781,N_13701,N_14344);
xor U14782 (N_14782,N_14257,N_13704);
nor U14783 (N_14783,N_14082,N_13907);
nor U14784 (N_14784,N_13655,N_14337);
xnor U14785 (N_14785,N_13638,N_14145);
nor U14786 (N_14786,N_14339,N_13880);
or U14787 (N_14787,N_14012,N_13686);
nor U14788 (N_14788,N_14108,N_13860);
nand U14789 (N_14789,N_14250,N_14288);
nand U14790 (N_14790,N_14155,N_13879);
nor U14791 (N_14791,N_14341,N_14196);
xnor U14792 (N_14792,N_14150,N_13661);
xnor U14793 (N_14793,N_13925,N_14227);
nor U14794 (N_14794,N_13642,N_13967);
xnor U14795 (N_14795,N_13644,N_13604);
xor U14796 (N_14796,N_13621,N_13877);
nor U14797 (N_14797,N_14249,N_13795);
nor U14798 (N_14798,N_13932,N_13975);
nor U14799 (N_14799,N_13807,N_14228);
nor U14800 (N_14800,N_13662,N_14115);
and U14801 (N_14801,N_13954,N_13816);
xor U14802 (N_14802,N_13993,N_14162);
nand U14803 (N_14803,N_14200,N_14351);
or U14804 (N_14804,N_14314,N_13882);
or U14805 (N_14805,N_14115,N_14039);
xor U14806 (N_14806,N_14333,N_14179);
and U14807 (N_14807,N_13967,N_14238);
or U14808 (N_14808,N_13816,N_13935);
or U14809 (N_14809,N_14115,N_13828);
nand U14810 (N_14810,N_14246,N_14389);
and U14811 (N_14811,N_13813,N_13789);
or U14812 (N_14812,N_14326,N_13901);
or U14813 (N_14813,N_14265,N_14105);
xor U14814 (N_14814,N_14325,N_14261);
nor U14815 (N_14815,N_14094,N_14325);
and U14816 (N_14816,N_13736,N_14235);
and U14817 (N_14817,N_13941,N_13943);
xnor U14818 (N_14818,N_13670,N_14004);
nand U14819 (N_14819,N_14289,N_14088);
or U14820 (N_14820,N_13752,N_13664);
nand U14821 (N_14821,N_13776,N_13779);
nor U14822 (N_14822,N_14275,N_13791);
xor U14823 (N_14823,N_13625,N_14109);
or U14824 (N_14824,N_14099,N_13733);
and U14825 (N_14825,N_13785,N_13946);
nor U14826 (N_14826,N_14144,N_14340);
nor U14827 (N_14827,N_14213,N_13839);
xor U14828 (N_14828,N_13915,N_14063);
xor U14829 (N_14829,N_13982,N_14003);
xor U14830 (N_14830,N_13844,N_13627);
xnor U14831 (N_14831,N_14368,N_14006);
and U14832 (N_14832,N_13856,N_13671);
xor U14833 (N_14833,N_13621,N_13874);
xnor U14834 (N_14834,N_13827,N_13611);
xnor U14835 (N_14835,N_13613,N_14355);
or U14836 (N_14836,N_13974,N_13866);
nand U14837 (N_14837,N_14215,N_14093);
and U14838 (N_14838,N_14146,N_13670);
xor U14839 (N_14839,N_14189,N_13848);
nor U14840 (N_14840,N_14142,N_14052);
nor U14841 (N_14841,N_13619,N_13873);
nand U14842 (N_14842,N_14189,N_13772);
xor U14843 (N_14843,N_14041,N_13988);
and U14844 (N_14844,N_14133,N_13787);
nand U14845 (N_14845,N_13844,N_14331);
nand U14846 (N_14846,N_13991,N_14183);
nand U14847 (N_14847,N_14375,N_13825);
or U14848 (N_14848,N_13637,N_14168);
or U14849 (N_14849,N_14345,N_14010);
nand U14850 (N_14850,N_13907,N_13722);
xnor U14851 (N_14851,N_14116,N_13655);
xnor U14852 (N_14852,N_13691,N_14247);
nand U14853 (N_14853,N_14259,N_13806);
nand U14854 (N_14854,N_13819,N_13873);
and U14855 (N_14855,N_13751,N_13953);
and U14856 (N_14856,N_14354,N_14340);
or U14857 (N_14857,N_14033,N_14072);
nor U14858 (N_14858,N_13600,N_14169);
or U14859 (N_14859,N_14305,N_13847);
and U14860 (N_14860,N_14363,N_14054);
and U14861 (N_14861,N_14011,N_14121);
nor U14862 (N_14862,N_13956,N_14159);
or U14863 (N_14863,N_14174,N_14289);
or U14864 (N_14864,N_13642,N_13858);
nand U14865 (N_14865,N_13633,N_14385);
and U14866 (N_14866,N_14343,N_14202);
or U14867 (N_14867,N_14317,N_13892);
xnor U14868 (N_14868,N_13611,N_14230);
and U14869 (N_14869,N_14108,N_14345);
or U14870 (N_14870,N_14004,N_13902);
nor U14871 (N_14871,N_13665,N_13699);
xor U14872 (N_14872,N_14363,N_14024);
xor U14873 (N_14873,N_13897,N_13947);
and U14874 (N_14874,N_13976,N_14115);
nand U14875 (N_14875,N_14185,N_14369);
xor U14876 (N_14876,N_13645,N_13981);
and U14877 (N_14877,N_13766,N_14064);
nor U14878 (N_14878,N_14104,N_13957);
nand U14879 (N_14879,N_14135,N_13945);
xnor U14880 (N_14880,N_13640,N_14355);
and U14881 (N_14881,N_13762,N_14016);
nor U14882 (N_14882,N_14391,N_14098);
or U14883 (N_14883,N_13770,N_13607);
nand U14884 (N_14884,N_13987,N_14222);
nand U14885 (N_14885,N_14153,N_14241);
xor U14886 (N_14886,N_13787,N_14362);
nand U14887 (N_14887,N_13726,N_14367);
nand U14888 (N_14888,N_13647,N_14015);
xor U14889 (N_14889,N_14169,N_13647);
or U14890 (N_14890,N_14010,N_13817);
and U14891 (N_14891,N_14253,N_13764);
xnor U14892 (N_14892,N_14338,N_14274);
nand U14893 (N_14893,N_13956,N_14042);
or U14894 (N_14894,N_13736,N_14027);
nand U14895 (N_14895,N_14142,N_14006);
and U14896 (N_14896,N_14018,N_13739);
nand U14897 (N_14897,N_14371,N_13632);
or U14898 (N_14898,N_14389,N_13688);
nand U14899 (N_14899,N_14380,N_14295);
and U14900 (N_14900,N_14247,N_13941);
or U14901 (N_14901,N_13603,N_14281);
and U14902 (N_14902,N_14317,N_13674);
or U14903 (N_14903,N_14123,N_14110);
nand U14904 (N_14904,N_13741,N_13948);
or U14905 (N_14905,N_14293,N_14076);
and U14906 (N_14906,N_13914,N_13632);
and U14907 (N_14907,N_14332,N_14314);
xor U14908 (N_14908,N_14046,N_14288);
xor U14909 (N_14909,N_13747,N_14280);
nor U14910 (N_14910,N_14305,N_14062);
xnor U14911 (N_14911,N_13845,N_14082);
nand U14912 (N_14912,N_14075,N_13792);
nor U14913 (N_14913,N_14204,N_14268);
nand U14914 (N_14914,N_13719,N_14009);
or U14915 (N_14915,N_14368,N_14366);
nor U14916 (N_14916,N_13634,N_14310);
nand U14917 (N_14917,N_13912,N_13861);
nand U14918 (N_14918,N_13799,N_14322);
nand U14919 (N_14919,N_13939,N_13967);
xor U14920 (N_14920,N_13785,N_14281);
nand U14921 (N_14921,N_14280,N_14021);
or U14922 (N_14922,N_13684,N_13959);
nor U14923 (N_14923,N_14320,N_14395);
or U14924 (N_14924,N_14389,N_14346);
nor U14925 (N_14925,N_13778,N_13848);
nor U14926 (N_14926,N_14327,N_13797);
xnor U14927 (N_14927,N_13626,N_14020);
xnor U14928 (N_14928,N_14350,N_14247);
and U14929 (N_14929,N_14369,N_14170);
xor U14930 (N_14930,N_14377,N_13880);
nor U14931 (N_14931,N_14292,N_13930);
nand U14932 (N_14932,N_14397,N_13749);
xor U14933 (N_14933,N_13830,N_13828);
xor U14934 (N_14934,N_13716,N_14233);
nor U14935 (N_14935,N_14256,N_14234);
nand U14936 (N_14936,N_14122,N_13894);
and U14937 (N_14937,N_13887,N_13967);
and U14938 (N_14938,N_13879,N_14112);
or U14939 (N_14939,N_13693,N_14098);
xor U14940 (N_14940,N_13766,N_14380);
and U14941 (N_14941,N_14241,N_13768);
nor U14942 (N_14942,N_14034,N_14275);
or U14943 (N_14943,N_14257,N_14112);
or U14944 (N_14944,N_13699,N_13747);
and U14945 (N_14945,N_14256,N_13776);
xnor U14946 (N_14946,N_14182,N_14199);
or U14947 (N_14947,N_14218,N_14034);
and U14948 (N_14948,N_13761,N_13635);
nand U14949 (N_14949,N_14245,N_14351);
xor U14950 (N_14950,N_14139,N_14255);
xnor U14951 (N_14951,N_13663,N_14255);
or U14952 (N_14952,N_13676,N_14232);
nor U14953 (N_14953,N_13790,N_13949);
and U14954 (N_14954,N_14018,N_13680);
nand U14955 (N_14955,N_14179,N_14285);
or U14956 (N_14956,N_14139,N_13731);
nor U14957 (N_14957,N_13731,N_13841);
xor U14958 (N_14958,N_13854,N_14338);
and U14959 (N_14959,N_13832,N_13840);
xnor U14960 (N_14960,N_14023,N_13723);
or U14961 (N_14961,N_14212,N_14192);
nor U14962 (N_14962,N_14034,N_13680);
or U14963 (N_14963,N_14030,N_14013);
xor U14964 (N_14964,N_13746,N_13772);
xnor U14965 (N_14965,N_14242,N_13682);
or U14966 (N_14966,N_14183,N_13830);
or U14967 (N_14967,N_13682,N_13968);
nand U14968 (N_14968,N_13944,N_14147);
nor U14969 (N_14969,N_14296,N_13727);
and U14970 (N_14970,N_14275,N_13666);
nand U14971 (N_14971,N_13930,N_13825);
nor U14972 (N_14972,N_14196,N_13943);
nand U14973 (N_14973,N_14298,N_13679);
nand U14974 (N_14974,N_14222,N_14153);
and U14975 (N_14975,N_14091,N_13958);
nand U14976 (N_14976,N_13679,N_14248);
xnor U14977 (N_14977,N_13886,N_13958);
xnor U14978 (N_14978,N_13820,N_13810);
xor U14979 (N_14979,N_14156,N_14183);
xor U14980 (N_14980,N_14240,N_13951);
or U14981 (N_14981,N_14056,N_13748);
nand U14982 (N_14982,N_14320,N_13831);
and U14983 (N_14983,N_13734,N_14250);
nand U14984 (N_14984,N_14232,N_13635);
nand U14985 (N_14985,N_14027,N_14335);
nor U14986 (N_14986,N_13701,N_14367);
nor U14987 (N_14987,N_13663,N_13751);
nand U14988 (N_14988,N_13645,N_13893);
nand U14989 (N_14989,N_14050,N_14382);
xnor U14990 (N_14990,N_13822,N_13604);
or U14991 (N_14991,N_14262,N_13863);
and U14992 (N_14992,N_13976,N_14208);
nor U14993 (N_14993,N_13678,N_14374);
nand U14994 (N_14994,N_14226,N_14348);
nand U14995 (N_14995,N_13860,N_13847);
or U14996 (N_14996,N_13726,N_14132);
nand U14997 (N_14997,N_14126,N_14259);
nor U14998 (N_14998,N_14108,N_13849);
nor U14999 (N_14999,N_13742,N_14086);
nand U15000 (N_15000,N_13786,N_14069);
or U15001 (N_15001,N_14095,N_14103);
or U15002 (N_15002,N_13770,N_14153);
and U15003 (N_15003,N_13941,N_13701);
xor U15004 (N_15004,N_13904,N_14338);
nand U15005 (N_15005,N_13631,N_14051);
xnor U15006 (N_15006,N_14004,N_14363);
and U15007 (N_15007,N_14281,N_14382);
nor U15008 (N_15008,N_14352,N_13848);
and U15009 (N_15009,N_14158,N_13797);
and U15010 (N_15010,N_14194,N_13901);
or U15011 (N_15011,N_13794,N_14309);
or U15012 (N_15012,N_13911,N_14284);
xor U15013 (N_15013,N_13937,N_13681);
and U15014 (N_15014,N_13609,N_13974);
and U15015 (N_15015,N_14005,N_13718);
or U15016 (N_15016,N_14250,N_14148);
nand U15017 (N_15017,N_13658,N_14114);
xnor U15018 (N_15018,N_14299,N_13848);
or U15019 (N_15019,N_13939,N_13893);
xnor U15020 (N_15020,N_13666,N_14157);
nor U15021 (N_15021,N_13667,N_13645);
xnor U15022 (N_15022,N_13783,N_13935);
or U15023 (N_15023,N_13767,N_14316);
nor U15024 (N_15024,N_13817,N_14020);
and U15025 (N_15025,N_14194,N_13620);
xor U15026 (N_15026,N_13768,N_13941);
nand U15027 (N_15027,N_14090,N_13615);
nor U15028 (N_15028,N_14084,N_14050);
and U15029 (N_15029,N_14395,N_14343);
nor U15030 (N_15030,N_13807,N_13653);
or U15031 (N_15031,N_14221,N_14361);
nand U15032 (N_15032,N_13677,N_14018);
xor U15033 (N_15033,N_14276,N_13810);
nor U15034 (N_15034,N_13643,N_14363);
nand U15035 (N_15035,N_13687,N_13982);
or U15036 (N_15036,N_14356,N_14097);
nand U15037 (N_15037,N_14203,N_14382);
and U15038 (N_15038,N_14107,N_13986);
nand U15039 (N_15039,N_14278,N_13662);
or U15040 (N_15040,N_13846,N_14223);
xor U15041 (N_15041,N_14207,N_14034);
or U15042 (N_15042,N_14176,N_14266);
xor U15043 (N_15043,N_14110,N_14214);
and U15044 (N_15044,N_13669,N_14110);
nor U15045 (N_15045,N_14199,N_14351);
nand U15046 (N_15046,N_13738,N_13801);
or U15047 (N_15047,N_13741,N_14092);
or U15048 (N_15048,N_13937,N_14136);
nor U15049 (N_15049,N_13955,N_14022);
or U15050 (N_15050,N_13717,N_13646);
nand U15051 (N_15051,N_13770,N_13978);
and U15052 (N_15052,N_14048,N_14397);
nand U15053 (N_15053,N_14383,N_13729);
or U15054 (N_15054,N_13920,N_13932);
or U15055 (N_15055,N_13983,N_14138);
xnor U15056 (N_15056,N_14316,N_13972);
xor U15057 (N_15057,N_14113,N_14390);
nor U15058 (N_15058,N_13966,N_13682);
or U15059 (N_15059,N_13608,N_13809);
and U15060 (N_15060,N_13877,N_13962);
and U15061 (N_15061,N_13669,N_13744);
and U15062 (N_15062,N_13977,N_14385);
nand U15063 (N_15063,N_13902,N_13971);
or U15064 (N_15064,N_14216,N_13869);
and U15065 (N_15065,N_14389,N_13648);
and U15066 (N_15066,N_14059,N_13914);
nor U15067 (N_15067,N_14060,N_13923);
or U15068 (N_15068,N_13986,N_14276);
or U15069 (N_15069,N_13833,N_14347);
and U15070 (N_15070,N_14365,N_13903);
and U15071 (N_15071,N_14226,N_14388);
or U15072 (N_15072,N_14026,N_14137);
nand U15073 (N_15073,N_13628,N_14121);
xor U15074 (N_15074,N_13982,N_13959);
nor U15075 (N_15075,N_14380,N_14017);
nand U15076 (N_15076,N_13628,N_13612);
and U15077 (N_15077,N_14022,N_14240);
and U15078 (N_15078,N_14259,N_14238);
or U15079 (N_15079,N_13775,N_13827);
nor U15080 (N_15080,N_14326,N_13919);
nor U15081 (N_15081,N_13646,N_14288);
xor U15082 (N_15082,N_14061,N_14349);
nor U15083 (N_15083,N_13896,N_14203);
and U15084 (N_15084,N_13747,N_14178);
xor U15085 (N_15085,N_14111,N_14170);
or U15086 (N_15086,N_14249,N_14334);
xnor U15087 (N_15087,N_14003,N_14196);
nand U15088 (N_15088,N_13935,N_13710);
nor U15089 (N_15089,N_14386,N_14167);
nor U15090 (N_15090,N_14065,N_14008);
nor U15091 (N_15091,N_13804,N_14381);
nand U15092 (N_15092,N_14287,N_14194);
nand U15093 (N_15093,N_14070,N_13819);
nand U15094 (N_15094,N_13751,N_14168);
nand U15095 (N_15095,N_13710,N_14113);
nor U15096 (N_15096,N_13967,N_14005);
and U15097 (N_15097,N_13700,N_14212);
or U15098 (N_15098,N_13869,N_14368);
and U15099 (N_15099,N_14053,N_14269);
xor U15100 (N_15100,N_14358,N_13938);
xor U15101 (N_15101,N_13884,N_14028);
and U15102 (N_15102,N_14007,N_13863);
nor U15103 (N_15103,N_14191,N_13938);
xnor U15104 (N_15104,N_14245,N_14391);
nand U15105 (N_15105,N_13652,N_14211);
nor U15106 (N_15106,N_13878,N_14259);
xor U15107 (N_15107,N_14135,N_14077);
or U15108 (N_15108,N_13734,N_14372);
nor U15109 (N_15109,N_13625,N_14246);
nor U15110 (N_15110,N_13853,N_13891);
nand U15111 (N_15111,N_14052,N_14216);
and U15112 (N_15112,N_14237,N_14313);
nor U15113 (N_15113,N_13840,N_14037);
or U15114 (N_15114,N_13765,N_14083);
and U15115 (N_15115,N_13871,N_14167);
nor U15116 (N_15116,N_14134,N_14071);
xnor U15117 (N_15117,N_14242,N_13635);
or U15118 (N_15118,N_14363,N_13619);
nand U15119 (N_15119,N_13958,N_14089);
and U15120 (N_15120,N_13727,N_13701);
or U15121 (N_15121,N_13890,N_14192);
or U15122 (N_15122,N_13720,N_14115);
or U15123 (N_15123,N_14247,N_13850);
or U15124 (N_15124,N_13721,N_14380);
xnor U15125 (N_15125,N_13889,N_14085);
nor U15126 (N_15126,N_13654,N_14223);
xnor U15127 (N_15127,N_13603,N_14096);
nor U15128 (N_15128,N_14370,N_13601);
xnor U15129 (N_15129,N_14033,N_13656);
xnor U15130 (N_15130,N_13936,N_13746);
nand U15131 (N_15131,N_13797,N_13726);
or U15132 (N_15132,N_14008,N_13823);
nor U15133 (N_15133,N_14382,N_13701);
nor U15134 (N_15134,N_14212,N_14138);
and U15135 (N_15135,N_13995,N_13612);
nand U15136 (N_15136,N_13801,N_13958);
xor U15137 (N_15137,N_14214,N_14241);
nor U15138 (N_15138,N_13962,N_14088);
or U15139 (N_15139,N_14239,N_13740);
nor U15140 (N_15140,N_13818,N_14296);
or U15141 (N_15141,N_14017,N_14178);
nand U15142 (N_15142,N_14166,N_13603);
xor U15143 (N_15143,N_13874,N_14148);
nand U15144 (N_15144,N_14366,N_14192);
or U15145 (N_15145,N_14153,N_13783);
or U15146 (N_15146,N_13727,N_13696);
and U15147 (N_15147,N_14136,N_14298);
or U15148 (N_15148,N_13810,N_13861);
and U15149 (N_15149,N_14340,N_13900);
or U15150 (N_15150,N_14292,N_13660);
or U15151 (N_15151,N_14032,N_13900);
or U15152 (N_15152,N_14086,N_13714);
xor U15153 (N_15153,N_14379,N_14312);
and U15154 (N_15154,N_13684,N_13810);
xor U15155 (N_15155,N_14106,N_14305);
xor U15156 (N_15156,N_13813,N_13654);
nor U15157 (N_15157,N_14254,N_13717);
nor U15158 (N_15158,N_14145,N_13610);
and U15159 (N_15159,N_14279,N_13920);
or U15160 (N_15160,N_13879,N_13958);
or U15161 (N_15161,N_14167,N_14215);
or U15162 (N_15162,N_13702,N_14323);
or U15163 (N_15163,N_14253,N_13926);
or U15164 (N_15164,N_13908,N_13901);
nor U15165 (N_15165,N_13624,N_14209);
and U15166 (N_15166,N_14254,N_13987);
nor U15167 (N_15167,N_13936,N_13978);
nor U15168 (N_15168,N_14169,N_13724);
or U15169 (N_15169,N_14265,N_13779);
or U15170 (N_15170,N_14024,N_13987);
or U15171 (N_15171,N_14237,N_13782);
or U15172 (N_15172,N_13834,N_14343);
and U15173 (N_15173,N_14254,N_13731);
or U15174 (N_15174,N_14103,N_14063);
xor U15175 (N_15175,N_14270,N_14314);
nor U15176 (N_15176,N_13837,N_14156);
nand U15177 (N_15177,N_14013,N_13723);
nor U15178 (N_15178,N_13805,N_14246);
and U15179 (N_15179,N_13615,N_14360);
or U15180 (N_15180,N_14183,N_13916);
nor U15181 (N_15181,N_13733,N_13797);
nand U15182 (N_15182,N_14360,N_14127);
or U15183 (N_15183,N_14319,N_13969);
and U15184 (N_15184,N_14098,N_13695);
nor U15185 (N_15185,N_14205,N_14301);
and U15186 (N_15186,N_14154,N_14215);
or U15187 (N_15187,N_13932,N_13736);
nand U15188 (N_15188,N_13915,N_13950);
and U15189 (N_15189,N_14014,N_14191);
nand U15190 (N_15190,N_13833,N_14363);
nand U15191 (N_15191,N_14354,N_13801);
nand U15192 (N_15192,N_14059,N_13831);
or U15193 (N_15193,N_13720,N_14274);
xnor U15194 (N_15194,N_13977,N_13806);
nor U15195 (N_15195,N_13799,N_14291);
nand U15196 (N_15196,N_14008,N_14019);
nand U15197 (N_15197,N_14026,N_14313);
or U15198 (N_15198,N_13601,N_13957);
or U15199 (N_15199,N_14145,N_14037);
xor U15200 (N_15200,N_14541,N_14940);
xnor U15201 (N_15201,N_14461,N_14968);
nor U15202 (N_15202,N_14855,N_14943);
nor U15203 (N_15203,N_14848,N_15133);
xnor U15204 (N_15204,N_14733,N_14813);
xnor U15205 (N_15205,N_14823,N_14729);
xor U15206 (N_15206,N_14866,N_15066);
xnor U15207 (N_15207,N_15039,N_15132);
nor U15208 (N_15208,N_14600,N_14479);
nor U15209 (N_15209,N_14981,N_15198);
and U15210 (N_15210,N_14913,N_15059);
or U15211 (N_15211,N_15197,N_15003);
xnor U15212 (N_15212,N_14402,N_14432);
and U15213 (N_15213,N_15121,N_14945);
or U15214 (N_15214,N_15137,N_14934);
nor U15215 (N_15215,N_14923,N_14587);
or U15216 (N_15216,N_14906,N_14840);
nand U15217 (N_15217,N_14686,N_14431);
xor U15218 (N_15218,N_15194,N_14803);
nor U15219 (N_15219,N_14928,N_15093);
xor U15220 (N_15220,N_14871,N_14498);
nand U15221 (N_15221,N_15038,N_15156);
or U15222 (N_15222,N_14671,N_15165);
nand U15223 (N_15223,N_14557,N_14895);
and U15224 (N_15224,N_14708,N_15042);
nand U15225 (N_15225,N_15120,N_14865);
and U15226 (N_15226,N_14944,N_14555);
xor U15227 (N_15227,N_15114,N_15124);
nor U15228 (N_15228,N_15142,N_14881);
nand U15229 (N_15229,N_14413,N_14536);
xnor U15230 (N_15230,N_14989,N_14509);
and U15231 (N_15231,N_15145,N_15177);
nor U15232 (N_15232,N_14878,N_14670);
xnor U15233 (N_15233,N_14453,N_14471);
or U15234 (N_15234,N_14506,N_14611);
nor U15235 (N_15235,N_14980,N_14910);
and U15236 (N_15236,N_14537,N_14789);
or U15237 (N_15237,N_14796,N_14914);
nor U15238 (N_15238,N_15049,N_14401);
nand U15239 (N_15239,N_15150,N_14510);
xnor U15240 (N_15240,N_14925,N_14668);
nor U15241 (N_15241,N_15018,N_14770);
nor U15242 (N_15242,N_14459,N_15080);
nor U15243 (N_15243,N_14596,N_14736);
or U15244 (N_15244,N_15036,N_14663);
and U15245 (N_15245,N_14825,N_14832);
nor U15246 (N_15246,N_14927,N_14893);
nand U15247 (N_15247,N_14674,N_14870);
and U15248 (N_15248,N_15123,N_14716);
xor U15249 (N_15249,N_14976,N_14751);
or U15250 (N_15250,N_14778,N_15166);
and U15251 (N_15251,N_14639,N_14853);
nor U15252 (N_15252,N_14451,N_14644);
nand U15253 (N_15253,N_14801,N_15108);
nor U15254 (N_15254,N_14588,N_14707);
or U15255 (N_15255,N_15033,N_14808);
or U15256 (N_15256,N_14548,N_14746);
and U15257 (N_15257,N_15106,N_14483);
nand U15258 (N_15258,N_14798,N_14858);
xnor U15259 (N_15259,N_14998,N_14754);
nand U15260 (N_15260,N_14423,N_15109);
or U15261 (N_15261,N_14810,N_14637);
xnor U15262 (N_15262,N_14669,N_14643);
xor U15263 (N_15263,N_14462,N_14558);
and U15264 (N_15264,N_15017,N_14966);
xnor U15265 (N_15265,N_15141,N_14655);
xor U15266 (N_15266,N_14486,N_14921);
or U15267 (N_15267,N_14983,N_15087);
nand U15268 (N_15268,N_14638,N_14955);
and U15269 (N_15269,N_14738,N_14666);
nand U15270 (N_15270,N_14884,N_14745);
xor U15271 (N_15271,N_14742,N_14922);
xor U15272 (N_15272,N_15117,N_15082);
nor U15273 (N_15273,N_15021,N_14783);
and U15274 (N_15274,N_14460,N_15182);
xnor U15275 (N_15275,N_14992,N_14433);
nor U15276 (N_15276,N_14814,N_14418);
or U15277 (N_15277,N_14752,N_15161);
and U15278 (N_15278,N_15027,N_14470);
or U15279 (N_15279,N_15164,N_14875);
nand U15280 (N_15280,N_14862,N_14522);
nand U15281 (N_15281,N_14930,N_15009);
or U15282 (N_15282,N_14718,N_15044);
and U15283 (N_15283,N_14723,N_15111);
xnor U15284 (N_15284,N_14873,N_14978);
xnor U15285 (N_15285,N_14542,N_14648);
or U15286 (N_15286,N_14775,N_14477);
xor U15287 (N_15287,N_14649,N_14597);
nand U15288 (N_15288,N_15012,N_14571);
xnor U15289 (N_15289,N_14436,N_14615);
xor U15290 (N_15290,N_14407,N_14891);
nor U15291 (N_15291,N_14838,N_14991);
nand U15292 (N_15292,N_14972,N_15035);
and U15293 (N_15293,N_15175,N_14816);
nand U15294 (N_15294,N_14476,N_14854);
nor U15295 (N_15295,N_14488,N_14835);
nor U15296 (N_15296,N_14846,N_14788);
or U15297 (N_15297,N_15006,N_15139);
nand U15298 (N_15298,N_14995,N_14647);
xor U15299 (N_15299,N_14852,N_14767);
and U15300 (N_15300,N_15174,N_14799);
xor U15301 (N_15301,N_14755,N_15160);
nor U15302 (N_15302,N_14688,N_14577);
or U15303 (N_15303,N_14888,N_14847);
nor U15304 (N_15304,N_14965,N_15187);
and U15305 (N_15305,N_14828,N_14714);
or U15306 (N_15306,N_15122,N_14740);
xor U15307 (N_15307,N_14699,N_14440);
or U15308 (N_15308,N_14826,N_14556);
nand U15309 (N_15309,N_14491,N_14566);
or U15310 (N_15310,N_14409,N_15115);
nand U15311 (N_15311,N_14503,N_14950);
nand U15312 (N_15312,N_14434,N_14812);
nand U15313 (N_15313,N_14497,N_15143);
or U15314 (N_15314,N_15045,N_15022);
xor U15315 (N_15315,N_15047,N_14758);
nor U15316 (N_15316,N_14684,N_15062);
or U15317 (N_15317,N_15015,N_14918);
or U15318 (N_15318,N_14784,N_14659);
xor U15319 (N_15319,N_14726,N_15056);
nand U15320 (N_15320,N_14539,N_14484);
xor U15321 (N_15321,N_14997,N_14986);
nand U15322 (N_15322,N_14926,N_14988);
nor U15323 (N_15323,N_14960,N_14843);
nor U15324 (N_15324,N_15181,N_15118);
and U15325 (N_15325,N_14710,N_14426);
or U15326 (N_15326,N_15172,N_14646);
or U15327 (N_15327,N_14869,N_15019);
xnor U15328 (N_15328,N_14719,N_14901);
and U15329 (N_15329,N_14482,N_14677);
xor U15330 (N_15330,N_14416,N_15020);
or U15331 (N_15331,N_14657,N_14593);
and U15332 (N_15332,N_15170,N_15040);
xnor U15333 (N_15333,N_14970,N_14595);
nor U15334 (N_15334,N_14636,N_14599);
and U15335 (N_15335,N_15070,N_14618);
and U15336 (N_15336,N_14867,N_14952);
xor U15337 (N_15337,N_15078,N_14552);
or U15338 (N_15338,N_14804,N_14908);
or U15339 (N_15339,N_14941,N_14525);
and U15340 (N_15340,N_14935,N_14642);
xnor U15341 (N_15341,N_15131,N_14792);
and U15342 (N_15342,N_14485,N_15067);
nor U15343 (N_15343,N_14757,N_14500);
or U15344 (N_15344,N_15178,N_15159);
nand U15345 (N_15345,N_14961,N_14653);
xnor U15346 (N_15346,N_14811,N_15058);
nand U15347 (N_15347,N_14516,N_14889);
or U15348 (N_15348,N_14517,N_14604);
xor U15349 (N_15349,N_15079,N_14463);
nand U15350 (N_15350,N_15179,N_14845);
xnor U15351 (N_15351,N_14468,N_15103);
or U15352 (N_15352,N_14779,N_14885);
xnor U15353 (N_15353,N_15104,N_14452);
nor U15354 (N_15354,N_15091,N_14549);
and U15355 (N_15355,N_14971,N_14731);
or U15356 (N_15356,N_15130,N_14495);
or U15357 (N_15357,N_14818,N_15180);
nand U15358 (N_15358,N_15051,N_14800);
nand U15359 (N_15359,N_14578,N_14912);
nor U15360 (N_15360,N_14520,N_14610);
or U15361 (N_15361,N_14762,N_15077);
nor U15362 (N_15362,N_14563,N_15025);
and U15363 (N_15363,N_15063,N_14609);
xor U15364 (N_15364,N_14598,N_14982);
or U15365 (N_15365,N_15007,N_14831);
or U15366 (N_15366,N_15129,N_14781);
xor U15367 (N_15367,N_14664,N_14446);
nand U15368 (N_15368,N_14861,N_15116);
xor U15369 (N_15369,N_14911,N_15026);
xor U15370 (N_15370,N_14447,N_14547);
or U15371 (N_15371,N_14999,N_14584);
nor U15372 (N_15372,N_15110,N_14905);
and U15373 (N_15373,N_14979,N_14732);
xnor U15374 (N_15374,N_15126,N_15053);
xor U15375 (N_15375,N_14737,N_14967);
nor U15376 (N_15376,N_14882,N_14951);
xnor U15377 (N_15377,N_15144,N_14857);
xor U15378 (N_15378,N_15119,N_14614);
nand U15379 (N_15379,N_14628,N_14675);
nand U15380 (N_15380,N_14466,N_15084);
nand U15381 (N_15381,N_14626,N_14984);
nor U15382 (N_15382,N_14896,N_15184);
and U15383 (N_15383,N_14819,N_14502);
and U15384 (N_15384,N_14937,N_14631);
nor U15385 (N_15385,N_14411,N_14730);
or U15386 (N_15386,N_15083,N_14420);
nand U15387 (N_15387,N_14765,N_14724);
and U15388 (N_15388,N_14836,N_14421);
or U15389 (N_15389,N_15016,N_15199);
and U15390 (N_15390,N_14620,N_14743);
and U15391 (N_15391,N_14877,N_14876);
xor U15392 (N_15392,N_14706,N_14464);
or U15393 (N_15393,N_14693,N_14851);
nand U15394 (N_15394,N_14443,N_14494);
xor U15395 (N_15395,N_14990,N_15125);
nor U15396 (N_15396,N_15005,N_15157);
xnor U15397 (N_15397,N_14985,N_15147);
nand U15398 (N_15398,N_14933,N_14640);
nand U15399 (N_15399,N_14932,N_15148);
xnor U15400 (N_15400,N_14424,N_14807);
or U15401 (N_15401,N_14568,N_15057);
or U15402 (N_15402,N_14475,N_14963);
nor U15403 (N_15403,N_15010,N_14809);
nor U15404 (N_15404,N_14709,N_14772);
nor U15405 (N_15405,N_15101,N_15081);
nand U15406 (N_15406,N_15191,N_14702);
nand U15407 (N_15407,N_15068,N_14410);
nand U15408 (N_15408,N_14805,N_14602);
nand U15409 (N_15409,N_15064,N_14430);
nor U15410 (N_15410,N_14533,N_15162);
nand U15411 (N_15411,N_14630,N_14903);
or U15412 (N_15412,N_14797,N_14713);
nand U15413 (N_15413,N_14996,N_14521);
xnor U15414 (N_15414,N_14607,N_14513);
xor U15415 (N_15415,N_14652,N_14863);
xor U15416 (N_15416,N_14512,N_14467);
nor U15417 (N_15417,N_14890,N_14658);
or U15418 (N_15418,N_14603,N_15023);
nand U15419 (N_15419,N_14472,N_15004);
nand U15420 (N_15420,N_14508,N_14728);
or U15421 (N_15421,N_14749,N_15193);
and U15422 (N_15422,N_14489,N_14592);
xnor U15423 (N_15423,N_14774,N_15102);
nand U15424 (N_15424,N_14705,N_14802);
xnor U15425 (N_15425,N_15168,N_14493);
or U15426 (N_15426,N_14821,N_14665);
nand U15427 (N_15427,N_14860,N_14616);
or U15428 (N_15428,N_15030,N_14404);
and U15429 (N_15429,N_14579,N_14573);
xor U15430 (N_15430,N_15008,N_15024);
nor U15431 (N_15431,N_14844,N_14524);
or U15432 (N_15432,N_15028,N_15043);
xor U15433 (N_15433,N_14872,N_14435);
or U15434 (N_15434,N_14920,N_14727);
nand U15435 (N_15435,N_14739,N_14575);
and U15436 (N_15436,N_14883,N_14696);
xnor U15437 (N_15437,N_14458,N_14564);
or U15438 (N_15438,N_14892,N_14793);
nand U15439 (N_15439,N_15183,N_14773);
or U15440 (N_15440,N_14829,N_14899);
xor U15441 (N_15441,N_14683,N_14776);
or U15442 (N_15442,N_14572,N_14629);
or U15443 (N_15443,N_14625,N_14504);
and U15444 (N_15444,N_14478,N_14581);
nor U15445 (N_15445,N_15032,N_14554);
nand U15446 (N_15446,N_15088,N_14422);
and U15447 (N_15447,N_15050,N_14529);
or U15448 (N_15448,N_14535,N_14787);
nor U15449 (N_15449,N_14824,N_14679);
nor U15450 (N_15450,N_14514,N_14790);
nor U15451 (N_15451,N_14689,N_14586);
and U15452 (N_15452,N_14957,N_15195);
xnor U15453 (N_15453,N_14850,N_15095);
or U15454 (N_15454,N_15011,N_14907);
and U15455 (N_15455,N_15085,N_14833);
and U15456 (N_15456,N_15135,N_14954);
and U15457 (N_15457,N_14938,N_14949);
and U15458 (N_15458,N_14769,N_15097);
or U15459 (N_15459,N_14766,N_14680);
nand U15460 (N_15460,N_15013,N_15075);
or U15461 (N_15461,N_15167,N_14676);
or U15462 (N_15462,N_14567,N_14806);
xor U15463 (N_15463,N_14627,N_14617);
xnor U15464 (N_15464,N_14859,N_14403);
nor U15465 (N_15465,N_14794,N_14904);
xnor U15466 (N_15466,N_14417,N_14842);
and U15467 (N_15467,N_15146,N_14527);
xnor U15468 (N_15468,N_14864,N_14785);
nor U15469 (N_15469,N_14887,N_14565);
or U15470 (N_15470,N_15190,N_14601);
nor U15471 (N_15471,N_14496,N_14448);
xnor U15472 (N_15472,N_14987,N_14656);
or U15473 (N_15473,N_14457,N_14544);
xnor U15474 (N_15474,N_14562,N_14694);
xnor U15475 (N_15475,N_14576,N_14969);
or U15476 (N_15476,N_14441,N_14419);
nor U15477 (N_15477,N_14771,N_14480);
nand U15478 (N_15478,N_14518,N_15014);
xor U15479 (N_15479,N_14849,N_15152);
xnor U15480 (N_15480,N_15151,N_14830);
or U15481 (N_15481,N_15099,N_14764);
and U15482 (N_15482,N_14760,N_14634);
and U15483 (N_15483,N_15112,N_14545);
or U15484 (N_15484,N_15140,N_14519);
nand U15485 (N_15485,N_14894,N_15192);
or U15486 (N_15486,N_14473,N_14550);
nor U15487 (N_15487,N_14942,N_14444);
and U15488 (N_15488,N_14605,N_14667);
xor U15489 (N_15489,N_15149,N_14837);
and U15490 (N_15490,N_14761,N_14791);
xor U15491 (N_15491,N_14469,N_14427);
xnor U15492 (N_15492,N_14662,N_14454);
nand U15493 (N_15493,N_15001,N_14582);
nor U15494 (N_15494,N_14487,N_14553);
nand U15495 (N_15495,N_14929,N_15173);
nand U15496 (N_15496,N_14777,N_14551);
and U15497 (N_15497,N_15054,N_14574);
xnor U15498 (N_15498,N_14449,N_14633);
nand U15499 (N_15499,N_14717,N_14622);
or U15500 (N_15500,N_15189,N_14975);
or U15501 (N_15501,N_14559,N_15031);
nor U15502 (N_15502,N_14585,N_14687);
nor U15503 (N_15503,N_14612,N_15052);
nor U15504 (N_15504,N_14915,N_14701);
or U15505 (N_15505,N_15098,N_14523);
or U15506 (N_15506,N_15138,N_14839);
nand U15507 (N_15507,N_14902,N_14492);
xor U15508 (N_15508,N_15073,N_14959);
and U15509 (N_15509,N_15096,N_15041);
and U15510 (N_15510,N_14993,N_14624);
or U15511 (N_15511,N_14583,N_14682);
or U15512 (N_15512,N_14569,N_14720);
nor U15513 (N_15513,N_14768,N_15090);
nand U15514 (N_15514,N_14532,N_15048);
nand U15515 (N_15515,N_15002,N_14704);
xor U15516 (N_15516,N_14763,N_15037);
xor U15517 (N_15517,N_14700,N_14712);
nand U15518 (N_15518,N_15196,N_14673);
nand U15519 (N_15519,N_14962,N_14827);
nor U15520 (N_15520,N_15071,N_14956);
nand U15521 (N_15521,N_15072,N_14543);
nand U15522 (N_15522,N_14546,N_14974);
nand U15523 (N_15523,N_14931,N_15185);
and U15524 (N_15524,N_14531,N_14408);
nand U15525 (N_15525,N_14822,N_14747);
nand U15526 (N_15526,N_14898,N_14400);
and U15527 (N_15527,N_15154,N_14499);
and U15528 (N_15528,N_15055,N_14507);
or U15529 (N_15529,N_14924,N_14994);
or U15530 (N_15530,N_14678,N_15000);
or U15531 (N_15531,N_14645,N_15094);
nor U15532 (N_15532,N_14953,N_14886);
or U15533 (N_15533,N_15061,N_14936);
nand U15534 (N_15534,N_14744,N_14455);
and U15535 (N_15535,N_14561,N_14672);
nor U15536 (N_15536,N_14589,N_14964);
nand U15537 (N_15537,N_14425,N_14759);
xor U15538 (N_15538,N_14834,N_14632);
nor U15539 (N_15539,N_14939,N_14958);
and U15540 (N_15540,N_15176,N_14868);
xor U15541 (N_15541,N_14526,N_14748);
nor U15542 (N_15542,N_15065,N_14654);
xnor U15543 (N_15543,N_14438,N_14621);
xnor U15544 (N_15544,N_14534,N_14721);
nand U15545 (N_15545,N_14490,N_14916);
xnor U15546 (N_15546,N_14900,N_14692);
nand U15547 (N_15547,N_14917,N_14623);
nand U15548 (N_15548,N_14697,N_14442);
nand U15549 (N_15549,N_14977,N_15113);
nand U15550 (N_15550,N_15171,N_14530);
and U15551 (N_15551,N_15153,N_14428);
nand U15552 (N_15552,N_15105,N_14560);
and U15553 (N_15553,N_14594,N_14780);
nand U15554 (N_15554,N_14651,N_14817);
nand U15555 (N_15555,N_14570,N_14456);
nor U15556 (N_15556,N_14820,N_15060);
and U15557 (N_15557,N_14481,N_14741);
nor U15558 (N_15558,N_14660,N_15074);
or U15559 (N_15559,N_14973,N_14715);
or U15560 (N_15560,N_14528,N_14946);
and U15561 (N_15561,N_14445,N_14879);
nand U15562 (N_15562,N_14691,N_14703);
and U15563 (N_15563,N_14606,N_14439);
and U15564 (N_15564,N_15107,N_15155);
nor U15565 (N_15565,N_14505,N_14756);
and U15566 (N_15566,N_14661,N_15127);
nor U15567 (N_15567,N_14880,N_14698);
xnor U15568 (N_15568,N_15163,N_15128);
nand U15569 (N_15569,N_14501,N_14815);
nand U15570 (N_15570,N_14608,N_14734);
nor U15571 (N_15571,N_14619,N_15076);
and U15572 (N_15572,N_14405,N_14415);
and U15573 (N_15573,N_14874,N_14750);
and U15574 (N_15574,N_14511,N_15086);
nor U15575 (N_15575,N_14782,N_14429);
nand U15576 (N_15576,N_14450,N_14474);
or U15577 (N_15577,N_14690,N_14711);
nand U15578 (N_15578,N_15158,N_14613);
xor U15579 (N_15579,N_14540,N_14909);
nor U15580 (N_15580,N_14735,N_14515);
nor U15581 (N_15581,N_15188,N_14685);
xnor U15582 (N_15582,N_15169,N_14650);
nand U15583 (N_15583,N_14580,N_15034);
xor U15584 (N_15584,N_14635,N_15134);
and U15585 (N_15585,N_15089,N_14856);
nor U15586 (N_15586,N_15092,N_15046);
or U15587 (N_15587,N_14681,N_14406);
and U15588 (N_15588,N_14795,N_14948);
and U15589 (N_15589,N_14641,N_14695);
xor U15590 (N_15590,N_15186,N_14786);
nor U15591 (N_15591,N_14947,N_15029);
or U15592 (N_15592,N_14412,N_14725);
and U15593 (N_15593,N_15100,N_14722);
nand U15594 (N_15594,N_15069,N_14753);
nand U15595 (N_15595,N_14591,N_14414);
nor U15596 (N_15596,N_14465,N_14538);
xor U15597 (N_15597,N_14897,N_14919);
and U15598 (N_15598,N_14437,N_14590);
xor U15599 (N_15599,N_15136,N_14841);
and U15600 (N_15600,N_15174,N_15099);
nand U15601 (N_15601,N_14516,N_14989);
nor U15602 (N_15602,N_15070,N_14462);
or U15603 (N_15603,N_14790,N_14438);
nand U15604 (N_15604,N_15001,N_14855);
xor U15605 (N_15605,N_15040,N_15114);
nand U15606 (N_15606,N_14674,N_14523);
xor U15607 (N_15607,N_14820,N_15008);
xor U15608 (N_15608,N_14747,N_14569);
nor U15609 (N_15609,N_14893,N_14547);
xnor U15610 (N_15610,N_14411,N_15051);
nor U15611 (N_15611,N_14818,N_15177);
or U15612 (N_15612,N_14761,N_14521);
and U15613 (N_15613,N_15054,N_15053);
nor U15614 (N_15614,N_14739,N_14980);
nand U15615 (N_15615,N_14540,N_14687);
or U15616 (N_15616,N_14942,N_14544);
xor U15617 (N_15617,N_14994,N_14707);
nand U15618 (N_15618,N_14936,N_14530);
and U15619 (N_15619,N_14486,N_15103);
or U15620 (N_15620,N_14614,N_14740);
xnor U15621 (N_15621,N_14865,N_14495);
xnor U15622 (N_15622,N_14462,N_15118);
xor U15623 (N_15623,N_15049,N_15023);
nand U15624 (N_15624,N_14889,N_14537);
xor U15625 (N_15625,N_14863,N_14776);
xor U15626 (N_15626,N_14960,N_14533);
and U15627 (N_15627,N_14986,N_14797);
nor U15628 (N_15628,N_15110,N_14958);
nand U15629 (N_15629,N_14950,N_14644);
nand U15630 (N_15630,N_14828,N_14510);
xnor U15631 (N_15631,N_14628,N_14796);
nor U15632 (N_15632,N_14440,N_14664);
or U15633 (N_15633,N_14860,N_14727);
nor U15634 (N_15634,N_14545,N_14421);
nor U15635 (N_15635,N_14824,N_14983);
and U15636 (N_15636,N_14963,N_14852);
nor U15637 (N_15637,N_14664,N_14508);
or U15638 (N_15638,N_14899,N_14743);
xnor U15639 (N_15639,N_14489,N_14708);
xor U15640 (N_15640,N_14651,N_14882);
nor U15641 (N_15641,N_14728,N_14447);
or U15642 (N_15642,N_14676,N_14464);
and U15643 (N_15643,N_14594,N_14798);
xnor U15644 (N_15644,N_14974,N_15008);
or U15645 (N_15645,N_14838,N_14779);
nor U15646 (N_15646,N_14911,N_14879);
and U15647 (N_15647,N_14698,N_14863);
nor U15648 (N_15648,N_14907,N_14687);
xor U15649 (N_15649,N_14816,N_14859);
or U15650 (N_15650,N_14901,N_14592);
nor U15651 (N_15651,N_14816,N_14554);
nand U15652 (N_15652,N_15046,N_15054);
nand U15653 (N_15653,N_14895,N_14846);
nor U15654 (N_15654,N_15193,N_14971);
nor U15655 (N_15655,N_15025,N_14459);
or U15656 (N_15656,N_14991,N_14921);
or U15657 (N_15657,N_14700,N_14452);
nand U15658 (N_15658,N_14677,N_14501);
nand U15659 (N_15659,N_15109,N_14462);
nor U15660 (N_15660,N_14850,N_15150);
nand U15661 (N_15661,N_14441,N_14826);
xnor U15662 (N_15662,N_14668,N_14604);
xor U15663 (N_15663,N_14445,N_14410);
nand U15664 (N_15664,N_14856,N_14404);
xor U15665 (N_15665,N_14916,N_14459);
nand U15666 (N_15666,N_14745,N_14596);
nand U15667 (N_15667,N_14550,N_14754);
nand U15668 (N_15668,N_15188,N_14862);
nor U15669 (N_15669,N_15096,N_14726);
or U15670 (N_15670,N_14685,N_14637);
xnor U15671 (N_15671,N_14741,N_14500);
xor U15672 (N_15672,N_14494,N_15008);
xor U15673 (N_15673,N_14552,N_15187);
or U15674 (N_15674,N_15030,N_15000);
or U15675 (N_15675,N_14581,N_14878);
and U15676 (N_15676,N_14652,N_14997);
xnor U15677 (N_15677,N_14862,N_14593);
or U15678 (N_15678,N_14695,N_14856);
nand U15679 (N_15679,N_15114,N_15093);
nor U15680 (N_15680,N_15101,N_15138);
nor U15681 (N_15681,N_14953,N_14450);
xnor U15682 (N_15682,N_14700,N_14839);
nor U15683 (N_15683,N_14569,N_14786);
or U15684 (N_15684,N_14854,N_14468);
nand U15685 (N_15685,N_14559,N_14647);
and U15686 (N_15686,N_15195,N_14709);
and U15687 (N_15687,N_14493,N_14761);
nand U15688 (N_15688,N_14541,N_14599);
or U15689 (N_15689,N_14583,N_14727);
and U15690 (N_15690,N_14762,N_15126);
nor U15691 (N_15691,N_14988,N_15077);
or U15692 (N_15692,N_14707,N_15025);
or U15693 (N_15693,N_15066,N_14569);
and U15694 (N_15694,N_14420,N_14815);
xor U15695 (N_15695,N_14653,N_14956);
nand U15696 (N_15696,N_14473,N_14726);
xor U15697 (N_15697,N_14966,N_14525);
xor U15698 (N_15698,N_15176,N_14838);
nor U15699 (N_15699,N_14879,N_14518);
or U15700 (N_15700,N_14977,N_14642);
or U15701 (N_15701,N_14623,N_14669);
or U15702 (N_15702,N_14479,N_15066);
xnor U15703 (N_15703,N_14811,N_14735);
nor U15704 (N_15704,N_14759,N_14763);
nor U15705 (N_15705,N_14580,N_14516);
xnor U15706 (N_15706,N_14527,N_14589);
nor U15707 (N_15707,N_14971,N_14677);
and U15708 (N_15708,N_15025,N_15055);
xor U15709 (N_15709,N_14899,N_14924);
xor U15710 (N_15710,N_14944,N_14926);
or U15711 (N_15711,N_14678,N_14834);
and U15712 (N_15712,N_14674,N_15081);
nand U15713 (N_15713,N_14409,N_14605);
or U15714 (N_15714,N_14424,N_14650);
xnor U15715 (N_15715,N_14629,N_14542);
xor U15716 (N_15716,N_15021,N_15087);
and U15717 (N_15717,N_14958,N_15179);
or U15718 (N_15718,N_14405,N_14892);
nand U15719 (N_15719,N_14499,N_14496);
nand U15720 (N_15720,N_14768,N_15021);
nor U15721 (N_15721,N_14616,N_15056);
nor U15722 (N_15722,N_14863,N_14631);
or U15723 (N_15723,N_14681,N_15195);
xor U15724 (N_15724,N_15139,N_15127);
xor U15725 (N_15725,N_15132,N_14856);
and U15726 (N_15726,N_15042,N_14844);
xor U15727 (N_15727,N_14449,N_14976);
or U15728 (N_15728,N_14964,N_14776);
and U15729 (N_15729,N_14980,N_14834);
nand U15730 (N_15730,N_14444,N_15036);
nor U15731 (N_15731,N_14545,N_15157);
xnor U15732 (N_15732,N_14862,N_14969);
nor U15733 (N_15733,N_14611,N_14409);
nand U15734 (N_15734,N_14999,N_15016);
and U15735 (N_15735,N_14627,N_14587);
nand U15736 (N_15736,N_14785,N_14421);
and U15737 (N_15737,N_14610,N_14682);
or U15738 (N_15738,N_14714,N_14664);
or U15739 (N_15739,N_14500,N_14781);
nand U15740 (N_15740,N_14445,N_14604);
nor U15741 (N_15741,N_14921,N_14406);
or U15742 (N_15742,N_14656,N_14409);
xor U15743 (N_15743,N_15131,N_14571);
and U15744 (N_15744,N_14647,N_14831);
nor U15745 (N_15745,N_14411,N_14732);
or U15746 (N_15746,N_14772,N_14473);
and U15747 (N_15747,N_14558,N_15048);
nand U15748 (N_15748,N_14630,N_14420);
or U15749 (N_15749,N_14613,N_15171);
and U15750 (N_15750,N_14691,N_14844);
xor U15751 (N_15751,N_14761,N_14971);
and U15752 (N_15752,N_15184,N_14699);
or U15753 (N_15753,N_14608,N_14988);
or U15754 (N_15754,N_14867,N_14917);
nor U15755 (N_15755,N_15155,N_15177);
and U15756 (N_15756,N_15091,N_14965);
xnor U15757 (N_15757,N_14813,N_14601);
or U15758 (N_15758,N_15138,N_14886);
nor U15759 (N_15759,N_14916,N_14787);
or U15760 (N_15760,N_14630,N_14445);
nor U15761 (N_15761,N_14761,N_14667);
nand U15762 (N_15762,N_14734,N_14973);
and U15763 (N_15763,N_15142,N_15075);
xor U15764 (N_15764,N_14650,N_14614);
xor U15765 (N_15765,N_14517,N_14805);
nand U15766 (N_15766,N_14503,N_14752);
or U15767 (N_15767,N_14794,N_14430);
and U15768 (N_15768,N_14515,N_15183);
or U15769 (N_15769,N_14443,N_14952);
and U15770 (N_15770,N_14664,N_14941);
or U15771 (N_15771,N_14892,N_14495);
or U15772 (N_15772,N_14774,N_14897);
nand U15773 (N_15773,N_14875,N_14542);
nand U15774 (N_15774,N_15100,N_14811);
nor U15775 (N_15775,N_14558,N_15127);
or U15776 (N_15776,N_14410,N_14889);
and U15777 (N_15777,N_15020,N_15027);
xor U15778 (N_15778,N_14470,N_14640);
xor U15779 (N_15779,N_14992,N_14756);
or U15780 (N_15780,N_14792,N_14974);
nor U15781 (N_15781,N_15075,N_14686);
nor U15782 (N_15782,N_14507,N_15017);
nand U15783 (N_15783,N_14412,N_14559);
or U15784 (N_15784,N_14850,N_14496);
nor U15785 (N_15785,N_14585,N_14990);
nand U15786 (N_15786,N_15147,N_14827);
nand U15787 (N_15787,N_15066,N_15048);
nand U15788 (N_15788,N_14987,N_14966);
nor U15789 (N_15789,N_14908,N_14958);
nor U15790 (N_15790,N_14573,N_15081);
xnor U15791 (N_15791,N_14924,N_15053);
nand U15792 (N_15792,N_15151,N_15175);
xor U15793 (N_15793,N_14475,N_14526);
xor U15794 (N_15794,N_14710,N_15164);
nand U15795 (N_15795,N_14564,N_15148);
nand U15796 (N_15796,N_14809,N_15125);
nand U15797 (N_15797,N_14854,N_14501);
and U15798 (N_15798,N_15061,N_14477);
xnor U15799 (N_15799,N_14676,N_14576);
nor U15800 (N_15800,N_15172,N_14818);
nand U15801 (N_15801,N_15132,N_14811);
and U15802 (N_15802,N_14802,N_14555);
nor U15803 (N_15803,N_14416,N_14814);
xor U15804 (N_15804,N_14927,N_15018);
nor U15805 (N_15805,N_14580,N_14794);
and U15806 (N_15806,N_14484,N_14692);
or U15807 (N_15807,N_14905,N_14751);
xor U15808 (N_15808,N_14522,N_14911);
nand U15809 (N_15809,N_14650,N_14902);
and U15810 (N_15810,N_15116,N_15166);
and U15811 (N_15811,N_15112,N_14938);
xnor U15812 (N_15812,N_14943,N_14723);
nor U15813 (N_15813,N_15105,N_15091);
nand U15814 (N_15814,N_14829,N_15100);
xor U15815 (N_15815,N_15013,N_14766);
nand U15816 (N_15816,N_15156,N_14987);
nor U15817 (N_15817,N_14689,N_14872);
nor U15818 (N_15818,N_14624,N_15174);
xor U15819 (N_15819,N_14946,N_14881);
or U15820 (N_15820,N_14869,N_14647);
nor U15821 (N_15821,N_15093,N_14808);
nand U15822 (N_15822,N_14464,N_14688);
nand U15823 (N_15823,N_15055,N_14732);
or U15824 (N_15824,N_15100,N_14954);
xor U15825 (N_15825,N_15127,N_14702);
xnor U15826 (N_15826,N_14973,N_14860);
and U15827 (N_15827,N_15013,N_14736);
nor U15828 (N_15828,N_15058,N_14906);
nor U15829 (N_15829,N_14601,N_14550);
or U15830 (N_15830,N_15177,N_14549);
nor U15831 (N_15831,N_14488,N_15014);
nor U15832 (N_15832,N_14510,N_15119);
xnor U15833 (N_15833,N_14634,N_14656);
and U15834 (N_15834,N_14888,N_14933);
nor U15835 (N_15835,N_15025,N_14804);
and U15836 (N_15836,N_14683,N_15041);
xnor U15837 (N_15837,N_15004,N_14845);
or U15838 (N_15838,N_14905,N_14681);
and U15839 (N_15839,N_14859,N_14553);
xnor U15840 (N_15840,N_14812,N_14697);
nor U15841 (N_15841,N_14779,N_14639);
and U15842 (N_15842,N_14693,N_14516);
and U15843 (N_15843,N_14418,N_14501);
or U15844 (N_15844,N_14679,N_14582);
and U15845 (N_15845,N_14924,N_14621);
nor U15846 (N_15846,N_14546,N_14472);
and U15847 (N_15847,N_15164,N_14599);
or U15848 (N_15848,N_14472,N_14513);
or U15849 (N_15849,N_15146,N_14506);
xor U15850 (N_15850,N_14960,N_14683);
nor U15851 (N_15851,N_14734,N_14777);
and U15852 (N_15852,N_14589,N_14410);
xnor U15853 (N_15853,N_14955,N_15073);
nand U15854 (N_15854,N_14720,N_14555);
nand U15855 (N_15855,N_15104,N_14760);
nor U15856 (N_15856,N_14550,N_14656);
and U15857 (N_15857,N_14736,N_14669);
or U15858 (N_15858,N_15060,N_15108);
or U15859 (N_15859,N_14834,N_15155);
and U15860 (N_15860,N_15173,N_15168);
nor U15861 (N_15861,N_14821,N_14980);
nor U15862 (N_15862,N_14997,N_14440);
nand U15863 (N_15863,N_15115,N_14583);
or U15864 (N_15864,N_15135,N_14698);
nor U15865 (N_15865,N_14889,N_15083);
xor U15866 (N_15866,N_14621,N_15019);
xnor U15867 (N_15867,N_15044,N_15126);
nor U15868 (N_15868,N_15038,N_14442);
nor U15869 (N_15869,N_15150,N_14551);
nor U15870 (N_15870,N_15099,N_14467);
or U15871 (N_15871,N_14891,N_14739);
nor U15872 (N_15872,N_14429,N_14646);
xor U15873 (N_15873,N_14954,N_14418);
and U15874 (N_15874,N_15138,N_15070);
nor U15875 (N_15875,N_14646,N_15043);
nor U15876 (N_15876,N_14422,N_14754);
xor U15877 (N_15877,N_14920,N_15127);
or U15878 (N_15878,N_14822,N_14880);
or U15879 (N_15879,N_14656,N_15083);
nand U15880 (N_15880,N_15143,N_15046);
nor U15881 (N_15881,N_14816,N_14851);
or U15882 (N_15882,N_15030,N_15090);
xnor U15883 (N_15883,N_14665,N_14524);
xor U15884 (N_15884,N_14900,N_14559);
nor U15885 (N_15885,N_14551,N_15180);
xor U15886 (N_15886,N_14701,N_14768);
nand U15887 (N_15887,N_14967,N_14518);
and U15888 (N_15888,N_14547,N_14445);
nor U15889 (N_15889,N_14818,N_14877);
xor U15890 (N_15890,N_14493,N_14487);
xnor U15891 (N_15891,N_14529,N_14975);
or U15892 (N_15892,N_15177,N_14960);
nand U15893 (N_15893,N_14749,N_14964);
or U15894 (N_15894,N_14423,N_14890);
and U15895 (N_15895,N_15188,N_15111);
nor U15896 (N_15896,N_14772,N_14992);
xnor U15897 (N_15897,N_15128,N_14821);
and U15898 (N_15898,N_15016,N_15008);
or U15899 (N_15899,N_14893,N_14668);
or U15900 (N_15900,N_14878,N_14824);
or U15901 (N_15901,N_14727,N_15024);
or U15902 (N_15902,N_14720,N_15106);
xor U15903 (N_15903,N_14673,N_14523);
xor U15904 (N_15904,N_14454,N_14876);
nand U15905 (N_15905,N_14841,N_14540);
nand U15906 (N_15906,N_15003,N_14714);
nand U15907 (N_15907,N_14553,N_14441);
nor U15908 (N_15908,N_15156,N_14651);
nor U15909 (N_15909,N_14795,N_14436);
nand U15910 (N_15910,N_14598,N_14764);
nand U15911 (N_15911,N_14684,N_14879);
nand U15912 (N_15912,N_15098,N_14628);
nor U15913 (N_15913,N_14425,N_14844);
xor U15914 (N_15914,N_14462,N_14992);
nor U15915 (N_15915,N_14717,N_14635);
and U15916 (N_15916,N_14471,N_14570);
nor U15917 (N_15917,N_14568,N_14708);
or U15918 (N_15918,N_14860,N_14918);
nor U15919 (N_15919,N_14527,N_14628);
nor U15920 (N_15920,N_14417,N_14574);
and U15921 (N_15921,N_15162,N_14638);
or U15922 (N_15922,N_14592,N_14983);
and U15923 (N_15923,N_14974,N_15139);
and U15924 (N_15924,N_15147,N_15028);
and U15925 (N_15925,N_14972,N_14786);
and U15926 (N_15926,N_14575,N_14687);
and U15927 (N_15927,N_14926,N_14746);
xnor U15928 (N_15928,N_15057,N_14755);
nand U15929 (N_15929,N_15186,N_14943);
xor U15930 (N_15930,N_14901,N_14550);
and U15931 (N_15931,N_14761,N_14908);
xor U15932 (N_15932,N_15165,N_15086);
nand U15933 (N_15933,N_14831,N_14480);
xnor U15934 (N_15934,N_14466,N_14874);
nor U15935 (N_15935,N_14791,N_14632);
and U15936 (N_15936,N_14438,N_14924);
xnor U15937 (N_15937,N_14665,N_14595);
xor U15938 (N_15938,N_14614,N_14845);
xnor U15939 (N_15939,N_14796,N_15138);
nand U15940 (N_15940,N_15106,N_14623);
nor U15941 (N_15941,N_14835,N_14419);
and U15942 (N_15942,N_14990,N_14760);
xor U15943 (N_15943,N_14687,N_15158);
or U15944 (N_15944,N_14434,N_14440);
nand U15945 (N_15945,N_14499,N_15169);
xor U15946 (N_15946,N_14627,N_15180);
or U15947 (N_15947,N_15177,N_14972);
nor U15948 (N_15948,N_14649,N_14454);
and U15949 (N_15949,N_14578,N_14865);
nand U15950 (N_15950,N_14870,N_15082);
nor U15951 (N_15951,N_14879,N_14634);
nor U15952 (N_15952,N_14429,N_14659);
and U15953 (N_15953,N_14473,N_14433);
and U15954 (N_15954,N_14452,N_15069);
nor U15955 (N_15955,N_14847,N_14659);
xor U15956 (N_15956,N_14628,N_14667);
and U15957 (N_15957,N_14656,N_14858);
xnor U15958 (N_15958,N_14605,N_15038);
and U15959 (N_15959,N_14681,N_14850);
or U15960 (N_15960,N_14483,N_15191);
and U15961 (N_15961,N_14984,N_14490);
nor U15962 (N_15962,N_14643,N_15042);
xor U15963 (N_15963,N_14904,N_14572);
nand U15964 (N_15964,N_14542,N_14934);
and U15965 (N_15965,N_15113,N_14908);
nand U15966 (N_15966,N_15057,N_14914);
or U15967 (N_15967,N_14545,N_14734);
nand U15968 (N_15968,N_14742,N_14731);
nor U15969 (N_15969,N_14902,N_14948);
xnor U15970 (N_15970,N_14825,N_14497);
and U15971 (N_15971,N_15008,N_14464);
nor U15972 (N_15972,N_14923,N_14980);
or U15973 (N_15973,N_14804,N_14916);
nand U15974 (N_15974,N_14453,N_15163);
or U15975 (N_15975,N_15097,N_14762);
and U15976 (N_15976,N_14851,N_14508);
xnor U15977 (N_15977,N_14531,N_14867);
nand U15978 (N_15978,N_14551,N_14864);
or U15979 (N_15979,N_15090,N_14563);
nor U15980 (N_15980,N_14725,N_14628);
xor U15981 (N_15981,N_14834,N_15123);
nand U15982 (N_15982,N_14629,N_14785);
nand U15983 (N_15983,N_14716,N_14803);
nand U15984 (N_15984,N_15105,N_14728);
xor U15985 (N_15985,N_14949,N_14593);
nor U15986 (N_15986,N_14736,N_14995);
nor U15987 (N_15987,N_15020,N_15067);
and U15988 (N_15988,N_14475,N_15115);
xnor U15989 (N_15989,N_14554,N_14580);
and U15990 (N_15990,N_15113,N_14443);
xor U15991 (N_15991,N_14665,N_15006);
nand U15992 (N_15992,N_14580,N_14410);
or U15993 (N_15993,N_15195,N_14403);
and U15994 (N_15994,N_14673,N_14440);
nand U15995 (N_15995,N_15118,N_14459);
and U15996 (N_15996,N_14823,N_14706);
nand U15997 (N_15997,N_14682,N_14477);
and U15998 (N_15998,N_14841,N_14931);
or U15999 (N_15999,N_14434,N_15025);
xor U16000 (N_16000,N_15382,N_15450);
or U16001 (N_16001,N_15324,N_15448);
nand U16002 (N_16002,N_15378,N_15720);
xor U16003 (N_16003,N_15276,N_15733);
or U16004 (N_16004,N_15941,N_15731);
nor U16005 (N_16005,N_15607,N_15546);
or U16006 (N_16006,N_15833,N_15309);
and U16007 (N_16007,N_15999,N_15839);
and U16008 (N_16008,N_15690,N_15203);
nor U16009 (N_16009,N_15680,N_15218);
or U16010 (N_16010,N_15869,N_15238);
xor U16011 (N_16011,N_15580,N_15722);
nor U16012 (N_16012,N_15704,N_15740);
or U16013 (N_16013,N_15861,N_15511);
nand U16014 (N_16014,N_15591,N_15481);
or U16015 (N_16015,N_15856,N_15452);
nand U16016 (N_16016,N_15706,N_15292);
and U16017 (N_16017,N_15441,N_15639);
xor U16018 (N_16018,N_15295,N_15512);
or U16019 (N_16019,N_15700,N_15391);
xor U16020 (N_16020,N_15887,N_15709);
nand U16021 (N_16021,N_15201,N_15249);
xnor U16022 (N_16022,N_15883,N_15601);
xnor U16023 (N_16023,N_15810,N_15552);
nor U16024 (N_16024,N_15393,N_15818);
xor U16025 (N_16025,N_15348,N_15302);
nor U16026 (N_16026,N_15461,N_15220);
and U16027 (N_16027,N_15853,N_15350);
nor U16028 (N_16028,N_15975,N_15590);
and U16029 (N_16029,N_15241,N_15300);
nor U16030 (N_16030,N_15911,N_15236);
xor U16031 (N_16031,N_15945,N_15354);
and U16032 (N_16032,N_15368,N_15223);
nor U16033 (N_16033,N_15436,N_15778);
and U16034 (N_16034,N_15625,N_15390);
and U16035 (N_16035,N_15409,N_15652);
or U16036 (N_16036,N_15454,N_15529);
nand U16037 (N_16037,N_15206,N_15769);
nand U16038 (N_16038,N_15864,N_15268);
and U16039 (N_16039,N_15245,N_15782);
and U16040 (N_16040,N_15797,N_15741);
and U16041 (N_16041,N_15403,N_15247);
and U16042 (N_16042,N_15996,N_15669);
nand U16043 (N_16043,N_15521,N_15629);
xnor U16044 (N_16044,N_15832,N_15963);
xnor U16045 (N_16045,N_15272,N_15237);
xor U16046 (N_16046,N_15408,N_15347);
or U16047 (N_16047,N_15484,N_15998);
xnor U16048 (N_16048,N_15496,N_15688);
and U16049 (N_16049,N_15508,N_15421);
xnor U16050 (N_16050,N_15344,N_15352);
nand U16051 (N_16051,N_15240,N_15449);
xnor U16052 (N_16052,N_15848,N_15889);
xnor U16053 (N_16053,N_15312,N_15277);
xor U16054 (N_16054,N_15574,N_15678);
or U16055 (N_16055,N_15858,N_15894);
or U16056 (N_16056,N_15375,N_15359);
or U16057 (N_16057,N_15799,N_15684);
and U16058 (N_16058,N_15524,N_15432);
and U16059 (N_16059,N_15761,N_15985);
and U16060 (N_16060,N_15407,N_15619);
and U16061 (N_16061,N_15993,N_15673);
nor U16062 (N_16062,N_15980,N_15798);
xor U16063 (N_16063,N_15248,N_15573);
nor U16064 (N_16064,N_15310,N_15918);
nand U16065 (N_16065,N_15760,N_15746);
nand U16066 (N_16066,N_15751,N_15341);
or U16067 (N_16067,N_15982,N_15318);
or U16068 (N_16068,N_15472,N_15239);
xor U16069 (N_16069,N_15732,N_15228);
nor U16070 (N_16070,N_15465,N_15369);
nor U16071 (N_16071,N_15846,N_15708);
xnor U16072 (N_16072,N_15986,N_15557);
nor U16073 (N_16073,N_15565,N_15715);
and U16074 (N_16074,N_15577,N_15583);
xnor U16075 (N_16075,N_15306,N_15876);
or U16076 (N_16076,N_15230,N_15242);
or U16077 (N_16077,N_15801,N_15602);
nand U16078 (N_16078,N_15756,N_15243);
xor U16079 (N_16079,N_15891,N_15947);
or U16080 (N_16080,N_15303,N_15335);
or U16081 (N_16081,N_15812,N_15665);
nor U16082 (N_16082,N_15613,N_15938);
or U16083 (N_16083,N_15576,N_15545);
and U16084 (N_16084,N_15559,N_15860);
xor U16085 (N_16085,N_15518,N_15367);
xnor U16086 (N_16086,N_15528,N_15374);
or U16087 (N_16087,N_15547,N_15457);
nand U16088 (N_16088,N_15517,N_15763);
and U16089 (N_16089,N_15298,N_15498);
nor U16090 (N_16090,N_15264,N_15486);
xnor U16091 (N_16091,N_15867,N_15422);
nand U16092 (N_16092,N_15427,N_15762);
or U16093 (N_16093,N_15568,N_15890);
and U16094 (N_16094,N_15610,N_15476);
xnor U16095 (N_16095,N_15364,N_15519);
nand U16096 (N_16096,N_15903,N_15596);
nand U16097 (N_16097,N_15424,N_15345);
nor U16098 (N_16098,N_15253,N_15495);
nor U16099 (N_16099,N_15389,N_15330);
or U16100 (N_16100,N_15214,N_15500);
or U16101 (N_16101,N_15595,N_15322);
and U16102 (N_16102,N_15719,N_15850);
or U16103 (N_16103,N_15217,N_15614);
and U16104 (N_16104,N_15262,N_15716);
xnor U16105 (N_16105,N_15585,N_15200);
nand U16106 (N_16106,N_15668,N_15828);
and U16107 (N_16107,N_15387,N_15926);
and U16108 (N_16108,N_15328,N_15824);
or U16109 (N_16109,N_15718,N_15396);
xor U16110 (N_16110,N_15428,N_15429);
and U16111 (N_16111,N_15453,N_15466);
nand U16112 (N_16112,N_15935,N_15315);
and U16113 (N_16113,N_15777,N_15445);
and U16114 (N_16114,N_15728,N_15480);
or U16115 (N_16115,N_15994,N_15925);
and U16116 (N_16116,N_15632,N_15872);
nor U16117 (N_16117,N_15388,N_15488);
nand U16118 (N_16118,N_15263,N_15397);
xnor U16119 (N_16119,N_15906,N_15394);
and U16120 (N_16120,N_15736,N_15748);
nor U16121 (N_16121,N_15725,N_15927);
nand U16122 (N_16122,N_15807,N_15342);
nor U16123 (N_16123,N_15744,N_15995);
or U16124 (N_16124,N_15962,N_15331);
or U16125 (N_16125,N_15551,N_15923);
or U16126 (N_16126,N_15522,N_15990);
xor U16127 (N_16127,N_15535,N_15587);
nor U16128 (N_16128,N_15329,N_15550);
nand U16129 (N_16129,N_15685,N_15415);
xor U16130 (N_16130,N_15285,N_15384);
or U16131 (N_16131,N_15666,N_15877);
nand U16132 (N_16132,N_15664,N_15361);
or U16133 (N_16133,N_15738,N_15930);
nor U16134 (N_16134,N_15297,N_15489);
or U16135 (N_16135,N_15443,N_15575);
xor U16136 (N_16136,N_15537,N_15477);
or U16137 (N_16137,N_15785,N_15615);
xnor U16138 (N_16138,N_15660,N_15229);
nand U16139 (N_16139,N_15490,N_15793);
and U16140 (N_16140,N_15234,N_15808);
nand U16141 (N_16141,N_15600,N_15635);
nor U16142 (N_16142,N_15905,N_15997);
and U16143 (N_16143,N_15520,N_15705);
xnor U16144 (N_16144,N_15843,N_15571);
or U16145 (N_16145,N_15819,N_15696);
xor U16146 (N_16146,N_15916,N_15623);
and U16147 (N_16147,N_15321,N_15663);
xnor U16148 (N_16148,N_15789,N_15971);
nor U16149 (N_16149,N_15627,N_15724);
and U16150 (N_16150,N_15758,N_15989);
xor U16151 (N_16151,N_15928,N_15815);
xnor U16152 (N_16152,N_15346,N_15544);
xnor U16153 (N_16153,N_15540,N_15425);
and U16154 (N_16154,N_15464,N_15270);
or U16155 (N_16155,N_15514,N_15435);
xnor U16156 (N_16156,N_15558,N_15594);
nor U16157 (N_16157,N_15672,N_15659);
nor U16158 (N_16158,N_15420,N_15654);
nor U16159 (N_16159,N_15358,N_15325);
xor U16160 (N_16160,N_15714,N_15811);
nand U16161 (N_16161,N_15473,N_15697);
or U16162 (N_16162,N_15806,N_15569);
xor U16163 (N_16163,N_15699,N_15854);
or U16164 (N_16164,N_15878,N_15874);
nor U16165 (N_16165,N_15305,N_15339);
xor U16166 (N_16166,N_15842,N_15503);
nor U16167 (N_16167,N_15866,N_15379);
and U16168 (N_16168,N_15337,N_15363);
or U16169 (N_16169,N_15549,N_15957);
nor U16170 (N_16170,N_15702,N_15543);
or U16171 (N_16171,N_15536,N_15353);
nor U16172 (N_16172,N_15981,N_15759);
xor U16173 (N_16173,N_15216,N_15226);
xnor U16174 (N_16174,N_15636,N_15531);
and U16175 (N_16175,N_15266,N_15437);
nor U16176 (N_16176,N_15749,N_15460);
xor U16177 (N_16177,N_15717,N_15506);
nor U16178 (N_16178,N_15598,N_15556);
nand U16179 (N_16179,N_15648,N_15875);
and U16180 (N_16180,N_15934,N_15804);
nand U16181 (N_16181,N_15745,N_15323);
nor U16182 (N_16182,N_15852,N_15712);
nand U16183 (N_16183,N_15308,N_15616);
or U16184 (N_16184,N_15606,N_15661);
or U16185 (N_16185,N_15795,N_15676);
xor U16186 (N_16186,N_15294,N_15735);
or U16187 (N_16187,N_15265,N_15752);
xor U16188 (N_16188,N_15340,N_15829);
nor U16189 (N_16189,N_15786,N_15739);
or U16190 (N_16190,N_15917,N_15467);
xor U16191 (N_16191,N_15649,N_15965);
nand U16192 (N_16192,N_15973,N_15838);
nand U16193 (N_16193,N_15796,N_15929);
nand U16194 (N_16194,N_15611,N_15968);
nand U16195 (N_16195,N_15640,N_15682);
nor U16196 (N_16196,N_15386,N_15210);
xor U16197 (N_16197,N_15566,N_15820);
or U16198 (N_16198,N_15527,N_15775);
nand U16199 (N_16199,N_15356,N_15770);
xor U16200 (N_16200,N_15456,N_15561);
xor U16201 (N_16201,N_15401,N_15455);
and U16202 (N_16202,N_15937,N_15753);
nand U16203 (N_16203,N_15880,N_15225);
nor U16204 (N_16204,N_15711,N_15827);
xnor U16205 (N_16205,N_15686,N_15948);
or U16206 (N_16206,N_15320,N_15978);
xor U16207 (N_16207,N_15400,N_15539);
xnor U16208 (N_16208,N_15653,N_15922);
or U16209 (N_16209,N_15771,N_15416);
and U16210 (N_16210,N_15992,N_15683);
nand U16211 (N_16211,N_15642,N_15491);
xor U16212 (N_16212,N_15444,N_15754);
and U16213 (N_16213,N_15534,N_15553);
and U16214 (N_16214,N_15991,N_15822);
and U16215 (N_16215,N_15772,N_15689);
nor U16216 (N_16216,N_15723,N_15250);
nor U16217 (N_16217,N_15944,N_15841);
nor U16218 (N_16218,N_15211,N_15936);
or U16219 (N_16219,N_15376,N_15383);
and U16220 (N_16220,N_15398,N_15727);
xor U16221 (N_16221,N_15414,N_15451);
xnor U16222 (N_16222,N_15964,N_15279);
nor U16223 (N_16223,N_15902,N_15423);
or U16224 (N_16224,N_15482,N_15316);
or U16225 (N_16225,N_15913,N_15343);
or U16226 (N_16226,N_15261,N_15794);
and U16227 (N_16227,N_15621,N_15780);
xnor U16228 (N_16228,N_15586,N_15882);
and U16229 (N_16229,N_15943,N_15845);
and U16230 (N_16230,N_15821,N_15679);
or U16231 (N_16231,N_15644,N_15509);
xnor U16232 (N_16232,N_15442,N_15317);
xor U16233 (N_16233,N_15560,N_15492);
nand U16234 (N_16234,N_15515,N_15497);
or U16235 (N_16235,N_15202,N_15784);
xnor U16236 (N_16236,N_15939,N_15283);
nor U16237 (N_16237,N_15224,N_15662);
xor U16238 (N_16238,N_15251,N_15617);
or U16239 (N_16239,N_15419,N_15355);
xnor U16240 (N_16240,N_15701,N_15899);
nor U16241 (N_16241,N_15510,N_15286);
and U16242 (N_16242,N_15956,N_15499);
nand U16243 (N_16243,N_15212,N_15677);
nand U16244 (N_16244,N_15764,N_15458);
nor U16245 (N_16245,N_15380,N_15333);
xor U16246 (N_16246,N_15670,N_15260);
or U16247 (N_16247,N_15908,N_15319);
or U16248 (N_16248,N_15651,N_15966);
nor U16249 (N_16249,N_15823,N_15609);
xnor U16250 (N_16250,N_15879,N_15570);
xor U16251 (N_16251,N_15470,N_15630);
xnor U16252 (N_16252,N_15703,N_15479);
nand U16253 (N_16253,N_15800,N_15650);
or U16254 (N_16254,N_15513,N_15221);
or U16255 (N_16255,N_15658,N_15681);
and U16256 (N_16256,N_15667,N_15385);
xor U16257 (N_16257,N_15231,N_15641);
nor U16258 (N_16258,N_15931,N_15983);
and U16259 (N_16259,N_15525,N_15494);
and U16260 (N_16260,N_15284,N_15381);
xnor U16261 (N_16261,N_15884,N_15693);
xor U16262 (N_16262,N_15791,N_15781);
and U16263 (N_16263,N_15834,N_15919);
nand U16264 (N_16264,N_15671,N_15768);
and U16265 (N_16265,N_15817,N_15896);
xnor U16266 (N_16266,N_15411,N_15532);
and U16267 (N_16267,N_15447,N_15988);
nand U16268 (N_16268,N_15825,N_15232);
xnor U16269 (N_16269,N_15256,N_15504);
nand U16270 (N_16270,N_15213,N_15471);
nand U16271 (N_16271,N_15338,N_15773);
xnor U16272 (N_16272,N_15254,N_15618);
xnor U16273 (N_16273,N_15729,N_15293);
nor U16274 (N_16274,N_15402,N_15392);
nand U16275 (N_16275,N_15314,N_15326);
xor U16276 (N_16276,N_15507,N_15886);
or U16277 (N_16277,N_15656,N_15205);
nor U16278 (N_16278,N_15430,N_15707);
and U16279 (N_16279,N_15307,N_15940);
xnor U16280 (N_16280,N_15603,N_15222);
and U16281 (N_16281,N_15269,N_15755);
xnor U16282 (N_16282,N_15438,N_15564);
nand U16283 (N_16283,N_15372,N_15984);
nand U16284 (N_16284,N_15855,N_15687);
or U16285 (N_16285,N_15439,N_15410);
nor U16286 (N_16286,N_15478,N_15579);
or U16287 (N_16287,N_15485,N_15357);
nand U16288 (N_16288,N_15204,N_15459);
and U16289 (N_16289,N_15892,N_15592);
xor U16290 (N_16290,N_15790,N_15960);
xnor U16291 (N_16291,N_15961,N_15933);
xnor U16292 (N_16292,N_15301,N_15967);
nand U16293 (N_16293,N_15267,N_15362);
or U16294 (N_16294,N_15446,N_15351);
nand U16295 (N_16295,N_15802,N_15502);
nand U16296 (N_16296,N_15788,N_15493);
nor U16297 (N_16297,N_15840,N_15949);
nor U16298 (N_16298,N_15207,N_15851);
and U16299 (N_16299,N_15914,N_15969);
and U16300 (N_16300,N_15275,N_15831);
nor U16301 (N_16301,N_15563,N_15730);
nor U16302 (N_16302,N_15313,N_15692);
nand U16303 (N_16303,N_15645,N_15377);
nor U16304 (N_16304,N_15244,N_15505);
xor U16305 (N_16305,N_15783,N_15258);
or U16306 (N_16306,N_15885,N_15721);
nand U16307 (N_16307,N_15849,N_15255);
nand U16308 (N_16308,N_15291,N_15516);
nor U16309 (N_16309,N_15288,N_15950);
xor U16310 (N_16310,N_15900,N_15897);
nor U16311 (N_16311,N_15920,N_15915);
or U16312 (N_16312,N_15501,N_15647);
or U16313 (N_16313,N_15826,N_15259);
xnor U16314 (N_16314,N_15646,N_15273);
nor U16315 (N_16315,N_15628,N_15593);
nand U16316 (N_16316,N_15582,N_15958);
nand U16317 (N_16317,N_15694,N_15541);
and U16318 (N_16318,N_15757,N_15208);
and U16319 (N_16319,N_15475,N_15624);
or U16320 (N_16320,N_15219,N_15526);
xnor U16321 (N_16321,N_15533,N_15530);
nand U16322 (N_16322,N_15280,N_15742);
xnor U16323 (N_16323,N_15743,N_15463);
and U16324 (N_16324,N_15979,N_15296);
and U16325 (N_16325,N_15898,N_15909);
and U16326 (N_16326,N_15835,N_15523);
and U16327 (N_16327,N_15830,N_15257);
or U16328 (N_16328,N_15572,N_15698);
nand U16329 (N_16329,N_15987,N_15578);
and U16330 (N_16330,N_15584,N_15946);
or U16331 (N_16331,N_15766,N_15637);
nor U16332 (N_16332,N_15332,N_15888);
and U16333 (N_16333,N_15299,N_15336);
and U16334 (N_16334,N_15589,N_15695);
or U16335 (N_16335,N_15859,N_15976);
nand U16336 (N_16336,N_15562,N_15538);
xor U16337 (N_16337,N_15863,N_15622);
or U16338 (N_16338,N_15774,N_15483);
and U16339 (N_16339,N_15893,N_15554);
nand U16340 (N_16340,N_15787,N_15281);
nand U16341 (N_16341,N_15462,N_15952);
nand U16342 (N_16342,N_15548,N_15765);
xnor U16343 (N_16343,N_15809,N_15776);
nor U16344 (N_16344,N_15881,N_15953);
and U16345 (N_16345,N_15921,N_15803);
nand U16346 (N_16346,N_15873,N_15816);
nor U16347 (N_16347,N_15311,N_15734);
nand U16348 (N_16348,N_15417,N_15404);
xnor U16349 (N_16349,N_15413,N_15371);
and U16350 (N_16350,N_15691,N_15779);
nand U16351 (N_16351,N_15370,N_15274);
nor U16352 (N_16352,N_15209,N_15418);
xor U16353 (N_16353,N_15895,N_15638);
nand U16354 (N_16354,N_15868,N_15278);
xor U16355 (N_16355,N_15227,N_15626);
nor U16356 (N_16356,N_15657,N_15542);
and U16357 (N_16357,N_15907,N_15327);
or U16358 (N_16358,N_15951,N_15431);
nor U16359 (N_16359,N_15862,N_15360);
xnor U16360 (N_16360,N_15633,N_15954);
nor U16361 (N_16361,N_15870,N_15282);
xnor U16362 (N_16362,N_15910,N_15289);
xnor U16363 (N_16363,N_15612,N_15631);
and U16364 (N_16364,N_15901,N_15912);
or U16365 (N_16365,N_15836,N_15567);
nand U16366 (N_16366,N_15674,N_15865);
xnor U16367 (N_16367,N_15252,N_15837);
nand U16368 (N_16368,N_15747,N_15487);
nand U16369 (N_16369,N_15290,N_15599);
xor U16370 (N_16370,N_15271,N_15871);
nor U16371 (N_16371,N_15365,N_15726);
nand U16372 (N_16372,N_15399,N_15334);
or U16373 (N_16373,N_15395,N_15970);
nor U16374 (N_16374,N_15959,N_15235);
nor U16375 (N_16375,N_15433,N_15434);
xnor U16376 (N_16376,N_15468,N_15844);
nor U16377 (N_16377,N_15366,N_15977);
nor U16378 (N_16378,N_15974,N_15608);
nand U16379 (N_16379,N_15942,N_15604);
nand U16380 (N_16380,N_15634,N_15737);
nor U16381 (N_16381,N_15955,N_15767);
or U16382 (N_16382,N_15373,N_15713);
nor U16383 (N_16383,N_15932,N_15847);
nand U16384 (N_16384,N_15405,N_15792);
and U16385 (N_16385,N_15233,N_15675);
and U16386 (N_16386,N_15426,N_15474);
nor U16387 (N_16387,N_15655,N_15750);
nand U16388 (N_16388,N_15620,N_15588);
and U16389 (N_16389,N_15246,N_15349);
or U16390 (N_16390,N_15924,N_15406);
nor U16391 (N_16391,N_15440,N_15814);
and U16392 (N_16392,N_15555,N_15972);
and U16393 (N_16393,N_15857,N_15581);
or U16394 (N_16394,N_15904,N_15469);
nor U16395 (N_16395,N_15412,N_15643);
xor U16396 (N_16396,N_15287,N_15605);
and U16397 (N_16397,N_15710,N_15597);
or U16398 (N_16398,N_15304,N_15813);
xor U16399 (N_16399,N_15215,N_15805);
nand U16400 (N_16400,N_15994,N_15744);
and U16401 (N_16401,N_15532,N_15387);
nand U16402 (N_16402,N_15420,N_15778);
xor U16403 (N_16403,N_15933,N_15712);
nor U16404 (N_16404,N_15760,N_15408);
or U16405 (N_16405,N_15433,N_15806);
nor U16406 (N_16406,N_15512,N_15814);
and U16407 (N_16407,N_15311,N_15342);
or U16408 (N_16408,N_15211,N_15360);
nor U16409 (N_16409,N_15695,N_15917);
xnor U16410 (N_16410,N_15409,N_15209);
xor U16411 (N_16411,N_15429,N_15462);
or U16412 (N_16412,N_15250,N_15714);
and U16413 (N_16413,N_15916,N_15430);
nor U16414 (N_16414,N_15381,N_15236);
xor U16415 (N_16415,N_15696,N_15475);
or U16416 (N_16416,N_15317,N_15444);
and U16417 (N_16417,N_15417,N_15739);
or U16418 (N_16418,N_15232,N_15569);
nand U16419 (N_16419,N_15842,N_15501);
and U16420 (N_16420,N_15725,N_15251);
and U16421 (N_16421,N_15387,N_15918);
nor U16422 (N_16422,N_15455,N_15309);
nor U16423 (N_16423,N_15533,N_15406);
and U16424 (N_16424,N_15563,N_15835);
and U16425 (N_16425,N_15400,N_15845);
nand U16426 (N_16426,N_15524,N_15310);
nor U16427 (N_16427,N_15740,N_15759);
nand U16428 (N_16428,N_15703,N_15869);
and U16429 (N_16429,N_15618,N_15837);
nor U16430 (N_16430,N_15865,N_15363);
nor U16431 (N_16431,N_15890,N_15864);
nor U16432 (N_16432,N_15611,N_15747);
or U16433 (N_16433,N_15447,N_15604);
nor U16434 (N_16434,N_15857,N_15646);
nor U16435 (N_16435,N_15921,N_15888);
and U16436 (N_16436,N_15290,N_15638);
xnor U16437 (N_16437,N_15768,N_15474);
nand U16438 (N_16438,N_15514,N_15468);
xor U16439 (N_16439,N_15596,N_15658);
xor U16440 (N_16440,N_15505,N_15939);
xnor U16441 (N_16441,N_15849,N_15566);
and U16442 (N_16442,N_15861,N_15365);
nand U16443 (N_16443,N_15578,N_15872);
nand U16444 (N_16444,N_15270,N_15616);
xor U16445 (N_16445,N_15864,N_15834);
or U16446 (N_16446,N_15278,N_15888);
nor U16447 (N_16447,N_15995,N_15316);
or U16448 (N_16448,N_15601,N_15957);
or U16449 (N_16449,N_15928,N_15235);
and U16450 (N_16450,N_15627,N_15546);
or U16451 (N_16451,N_15813,N_15689);
and U16452 (N_16452,N_15460,N_15259);
xor U16453 (N_16453,N_15653,N_15345);
xor U16454 (N_16454,N_15368,N_15651);
xnor U16455 (N_16455,N_15986,N_15569);
or U16456 (N_16456,N_15792,N_15723);
nand U16457 (N_16457,N_15434,N_15472);
nand U16458 (N_16458,N_15611,N_15356);
nand U16459 (N_16459,N_15644,N_15976);
xnor U16460 (N_16460,N_15774,N_15279);
xnor U16461 (N_16461,N_15535,N_15335);
xor U16462 (N_16462,N_15255,N_15446);
xnor U16463 (N_16463,N_15705,N_15788);
nor U16464 (N_16464,N_15873,N_15326);
nor U16465 (N_16465,N_15333,N_15727);
xnor U16466 (N_16466,N_15928,N_15370);
or U16467 (N_16467,N_15783,N_15238);
nor U16468 (N_16468,N_15674,N_15510);
or U16469 (N_16469,N_15331,N_15604);
and U16470 (N_16470,N_15585,N_15586);
nor U16471 (N_16471,N_15998,N_15669);
nand U16472 (N_16472,N_15565,N_15532);
or U16473 (N_16473,N_15270,N_15501);
and U16474 (N_16474,N_15601,N_15941);
nand U16475 (N_16475,N_15607,N_15389);
or U16476 (N_16476,N_15571,N_15896);
nand U16477 (N_16477,N_15418,N_15837);
and U16478 (N_16478,N_15455,N_15808);
nand U16479 (N_16479,N_15225,N_15399);
nand U16480 (N_16480,N_15940,N_15924);
and U16481 (N_16481,N_15994,N_15364);
nor U16482 (N_16482,N_15941,N_15690);
nor U16483 (N_16483,N_15974,N_15630);
nand U16484 (N_16484,N_15555,N_15934);
or U16485 (N_16485,N_15676,N_15864);
nor U16486 (N_16486,N_15296,N_15358);
or U16487 (N_16487,N_15277,N_15789);
nand U16488 (N_16488,N_15336,N_15982);
nor U16489 (N_16489,N_15697,N_15226);
and U16490 (N_16490,N_15248,N_15220);
or U16491 (N_16491,N_15747,N_15431);
nor U16492 (N_16492,N_15292,N_15626);
nor U16493 (N_16493,N_15996,N_15210);
or U16494 (N_16494,N_15508,N_15446);
xor U16495 (N_16495,N_15533,N_15719);
nor U16496 (N_16496,N_15518,N_15979);
nor U16497 (N_16497,N_15203,N_15968);
nand U16498 (N_16498,N_15222,N_15908);
nand U16499 (N_16499,N_15709,N_15863);
and U16500 (N_16500,N_15563,N_15296);
nand U16501 (N_16501,N_15235,N_15776);
nand U16502 (N_16502,N_15297,N_15528);
nand U16503 (N_16503,N_15615,N_15319);
nor U16504 (N_16504,N_15752,N_15528);
nor U16505 (N_16505,N_15519,N_15295);
and U16506 (N_16506,N_15895,N_15371);
nor U16507 (N_16507,N_15435,N_15971);
and U16508 (N_16508,N_15695,N_15997);
nand U16509 (N_16509,N_15776,N_15908);
and U16510 (N_16510,N_15759,N_15723);
and U16511 (N_16511,N_15646,N_15673);
and U16512 (N_16512,N_15627,N_15642);
nor U16513 (N_16513,N_15624,N_15416);
and U16514 (N_16514,N_15200,N_15657);
nor U16515 (N_16515,N_15308,N_15203);
nor U16516 (N_16516,N_15683,N_15928);
or U16517 (N_16517,N_15844,N_15288);
nand U16518 (N_16518,N_15745,N_15789);
nand U16519 (N_16519,N_15413,N_15745);
nand U16520 (N_16520,N_15441,N_15323);
nor U16521 (N_16521,N_15611,N_15344);
or U16522 (N_16522,N_15877,N_15584);
nand U16523 (N_16523,N_15341,N_15806);
xnor U16524 (N_16524,N_15626,N_15271);
and U16525 (N_16525,N_15394,N_15946);
and U16526 (N_16526,N_15690,N_15202);
nor U16527 (N_16527,N_15748,N_15593);
nand U16528 (N_16528,N_15646,N_15950);
or U16529 (N_16529,N_15228,N_15734);
nor U16530 (N_16530,N_15780,N_15326);
nor U16531 (N_16531,N_15357,N_15403);
nand U16532 (N_16532,N_15769,N_15763);
nand U16533 (N_16533,N_15886,N_15822);
nor U16534 (N_16534,N_15745,N_15687);
nand U16535 (N_16535,N_15882,N_15754);
nand U16536 (N_16536,N_15634,N_15340);
nand U16537 (N_16537,N_15497,N_15580);
xnor U16538 (N_16538,N_15966,N_15617);
and U16539 (N_16539,N_15653,N_15271);
nor U16540 (N_16540,N_15475,N_15201);
nand U16541 (N_16541,N_15561,N_15424);
nand U16542 (N_16542,N_15798,N_15822);
or U16543 (N_16543,N_15280,N_15677);
or U16544 (N_16544,N_15630,N_15666);
nor U16545 (N_16545,N_15233,N_15973);
nand U16546 (N_16546,N_15370,N_15987);
and U16547 (N_16547,N_15990,N_15498);
xor U16548 (N_16548,N_15592,N_15828);
xor U16549 (N_16549,N_15807,N_15754);
nand U16550 (N_16550,N_15553,N_15219);
xor U16551 (N_16551,N_15490,N_15702);
nand U16552 (N_16552,N_15485,N_15920);
or U16553 (N_16553,N_15649,N_15714);
nor U16554 (N_16554,N_15655,N_15722);
or U16555 (N_16555,N_15998,N_15961);
xnor U16556 (N_16556,N_15668,N_15872);
nand U16557 (N_16557,N_15507,N_15268);
nand U16558 (N_16558,N_15804,N_15328);
xnor U16559 (N_16559,N_15684,N_15613);
nor U16560 (N_16560,N_15713,N_15798);
nand U16561 (N_16561,N_15497,N_15662);
nand U16562 (N_16562,N_15417,N_15440);
or U16563 (N_16563,N_15559,N_15479);
nand U16564 (N_16564,N_15952,N_15903);
and U16565 (N_16565,N_15755,N_15495);
nor U16566 (N_16566,N_15467,N_15794);
or U16567 (N_16567,N_15946,N_15314);
nor U16568 (N_16568,N_15643,N_15910);
or U16569 (N_16569,N_15367,N_15666);
or U16570 (N_16570,N_15717,N_15551);
nor U16571 (N_16571,N_15463,N_15594);
nor U16572 (N_16572,N_15813,N_15355);
nand U16573 (N_16573,N_15979,N_15779);
xnor U16574 (N_16574,N_15538,N_15919);
xor U16575 (N_16575,N_15816,N_15741);
nand U16576 (N_16576,N_15643,N_15447);
nand U16577 (N_16577,N_15373,N_15210);
nor U16578 (N_16578,N_15674,N_15411);
and U16579 (N_16579,N_15249,N_15213);
or U16580 (N_16580,N_15654,N_15505);
xnor U16581 (N_16581,N_15792,N_15452);
and U16582 (N_16582,N_15631,N_15960);
nor U16583 (N_16583,N_15329,N_15774);
nor U16584 (N_16584,N_15927,N_15916);
xnor U16585 (N_16585,N_15261,N_15658);
xor U16586 (N_16586,N_15989,N_15486);
nor U16587 (N_16587,N_15754,N_15287);
nor U16588 (N_16588,N_15570,N_15351);
nand U16589 (N_16589,N_15375,N_15704);
nand U16590 (N_16590,N_15350,N_15767);
or U16591 (N_16591,N_15465,N_15989);
xor U16592 (N_16592,N_15643,N_15956);
xnor U16593 (N_16593,N_15627,N_15445);
and U16594 (N_16594,N_15504,N_15870);
xnor U16595 (N_16595,N_15888,N_15480);
nand U16596 (N_16596,N_15965,N_15567);
nor U16597 (N_16597,N_15798,N_15363);
nor U16598 (N_16598,N_15319,N_15691);
or U16599 (N_16599,N_15806,N_15729);
xor U16600 (N_16600,N_15315,N_15733);
or U16601 (N_16601,N_15460,N_15805);
nand U16602 (N_16602,N_15437,N_15713);
or U16603 (N_16603,N_15490,N_15303);
nor U16604 (N_16604,N_15761,N_15436);
or U16605 (N_16605,N_15547,N_15842);
xor U16606 (N_16606,N_15835,N_15689);
nor U16607 (N_16607,N_15582,N_15609);
and U16608 (N_16608,N_15244,N_15243);
or U16609 (N_16609,N_15680,N_15543);
or U16610 (N_16610,N_15348,N_15583);
nor U16611 (N_16611,N_15902,N_15722);
xor U16612 (N_16612,N_15875,N_15659);
xnor U16613 (N_16613,N_15365,N_15882);
xor U16614 (N_16614,N_15697,N_15901);
or U16615 (N_16615,N_15271,N_15999);
nor U16616 (N_16616,N_15858,N_15721);
nor U16617 (N_16617,N_15213,N_15528);
nor U16618 (N_16618,N_15846,N_15285);
xnor U16619 (N_16619,N_15815,N_15937);
nand U16620 (N_16620,N_15955,N_15303);
nand U16621 (N_16621,N_15782,N_15361);
nand U16622 (N_16622,N_15338,N_15388);
xor U16623 (N_16623,N_15617,N_15242);
or U16624 (N_16624,N_15901,N_15395);
nand U16625 (N_16625,N_15304,N_15544);
and U16626 (N_16626,N_15226,N_15868);
xor U16627 (N_16627,N_15720,N_15218);
nand U16628 (N_16628,N_15469,N_15934);
nand U16629 (N_16629,N_15692,N_15761);
xnor U16630 (N_16630,N_15952,N_15586);
or U16631 (N_16631,N_15351,N_15461);
nand U16632 (N_16632,N_15897,N_15378);
and U16633 (N_16633,N_15923,N_15957);
nor U16634 (N_16634,N_15318,N_15495);
and U16635 (N_16635,N_15459,N_15429);
xnor U16636 (N_16636,N_15456,N_15892);
or U16637 (N_16637,N_15780,N_15338);
nor U16638 (N_16638,N_15254,N_15294);
or U16639 (N_16639,N_15638,N_15855);
nand U16640 (N_16640,N_15982,N_15225);
xor U16641 (N_16641,N_15723,N_15529);
or U16642 (N_16642,N_15762,N_15701);
xnor U16643 (N_16643,N_15931,N_15234);
xnor U16644 (N_16644,N_15760,N_15634);
or U16645 (N_16645,N_15226,N_15361);
and U16646 (N_16646,N_15830,N_15498);
nor U16647 (N_16647,N_15499,N_15774);
or U16648 (N_16648,N_15881,N_15566);
and U16649 (N_16649,N_15992,N_15448);
nor U16650 (N_16650,N_15283,N_15989);
xor U16651 (N_16651,N_15400,N_15755);
and U16652 (N_16652,N_15858,N_15421);
nand U16653 (N_16653,N_15251,N_15230);
nor U16654 (N_16654,N_15573,N_15581);
or U16655 (N_16655,N_15848,N_15264);
or U16656 (N_16656,N_15217,N_15372);
nand U16657 (N_16657,N_15852,N_15918);
or U16658 (N_16658,N_15260,N_15846);
nor U16659 (N_16659,N_15549,N_15582);
nand U16660 (N_16660,N_15756,N_15352);
nand U16661 (N_16661,N_15239,N_15431);
or U16662 (N_16662,N_15983,N_15627);
nor U16663 (N_16663,N_15913,N_15856);
and U16664 (N_16664,N_15289,N_15858);
nor U16665 (N_16665,N_15594,N_15879);
or U16666 (N_16666,N_15233,N_15470);
nand U16667 (N_16667,N_15412,N_15799);
xnor U16668 (N_16668,N_15946,N_15638);
nor U16669 (N_16669,N_15311,N_15531);
nand U16670 (N_16670,N_15619,N_15712);
nor U16671 (N_16671,N_15260,N_15698);
nand U16672 (N_16672,N_15329,N_15622);
and U16673 (N_16673,N_15301,N_15239);
xnor U16674 (N_16674,N_15449,N_15760);
nand U16675 (N_16675,N_15593,N_15333);
or U16676 (N_16676,N_15336,N_15922);
and U16677 (N_16677,N_15250,N_15654);
or U16678 (N_16678,N_15394,N_15308);
xnor U16679 (N_16679,N_15888,N_15719);
or U16680 (N_16680,N_15321,N_15312);
nor U16681 (N_16681,N_15681,N_15952);
or U16682 (N_16682,N_15981,N_15574);
and U16683 (N_16683,N_15684,N_15756);
xnor U16684 (N_16684,N_15410,N_15340);
nand U16685 (N_16685,N_15764,N_15584);
xor U16686 (N_16686,N_15844,N_15933);
and U16687 (N_16687,N_15887,N_15427);
nor U16688 (N_16688,N_15574,N_15757);
nand U16689 (N_16689,N_15314,N_15954);
xnor U16690 (N_16690,N_15447,N_15945);
xor U16691 (N_16691,N_15907,N_15670);
nand U16692 (N_16692,N_15395,N_15411);
nand U16693 (N_16693,N_15362,N_15403);
nand U16694 (N_16694,N_15568,N_15955);
nor U16695 (N_16695,N_15321,N_15262);
nand U16696 (N_16696,N_15238,N_15735);
or U16697 (N_16697,N_15983,N_15279);
and U16698 (N_16698,N_15859,N_15675);
nand U16699 (N_16699,N_15884,N_15711);
nand U16700 (N_16700,N_15840,N_15315);
and U16701 (N_16701,N_15451,N_15924);
xnor U16702 (N_16702,N_15986,N_15647);
nand U16703 (N_16703,N_15631,N_15785);
and U16704 (N_16704,N_15337,N_15410);
and U16705 (N_16705,N_15759,N_15755);
nand U16706 (N_16706,N_15693,N_15315);
nand U16707 (N_16707,N_15472,N_15683);
nor U16708 (N_16708,N_15661,N_15968);
nand U16709 (N_16709,N_15554,N_15453);
nor U16710 (N_16710,N_15854,N_15883);
xnor U16711 (N_16711,N_15604,N_15842);
nor U16712 (N_16712,N_15496,N_15415);
or U16713 (N_16713,N_15682,N_15282);
xnor U16714 (N_16714,N_15355,N_15627);
xor U16715 (N_16715,N_15736,N_15344);
nor U16716 (N_16716,N_15502,N_15788);
or U16717 (N_16717,N_15371,N_15329);
or U16718 (N_16718,N_15285,N_15359);
nand U16719 (N_16719,N_15952,N_15208);
nor U16720 (N_16720,N_15690,N_15877);
and U16721 (N_16721,N_15321,N_15648);
nor U16722 (N_16722,N_15554,N_15219);
nor U16723 (N_16723,N_15576,N_15420);
and U16724 (N_16724,N_15820,N_15362);
xnor U16725 (N_16725,N_15674,N_15445);
and U16726 (N_16726,N_15521,N_15216);
xnor U16727 (N_16727,N_15742,N_15484);
and U16728 (N_16728,N_15233,N_15731);
and U16729 (N_16729,N_15629,N_15766);
or U16730 (N_16730,N_15771,N_15800);
xor U16731 (N_16731,N_15599,N_15472);
xor U16732 (N_16732,N_15720,N_15437);
xor U16733 (N_16733,N_15889,N_15271);
nor U16734 (N_16734,N_15933,N_15344);
nand U16735 (N_16735,N_15665,N_15467);
xnor U16736 (N_16736,N_15683,N_15457);
and U16737 (N_16737,N_15967,N_15820);
or U16738 (N_16738,N_15750,N_15854);
xnor U16739 (N_16739,N_15457,N_15969);
xor U16740 (N_16740,N_15918,N_15780);
nor U16741 (N_16741,N_15870,N_15871);
xor U16742 (N_16742,N_15343,N_15357);
xor U16743 (N_16743,N_15731,N_15865);
nor U16744 (N_16744,N_15558,N_15525);
and U16745 (N_16745,N_15517,N_15925);
xor U16746 (N_16746,N_15525,N_15446);
nand U16747 (N_16747,N_15654,N_15226);
nand U16748 (N_16748,N_15601,N_15367);
xnor U16749 (N_16749,N_15466,N_15292);
nor U16750 (N_16750,N_15309,N_15708);
nor U16751 (N_16751,N_15334,N_15733);
or U16752 (N_16752,N_15427,N_15496);
nand U16753 (N_16753,N_15368,N_15676);
or U16754 (N_16754,N_15543,N_15341);
xor U16755 (N_16755,N_15957,N_15848);
and U16756 (N_16756,N_15235,N_15428);
xnor U16757 (N_16757,N_15737,N_15694);
xnor U16758 (N_16758,N_15305,N_15872);
nand U16759 (N_16759,N_15230,N_15572);
nor U16760 (N_16760,N_15892,N_15653);
or U16761 (N_16761,N_15341,N_15650);
nand U16762 (N_16762,N_15720,N_15739);
nor U16763 (N_16763,N_15868,N_15780);
xnor U16764 (N_16764,N_15824,N_15878);
nor U16765 (N_16765,N_15338,N_15799);
nor U16766 (N_16766,N_15726,N_15292);
nor U16767 (N_16767,N_15599,N_15380);
or U16768 (N_16768,N_15600,N_15529);
xnor U16769 (N_16769,N_15641,N_15794);
and U16770 (N_16770,N_15777,N_15441);
xnor U16771 (N_16771,N_15601,N_15536);
nand U16772 (N_16772,N_15634,N_15369);
or U16773 (N_16773,N_15291,N_15844);
or U16774 (N_16774,N_15862,N_15890);
and U16775 (N_16775,N_15441,N_15517);
xor U16776 (N_16776,N_15363,N_15284);
xor U16777 (N_16777,N_15341,N_15251);
nor U16778 (N_16778,N_15397,N_15784);
and U16779 (N_16779,N_15847,N_15828);
nand U16780 (N_16780,N_15538,N_15443);
nor U16781 (N_16781,N_15782,N_15648);
or U16782 (N_16782,N_15502,N_15406);
nor U16783 (N_16783,N_15668,N_15927);
and U16784 (N_16784,N_15962,N_15407);
xnor U16785 (N_16785,N_15645,N_15927);
or U16786 (N_16786,N_15660,N_15272);
nand U16787 (N_16787,N_15413,N_15469);
xor U16788 (N_16788,N_15873,N_15897);
nor U16789 (N_16789,N_15439,N_15583);
xor U16790 (N_16790,N_15489,N_15277);
or U16791 (N_16791,N_15486,N_15752);
nor U16792 (N_16792,N_15238,N_15911);
xor U16793 (N_16793,N_15633,N_15419);
nor U16794 (N_16794,N_15650,N_15248);
xor U16795 (N_16795,N_15988,N_15395);
nand U16796 (N_16796,N_15394,N_15583);
nor U16797 (N_16797,N_15947,N_15612);
or U16798 (N_16798,N_15995,N_15757);
and U16799 (N_16799,N_15365,N_15684);
nand U16800 (N_16800,N_16360,N_16567);
xor U16801 (N_16801,N_16749,N_16337);
nor U16802 (N_16802,N_16027,N_16153);
xnor U16803 (N_16803,N_16720,N_16335);
nor U16804 (N_16804,N_16293,N_16223);
nor U16805 (N_16805,N_16588,N_16002);
xor U16806 (N_16806,N_16592,N_16517);
nand U16807 (N_16807,N_16549,N_16776);
xnor U16808 (N_16808,N_16375,N_16751);
nand U16809 (N_16809,N_16119,N_16650);
or U16810 (N_16810,N_16186,N_16409);
nor U16811 (N_16811,N_16563,N_16421);
nand U16812 (N_16812,N_16265,N_16458);
nor U16813 (N_16813,N_16077,N_16114);
and U16814 (N_16814,N_16759,N_16757);
nand U16815 (N_16815,N_16767,N_16454);
nand U16816 (N_16816,N_16770,N_16343);
nand U16817 (N_16817,N_16593,N_16516);
or U16818 (N_16818,N_16134,N_16161);
or U16819 (N_16819,N_16124,N_16699);
or U16820 (N_16820,N_16345,N_16208);
and U16821 (N_16821,N_16664,N_16475);
or U16822 (N_16822,N_16457,N_16294);
nand U16823 (N_16823,N_16729,N_16175);
nor U16824 (N_16824,N_16012,N_16507);
and U16825 (N_16825,N_16427,N_16222);
or U16826 (N_16826,N_16255,N_16308);
nor U16827 (N_16827,N_16341,N_16403);
nor U16828 (N_16828,N_16607,N_16067);
nand U16829 (N_16829,N_16252,N_16756);
and U16830 (N_16830,N_16399,N_16116);
or U16831 (N_16831,N_16526,N_16111);
nor U16832 (N_16832,N_16416,N_16383);
nand U16833 (N_16833,N_16750,N_16311);
and U16834 (N_16834,N_16589,N_16371);
or U16835 (N_16835,N_16629,N_16227);
or U16836 (N_16836,N_16211,N_16347);
xor U16837 (N_16837,N_16667,N_16071);
or U16838 (N_16838,N_16774,N_16064);
xnor U16839 (N_16839,N_16641,N_16519);
nand U16840 (N_16840,N_16103,N_16669);
or U16841 (N_16841,N_16238,N_16673);
nand U16842 (N_16842,N_16556,N_16105);
nor U16843 (N_16843,N_16418,N_16039);
xor U16844 (N_16844,N_16697,N_16781);
and U16845 (N_16845,N_16069,N_16397);
nand U16846 (N_16846,N_16166,N_16484);
nand U16847 (N_16847,N_16497,N_16769);
and U16848 (N_16848,N_16730,N_16796);
xor U16849 (N_16849,N_16483,N_16711);
xor U16850 (N_16850,N_16180,N_16553);
xnor U16851 (N_16851,N_16561,N_16679);
nand U16852 (N_16852,N_16368,N_16083);
nor U16853 (N_16853,N_16339,N_16110);
or U16854 (N_16854,N_16286,N_16163);
nand U16855 (N_16855,N_16572,N_16499);
or U16856 (N_16856,N_16511,N_16419);
nand U16857 (N_16857,N_16194,N_16538);
nand U16858 (N_16858,N_16634,N_16537);
xnor U16859 (N_16859,N_16018,N_16192);
xnor U16860 (N_16860,N_16213,N_16173);
and U16861 (N_16861,N_16212,N_16521);
and U16862 (N_16862,N_16266,N_16564);
and U16863 (N_16863,N_16098,N_16178);
nor U16864 (N_16864,N_16491,N_16530);
nand U16865 (N_16865,N_16414,N_16482);
or U16866 (N_16866,N_16702,N_16113);
nor U16867 (N_16867,N_16696,N_16102);
or U16868 (N_16868,N_16226,N_16628);
and U16869 (N_16869,N_16554,N_16658);
xnor U16870 (N_16870,N_16682,N_16181);
nand U16871 (N_16871,N_16787,N_16406);
nor U16872 (N_16872,N_16512,N_16498);
nand U16873 (N_16873,N_16108,N_16599);
xor U16874 (N_16874,N_16202,N_16616);
or U16875 (N_16875,N_16237,N_16468);
nand U16876 (N_16876,N_16434,N_16043);
and U16877 (N_16877,N_16026,N_16063);
nor U16878 (N_16878,N_16597,N_16036);
nand U16879 (N_16879,N_16566,N_16154);
and U16880 (N_16880,N_16687,N_16084);
nand U16881 (N_16881,N_16269,N_16066);
nand U16882 (N_16882,N_16019,N_16765);
nor U16883 (N_16883,N_16303,N_16524);
nor U16884 (N_16884,N_16032,N_16410);
or U16885 (N_16885,N_16480,N_16356);
nor U16886 (N_16886,N_16671,N_16578);
and U16887 (N_16887,N_16612,N_16353);
nor U16888 (N_16888,N_16695,N_16300);
xor U16889 (N_16889,N_16056,N_16239);
xnor U16890 (N_16890,N_16059,N_16678);
or U16891 (N_16891,N_16726,N_16253);
xnor U16892 (N_16892,N_16555,N_16327);
xnor U16893 (N_16893,N_16144,N_16241);
nand U16894 (N_16894,N_16030,N_16734);
nand U16895 (N_16895,N_16263,N_16460);
xnor U16896 (N_16896,N_16630,N_16305);
nand U16897 (N_16897,N_16006,N_16319);
and U16898 (N_16898,N_16306,N_16686);
or U16899 (N_16899,N_16118,N_16463);
or U16900 (N_16900,N_16714,N_16389);
nor U16901 (N_16901,N_16047,N_16617);
nor U16902 (N_16902,N_16433,N_16557);
or U16903 (N_16903,N_16179,N_16704);
xor U16904 (N_16904,N_16025,N_16011);
nor U16905 (N_16905,N_16171,N_16577);
nor U16906 (N_16906,N_16284,N_16708);
nor U16907 (N_16907,N_16590,N_16768);
or U16908 (N_16908,N_16296,N_16292);
or U16909 (N_16909,N_16689,N_16159);
or U16910 (N_16910,N_16694,N_16349);
nor U16911 (N_16911,N_16231,N_16070);
xnor U16912 (N_16912,N_16545,N_16660);
xnor U16913 (N_16913,N_16388,N_16274);
xnor U16914 (N_16914,N_16243,N_16568);
nor U16915 (N_16915,N_16261,N_16271);
nor U16916 (N_16916,N_16580,N_16031);
xor U16917 (N_16917,N_16753,N_16605);
and U16918 (N_16918,N_16086,N_16050);
and U16919 (N_16919,N_16394,N_16752);
nor U16920 (N_16920,N_16579,N_16533);
and U16921 (N_16921,N_16426,N_16624);
and U16922 (N_16922,N_16444,N_16646);
or U16923 (N_16923,N_16065,N_16438);
xnor U16924 (N_16924,N_16675,N_16520);
and U16925 (N_16925,N_16772,N_16120);
nand U16926 (N_16926,N_16326,N_16038);
nand U16927 (N_16927,N_16719,N_16312);
or U16928 (N_16928,N_16277,N_16143);
nand U16929 (N_16929,N_16355,N_16425);
nor U16930 (N_16930,N_16374,N_16022);
and U16931 (N_16931,N_16775,N_16574);
nor U16932 (N_16932,N_16127,N_16273);
and U16933 (N_16933,N_16654,N_16352);
and U16934 (N_16934,N_16464,N_16373);
nand U16935 (N_16935,N_16090,N_16150);
nand U16936 (N_16936,N_16453,N_16112);
nand U16937 (N_16937,N_16029,N_16569);
nor U16938 (N_16938,N_16158,N_16104);
and U16939 (N_16939,N_16053,N_16792);
and U16940 (N_16940,N_16623,N_16783);
or U16941 (N_16941,N_16417,N_16191);
and U16942 (N_16942,N_16363,N_16637);
nand U16943 (N_16943,N_16741,N_16270);
nand U16944 (N_16944,N_16185,N_16754);
nor U16945 (N_16945,N_16042,N_16320);
nor U16946 (N_16946,N_16722,N_16076);
and U16947 (N_16947,N_16254,N_16583);
or U16948 (N_16948,N_16493,N_16651);
and U16949 (N_16949,N_16365,N_16610);
or U16950 (N_16950,N_16182,N_16221);
nor U16951 (N_16951,N_16404,N_16174);
nand U16952 (N_16952,N_16299,N_16502);
nor U16953 (N_16953,N_16706,N_16302);
nor U16954 (N_16954,N_16256,N_16717);
and U16955 (N_16955,N_16338,N_16172);
or U16956 (N_16956,N_16587,N_16534);
or U16957 (N_16957,N_16663,N_16354);
nor U16958 (N_16958,N_16074,N_16200);
nand U16959 (N_16959,N_16441,N_16121);
nand U16960 (N_16960,N_16412,N_16529);
nand U16961 (N_16961,N_16715,N_16448);
xor U16962 (N_16962,N_16681,N_16662);
nand U16963 (N_16963,N_16198,N_16473);
and U16964 (N_16964,N_16034,N_16423);
or U16965 (N_16965,N_16122,N_16461);
xnor U16966 (N_16966,N_16495,N_16236);
xnor U16967 (N_16967,N_16633,N_16496);
nand U16968 (N_16968,N_16206,N_16744);
and U16969 (N_16969,N_16209,N_16073);
and U16970 (N_16970,N_16531,N_16435);
nand U16971 (N_16971,N_16009,N_16700);
or U16972 (N_16972,N_16558,N_16401);
and U16973 (N_16973,N_16193,N_16291);
or U16974 (N_16974,N_16248,N_16547);
nand U16975 (N_16975,N_16137,N_16297);
xnor U16976 (N_16976,N_16405,N_16196);
and U16977 (N_16977,N_16328,N_16723);
xor U16978 (N_16978,N_16797,N_16400);
and U16979 (N_16979,N_16692,N_16298);
nand U16980 (N_16980,N_16259,N_16142);
or U16981 (N_16981,N_16245,N_16528);
nor U16982 (N_16982,N_16505,N_16275);
and U16983 (N_16983,N_16010,N_16201);
and U16984 (N_16984,N_16677,N_16078);
xor U16985 (N_16985,N_16535,N_16123);
xor U16986 (N_16986,N_16489,N_16411);
nor U16987 (N_16987,N_16081,N_16408);
nand U16988 (N_16988,N_16546,N_16344);
xor U16989 (N_16989,N_16332,N_16737);
nand U16990 (N_16990,N_16325,N_16443);
nor U16991 (N_16991,N_16469,N_16015);
xnor U16992 (N_16992,N_16415,N_16100);
and U16993 (N_16993,N_16422,N_16685);
xor U16994 (N_16994,N_16350,N_16523);
nand U16995 (N_16995,N_16640,N_16016);
nand U16996 (N_16996,N_16346,N_16364);
nand U16997 (N_16997,N_16614,N_16514);
xor U16998 (N_16998,N_16348,N_16515);
or U16999 (N_16999,N_16620,N_16004);
nand U17000 (N_17000,N_16764,N_16246);
nor U17001 (N_17001,N_16479,N_16283);
nor U17002 (N_17002,N_16653,N_16342);
xnor U17003 (N_17003,N_16135,N_16440);
and U17004 (N_17004,N_16632,N_16591);
nand U17005 (N_17005,N_16232,N_16329);
xor U17006 (N_17006,N_16771,N_16540);
nand U17007 (N_17007,N_16366,N_16462);
nor U17008 (N_17008,N_16490,N_16684);
nand U17009 (N_17009,N_16760,N_16385);
and U17010 (N_17010,N_16258,N_16168);
or U17011 (N_17011,N_16655,N_16207);
nor U17012 (N_17012,N_16581,N_16518);
and U17013 (N_17013,N_16014,N_16289);
and U17014 (N_17014,N_16778,N_16508);
nand U17015 (N_17015,N_16096,N_16099);
nand U17016 (N_17016,N_16645,N_16377);
xnor U17017 (N_17017,N_16683,N_16659);
nand U17018 (N_17018,N_16205,N_16260);
or U17019 (N_17019,N_16233,N_16177);
and U17020 (N_17020,N_16310,N_16219);
and U17021 (N_17021,N_16131,N_16657);
nand U17022 (N_17022,N_16690,N_16527);
xor U17023 (N_17023,N_16281,N_16228);
nand U17024 (N_17024,N_16167,N_16710);
or U17025 (N_17025,N_16647,N_16392);
xnor U17026 (N_17026,N_16054,N_16522);
nor U17027 (N_17027,N_16627,N_16267);
nor U17028 (N_17028,N_16777,N_16625);
nand U17029 (N_17029,N_16550,N_16727);
and U17030 (N_17030,N_16148,N_16324);
or U17031 (N_17031,N_16393,N_16264);
or U17032 (N_17032,N_16691,N_16552);
nor U17033 (N_17033,N_16506,N_16323);
or U17034 (N_17034,N_16576,N_16045);
nand U17035 (N_17035,N_16075,N_16739);
nor U17036 (N_17036,N_16301,N_16176);
nor U17037 (N_17037,N_16733,N_16539);
nor U17038 (N_17038,N_16509,N_16485);
or U17039 (N_17039,N_16442,N_16378);
xor U17040 (N_17040,N_16109,N_16060);
nand U17041 (N_17041,N_16477,N_16188);
or U17042 (N_17042,N_16382,N_16456);
nand U17043 (N_17043,N_16079,N_16562);
or U17044 (N_17044,N_16676,N_16280);
nand U17045 (N_17045,N_16052,N_16474);
and U17046 (N_17046,N_16656,N_16707);
nor U17047 (N_17047,N_16340,N_16668);
xnor U17048 (N_17048,N_16017,N_16115);
xnor U17049 (N_17049,N_16062,N_16369);
and U17050 (N_17050,N_16013,N_16133);
and U17051 (N_17051,N_16471,N_16565);
or U17052 (N_17052,N_16304,N_16407);
and U17053 (N_17053,N_16745,N_16139);
nand U17054 (N_17054,N_16244,N_16156);
nor U17055 (N_17055,N_16055,N_16218);
nand U17056 (N_17056,N_16234,N_16216);
or U17057 (N_17057,N_16513,N_16398);
or U17058 (N_17058,N_16204,N_16082);
nor U17059 (N_17059,N_16608,N_16169);
nor U17060 (N_17060,N_16041,N_16445);
or U17061 (N_17061,N_16307,N_16007);
xnor U17062 (N_17062,N_16210,N_16250);
nor U17063 (N_17063,N_16085,N_16318);
nand U17064 (N_17064,N_16780,N_16165);
xnor U17065 (N_17065,N_16680,N_16542);
nand U17066 (N_17066,N_16097,N_16317);
xnor U17067 (N_17067,N_16170,N_16197);
nor U17068 (N_17068,N_16709,N_16141);
xnor U17069 (N_17069,N_16278,N_16068);
nand U17070 (N_17070,N_16431,N_16359);
and U17071 (N_17071,N_16376,N_16187);
nor U17072 (N_17072,N_16088,N_16449);
or U17073 (N_17073,N_16020,N_16609);
xnor U17074 (N_17074,N_16451,N_16510);
nor U17075 (N_17075,N_16785,N_16432);
nand U17076 (N_17076,N_16282,N_16779);
nand U17077 (N_17077,N_16747,N_16358);
nand U17078 (N_17078,N_16439,N_16459);
nor U17079 (N_17079,N_16035,N_16008);
and U17080 (N_17080,N_16688,N_16229);
and U17081 (N_17081,N_16000,N_16402);
nor U17082 (N_17082,N_16257,N_16452);
and U17083 (N_17083,N_16136,N_16330);
and U17084 (N_17084,N_16199,N_16138);
xor U17085 (N_17085,N_16586,N_16638);
nand U17086 (N_17086,N_16146,N_16386);
nor U17087 (N_17087,N_16420,N_16024);
xnor U17088 (N_17088,N_16598,N_16295);
nor U17089 (N_17089,N_16560,N_16661);
and U17090 (N_17090,N_16786,N_16429);
xnor U17091 (N_17091,N_16057,N_16094);
and U17092 (N_17092,N_16331,N_16370);
xnor U17093 (N_17093,N_16486,N_16333);
or U17094 (N_17094,N_16321,N_16089);
nand U17095 (N_17095,N_16093,N_16666);
and U17096 (N_17096,N_16773,N_16582);
nand U17097 (N_17097,N_16743,N_16230);
nor U17098 (N_17098,N_16559,N_16606);
and U17099 (N_17099,N_16543,N_16643);
nand U17100 (N_17100,N_16698,N_16467);
and U17101 (N_17101,N_16602,N_16611);
or U17102 (N_17102,N_16642,N_16396);
xnor U17103 (N_17103,N_16476,N_16648);
xnor U17104 (N_17104,N_16087,N_16631);
nor U17105 (N_17105,N_16532,N_16789);
or U17106 (N_17106,N_16570,N_16424);
nor U17107 (N_17107,N_16446,N_16080);
nand U17108 (N_17108,N_16622,N_16447);
nand U17109 (N_17109,N_16652,N_16128);
nand U17110 (N_17110,N_16740,N_16336);
or U17111 (N_17111,N_16470,N_16626);
and U17112 (N_17112,N_16314,N_16674);
and U17113 (N_17113,N_16736,N_16548);
and U17114 (N_17114,N_16037,N_16040);
nand U17115 (N_17115,N_16791,N_16573);
or U17116 (N_17116,N_16746,N_16203);
or U17117 (N_17117,N_16639,N_16672);
nor U17118 (N_17118,N_16367,N_16313);
or U17119 (N_17119,N_16130,N_16287);
and U17120 (N_17120,N_16285,N_16240);
nand U17121 (N_17121,N_16718,N_16615);
nor U17122 (N_17122,N_16162,N_16224);
nor U17123 (N_17123,N_16701,N_16106);
nand U17124 (N_17124,N_16001,N_16276);
xor U17125 (N_17125,N_16091,N_16450);
and U17126 (N_17126,N_16379,N_16584);
or U17127 (N_17127,N_16413,N_16735);
and U17128 (N_17128,N_16790,N_16021);
nor U17129 (N_17129,N_16455,N_16600);
nor U17130 (N_17130,N_16003,N_16763);
and U17131 (N_17131,N_16536,N_16636);
nand U17132 (N_17132,N_16541,N_16784);
xor U17133 (N_17133,N_16613,N_16334);
nand U17134 (N_17134,N_16544,N_16799);
xnor U17135 (N_17135,N_16157,N_16488);
and U17136 (N_17136,N_16129,N_16703);
xor U17137 (N_17137,N_16217,N_16713);
or U17138 (N_17138,N_16072,N_16604);
nand U17139 (N_17139,N_16242,N_16322);
nand U17140 (N_17140,N_16788,N_16782);
nor U17141 (N_17141,N_16428,N_16738);
or U17142 (N_17142,N_16793,N_16748);
and U17143 (N_17143,N_16381,N_16235);
and U17144 (N_17144,N_16478,N_16742);
xor U17145 (N_17145,N_16436,N_16140);
xnor U17146 (N_17146,N_16145,N_16351);
or U17147 (N_17147,N_16761,N_16390);
xnor U17148 (N_17148,N_16575,N_16272);
nand U17149 (N_17149,N_16362,N_16731);
or U17150 (N_17150,N_16044,N_16184);
or U17151 (N_17151,N_16126,N_16487);
nand U17152 (N_17152,N_16494,N_16149);
nor U17153 (N_17153,N_16247,N_16262);
nor U17154 (N_17154,N_16665,N_16095);
or U17155 (N_17155,N_16249,N_16005);
or U17156 (N_17156,N_16732,N_16670);
xor U17157 (N_17157,N_16189,N_16164);
nand U17158 (N_17158,N_16058,N_16051);
or U17159 (N_17159,N_16387,N_16147);
nor U17160 (N_17160,N_16721,N_16048);
and U17161 (N_17161,N_16492,N_16290);
xor U17162 (N_17162,N_16649,N_16195);
nor U17163 (N_17163,N_16465,N_16603);
and U17164 (N_17164,N_16466,N_16728);
nor U17165 (N_17165,N_16315,N_16288);
or U17166 (N_17166,N_16214,N_16635);
and U17167 (N_17167,N_16391,N_16220);
nor U17168 (N_17168,N_16316,N_16481);
xnor U17169 (N_17169,N_16755,N_16160);
or U17170 (N_17170,N_16107,N_16716);
xnor U17171 (N_17171,N_16798,N_16380);
xnor U17172 (N_17172,N_16724,N_16117);
xor U17173 (N_17173,N_16571,N_16596);
nor U17174 (N_17174,N_16132,N_16152);
and U17175 (N_17175,N_16501,N_16725);
xnor U17176 (N_17176,N_16758,N_16049);
nor U17177 (N_17177,N_16309,N_16762);
xor U17178 (N_17178,N_16500,N_16766);
xnor U17179 (N_17179,N_16504,N_16215);
or U17180 (N_17180,N_16503,N_16225);
or U17181 (N_17181,N_16023,N_16595);
or U17182 (N_17182,N_16795,N_16061);
xnor U17183 (N_17183,N_16618,N_16712);
xor U17184 (N_17184,N_16472,N_16268);
nand U17185 (N_17185,N_16357,N_16125);
nand U17186 (N_17186,N_16551,N_16585);
xnor U17187 (N_17187,N_16705,N_16621);
xor U17188 (N_17188,N_16183,N_16693);
nor U17189 (N_17189,N_16190,N_16644);
xor U17190 (N_17190,N_16101,N_16525);
or U17191 (N_17191,N_16794,N_16151);
and U17192 (N_17192,N_16361,N_16601);
xnor U17193 (N_17193,N_16046,N_16619);
xor U17194 (N_17194,N_16155,N_16372);
nor U17195 (N_17195,N_16594,N_16028);
nand U17196 (N_17196,N_16384,N_16251);
or U17197 (N_17197,N_16033,N_16092);
xnor U17198 (N_17198,N_16437,N_16279);
or U17199 (N_17199,N_16430,N_16395);
nor U17200 (N_17200,N_16345,N_16328);
or U17201 (N_17201,N_16502,N_16501);
nand U17202 (N_17202,N_16748,N_16433);
nand U17203 (N_17203,N_16323,N_16067);
and U17204 (N_17204,N_16533,N_16496);
and U17205 (N_17205,N_16459,N_16623);
xnor U17206 (N_17206,N_16082,N_16065);
nand U17207 (N_17207,N_16309,N_16354);
xor U17208 (N_17208,N_16323,N_16213);
xnor U17209 (N_17209,N_16657,N_16394);
xor U17210 (N_17210,N_16750,N_16014);
nand U17211 (N_17211,N_16669,N_16045);
and U17212 (N_17212,N_16736,N_16475);
nand U17213 (N_17213,N_16213,N_16574);
or U17214 (N_17214,N_16653,N_16293);
nor U17215 (N_17215,N_16171,N_16634);
and U17216 (N_17216,N_16288,N_16181);
or U17217 (N_17217,N_16338,N_16421);
xor U17218 (N_17218,N_16278,N_16698);
and U17219 (N_17219,N_16483,N_16510);
xnor U17220 (N_17220,N_16275,N_16404);
nor U17221 (N_17221,N_16498,N_16694);
or U17222 (N_17222,N_16613,N_16077);
nor U17223 (N_17223,N_16489,N_16026);
or U17224 (N_17224,N_16130,N_16764);
or U17225 (N_17225,N_16423,N_16627);
or U17226 (N_17226,N_16496,N_16048);
and U17227 (N_17227,N_16369,N_16273);
or U17228 (N_17228,N_16179,N_16712);
or U17229 (N_17229,N_16568,N_16767);
and U17230 (N_17230,N_16057,N_16230);
or U17231 (N_17231,N_16512,N_16469);
xnor U17232 (N_17232,N_16128,N_16621);
nor U17233 (N_17233,N_16293,N_16670);
or U17234 (N_17234,N_16666,N_16730);
xor U17235 (N_17235,N_16371,N_16714);
nor U17236 (N_17236,N_16049,N_16757);
nor U17237 (N_17237,N_16709,N_16106);
nor U17238 (N_17238,N_16164,N_16010);
or U17239 (N_17239,N_16092,N_16689);
nor U17240 (N_17240,N_16215,N_16054);
xor U17241 (N_17241,N_16508,N_16355);
and U17242 (N_17242,N_16795,N_16789);
and U17243 (N_17243,N_16292,N_16608);
or U17244 (N_17244,N_16072,N_16051);
nor U17245 (N_17245,N_16312,N_16766);
nor U17246 (N_17246,N_16200,N_16285);
or U17247 (N_17247,N_16197,N_16112);
nand U17248 (N_17248,N_16236,N_16683);
and U17249 (N_17249,N_16646,N_16265);
xor U17250 (N_17250,N_16177,N_16686);
or U17251 (N_17251,N_16667,N_16233);
and U17252 (N_17252,N_16216,N_16096);
xor U17253 (N_17253,N_16673,N_16796);
nand U17254 (N_17254,N_16237,N_16365);
or U17255 (N_17255,N_16153,N_16767);
xnor U17256 (N_17256,N_16284,N_16751);
and U17257 (N_17257,N_16216,N_16137);
and U17258 (N_17258,N_16026,N_16735);
nand U17259 (N_17259,N_16263,N_16597);
and U17260 (N_17260,N_16371,N_16329);
xor U17261 (N_17261,N_16731,N_16070);
nand U17262 (N_17262,N_16423,N_16440);
and U17263 (N_17263,N_16277,N_16506);
xnor U17264 (N_17264,N_16450,N_16778);
or U17265 (N_17265,N_16529,N_16247);
nor U17266 (N_17266,N_16108,N_16655);
and U17267 (N_17267,N_16365,N_16594);
xor U17268 (N_17268,N_16197,N_16327);
nor U17269 (N_17269,N_16563,N_16078);
and U17270 (N_17270,N_16255,N_16004);
xor U17271 (N_17271,N_16404,N_16495);
nor U17272 (N_17272,N_16201,N_16706);
or U17273 (N_17273,N_16318,N_16425);
or U17274 (N_17274,N_16362,N_16027);
or U17275 (N_17275,N_16357,N_16204);
or U17276 (N_17276,N_16583,N_16300);
and U17277 (N_17277,N_16429,N_16034);
or U17278 (N_17278,N_16410,N_16216);
nor U17279 (N_17279,N_16361,N_16199);
xnor U17280 (N_17280,N_16353,N_16384);
nor U17281 (N_17281,N_16349,N_16625);
nand U17282 (N_17282,N_16302,N_16646);
nor U17283 (N_17283,N_16445,N_16178);
and U17284 (N_17284,N_16188,N_16410);
nor U17285 (N_17285,N_16725,N_16706);
or U17286 (N_17286,N_16311,N_16399);
nor U17287 (N_17287,N_16563,N_16759);
and U17288 (N_17288,N_16515,N_16438);
nand U17289 (N_17289,N_16631,N_16247);
or U17290 (N_17290,N_16126,N_16238);
and U17291 (N_17291,N_16086,N_16216);
nor U17292 (N_17292,N_16439,N_16295);
or U17293 (N_17293,N_16389,N_16136);
xor U17294 (N_17294,N_16501,N_16432);
and U17295 (N_17295,N_16060,N_16306);
and U17296 (N_17296,N_16711,N_16582);
or U17297 (N_17297,N_16390,N_16028);
xnor U17298 (N_17298,N_16501,N_16396);
nand U17299 (N_17299,N_16650,N_16619);
nand U17300 (N_17300,N_16413,N_16742);
nand U17301 (N_17301,N_16538,N_16755);
xnor U17302 (N_17302,N_16504,N_16358);
and U17303 (N_17303,N_16738,N_16270);
nand U17304 (N_17304,N_16629,N_16515);
or U17305 (N_17305,N_16289,N_16544);
xor U17306 (N_17306,N_16261,N_16549);
nand U17307 (N_17307,N_16766,N_16057);
nor U17308 (N_17308,N_16256,N_16177);
xor U17309 (N_17309,N_16205,N_16049);
and U17310 (N_17310,N_16694,N_16538);
xor U17311 (N_17311,N_16727,N_16291);
nand U17312 (N_17312,N_16395,N_16245);
and U17313 (N_17313,N_16696,N_16292);
xnor U17314 (N_17314,N_16182,N_16348);
nand U17315 (N_17315,N_16415,N_16154);
xor U17316 (N_17316,N_16641,N_16020);
or U17317 (N_17317,N_16625,N_16797);
xor U17318 (N_17318,N_16594,N_16132);
or U17319 (N_17319,N_16156,N_16074);
or U17320 (N_17320,N_16610,N_16294);
nor U17321 (N_17321,N_16672,N_16372);
and U17322 (N_17322,N_16505,N_16428);
or U17323 (N_17323,N_16736,N_16457);
nor U17324 (N_17324,N_16468,N_16092);
nand U17325 (N_17325,N_16025,N_16778);
nor U17326 (N_17326,N_16575,N_16264);
nand U17327 (N_17327,N_16553,N_16702);
nor U17328 (N_17328,N_16552,N_16484);
or U17329 (N_17329,N_16206,N_16115);
or U17330 (N_17330,N_16568,N_16173);
xor U17331 (N_17331,N_16646,N_16541);
xor U17332 (N_17332,N_16523,N_16341);
nor U17333 (N_17333,N_16260,N_16185);
and U17334 (N_17334,N_16105,N_16061);
or U17335 (N_17335,N_16757,N_16641);
nor U17336 (N_17336,N_16536,N_16344);
and U17337 (N_17337,N_16040,N_16524);
nand U17338 (N_17338,N_16642,N_16002);
nand U17339 (N_17339,N_16182,N_16420);
or U17340 (N_17340,N_16088,N_16131);
nand U17341 (N_17341,N_16393,N_16353);
nor U17342 (N_17342,N_16638,N_16281);
xor U17343 (N_17343,N_16293,N_16427);
or U17344 (N_17344,N_16614,N_16295);
nor U17345 (N_17345,N_16255,N_16515);
nand U17346 (N_17346,N_16191,N_16152);
or U17347 (N_17347,N_16318,N_16574);
nand U17348 (N_17348,N_16282,N_16383);
xnor U17349 (N_17349,N_16107,N_16187);
and U17350 (N_17350,N_16679,N_16047);
xor U17351 (N_17351,N_16488,N_16666);
xor U17352 (N_17352,N_16757,N_16393);
xnor U17353 (N_17353,N_16365,N_16622);
or U17354 (N_17354,N_16589,N_16284);
nor U17355 (N_17355,N_16258,N_16405);
and U17356 (N_17356,N_16111,N_16002);
and U17357 (N_17357,N_16541,N_16716);
and U17358 (N_17358,N_16078,N_16162);
nand U17359 (N_17359,N_16356,N_16545);
xor U17360 (N_17360,N_16492,N_16685);
nand U17361 (N_17361,N_16066,N_16136);
and U17362 (N_17362,N_16590,N_16550);
xor U17363 (N_17363,N_16272,N_16020);
and U17364 (N_17364,N_16013,N_16292);
nand U17365 (N_17365,N_16461,N_16538);
or U17366 (N_17366,N_16408,N_16332);
and U17367 (N_17367,N_16127,N_16510);
nand U17368 (N_17368,N_16018,N_16031);
nor U17369 (N_17369,N_16124,N_16512);
and U17370 (N_17370,N_16290,N_16657);
nor U17371 (N_17371,N_16546,N_16185);
or U17372 (N_17372,N_16312,N_16567);
xnor U17373 (N_17373,N_16582,N_16538);
nand U17374 (N_17374,N_16316,N_16725);
or U17375 (N_17375,N_16026,N_16024);
nand U17376 (N_17376,N_16637,N_16069);
and U17377 (N_17377,N_16443,N_16240);
or U17378 (N_17378,N_16734,N_16096);
or U17379 (N_17379,N_16488,N_16714);
nor U17380 (N_17380,N_16394,N_16115);
and U17381 (N_17381,N_16755,N_16018);
or U17382 (N_17382,N_16153,N_16097);
and U17383 (N_17383,N_16298,N_16739);
nor U17384 (N_17384,N_16140,N_16549);
nand U17385 (N_17385,N_16107,N_16393);
nor U17386 (N_17386,N_16770,N_16472);
nor U17387 (N_17387,N_16055,N_16275);
nand U17388 (N_17388,N_16359,N_16146);
and U17389 (N_17389,N_16356,N_16611);
xor U17390 (N_17390,N_16023,N_16781);
or U17391 (N_17391,N_16541,N_16612);
nand U17392 (N_17392,N_16780,N_16523);
nor U17393 (N_17393,N_16022,N_16621);
xnor U17394 (N_17394,N_16541,N_16768);
or U17395 (N_17395,N_16606,N_16487);
or U17396 (N_17396,N_16281,N_16368);
nor U17397 (N_17397,N_16590,N_16161);
and U17398 (N_17398,N_16612,N_16517);
xnor U17399 (N_17399,N_16141,N_16594);
xor U17400 (N_17400,N_16498,N_16677);
nand U17401 (N_17401,N_16558,N_16729);
xor U17402 (N_17402,N_16686,N_16582);
nand U17403 (N_17403,N_16503,N_16128);
nand U17404 (N_17404,N_16554,N_16266);
and U17405 (N_17405,N_16084,N_16735);
nor U17406 (N_17406,N_16281,N_16188);
and U17407 (N_17407,N_16744,N_16428);
xnor U17408 (N_17408,N_16454,N_16042);
and U17409 (N_17409,N_16599,N_16732);
and U17410 (N_17410,N_16356,N_16691);
and U17411 (N_17411,N_16583,N_16679);
and U17412 (N_17412,N_16173,N_16079);
or U17413 (N_17413,N_16258,N_16123);
xnor U17414 (N_17414,N_16523,N_16752);
or U17415 (N_17415,N_16458,N_16075);
and U17416 (N_17416,N_16557,N_16014);
nor U17417 (N_17417,N_16128,N_16394);
and U17418 (N_17418,N_16506,N_16036);
xor U17419 (N_17419,N_16431,N_16099);
or U17420 (N_17420,N_16795,N_16505);
nor U17421 (N_17421,N_16404,N_16612);
nor U17422 (N_17422,N_16459,N_16251);
nor U17423 (N_17423,N_16750,N_16371);
nand U17424 (N_17424,N_16780,N_16612);
nor U17425 (N_17425,N_16285,N_16464);
or U17426 (N_17426,N_16377,N_16333);
or U17427 (N_17427,N_16103,N_16058);
and U17428 (N_17428,N_16077,N_16196);
xnor U17429 (N_17429,N_16457,N_16474);
nand U17430 (N_17430,N_16458,N_16699);
xnor U17431 (N_17431,N_16277,N_16625);
or U17432 (N_17432,N_16637,N_16350);
or U17433 (N_17433,N_16308,N_16145);
xnor U17434 (N_17434,N_16059,N_16047);
and U17435 (N_17435,N_16057,N_16184);
nor U17436 (N_17436,N_16481,N_16115);
nor U17437 (N_17437,N_16000,N_16205);
xnor U17438 (N_17438,N_16563,N_16056);
and U17439 (N_17439,N_16087,N_16008);
xnor U17440 (N_17440,N_16345,N_16420);
and U17441 (N_17441,N_16539,N_16070);
or U17442 (N_17442,N_16633,N_16352);
nand U17443 (N_17443,N_16615,N_16329);
and U17444 (N_17444,N_16736,N_16160);
and U17445 (N_17445,N_16721,N_16492);
or U17446 (N_17446,N_16395,N_16210);
and U17447 (N_17447,N_16417,N_16304);
and U17448 (N_17448,N_16627,N_16147);
or U17449 (N_17449,N_16338,N_16013);
or U17450 (N_17450,N_16034,N_16548);
nand U17451 (N_17451,N_16050,N_16101);
xor U17452 (N_17452,N_16546,N_16069);
nand U17453 (N_17453,N_16244,N_16217);
nor U17454 (N_17454,N_16738,N_16586);
nor U17455 (N_17455,N_16200,N_16682);
and U17456 (N_17456,N_16667,N_16776);
xnor U17457 (N_17457,N_16136,N_16211);
and U17458 (N_17458,N_16055,N_16338);
xor U17459 (N_17459,N_16718,N_16728);
xor U17460 (N_17460,N_16260,N_16601);
nand U17461 (N_17461,N_16218,N_16344);
nor U17462 (N_17462,N_16203,N_16338);
or U17463 (N_17463,N_16765,N_16642);
nand U17464 (N_17464,N_16430,N_16626);
xnor U17465 (N_17465,N_16304,N_16115);
and U17466 (N_17466,N_16067,N_16496);
nand U17467 (N_17467,N_16442,N_16510);
xnor U17468 (N_17468,N_16546,N_16745);
nand U17469 (N_17469,N_16701,N_16160);
or U17470 (N_17470,N_16125,N_16534);
and U17471 (N_17471,N_16752,N_16746);
xnor U17472 (N_17472,N_16386,N_16140);
xnor U17473 (N_17473,N_16682,N_16592);
xnor U17474 (N_17474,N_16605,N_16249);
and U17475 (N_17475,N_16663,N_16201);
nand U17476 (N_17476,N_16576,N_16606);
or U17477 (N_17477,N_16629,N_16164);
nand U17478 (N_17478,N_16581,N_16521);
xor U17479 (N_17479,N_16651,N_16229);
nand U17480 (N_17480,N_16384,N_16748);
nand U17481 (N_17481,N_16615,N_16416);
and U17482 (N_17482,N_16535,N_16612);
or U17483 (N_17483,N_16779,N_16508);
or U17484 (N_17484,N_16133,N_16494);
nand U17485 (N_17485,N_16399,N_16071);
nor U17486 (N_17486,N_16575,N_16336);
xnor U17487 (N_17487,N_16281,N_16458);
and U17488 (N_17488,N_16159,N_16291);
nor U17489 (N_17489,N_16776,N_16053);
nand U17490 (N_17490,N_16244,N_16646);
nor U17491 (N_17491,N_16772,N_16664);
nand U17492 (N_17492,N_16539,N_16610);
or U17493 (N_17493,N_16585,N_16492);
or U17494 (N_17494,N_16230,N_16290);
and U17495 (N_17495,N_16534,N_16551);
nor U17496 (N_17496,N_16647,N_16071);
or U17497 (N_17497,N_16194,N_16020);
nand U17498 (N_17498,N_16498,N_16433);
nor U17499 (N_17499,N_16380,N_16576);
and U17500 (N_17500,N_16162,N_16591);
nand U17501 (N_17501,N_16261,N_16673);
nand U17502 (N_17502,N_16032,N_16378);
xor U17503 (N_17503,N_16139,N_16612);
or U17504 (N_17504,N_16150,N_16204);
and U17505 (N_17505,N_16178,N_16012);
or U17506 (N_17506,N_16369,N_16282);
nand U17507 (N_17507,N_16586,N_16309);
or U17508 (N_17508,N_16491,N_16355);
nor U17509 (N_17509,N_16102,N_16779);
or U17510 (N_17510,N_16543,N_16499);
nor U17511 (N_17511,N_16449,N_16397);
and U17512 (N_17512,N_16039,N_16370);
xnor U17513 (N_17513,N_16178,N_16711);
and U17514 (N_17514,N_16552,N_16642);
nand U17515 (N_17515,N_16222,N_16023);
nor U17516 (N_17516,N_16567,N_16146);
and U17517 (N_17517,N_16135,N_16603);
xor U17518 (N_17518,N_16732,N_16726);
xor U17519 (N_17519,N_16078,N_16597);
and U17520 (N_17520,N_16382,N_16753);
nand U17521 (N_17521,N_16432,N_16142);
xnor U17522 (N_17522,N_16120,N_16572);
nand U17523 (N_17523,N_16335,N_16107);
and U17524 (N_17524,N_16227,N_16280);
nor U17525 (N_17525,N_16621,N_16058);
nor U17526 (N_17526,N_16659,N_16610);
or U17527 (N_17527,N_16676,N_16062);
and U17528 (N_17528,N_16051,N_16729);
nor U17529 (N_17529,N_16567,N_16040);
and U17530 (N_17530,N_16035,N_16184);
nor U17531 (N_17531,N_16693,N_16636);
nor U17532 (N_17532,N_16349,N_16768);
nor U17533 (N_17533,N_16691,N_16605);
or U17534 (N_17534,N_16280,N_16142);
nand U17535 (N_17535,N_16496,N_16599);
or U17536 (N_17536,N_16184,N_16592);
and U17537 (N_17537,N_16042,N_16411);
nand U17538 (N_17538,N_16791,N_16777);
nand U17539 (N_17539,N_16482,N_16294);
xnor U17540 (N_17540,N_16209,N_16378);
nand U17541 (N_17541,N_16473,N_16632);
nor U17542 (N_17542,N_16758,N_16308);
xnor U17543 (N_17543,N_16564,N_16351);
nor U17544 (N_17544,N_16266,N_16711);
or U17545 (N_17545,N_16101,N_16410);
nand U17546 (N_17546,N_16552,N_16545);
nor U17547 (N_17547,N_16335,N_16584);
and U17548 (N_17548,N_16129,N_16389);
xor U17549 (N_17549,N_16068,N_16223);
nand U17550 (N_17550,N_16604,N_16649);
and U17551 (N_17551,N_16767,N_16240);
nand U17552 (N_17552,N_16020,N_16458);
or U17553 (N_17553,N_16073,N_16670);
xor U17554 (N_17554,N_16783,N_16531);
nand U17555 (N_17555,N_16309,N_16302);
nand U17556 (N_17556,N_16701,N_16363);
or U17557 (N_17557,N_16126,N_16520);
and U17558 (N_17558,N_16296,N_16526);
nor U17559 (N_17559,N_16731,N_16706);
xnor U17560 (N_17560,N_16014,N_16033);
xor U17561 (N_17561,N_16715,N_16175);
xor U17562 (N_17562,N_16500,N_16539);
nor U17563 (N_17563,N_16767,N_16482);
xnor U17564 (N_17564,N_16160,N_16502);
or U17565 (N_17565,N_16434,N_16407);
xnor U17566 (N_17566,N_16118,N_16714);
xor U17567 (N_17567,N_16348,N_16359);
and U17568 (N_17568,N_16177,N_16009);
or U17569 (N_17569,N_16470,N_16128);
xnor U17570 (N_17570,N_16227,N_16538);
nand U17571 (N_17571,N_16268,N_16077);
or U17572 (N_17572,N_16774,N_16664);
nand U17573 (N_17573,N_16220,N_16575);
xnor U17574 (N_17574,N_16573,N_16372);
or U17575 (N_17575,N_16559,N_16755);
xor U17576 (N_17576,N_16138,N_16327);
and U17577 (N_17577,N_16502,N_16676);
or U17578 (N_17578,N_16020,N_16490);
nor U17579 (N_17579,N_16452,N_16323);
xor U17580 (N_17580,N_16097,N_16469);
nor U17581 (N_17581,N_16014,N_16376);
nor U17582 (N_17582,N_16530,N_16234);
and U17583 (N_17583,N_16632,N_16325);
nand U17584 (N_17584,N_16134,N_16524);
xnor U17585 (N_17585,N_16376,N_16220);
or U17586 (N_17586,N_16355,N_16591);
and U17587 (N_17587,N_16192,N_16183);
and U17588 (N_17588,N_16307,N_16515);
xnor U17589 (N_17589,N_16180,N_16382);
xor U17590 (N_17590,N_16596,N_16462);
and U17591 (N_17591,N_16119,N_16411);
and U17592 (N_17592,N_16143,N_16070);
or U17593 (N_17593,N_16714,N_16565);
and U17594 (N_17594,N_16788,N_16402);
nand U17595 (N_17595,N_16284,N_16288);
nor U17596 (N_17596,N_16748,N_16415);
nor U17597 (N_17597,N_16568,N_16038);
and U17598 (N_17598,N_16199,N_16148);
xor U17599 (N_17599,N_16709,N_16731);
nand U17600 (N_17600,N_16885,N_17330);
and U17601 (N_17601,N_17242,N_17306);
and U17602 (N_17602,N_17346,N_17019);
xnor U17603 (N_17603,N_16863,N_17406);
nand U17604 (N_17604,N_17590,N_17085);
nand U17605 (N_17605,N_17294,N_17484);
nand U17606 (N_17606,N_17094,N_17175);
nand U17607 (N_17607,N_16988,N_17587);
nand U17608 (N_17608,N_17221,N_17064);
nand U17609 (N_17609,N_17383,N_17349);
nand U17610 (N_17610,N_16913,N_17488);
nor U17611 (N_17611,N_17328,N_16827);
nand U17612 (N_17612,N_16860,N_16881);
and U17613 (N_17613,N_17438,N_17030);
or U17614 (N_17614,N_17451,N_17117);
and U17615 (N_17615,N_16891,N_17354);
or U17616 (N_17616,N_16907,N_16877);
and U17617 (N_17617,N_17408,N_17059);
xor U17618 (N_17618,N_17455,N_17417);
nand U17619 (N_17619,N_17022,N_16916);
nand U17620 (N_17620,N_17017,N_17462);
and U17621 (N_17621,N_16861,N_17382);
nor U17622 (N_17622,N_17142,N_17478);
or U17623 (N_17623,N_17139,N_17191);
xnor U17624 (N_17624,N_17497,N_17146);
nor U17625 (N_17625,N_16899,N_17461);
or U17626 (N_17626,N_16992,N_17166);
nor U17627 (N_17627,N_17169,N_17419);
nand U17628 (N_17628,N_17174,N_17095);
xnor U17629 (N_17629,N_17144,N_16832);
nand U17630 (N_17630,N_17519,N_16925);
nand U17631 (N_17631,N_17183,N_16928);
nand U17632 (N_17632,N_17155,N_17375);
or U17633 (N_17633,N_16846,N_17263);
nor U17634 (N_17634,N_16973,N_17534);
or U17635 (N_17635,N_16840,N_16966);
xnor U17636 (N_17636,N_17343,N_17141);
nor U17637 (N_17637,N_16857,N_17345);
and U17638 (N_17638,N_17543,N_17333);
nor U17639 (N_17639,N_17062,N_17122);
and U17640 (N_17640,N_16829,N_17479);
xor U17641 (N_17641,N_16964,N_17197);
nor U17642 (N_17642,N_17229,N_17036);
or U17643 (N_17643,N_17381,N_17222);
xnor U17644 (N_17644,N_17070,N_17244);
nand U17645 (N_17645,N_16883,N_17318);
nand U17646 (N_17646,N_17416,N_17131);
and U17647 (N_17647,N_17362,N_17501);
or U17648 (N_17648,N_17291,N_17482);
or U17649 (N_17649,N_17151,N_17551);
and U17650 (N_17650,N_17329,N_17153);
nand U17651 (N_17651,N_17110,N_17031);
or U17652 (N_17652,N_17215,N_17317);
nand U17653 (N_17653,N_17218,N_17292);
xnor U17654 (N_17654,N_17554,N_16956);
xnor U17655 (N_17655,N_17530,N_16972);
nor U17656 (N_17656,N_16869,N_17258);
or U17657 (N_17657,N_17261,N_16971);
nand U17658 (N_17658,N_16921,N_17477);
and U17659 (N_17659,N_17537,N_17570);
or U17660 (N_17660,N_16882,N_16989);
and U17661 (N_17661,N_17264,N_16823);
and U17662 (N_17662,N_17377,N_17252);
nor U17663 (N_17663,N_17213,N_17268);
nor U17664 (N_17664,N_17054,N_16876);
xnor U17665 (N_17665,N_17160,N_17104);
xor U17666 (N_17666,N_16984,N_16957);
nand U17667 (N_17667,N_17340,N_17067);
xnor U17668 (N_17668,N_16959,N_17165);
and U17669 (N_17669,N_17023,N_17108);
nand U17670 (N_17670,N_17116,N_17386);
and U17671 (N_17671,N_17506,N_17531);
nand U17672 (N_17672,N_17392,N_17090);
and U17673 (N_17673,N_16960,N_17597);
xnor U17674 (N_17674,N_17063,N_17405);
nor U17675 (N_17675,N_17557,N_17047);
and U17676 (N_17676,N_16810,N_17336);
or U17677 (N_17677,N_16894,N_16815);
nor U17678 (N_17678,N_17508,N_16849);
and U17679 (N_17679,N_17500,N_17300);
nand U17680 (N_17680,N_17367,N_17172);
nand U17681 (N_17681,N_17331,N_17372);
and U17682 (N_17682,N_17210,N_17295);
nand U17683 (N_17683,N_16900,N_17514);
xnor U17684 (N_17684,N_17260,N_17236);
or U17685 (N_17685,N_17135,N_17020);
nor U17686 (N_17686,N_16886,N_16932);
or U17687 (N_17687,N_17401,N_16938);
or U17688 (N_17688,N_17496,N_17460);
and U17689 (N_17689,N_17250,N_17008);
nand U17690 (N_17690,N_16858,N_17180);
nand U17691 (N_17691,N_17398,N_17071);
xor U17692 (N_17692,N_16843,N_17399);
nor U17693 (N_17693,N_16830,N_17220);
or U17694 (N_17694,N_17536,N_16835);
nand U17695 (N_17695,N_16987,N_17505);
xnor U17696 (N_17696,N_17523,N_17209);
nand U17697 (N_17697,N_17545,N_17446);
xor U17698 (N_17698,N_17303,N_17353);
or U17699 (N_17699,N_17055,N_16933);
xnor U17700 (N_17700,N_17088,N_16834);
nor U17701 (N_17701,N_17302,N_17288);
nand U17702 (N_17702,N_16930,N_16852);
or U17703 (N_17703,N_16980,N_17509);
nor U17704 (N_17704,N_17569,N_17384);
and U17705 (N_17705,N_16888,N_16944);
nor U17706 (N_17706,N_16948,N_16958);
and U17707 (N_17707,N_16802,N_17048);
nand U17708 (N_17708,N_17276,N_17352);
or U17709 (N_17709,N_17112,N_17511);
nand U17710 (N_17710,N_17301,N_16870);
nand U17711 (N_17711,N_17498,N_17173);
and U17712 (N_17712,N_16914,N_17259);
xor U17713 (N_17713,N_16906,N_16873);
and U17714 (N_17714,N_17470,N_16854);
xor U17715 (N_17715,N_17513,N_17271);
nand U17716 (N_17716,N_17177,N_17573);
xor U17717 (N_17717,N_16917,N_17237);
nand U17718 (N_17718,N_17240,N_17439);
xnor U17719 (N_17719,N_17583,N_17243);
nor U17720 (N_17720,N_17521,N_17136);
and U17721 (N_17721,N_17368,N_16826);
and U17722 (N_17722,N_17212,N_17253);
nor U17723 (N_17723,N_16892,N_16879);
or U17724 (N_17724,N_17380,N_17045);
nand U17725 (N_17725,N_17158,N_17457);
or U17726 (N_17726,N_16818,N_17574);
nand U17727 (N_17727,N_17357,N_16983);
or U17728 (N_17728,N_17159,N_17546);
and U17729 (N_17729,N_17121,N_17058);
or U17730 (N_17730,N_17378,N_17200);
nor U17731 (N_17731,N_17099,N_17167);
and U17732 (N_17732,N_17075,N_17388);
and U17733 (N_17733,N_17185,N_17491);
xor U17734 (N_17734,N_17422,N_17369);
xor U17735 (N_17735,N_17517,N_17114);
nor U17736 (N_17736,N_17395,N_17480);
and U17737 (N_17737,N_17011,N_17046);
xor U17738 (N_17738,N_17415,N_17339);
nor U17739 (N_17739,N_17450,N_17168);
xnor U17740 (N_17740,N_16844,N_16874);
nand U17741 (N_17741,N_17015,N_17418);
or U17742 (N_17742,N_17434,N_17356);
and U17743 (N_17743,N_17178,N_17321);
nor U17744 (N_17744,N_16871,N_17309);
or U17745 (N_17745,N_17072,N_17098);
nand U17746 (N_17746,N_17262,N_17133);
or U17747 (N_17747,N_17425,N_17016);
xor U17748 (N_17748,N_17421,N_17000);
nand U17749 (N_17749,N_17181,N_16967);
nor U17750 (N_17750,N_17194,N_17565);
xnor U17751 (N_17751,N_17563,N_17476);
xnor U17752 (N_17752,N_16847,N_17105);
and U17753 (N_17753,N_16998,N_17586);
xnor U17754 (N_17754,N_17225,N_17006);
or U17755 (N_17755,N_17083,N_17371);
nor U17756 (N_17756,N_17324,N_16982);
xnor U17757 (N_17757,N_17246,N_16954);
nand U17758 (N_17758,N_17429,N_16813);
nand U17759 (N_17759,N_16821,N_16911);
and U17760 (N_17760,N_17113,N_17073);
nand U17761 (N_17761,N_17009,N_17293);
nand U17762 (N_17762,N_16922,N_16946);
nor U17763 (N_17763,N_16878,N_17548);
xnor U17764 (N_17764,N_17107,N_17111);
nor U17765 (N_17765,N_17475,N_17494);
or U17766 (N_17766,N_17486,N_17156);
xor U17767 (N_17767,N_16996,N_17049);
xor U17768 (N_17768,N_17270,N_17118);
nand U17769 (N_17769,N_16994,N_16985);
or U17770 (N_17770,N_16819,N_17255);
xnor U17771 (N_17771,N_17091,N_17124);
nand U17772 (N_17772,N_16997,N_17404);
or U17773 (N_17773,N_17483,N_16993);
xnor U17774 (N_17774,N_17029,N_17510);
or U17775 (N_17775,N_17305,N_17502);
xor U17776 (N_17776,N_17143,N_17005);
or U17777 (N_17777,N_17039,N_16908);
and U17778 (N_17778,N_17089,N_17192);
or U17779 (N_17779,N_17572,N_17092);
nand U17780 (N_17780,N_17130,N_17216);
xor U17781 (N_17781,N_17096,N_17231);
nand U17782 (N_17782,N_17199,N_17472);
nand U17783 (N_17783,N_16920,N_17577);
nor U17784 (N_17784,N_17120,N_17391);
or U17785 (N_17785,N_17580,N_16942);
and U17786 (N_17786,N_16848,N_17424);
and U17787 (N_17787,N_17564,N_17524);
xor U17788 (N_17788,N_17444,N_17297);
and U17789 (N_17789,N_17445,N_17355);
nor U17790 (N_17790,N_17440,N_17018);
nor U17791 (N_17791,N_17481,N_16865);
nand U17792 (N_17792,N_17069,N_16817);
nor U17793 (N_17793,N_16962,N_17525);
or U17794 (N_17794,N_17539,N_17208);
or U17795 (N_17795,N_17423,N_16902);
or U17796 (N_17796,N_17235,N_17584);
nand U17797 (N_17797,N_16923,N_16880);
nand U17798 (N_17798,N_17273,N_16918);
or U17799 (N_17799,N_16872,N_17432);
nor U17800 (N_17800,N_17533,N_16935);
or U17801 (N_17801,N_17335,N_16945);
and U17802 (N_17802,N_17256,N_17061);
xor U17803 (N_17803,N_17241,N_17076);
nand U17804 (N_17804,N_17190,N_17161);
xor U17805 (N_17805,N_17430,N_17585);
xor U17806 (N_17806,N_17021,N_17447);
nor U17807 (N_17807,N_17203,N_17561);
nand U17808 (N_17808,N_16963,N_17082);
or U17809 (N_17809,N_16934,N_16952);
xor U17810 (N_17810,N_16841,N_17041);
nor U17811 (N_17811,N_16941,N_17540);
or U17812 (N_17812,N_17038,N_17201);
or U17813 (N_17813,N_17079,N_17576);
xor U17814 (N_17814,N_17269,N_16875);
or U17815 (N_17815,N_17487,N_17275);
and U17816 (N_17816,N_17024,N_17591);
nor U17817 (N_17817,N_17176,N_17374);
or U17818 (N_17818,N_17050,N_17467);
xnor U17819 (N_17819,N_17459,N_17164);
nand U17820 (N_17820,N_17065,N_17184);
and U17821 (N_17821,N_17449,N_16955);
and U17822 (N_17822,N_16931,N_16868);
nand U17823 (N_17823,N_17552,N_16969);
xor U17824 (N_17824,N_17097,N_17214);
or U17825 (N_17825,N_16884,N_17397);
and U17826 (N_17826,N_16893,N_17219);
nand U17827 (N_17827,N_17140,N_17313);
nand U17828 (N_17828,N_17385,N_17289);
and U17829 (N_17829,N_16929,N_17535);
xnor U17830 (N_17830,N_17581,N_16897);
nand U17831 (N_17831,N_17347,N_17589);
and U17832 (N_17832,N_17248,N_16831);
xor U17833 (N_17833,N_17403,N_17550);
or U17834 (N_17834,N_17342,N_17393);
or U17835 (N_17835,N_17549,N_17427);
nand U17836 (N_17836,N_16828,N_17492);
or U17837 (N_17837,N_17341,N_17448);
xnor U17838 (N_17838,N_17034,N_16990);
or U17839 (N_17839,N_17251,N_17542);
nor U17840 (N_17840,N_17559,N_17358);
xor U17841 (N_17841,N_16867,N_16995);
and U17842 (N_17842,N_17431,N_16845);
and U17843 (N_17843,N_16905,N_17232);
or U17844 (N_17844,N_17426,N_17053);
nor U17845 (N_17845,N_17081,N_17026);
nor U17846 (N_17846,N_16968,N_17280);
nand U17847 (N_17847,N_17512,N_17101);
nand U17848 (N_17848,N_17588,N_17051);
nand U17849 (N_17849,N_17566,N_17522);
nor U17850 (N_17850,N_17170,N_16979);
or U17851 (N_17851,N_17411,N_16949);
or U17852 (N_17852,N_17102,N_17490);
xnor U17853 (N_17853,N_17507,N_17007);
and U17854 (N_17854,N_17435,N_17066);
or U17855 (N_17855,N_17226,N_16842);
nor U17856 (N_17856,N_17532,N_17413);
and U17857 (N_17857,N_16950,N_16889);
nand U17858 (N_17858,N_17334,N_17217);
and U17859 (N_17859,N_16975,N_16937);
and U17860 (N_17860,N_17189,N_17314);
xnor U17861 (N_17861,N_17553,N_17125);
and U17862 (N_17862,N_17351,N_17468);
and U17863 (N_17863,N_16974,N_16981);
nor U17864 (N_17864,N_16850,N_17282);
or U17865 (N_17865,N_16804,N_17515);
nor U17866 (N_17866,N_17086,N_17115);
and U17867 (N_17867,N_16800,N_16809);
or U17868 (N_17868,N_17323,N_17465);
xnor U17869 (N_17869,N_17312,N_16940);
nand U17870 (N_17870,N_17361,N_17503);
nor U17871 (N_17871,N_17348,N_17578);
xnor U17872 (N_17872,N_17366,N_17469);
nand U17873 (N_17873,N_17127,N_17555);
nand U17874 (N_17874,N_17037,N_17454);
and U17875 (N_17875,N_17012,N_17272);
or U17876 (N_17876,N_17148,N_17456);
xnor U17877 (N_17877,N_16825,N_17409);
nand U17878 (N_17878,N_17238,N_16910);
xor U17879 (N_17879,N_17596,N_17410);
nand U17880 (N_17880,N_17182,N_16965);
or U17881 (N_17881,N_17149,N_16812);
nor U17882 (N_17882,N_17338,N_16986);
and U17883 (N_17883,N_17206,N_17123);
and U17884 (N_17884,N_17068,N_17157);
nor U17885 (N_17885,N_17598,N_17254);
nor U17886 (N_17886,N_17211,N_16839);
or U17887 (N_17887,N_17595,N_17057);
nor U17888 (N_17888,N_16803,N_16862);
and U17889 (N_17889,N_17400,N_16898);
and U17890 (N_17890,N_17284,N_16951);
nand U17891 (N_17891,N_17171,N_17376);
nor U17892 (N_17892,N_17290,N_17287);
nor U17893 (N_17893,N_17593,N_16943);
and U17894 (N_17894,N_17520,N_17360);
or U17895 (N_17895,N_17594,N_17499);
or U17896 (N_17896,N_17308,N_17528);
xor U17897 (N_17897,N_16939,N_17359);
or U17898 (N_17898,N_16976,N_17265);
xnor U17899 (N_17899,N_17202,N_17223);
nand U17900 (N_17900,N_17373,N_17224);
xnor U17901 (N_17901,N_17186,N_16924);
or U17902 (N_17902,N_17370,N_17103);
nand U17903 (N_17903,N_16853,N_17003);
nor U17904 (N_17904,N_17060,N_17529);
or U17905 (N_17905,N_17402,N_16919);
nor U17906 (N_17906,N_17147,N_17504);
xnor U17907 (N_17907,N_16909,N_17562);
or U17908 (N_17908,N_17389,N_16901);
or U17909 (N_17909,N_17541,N_17002);
or U17910 (N_17910,N_17547,N_16822);
xnor U17911 (N_17911,N_17152,N_17257);
nor U17912 (N_17912,N_17452,N_17379);
nor U17913 (N_17913,N_17198,N_17249);
nand U17914 (N_17914,N_17433,N_17350);
nand U17915 (N_17915,N_16912,N_17516);
and U17916 (N_17916,N_17077,N_17285);
and U17917 (N_17917,N_17150,N_16824);
nand U17918 (N_17918,N_16808,N_16936);
and U17919 (N_17919,N_17365,N_17327);
or U17920 (N_17920,N_17556,N_16814);
or U17921 (N_17921,N_17138,N_16864);
and U17922 (N_17922,N_17316,N_17326);
xnor U17923 (N_17923,N_17001,N_17032);
and U17924 (N_17924,N_16859,N_17286);
or U17925 (N_17925,N_17010,N_16926);
and U17926 (N_17926,N_16927,N_17599);
nor U17927 (N_17927,N_17044,N_17568);
or U17928 (N_17928,N_17310,N_16896);
or U17929 (N_17929,N_17093,N_17106);
or U17930 (N_17930,N_17320,N_16833);
or U17931 (N_17931,N_16816,N_17567);
xnor U17932 (N_17932,N_17109,N_17441);
nand U17933 (N_17933,N_16953,N_17234);
or U17934 (N_17934,N_17560,N_17337);
nand U17935 (N_17935,N_16961,N_17195);
or U17936 (N_17936,N_17311,N_17387);
nor U17937 (N_17937,N_17128,N_17162);
and U17938 (N_17938,N_17154,N_17233);
xor U17939 (N_17939,N_17196,N_17298);
nor U17940 (N_17940,N_17414,N_17126);
nand U17941 (N_17941,N_17042,N_17319);
nand U17942 (N_17942,N_17538,N_16806);
and U17943 (N_17943,N_17230,N_16947);
and U17944 (N_17944,N_17207,N_16970);
nor U17945 (N_17945,N_17363,N_16903);
and U17946 (N_17946,N_17453,N_17582);
xnor U17947 (N_17947,N_17575,N_17493);
nor U17948 (N_17948,N_17544,N_17390);
and U17949 (N_17949,N_17412,N_16805);
or U17950 (N_17950,N_17518,N_17558);
xnor U17951 (N_17951,N_17283,N_17471);
xnor U17952 (N_17952,N_16978,N_17028);
xnor U17953 (N_17953,N_17526,N_16890);
nand U17954 (N_17954,N_17056,N_16866);
or U17955 (N_17955,N_17458,N_16895);
or U17956 (N_17956,N_17420,N_17043);
nor U17957 (N_17957,N_17187,N_17193);
or U17958 (N_17958,N_17132,N_16856);
nand U17959 (N_17959,N_16915,N_17489);
or U17960 (N_17960,N_16887,N_17078);
nand U17961 (N_17961,N_17228,N_17466);
nand U17962 (N_17962,N_17495,N_17052);
nor U17963 (N_17963,N_17307,N_17464);
and U17964 (N_17964,N_17443,N_17267);
or U17965 (N_17965,N_17239,N_17027);
and U17966 (N_17966,N_17296,N_17442);
or U17967 (N_17967,N_17100,N_17407);
nor U17968 (N_17968,N_16838,N_17485);
nand U17969 (N_17969,N_17299,N_17137);
nand U17970 (N_17970,N_16820,N_16807);
nand U17971 (N_17971,N_17315,N_17074);
or U17972 (N_17972,N_17013,N_17040);
xor U17973 (N_17973,N_17204,N_17592);
or U17974 (N_17974,N_17396,N_17322);
xnor U17975 (N_17975,N_17474,N_16801);
nor U17976 (N_17976,N_17571,N_17277);
nor U17977 (N_17977,N_16837,N_17463);
nor U17978 (N_17978,N_17527,N_17332);
or U17979 (N_17979,N_17025,N_16904);
nor U17980 (N_17980,N_17227,N_17304);
nor U17981 (N_17981,N_17119,N_17266);
xnor U17982 (N_17982,N_16999,N_17247);
nor U17983 (N_17983,N_16977,N_17163);
xor U17984 (N_17984,N_17344,N_17035);
nor U17985 (N_17985,N_16811,N_17080);
nor U17986 (N_17986,N_17245,N_17179);
nand U17987 (N_17987,N_17129,N_17437);
nand U17988 (N_17988,N_17274,N_17278);
and U17989 (N_17989,N_17084,N_17033);
and U17990 (N_17990,N_17281,N_17134);
nand U17991 (N_17991,N_16991,N_17087);
and U17992 (N_17992,N_17364,N_17004);
or U17993 (N_17993,N_17436,N_16836);
nor U17994 (N_17994,N_17394,N_17014);
and U17995 (N_17995,N_16855,N_17188);
nor U17996 (N_17996,N_17428,N_17145);
nand U17997 (N_17997,N_17279,N_17205);
or U17998 (N_17998,N_17325,N_17473);
and U17999 (N_17999,N_16851,N_17579);
nor U18000 (N_18000,N_16892,N_17098);
and U18001 (N_18001,N_17042,N_17525);
nor U18002 (N_18002,N_17326,N_17148);
and U18003 (N_18003,N_16936,N_16917);
xnor U18004 (N_18004,N_17404,N_17441);
and U18005 (N_18005,N_17344,N_17229);
nor U18006 (N_18006,N_17349,N_17551);
or U18007 (N_18007,N_16859,N_17143);
or U18008 (N_18008,N_17038,N_17168);
xnor U18009 (N_18009,N_17062,N_17035);
or U18010 (N_18010,N_17149,N_17158);
or U18011 (N_18011,N_17283,N_16864);
or U18012 (N_18012,N_17151,N_17202);
nand U18013 (N_18013,N_17589,N_17344);
or U18014 (N_18014,N_17053,N_16878);
or U18015 (N_18015,N_17038,N_17337);
or U18016 (N_18016,N_17209,N_17105);
and U18017 (N_18017,N_17482,N_16833);
xor U18018 (N_18018,N_17326,N_17115);
or U18019 (N_18019,N_17337,N_17198);
xor U18020 (N_18020,N_17505,N_16907);
and U18021 (N_18021,N_17110,N_17457);
nor U18022 (N_18022,N_17579,N_17507);
xnor U18023 (N_18023,N_17201,N_17485);
and U18024 (N_18024,N_17410,N_17575);
xor U18025 (N_18025,N_16938,N_17309);
and U18026 (N_18026,N_16886,N_16877);
or U18027 (N_18027,N_17004,N_17149);
nor U18028 (N_18028,N_17254,N_17084);
and U18029 (N_18029,N_17067,N_17475);
and U18030 (N_18030,N_17187,N_17366);
or U18031 (N_18031,N_17195,N_17498);
or U18032 (N_18032,N_17547,N_16874);
xnor U18033 (N_18033,N_17287,N_17130);
and U18034 (N_18034,N_16975,N_16827);
xnor U18035 (N_18035,N_16873,N_17308);
nor U18036 (N_18036,N_17206,N_17038);
xor U18037 (N_18037,N_16996,N_17548);
nand U18038 (N_18038,N_16901,N_16943);
xor U18039 (N_18039,N_17264,N_17545);
nor U18040 (N_18040,N_16902,N_17043);
xnor U18041 (N_18041,N_17527,N_16863);
nor U18042 (N_18042,N_17282,N_16893);
nand U18043 (N_18043,N_17343,N_17427);
or U18044 (N_18044,N_17587,N_17554);
and U18045 (N_18045,N_17521,N_17280);
nor U18046 (N_18046,N_16904,N_17460);
or U18047 (N_18047,N_17308,N_17291);
or U18048 (N_18048,N_17399,N_16875);
nor U18049 (N_18049,N_17319,N_17061);
nand U18050 (N_18050,N_17149,N_16848);
and U18051 (N_18051,N_17451,N_16918);
nor U18052 (N_18052,N_16956,N_17268);
xnor U18053 (N_18053,N_17155,N_17358);
and U18054 (N_18054,N_16943,N_17158);
nand U18055 (N_18055,N_17100,N_16994);
nor U18056 (N_18056,N_17396,N_16962);
and U18057 (N_18057,N_17265,N_17262);
xnor U18058 (N_18058,N_17011,N_16912);
xor U18059 (N_18059,N_16876,N_17243);
nor U18060 (N_18060,N_17441,N_17035);
and U18061 (N_18061,N_17099,N_17585);
and U18062 (N_18062,N_17460,N_17572);
nor U18063 (N_18063,N_16826,N_17037);
nand U18064 (N_18064,N_17150,N_17340);
and U18065 (N_18065,N_16986,N_16935);
nand U18066 (N_18066,N_17525,N_17250);
nor U18067 (N_18067,N_17468,N_17143);
xor U18068 (N_18068,N_16937,N_16819);
and U18069 (N_18069,N_16914,N_17302);
nand U18070 (N_18070,N_17050,N_17566);
nor U18071 (N_18071,N_17120,N_17088);
nand U18072 (N_18072,N_16920,N_17585);
xnor U18073 (N_18073,N_17511,N_17188);
and U18074 (N_18074,N_17549,N_17409);
xor U18075 (N_18075,N_17475,N_17124);
nand U18076 (N_18076,N_17001,N_16923);
or U18077 (N_18077,N_16833,N_16805);
nor U18078 (N_18078,N_17342,N_17190);
and U18079 (N_18079,N_17494,N_17500);
and U18080 (N_18080,N_16998,N_17523);
nor U18081 (N_18081,N_17516,N_17265);
nor U18082 (N_18082,N_17046,N_17423);
nand U18083 (N_18083,N_16998,N_16949);
and U18084 (N_18084,N_17130,N_16813);
nor U18085 (N_18085,N_17283,N_17066);
xnor U18086 (N_18086,N_16938,N_17035);
nor U18087 (N_18087,N_16934,N_17578);
xnor U18088 (N_18088,N_17589,N_17436);
or U18089 (N_18089,N_17558,N_17498);
and U18090 (N_18090,N_17200,N_17001);
xnor U18091 (N_18091,N_17272,N_17101);
xor U18092 (N_18092,N_17144,N_17411);
or U18093 (N_18093,N_17375,N_16876);
and U18094 (N_18094,N_17129,N_17508);
xor U18095 (N_18095,N_17260,N_16898);
or U18096 (N_18096,N_17569,N_17249);
nand U18097 (N_18097,N_17279,N_16948);
xnor U18098 (N_18098,N_16999,N_17437);
nand U18099 (N_18099,N_16886,N_17143);
and U18100 (N_18100,N_17047,N_16934);
nand U18101 (N_18101,N_17116,N_16898);
nor U18102 (N_18102,N_17367,N_16923);
or U18103 (N_18103,N_17240,N_16957);
or U18104 (N_18104,N_16829,N_17084);
and U18105 (N_18105,N_16992,N_17183);
xnor U18106 (N_18106,N_17170,N_17289);
and U18107 (N_18107,N_17291,N_17338);
nor U18108 (N_18108,N_17253,N_16903);
nor U18109 (N_18109,N_17272,N_17455);
nand U18110 (N_18110,N_16810,N_17573);
xnor U18111 (N_18111,N_17405,N_17365);
or U18112 (N_18112,N_17100,N_17000);
nand U18113 (N_18113,N_17162,N_17268);
and U18114 (N_18114,N_17076,N_17230);
xor U18115 (N_18115,N_17408,N_17206);
or U18116 (N_18116,N_17531,N_17580);
and U18117 (N_18117,N_17399,N_16977);
and U18118 (N_18118,N_17226,N_17576);
xor U18119 (N_18119,N_17568,N_16997);
nor U18120 (N_18120,N_17569,N_17544);
or U18121 (N_18121,N_16889,N_16971);
xor U18122 (N_18122,N_17510,N_17390);
nand U18123 (N_18123,N_16983,N_17004);
nor U18124 (N_18124,N_16809,N_17049);
nand U18125 (N_18125,N_16832,N_17425);
or U18126 (N_18126,N_17095,N_16998);
or U18127 (N_18127,N_17434,N_17189);
nand U18128 (N_18128,N_17147,N_17411);
nor U18129 (N_18129,N_17218,N_17127);
nand U18130 (N_18130,N_16918,N_17403);
or U18131 (N_18131,N_17411,N_16990);
or U18132 (N_18132,N_17262,N_17268);
and U18133 (N_18133,N_17467,N_17230);
or U18134 (N_18134,N_16891,N_17327);
nor U18135 (N_18135,N_17537,N_17543);
or U18136 (N_18136,N_17232,N_17137);
and U18137 (N_18137,N_17304,N_16883);
and U18138 (N_18138,N_17412,N_16868);
and U18139 (N_18139,N_17118,N_17572);
and U18140 (N_18140,N_17522,N_16815);
or U18141 (N_18141,N_17339,N_17373);
nand U18142 (N_18142,N_17125,N_17446);
xor U18143 (N_18143,N_16923,N_17572);
nor U18144 (N_18144,N_17260,N_16905);
nor U18145 (N_18145,N_17161,N_17512);
or U18146 (N_18146,N_16857,N_17080);
and U18147 (N_18147,N_17032,N_17332);
or U18148 (N_18148,N_17217,N_17273);
nor U18149 (N_18149,N_17559,N_16966);
nor U18150 (N_18150,N_17235,N_17534);
nand U18151 (N_18151,N_17399,N_17155);
nor U18152 (N_18152,N_16862,N_17271);
and U18153 (N_18153,N_16844,N_17038);
or U18154 (N_18154,N_17252,N_16921);
or U18155 (N_18155,N_17483,N_17035);
and U18156 (N_18156,N_17354,N_17007);
or U18157 (N_18157,N_16855,N_17590);
nor U18158 (N_18158,N_16975,N_17544);
or U18159 (N_18159,N_17353,N_17231);
xor U18160 (N_18160,N_17155,N_17261);
or U18161 (N_18161,N_17095,N_17276);
xor U18162 (N_18162,N_17198,N_16876);
and U18163 (N_18163,N_17307,N_17021);
nor U18164 (N_18164,N_17326,N_17342);
xor U18165 (N_18165,N_17142,N_17418);
nand U18166 (N_18166,N_16920,N_17292);
and U18167 (N_18167,N_17350,N_16828);
and U18168 (N_18168,N_17558,N_17430);
and U18169 (N_18169,N_17546,N_17514);
nor U18170 (N_18170,N_17019,N_16903);
or U18171 (N_18171,N_17219,N_16984);
nand U18172 (N_18172,N_17068,N_16849);
or U18173 (N_18173,N_17544,N_17124);
or U18174 (N_18174,N_17100,N_16940);
xnor U18175 (N_18175,N_17132,N_17567);
or U18176 (N_18176,N_17157,N_17257);
nor U18177 (N_18177,N_17024,N_17494);
and U18178 (N_18178,N_17223,N_17483);
and U18179 (N_18179,N_17541,N_17568);
nand U18180 (N_18180,N_17417,N_16820);
or U18181 (N_18181,N_17030,N_17024);
nor U18182 (N_18182,N_17138,N_17227);
xor U18183 (N_18183,N_16941,N_17558);
or U18184 (N_18184,N_17318,N_17365);
or U18185 (N_18185,N_17578,N_16897);
and U18186 (N_18186,N_17119,N_17593);
nand U18187 (N_18187,N_17097,N_17538);
nor U18188 (N_18188,N_17509,N_17336);
xor U18189 (N_18189,N_17392,N_17412);
nand U18190 (N_18190,N_17478,N_17277);
nor U18191 (N_18191,N_16965,N_17098);
or U18192 (N_18192,N_16919,N_16928);
nand U18193 (N_18193,N_17413,N_16951);
and U18194 (N_18194,N_17594,N_17001);
nor U18195 (N_18195,N_16884,N_16802);
xnor U18196 (N_18196,N_17465,N_17195);
nand U18197 (N_18197,N_16922,N_17374);
nor U18198 (N_18198,N_17021,N_16816);
xnor U18199 (N_18199,N_17019,N_16957);
or U18200 (N_18200,N_17076,N_17592);
nor U18201 (N_18201,N_17329,N_17577);
nand U18202 (N_18202,N_16941,N_16819);
or U18203 (N_18203,N_17553,N_17259);
or U18204 (N_18204,N_17356,N_17415);
and U18205 (N_18205,N_17599,N_17283);
nand U18206 (N_18206,N_17400,N_16862);
and U18207 (N_18207,N_17511,N_17573);
or U18208 (N_18208,N_16990,N_17047);
or U18209 (N_18209,N_17347,N_17346);
and U18210 (N_18210,N_17092,N_17509);
xnor U18211 (N_18211,N_17131,N_17434);
nor U18212 (N_18212,N_17425,N_16829);
xor U18213 (N_18213,N_17344,N_17034);
and U18214 (N_18214,N_17491,N_16878);
and U18215 (N_18215,N_16863,N_16878);
nor U18216 (N_18216,N_17591,N_17488);
and U18217 (N_18217,N_17159,N_17238);
or U18218 (N_18218,N_16981,N_17437);
and U18219 (N_18219,N_17337,N_16880);
nor U18220 (N_18220,N_17483,N_17207);
nor U18221 (N_18221,N_17282,N_16951);
or U18222 (N_18222,N_17051,N_17395);
nand U18223 (N_18223,N_17286,N_17002);
or U18224 (N_18224,N_17296,N_17255);
and U18225 (N_18225,N_16896,N_16933);
nor U18226 (N_18226,N_17209,N_17185);
xnor U18227 (N_18227,N_17019,N_17570);
and U18228 (N_18228,N_17107,N_17494);
xnor U18229 (N_18229,N_17297,N_17503);
or U18230 (N_18230,N_17594,N_17179);
xnor U18231 (N_18231,N_16922,N_17082);
and U18232 (N_18232,N_17383,N_16926);
xor U18233 (N_18233,N_17293,N_17423);
and U18234 (N_18234,N_17597,N_16950);
nor U18235 (N_18235,N_17284,N_17185);
nand U18236 (N_18236,N_17017,N_16904);
and U18237 (N_18237,N_17034,N_16833);
and U18238 (N_18238,N_17410,N_17178);
or U18239 (N_18239,N_17151,N_17494);
and U18240 (N_18240,N_17515,N_17182);
or U18241 (N_18241,N_17100,N_16885);
nor U18242 (N_18242,N_17058,N_16939);
nor U18243 (N_18243,N_17171,N_17086);
and U18244 (N_18244,N_16963,N_17090);
nor U18245 (N_18245,N_16840,N_17421);
nor U18246 (N_18246,N_16838,N_16921);
nor U18247 (N_18247,N_17377,N_17541);
xor U18248 (N_18248,N_16938,N_16978);
nor U18249 (N_18249,N_17241,N_17249);
and U18250 (N_18250,N_17155,N_17263);
and U18251 (N_18251,N_17444,N_17283);
nor U18252 (N_18252,N_16846,N_16938);
and U18253 (N_18253,N_16817,N_17130);
and U18254 (N_18254,N_17226,N_17354);
nand U18255 (N_18255,N_16830,N_17223);
and U18256 (N_18256,N_17259,N_17544);
xor U18257 (N_18257,N_17598,N_17307);
or U18258 (N_18258,N_17019,N_17591);
xnor U18259 (N_18259,N_17028,N_16807);
xor U18260 (N_18260,N_16828,N_16956);
nand U18261 (N_18261,N_16861,N_17349);
nand U18262 (N_18262,N_17397,N_16863);
nor U18263 (N_18263,N_16803,N_17031);
or U18264 (N_18264,N_17469,N_17321);
and U18265 (N_18265,N_17257,N_17141);
nand U18266 (N_18266,N_17186,N_17347);
xnor U18267 (N_18267,N_17478,N_17187);
and U18268 (N_18268,N_17020,N_17109);
and U18269 (N_18269,N_16917,N_16882);
nand U18270 (N_18270,N_17589,N_16925);
or U18271 (N_18271,N_16972,N_16818);
nand U18272 (N_18272,N_17151,N_17313);
nand U18273 (N_18273,N_16832,N_17072);
nand U18274 (N_18274,N_17153,N_16979);
and U18275 (N_18275,N_17106,N_17568);
xnor U18276 (N_18276,N_16887,N_17449);
or U18277 (N_18277,N_16924,N_17281);
xnor U18278 (N_18278,N_17071,N_17307);
or U18279 (N_18279,N_16877,N_17309);
or U18280 (N_18280,N_17047,N_17066);
nand U18281 (N_18281,N_17343,N_16863);
nand U18282 (N_18282,N_17333,N_17203);
or U18283 (N_18283,N_17455,N_17120);
nand U18284 (N_18284,N_17001,N_17380);
xor U18285 (N_18285,N_17235,N_17163);
nand U18286 (N_18286,N_17413,N_16918);
nand U18287 (N_18287,N_17080,N_17435);
nor U18288 (N_18288,N_17530,N_17523);
or U18289 (N_18289,N_17570,N_17180);
or U18290 (N_18290,N_17282,N_17005);
nand U18291 (N_18291,N_17550,N_17216);
or U18292 (N_18292,N_16864,N_17503);
nand U18293 (N_18293,N_16878,N_17222);
and U18294 (N_18294,N_17239,N_16935);
or U18295 (N_18295,N_17500,N_17575);
nand U18296 (N_18296,N_17205,N_17344);
nand U18297 (N_18297,N_16829,N_16977);
xnor U18298 (N_18298,N_17296,N_17444);
nand U18299 (N_18299,N_16860,N_16978);
nand U18300 (N_18300,N_17200,N_17053);
and U18301 (N_18301,N_17346,N_17466);
nand U18302 (N_18302,N_17394,N_17575);
nand U18303 (N_18303,N_16820,N_17488);
nor U18304 (N_18304,N_16924,N_17158);
nor U18305 (N_18305,N_17517,N_17026);
nand U18306 (N_18306,N_17043,N_17233);
xor U18307 (N_18307,N_17545,N_17224);
and U18308 (N_18308,N_17062,N_17194);
xnor U18309 (N_18309,N_17481,N_17512);
nor U18310 (N_18310,N_16975,N_17381);
and U18311 (N_18311,N_17034,N_17107);
nor U18312 (N_18312,N_17456,N_16906);
nor U18313 (N_18313,N_17479,N_17447);
nand U18314 (N_18314,N_17508,N_17229);
and U18315 (N_18315,N_17556,N_17548);
nor U18316 (N_18316,N_17243,N_16822);
xor U18317 (N_18317,N_17186,N_17559);
nor U18318 (N_18318,N_17080,N_17231);
xor U18319 (N_18319,N_17119,N_17165);
xnor U18320 (N_18320,N_16976,N_17521);
nor U18321 (N_18321,N_17348,N_17261);
and U18322 (N_18322,N_16826,N_17061);
nand U18323 (N_18323,N_16885,N_16884);
or U18324 (N_18324,N_16937,N_17099);
nor U18325 (N_18325,N_17192,N_17294);
or U18326 (N_18326,N_17212,N_16856);
and U18327 (N_18327,N_17238,N_16957);
and U18328 (N_18328,N_17198,N_17522);
xnor U18329 (N_18329,N_16950,N_17592);
xor U18330 (N_18330,N_17064,N_17039);
nor U18331 (N_18331,N_17051,N_17090);
xnor U18332 (N_18332,N_17573,N_17312);
nor U18333 (N_18333,N_17445,N_16851);
or U18334 (N_18334,N_17167,N_17034);
and U18335 (N_18335,N_17192,N_17156);
xor U18336 (N_18336,N_17176,N_17164);
nor U18337 (N_18337,N_17593,N_16980);
or U18338 (N_18338,N_17347,N_17277);
xnor U18339 (N_18339,N_17553,N_16825);
nor U18340 (N_18340,N_17467,N_17580);
and U18341 (N_18341,N_17557,N_17465);
nor U18342 (N_18342,N_17165,N_16863);
xnor U18343 (N_18343,N_17559,N_16864);
xnor U18344 (N_18344,N_17148,N_16953);
nand U18345 (N_18345,N_17104,N_17043);
nor U18346 (N_18346,N_16939,N_17442);
nor U18347 (N_18347,N_17518,N_16928);
xor U18348 (N_18348,N_17015,N_17125);
nor U18349 (N_18349,N_17356,N_17076);
and U18350 (N_18350,N_17248,N_17545);
xor U18351 (N_18351,N_17261,N_17360);
xor U18352 (N_18352,N_16881,N_17069);
and U18353 (N_18353,N_17026,N_17050);
and U18354 (N_18354,N_16920,N_17207);
or U18355 (N_18355,N_17553,N_16975);
xnor U18356 (N_18356,N_17127,N_17123);
and U18357 (N_18357,N_17481,N_16994);
nor U18358 (N_18358,N_17486,N_17244);
and U18359 (N_18359,N_17080,N_17114);
xor U18360 (N_18360,N_17539,N_17251);
and U18361 (N_18361,N_17192,N_16829);
or U18362 (N_18362,N_17383,N_17573);
nor U18363 (N_18363,N_17428,N_16869);
xnor U18364 (N_18364,N_17492,N_17525);
nand U18365 (N_18365,N_17189,N_16923);
or U18366 (N_18366,N_16818,N_17331);
nand U18367 (N_18367,N_17084,N_16990);
nor U18368 (N_18368,N_17295,N_17424);
nand U18369 (N_18369,N_17534,N_17239);
xnor U18370 (N_18370,N_17561,N_17327);
nor U18371 (N_18371,N_17123,N_17255);
and U18372 (N_18372,N_16918,N_17130);
nor U18373 (N_18373,N_17580,N_17371);
and U18374 (N_18374,N_16956,N_16906);
and U18375 (N_18375,N_17257,N_17109);
xnor U18376 (N_18376,N_17046,N_17488);
or U18377 (N_18377,N_17164,N_17448);
nand U18378 (N_18378,N_17500,N_17501);
nand U18379 (N_18379,N_17485,N_16901);
nand U18380 (N_18380,N_17177,N_17076);
and U18381 (N_18381,N_17577,N_17145);
and U18382 (N_18382,N_17469,N_17551);
nand U18383 (N_18383,N_16834,N_16930);
xnor U18384 (N_18384,N_16934,N_16829);
or U18385 (N_18385,N_16914,N_16988);
nand U18386 (N_18386,N_17475,N_17421);
nand U18387 (N_18387,N_17060,N_17146);
or U18388 (N_18388,N_17175,N_17259);
and U18389 (N_18389,N_17186,N_17304);
and U18390 (N_18390,N_16847,N_17386);
nand U18391 (N_18391,N_17504,N_17293);
nor U18392 (N_18392,N_17544,N_16972);
nor U18393 (N_18393,N_17066,N_17477);
xor U18394 (N_18394,N_17202,N_17337);
or U18395 (N_18395,N_17134,N_17189);
and U18396 (N_18396,N_17465,N_16903);
xnor U18397 (N_18397,N_17217,N_16801);
or U18398 (N_18398,N_17249,N_17335);
xor U18399 (N_18399,N_16934,N_17128);
and U18400 (N_18400,N_17808,N_18105);
xnor U18401 (N_18401,N_17795,N_17753);
xnor U18402 (N_18402,N_17740,N_17998);
nor U18403 (N_18403,N_18117,N_18092);
nand U18404 (N_18404,N_18292,N_18139);
nor U18405 (N_18405,N_17786,N_17922);
nor U18406 (N_18406,N_17966,N_18041);
and U18407 (N_18407,N_17777,N_17709);
and U18408 (N_18408,N_18118,N_18328);
or U18409 (N_18409,N_17833,N_17654);
nor U18410 (N_18410,N_17695,N_17863);
xnor U18411 (N_18411,N_17982,N_17947);
nand U18412 (N_18412,N_18355,N_18007);
xnor U18413 (N_18413,N_18182,N_17890);
and U18414 (N_18414,N_18124,N_17679);
nor U18415 (N_18415,N_18214,N_17979);
nor U18416 (N_18416,N_18131,N_18350);
or U18417 (N_18417,N_18019,N_18337);
and U18418 (N_18418,N_18033,N_17694);
or U18419 (N_18419,N_18157,N_18209);
nor U18420 (N_18420,N_18104,N_17938);
nor U18421 (N_18421,N_18070,N_17705);
nand U18422 (N_18422,N_18225,N_18314);
nand U18423 (N_18423,N_17633,N_18243);
nand U18424 (N_18424,N_17731,N_18126);
and U18425 (N_18425,N_18344,N_18060);
nand U18426 (N_18426,N_18330,N_18221);
nor U18427 (N_18427,N_18080,N_18291);
or U18428 (N_18428,N_18385,N_18322);
nand U18429 (N_18429,N_18374,N_18062);
or U18430 (N_18430,N_17734,N_17603);
nand U18431 (N_18431,N_18015,N_18269);
or U18432 (N_18432,N_18300,N_18217);
or U18433 (N_18433,N_17675,N_17946);
and U18434 (N_18434,N_17672,N_18030);
nand U18435 (N_18435,N_17907,N_17847);
nor U18436 (N_18436,N_17832,N_18232);
xor U18437 (N_18437,N_17949,N_17976);
xnor U18438 (N_18438,N_17671,N_18333);
or U18439 (N_18439,N_18055,N_17886);
or U18440 (N_18440,N_17700,N_17919);
nor U18441 (N_18441,N_18081,N_18321);
or U18442 (N_18442,N_18053,N_18318);
xnor U18443 (N_18443,N_18133,N_18307);
nor U18444 (N_18444,N_17676,N_17960);
or U18445 (N_18445,N_18230,N_18010);
nor U18446 (N_18446,N_17877,N_17750);
and U18447 (N_18447,N_18151,N_18096);
or U18448 (N_18448,N_17984,N_18359);
nor U18449 (N_18449,N_18311,N_18305);
nor U18450 (N_18450,N_18177,N_18128);
xor U18451 (N_18451,N_17882,N_18399);
nor U18452 (N_18452,N_17992,N_17666);
or U18453 (N_18453,N_18373,N_17606);
nor U18454 (N_18454,N_17751,N_17878);
and U18455 (N_18455,N_18263,N_18331);
and U18456 (N_18456,N_18150,N_17715);
nand U18457 (N_18457,N_17687,N_17796);
and U18458 (N_18458,N_18332,N_17798);
and U18459 (N_18459,N_18021,N_18073);
or U18460 (N_18460,N_17683,N_18259);
xor U18461 (N_18461,N_18265,N_18034);
or U18462 (N_18462,N_18024,N_18247);
or U18463 (N_18463,N_18368,N_18327);
or U18464 (N_18464,N_18098,N_18160);
xor U18465 (N_18465,N_17814,N_18203);
nand U18466 (N_18466,N_17885,N_17622);
nand U18467 (N_18467,N_18339,N_18186);
or U18468 (N_18468,N_18082,N_17648);
nand U18469 (N_18469,N_17988,N_18086);
or U18470 (N_18470,N_17895,N_17996);
xnor U18471 (N_18471,N_18100,N_17875);
or U18472 (N_18472,N_17754,N_18165);
and U18473 (N_18473,N_18116,N_18195);
xor U18474 (N_18474,N_18037,N_17841);
xnor U18475 (N_18475,N_17978,N_17821);
nand U18476 (N_18476,N_17692,N_17968);
nand U18477 (N_18477,N_18046,N_18155);
and U18478 (N_18478,N_18085,N_17755);
nor U18479 (N_18479,N_17839,N_17824);
nor U18480 (N_18480,N_17869,N_17723);
nor U18481 (N_18481,N_17756,N_17725);
xnor U18482 (N_18482,N_17763,N_18397);
nor U18483 (N_18483,N_18083,N_17899);
xor U18484 (N_18484,N_18145,N_17858);
and U18485 (N_18485,N_18043,N_17720);
and U18486 (N_18486,N_18285,N_18237);
and U18487 (N_18487,N_17933,N_17733);
xnor U18488 (N_18488,N_18168,N_17952);
nor U18489 (N_18489,N_18241,N_18233);
nor U18490 (N_18490,N_18121,N_17879);
xor U18491 (N_18491,N_18347,N_18384);
or U18492 (N_18492,N_18044,N_17930);
or U18493 (N_18493,N_17881,N_17953);
and U18494 (N_18494,N_18246,N_17985);
xor U18495 (N_18495,N_17950,N_17776);
nor U18496 (N_18496,N_18306,N_18271);
and U18497 (N_18497,N_18293,N_18357);
nand U18498 (N_18498,N_18058,N_18308);
nand U18499 (N_18499,N_17771,N_18180);
xnor U18500 (N_18500,N_18023,N_18147);
nand U18501 (N_18501,N_17663,N_18262);
or U18502 (N_18502,N_18141,N_17722);
and U18503 (N_18503,N_17975,N_17790);
nor U18504 (N_18504,N_18252,N_17713);
nor U18505 (N_18505,N_18094,N_17853);
and U18506 (N_18506,N_17717,N_18334);
xnor U18507 (N_18507,N_18395,N_18301);
nor U18508 (N_18508,N_18272,N_17629);
nand U18509 (N_18509,N_17956,N_17703);
or U18510 (N_18510,N_18009,N_18335);
nand U18511 (N_18511,N_17806,N_18051);
nand U18512 (N_18512,N_17941,N_18266);
nor U18513 (N_18513,N_17641,N_17920);
and U18514 (N_18514,N_18224,N_17859);
or U18515 (N_18515,N_18063,N_18178);
nor U18516 (N_18516,N_18380,N_18362);
and U18517 (N_18517,N_18173,N_17974);
or U18518 (N_18518,N_17924,N_18202);
nand U18519 (N_18519,N_17757,N_18302);
nor U18520 (N_18520,N_18371,N_17927);
nor U18521 (N_18521,N_18206,N_18066);
and U18522 (N_18522,N_18227,N_18002);
nor U18523 (N_18523,N_18277,N_18281);
nand U18524 (N_18524,N_17785,N_17864);
and U18525 (N_18525,N_17916,N_18356);
nor U18526 (N_18526,N_18336,N_17768);
or U18527 (N_18527,N_17772,N_17707);
and U18528 (N_18528,N_18363,N_17904);
xnor U18529 (N_18529,N_17873,N_17741);
xnor U18530 (N_18530,N_18201,N_17967);
xnor U18531 (N_18531,N_17604,N_18025);
or U18532 (N_18532,N_18235,N_17787);
or U18533 (N_18533,N_18240,N_18372);
nand U18534 (N_18534,N_18383,N_17970);
and U18535 (N_18535,N_18011,N_17690);
xnor U18536 (N_18536,N_18215,N_18289);
nor U18537 (N_18537,N_17926,N_18138);
nor U18538 (N_18538,N_18008,N_17632);
and U18539 (N_18539,N_17862,N_17719);
xnor U18540 (N_18540,N_18342,N_17818);
and U18541 (N_18541,N_18387,N_18148);
nand U18542 (N_18542,N_17830,N_18052);
and U18543 (N_18543,N_17804,N_17827);
nand U18544 (N_18544,N_17834,N_18273);
nand U18545 (N_18545,N_18244,N_17943);
nor U18546 (N_18546,N_18276,N_17749);
nand U18547 (N_18547,N_17857,N_17860);
or U18548 (N_18548,N_18067,N_18068);
nand U18549 (N_18549,N_18048,N_17912);
or U18550 (N_18550,N_17630,N_17793);
xor U18551 (N_18551,N_17842,N_17764);
or U18552 (N_18552,N_17961,N_17716);
and U18553 (N_18553,N_17684,N_17893);
xnor U18554 (N_18554,N_18249,N_17743);
nand U18555 (N_18555,N_17959,N_17752);
and U18556 (N_18556,N_18078,N_18018);
or U18557 (N_18557,N_18323,N_18340);
or U18558 (N_18558,N_18346,N_18135);
xor U18559 (N_18559,N_17929,N_18170);
nor U18560 (N_18560,N_18375,N_18156);
nand U18561 (N_18561,N_18250,N_18358);
or U18562 (N_18562,N_18123,N_18379);
or U18563 (N_18563,N_18114,N_17908);
nor U18564 (N_18564,N_18125,N_17736);
xor U18565 (N_18565,N_18386,N_17655);
or U18566 (N_18566,N_17681,N_18392);
nor U18567 (N_18567,N_18120,N_17625);
nand U18568 (N_18568,N_17657,N_17738);
xnor U18569 (N_18569,N_18196,N_17989);
or U18570 (N_18570,N_18090,N_18057);
and U18571 (N_18571,N_18187,N_17923);
nand U18572 (N_18572,N_17925,N_18315);
nor U18573 (N_18573,N_18158,N_18261);
xnor U18574 (N_18574,N_17600,N_17619);
nor U18575 (N_18575,N_17650,N_17658);
xnor U18576 (N_18576,N_18102,N_17610);
xor U18577 (N_18577,N_18376,N_17963);
xnor U18578 (N_18578,N_18309,N_17708);
nor U18579 (N_18579,N_17789,N_17816);
and U18580 (N_18580,N_18260,N_17706);
or U18581 (N_18581,N_18297,N_18212);
nand U18582 (N_18582,N_17746,N_17739);
xnor U18583 (N_18583,N_18199,N_17880);
nand U18584 (N_18584,N_18097,N_17987);
or U18585 (N_18585,N_18324,N_18320);
nand U18586 (N_18586,N_17732,N_18231);
or U18587 (N_18587,N_17727,N_17653);
xnor U18588 (N_18588,N_17794,N_18061);
nand U18589 (N_18589,N_18312,N_18394);
nor U18590 (N_18590,N_17640,N_17673);
or U18591 (N_18591,N_17822,N_18299);
nand U18592 (N_18592,N_17621,N_18258);
nor U18593 (N_18593,N_17730,N_17712);
nand U18594 (N_18594,N_17767,N_17981);
nand U18595 (N_18595,N_18349,N_18108);
nand U18596 (N_18596,N_17791,N_17797);
or U18597 (N_18597,N_17783,N_18369);
or U18598 (N_18598,N_17686,N_18219);
xnor U18599 (N_18599,N_18248,N_18056);
nand U18600 (N_18600,N_18255,N_17866);
or U18601 (N_18601,N_17674,N_17773);
or U18602 (N_18602,N_17747,N_18091);
or U18603 (N_18603,N_18036,N_17761);
nand U18604 (N_18604,N_17784,N_18282);
and U18605 (N_18605,N_17903,N_18031);
or U18606 (N_18606,N_17759,N_18205);
and U18607 (N_18607,N_18175,N_18191);
xnor U18608 (N_18608,N_17710,N_18207);
nand U18609 (N_18609,N_17615,N_18366);
or U18610 (N_18610,N_17628,N_18185);
nand U18611 (N_18611,N_18242,N_18190);
xnor U18612 (N_18612,N_17744,N_17646);
or U18613 (N_18613,N_18174,N_18211);
or U18614 (N_18614,N_17910,N_18088);
nor U18615 (N_18615,N_17909,N_18099);
or U18616 (N_18616,N_17608,N_18218);
or U18617 (N_18617,N_18198,N_18251);
xnor U18618 (N_18618,N_17677,N_17845);
nand U18619 (N_18619,N_18172,N_17931);
xor U18620 (N_18620,N_18163,N_18213);
and U18621 (N_18621,N_17894,N_18181);
nand U18622 (N_18622,N_17721,N_18129);
nand U18623 (N_18623,N_18176,N_18154);
or U18624 (N_18624,N_18003,N_17788);
xor U18625 (N_18625,N_18310,N_18093);
or U18626 (N_18626,N_18278,N_17851);
nor U18627 (N_18627,N_18210,N_18069);
or U18628 (N_18628,N_17993,N_18075);
nand U18629 (N_18629,N_17680,N_17983);
and U18630 (N_18630,N_17843,N_17940);
or U18631 (N_18631,N_17889,N_18345);
and U18632 (N_18632,N_17637,N_17918);
nor U18633 (N_18633,N_17765,N_17607);
nor U18634 (N_18634,N_18353,N_18040);
xnor U18635 (N_18635,N_18390,N_17627);
and U18636 (N_18636,N_17670,N_18159);
nor U18637 (N_18637,N_17826,N_18200);
or U18638 (N_18638,N_17972,N_17884);
xnor U18639 (N_18639,N_17699,N_17928);
and U18640 (N_18640,N_18194,N_17942);
and U18641 (N_18641,N_18140,N_17965);
nor U18642 (N_18642,N_18381,N_18054);
nor U18643 (N_18643,N_18064,N_17829);
nand U18644 (N_18644,N_17626,N_17802);
nor U18645 (N_18645,N_17865,N_18326);
and U18646 (N_18646,N_17601,N_18050);
and U18647 (N_18647,N_17986,N_18377);
or U18648 (N_18648,N_17867,N_17999);
nor U18649 (N_18649,N_18351,N_18136);
or U18650 (N_18650,N_18005,N_17769);
or U18651 (N_18651,N_17726,N_17871);
xor U18652 (N_18652,N_17825,N_18006);
or U18653 (N_18653,N_17915,N_18283);
xor U18654 (N_18654,N_17977,N_17911);
nand U18655 (N_18655,N_18027,N_17799);
or U18656 (N_18656,N_18071,N_17635);
nor U18657 (N_18657,N_18317,N_17696);
xnor U18658 (N_18658,N_17724,N_17902);
nor U18659 (N_18659,N_18072,N_18014);
nor U18660 (N_18660,N_17770,N_18396);
nand U18661 (N_18661,N_18076,N_17897);
nand U18662 (N_18662,N_18226,N_18119);
or U18663 (N_18663,N_18267,N_18000);
nand U18664 (N_18664,N_18341,N_18229);
nand U18665 (N_18665,N_18013,N_18268);
xor U18666 (N_18666,N_17945,N_17921);
or U18667 (N_18667,N_17614,N_18313);
nand U18668 (N_18668,N_17874,N_17813);
xnor U18669 (N_18669,N_18280,N_17661);
nand U18670 (N_18670,N_18049,N_18389);
or U18671 (N_18671,N_17701,N_18004);
nand U18672 (N_18672,N_18074,N_18039);
xor U18673 (N_18673,N_17643,N_17819);
or U18674 (N_18674,N_18253,N_18109);
and U18675 (N_18675,N_17639,N_17861);
nor U18676 (N_18676,N_18228,N_18348);
xor U18677 (N_18677,N_18329,N_17617);
nand U18678 (N_18678,N_18047,N_17623);
xor U18679 (N_18679,N_17991,N_17647);
xor U18680 (N_18680,N_17831,N_18288);
and U18681 (N_18681,N_18038,N_17737);
nor U18682 (N_18682,N_17691,N_17735);
nor U18683 (N_18683,N_17669,N_17914);
nand U18684 (N_18684,N_17951,N_17651);
xnor U18685 (N_18685,N_18290,N_18112);
nand U18686 (N_18686,N_18294,N_18343);
nor U18687 (N_18687,N_18254,N_18236);
and U18688 (N_18688,N_17702,N_17964);
xnor U18689 (N_18689,N_17652,N_18103);
xnor U18690 (N_18690,N_18084,N_18179);
nand U18691 (N_18691,N_17955,N_18026);
nand U18692 (N_18692,N_17896,N_18220);
nor U18693 (N_18693,N_18137,N_18127);
and U18694 (N_18694,N_18378,N_17917);
or U18695 (N_18695,N_17848,N_18298);
xor U18696 (N_18696,N_18001,N_18012);
nand U18697 (N_18697,N_17846,N_17932);
or U18698 (N_18698,N_17689,N_18020);
nand U18699 (N_18699,N_17642,N_17728);
and U18700 (N_18700,N_17828,N_17711);
nand U18701 (N_18701,N_18059,N_18153);
xor U18702 (N_18702,N_18089,N_17613);
or U18703 (N_18703,N_18166,N_17748);
and U18704 (N_18704,N_17855,N_18367);
nand U18705 (N_18705,N_17913,N_17990);
nor U18706 (N_18706,N_18130,N_17778);
and U18707 (N_18707,N_18319,N_17849);
nor U18708 (N_18708,N_18087,N_18245);
nand U18709 (N_18709,N_17616,N_17854);
or U18710 (N_18710,N_17948,N_18208);
nand U18711 (N_18711,N_18398,N_17668);
nand U18712 (N_18712,N_18101,N_18042);
xor U18713 (N_18713,N_17662,N_18164);
and U18714 (N_18714,N_18193,N_18107);
and U18715 (N_18715,N_17876,N_18095);
nand U18716 (N_18716,N_17971,N_17638);
xnor U18717 (N_18717,N_17774,N_18274);
nor U18718 (N_18718,N_18115,N_17611);
nor U18719 (N_18719,N_18077,N_18393);
or U18720 (N_18720,N_18325,N_17800);
nor U18721 (N_18721,N_17815,N_17823);
nor U18722 (N_18722,N_18370,N_17969);
and U18723 (N_18723,N_18388,N_17870);
nor U18724 (N_18724,N_17939,N_17644);
or U18725 (N_18725,N_17704,N_17934);
nor U18726 (N_18726,N_17835,N_17888);
nor U18727 (N_18727,N_17836,N_18189);
nand U18728 (N_18728,N_18113,N_18295);
xor U18729 (N_18729,N_18279,N_17944);
or U18730 (N_18730,N_18184,N_18162);
and U18731 (N_18731,N_18361,N_17820);
xnor U18732 (N_18732,N_18152,N_18316);
and U18733 (N_18733,N_18360,N_18270);
nor U18734 (N_18734,N_18161,N_18264);
xor U18735 (N_18735,N_17883,N_18146);
or U18736 (N_18736,N_17631,N_18017);
xnor U18737 (N_18737,N_17636,N_18029);
or U18738 (N_18738,N_18022,N_17781);
and U18739 (N_18739,N_18352,N_17685);
and U18740 (N_18740,N_18338,N_17612);
or U18741 (N_18741,N_17805,N_18382);
and U18742 (N_18742,N_17775,N_17892);
xor U18743 (N_18743,N_18142,N_18284);
nand U18744 (N_18744,N_18275,N_18188);
nand U18745 (N_18745,N_17745,N_17665);
nor U18746 (N_18746,N_17837,N_17742);
and U18747 (N_18747,N_18296,N_17840);
nor U18748 (N_18748,N_17780,N_17973);
nand U18749 (N_18749,N_18391,N_18222);
xnor U18750 (N_18750,N_17792,N_17936);
nand U18751 (N_18751,N_18364,N_17954);
or U18752 (N_18752,N_18183,N_17906);
xnor U18753 (N_18753,N_17980,N_18143);
and U18754 (N_18754,N_18171,N_18286);
and U18755 (N_18755,N_17624,N_17620);
xnor U18756 (N_18756,N_17868,N_17810);
nand U18757 (N_18757,N_18365,N_18106);
or U18758 (N_18758,N_17664,N_17803);
xnor U18759 (N_18759,N_18223,N_17602);
nand U18760 (N_18760,N_18167,N_17838);
nor U18761 (N_18761,N_17898,N_18035);
nor U18762 (N_18762,N_17900,N_17994);
and U18763 (N_18763,N_17688,N_17779);
and U18764 (N_18764,N_17807,N_17667);
nor U18765 (N_18765,N_18045,N_17660);
or U18766 (N_18766,N_17649,N_18016);
or U18767 (N_18767,N_17714,N_17887);
nand U18768 (N_18768,N_18079,N_17645);
nor U18769 (N_18769,N_17957,N_17891);
nand U18770 (N_18770,N_17656,N_17697);
nand U18771 (N_18771,N_18287,N_17872);
nand U18772 (N_18772,N_17812,N_18028);
or U18773 (N_18773,N_17809,N_18134);
xor U18774 (N_18774,N_17817,N_18197);
xor U18775 (N_18775,N_18144,N_18257);
or U18776 (N_18776,N_18032,N_18132);
nor U18777 (N_18777,N_17760,N_17850);
xor U18778 (N_18778,N_18216,N_18169);
nor U18779 (N_18779,N_17693,N_18239);
or U18780 (N_18780,N_17678,N_17634);
and U18781 (N_18781,N_17618,N_17609);
nand U18782 (N_18782,N_18303,N_18149);
xor U18783 (N_18783,N_18122,N_17801);
nor U18784 (N_18784,N_17852,N_17698);
or U18785 (N_18785,N_18234,N_18065);
nand U18786 (N_18786,N_17901,N_17905);
xor U18787 (N_18787,N_17997,N_17995);
nand U18788 (N_18788,N_17758,N_17762);
and U18789 (N_18789,N_17935,N_18238);
nor U18790 (N_18790,N_17605,N_17729);
and U18791 (N_18791,N_18204,N_17856);
or U18792 (N_18792,N_17782,N_18354);
nand U18793 (N_18793,N_17937,N_17682);
nor U18794 (N_18794,N_18110,N_18192);
nor U18795 (N_18795,N_18304,N_17811);
nand U18796 (N_18796,N_17718,N_17958);
nor U18797 (N_18797,N_17659,N_17962);
or U18798 (N_18798,N_18256,N_17844);
or U18799 (N_18799,N_17766,N_18111);
nor U18800 (N_18800,N_18036,N_17831);
or U18801 (N_18801,N_17921,N_17769);
or U18802 (N_18802,N_18238,N_17898);
xnor U18803 (N_18803,N_18196,N_17968);
or U18804 (N_18804,N_18354,N_18048);
nor U18805 (N_18805,N_18361,N_18327);
nor U18806 (N_18806,N_18136,N_17919);
and U18807 (N_18807,N_18375,N_17648);
or U18808 (N_18808,N_18376,N_17934);
xor U18809 (N_18809,N_17761,N_18332);
nor U18810 (N_18810,N_17960,N_17897);
nand U18811 (N_18811,N_18303,N_17759);
or U18812 (N_18812,N_17719,N_18049);
xor U18813 (N_18813,N_18288,N_17828);
or U18814 (N_18814,N_17944,N_18255);
xnor U18815 (N_18815,N_18262,N_17900);
or U18816 (N_18816,N_18263,N_18201);
and U18817 (N_18817,N_18155,N_17879);
and U18818 (N_18818,N_18305,N_18239);
xnor U18819 (N_18819,N_17766,N_17641);
xnor U18820 (N_18820,N_17949,N_17889);
nor U18821 (N_18821,N_17985,N_18153);
and U18822 (N_18822,N_18308,N_17991);
nor U18823 (N_18823,N_17890,N_17759);
nand U18824 (N_18824,N_17997,N_18294);
or U18825 (N_18825,N_17732,N_17969);
xnor U18826 (N_18826,N_18068,N_17769);
xnor U18827 (N_18827,N_17674,N_17749);
nor U18828 (N_18828,N_17881,N_17862);
xor U18829 (N_18829,N_17667,N_17944);
and U18830 (N_18830,N_17675,N_17900);
xor U18831 (N_18831,N_17732,N_17795);
xor U18832 (N_18832,N_18081,N_18092);
xnor U18833 (N_18833,N_17936,N_17628);
nor U18834 (N_18834,N_17742,N_18088);
nand U18835 (N_18835,N_18116,N_18055);
nor U18836 (N_18836,N_18391,N_18293);
and U18837 (N_18837,N_17933,N_18149);
xor U18838 (N_18838,N_17957,N_17956);
and U18839 (N_18839,N_17668,N_17931);
nand U18840 (N_18840,N_17749,N_17954);
nor U18841 (N_18841,N_18020,N_18209);
or U18842 (N_18842,N_17936,N_18033);
and U18843 (N_18843,N_18293,N_18222);
or U18844 (N_18844,N_17602,N_17984);
xor U18845 (N_18845,N_17663,N_17769);
nor U18846 (N_18846,N_18290,N_18380);
xnor U18847 (N_18847,N_18395,N_17729);
or U18848 (N_18848,N_18192,N_18020);
xor U18849 (N_18849,N_17695,N_18270);
or U18850 (N_18850,N_18254,N_18368);
nand U18851 (N_18851,N_18113,N_17826);
and U18852 (N_18852,N_18194,N_17816);
xnor U18853 (N_18853,N_17858,N_17735);
nor U18854 (N_18854,N_17633,N_18068);
or U18855 (N_18855,N_18017,N_18012);
and U18856 (N_18856,N_17640,N_17895);
and U18857 (N_18857,N_18379,N_17880);
nor U18858 (N_18858,N_18088,N_17836);
or U18859 (N_18859,N_17842,N_18017);
nand U18860 (N_18860,N_17840,N_18280);
and U18861 (N_18861,N_18032,N_18020);
or U18862 (N_18862,N_17898,N_17962);
and U18863 (N_18863,N_18176,N_18201);
or U18864 (N_18864,N_18249,N_18190);
and U18865 (N_18865,N_18391,N_18171);
and U18866 (N_18866,N_17679,N_18206);
xnor U18867 (N_18867,N_18299,N_18100);
or U18868 (N_18868,N_17692,N_18081);
or U18869 (N_18869,N_18157,N_17629);
nand U18870 (N_18870,N_17926,N_17676);
nor U18871 (N_18871,N_17743,N_17933);
or U18872 (N_18872,N_17806,N_17912);
nor U18873 (N_18873,N_18369,N_17886);
nor U18874 (N_18874,N_17683,N_18037);
nor U18875 (N_18875,N_17979,N_17755);
nor U18876 (N_18876,N_18101,N_18071);
nand U18877 (N_18877,N_18042,N_18367);
xnor U18878 (N_18878,N_18397,N_17646);
nor U18879 (N_18879,N_18026,N_17665);
and U18880 (N_18880,N_17877,N_18306);
or U18881 (N_18881,N_18235,N_17847);
xor U18882 (N_18882,N_18135,N_17986);
and U18883 (N_18883,N_18229,N_18235);
nand U18884 (N_18884,N_18156,N_18225);
and U18885 (N_18885,N_17652,N_17789);
xor U18886 (N_18886,N_17877,N_17831);
and U18887 (N_18887,N_18055,N_17975);
xor U18888 (N_18888,N_17984,N_18042);
and U18889 (N_18889,N_17855,N_18041);
nor U18890 (N_18890,N_18374,N_18316);
xor U18891 (N_18891,N_17943,N_18286);
and U18892 (N_18892,N_17811,N_18224);
xnor U18893 (N_18893,N_18399,N_17698);
nor U18894 (N_18894,N_17722,N_17735);
nor U18895 (N_18895,N_18102,N_18307);
nor U18896 (N_18896,N_17697,N_17847);
xnor U18897 (N_18897,N_18156,N_17725);
nand U18898 (N_18898,N_18167,N_17722);
nand U18899 (N_18899,N_18345,N_17609);
or U18900 (N_18900,N_18200,N_17651);
nand U18901 (N_18901,N_17704,N_18308);
or U18902 (N_18902,N_18104,N_18194);
nand U18903 (N_18903,N_17814,N_18229);
xor U18904 (N_18904,N_17680,N_17842);
or U18905 (N_18905,N_18265,N_18015);
and U18906 (N_18906,N_18200,N_18158);
xor U18907 (N_18907,N_18135,N_18342);
nand U18908 (N_18908,N_18024,N_18260);
xor U18909 (N_18909,N_17609,N_18157);
xnor U18910 (N_18910,N_17858,N_17602);
nand U18911 (N_18911,N_18140,N_17909);
and U18912 (N_18912,N_17985,N_18364);
or U18913 (N_18913,N_17677,N_18398);
and U18914 (N_18914,N_17741,N_17882);
nor U18915 (N_18915,N_18283,N_18314);
nand U18916 (N_18916,N_18243,N_18297);
and U18917 (N_18917,N_18186,N_18085);
xor U18918 (N_18918,N_18182,N_18245);
and U18919 (N_18919,N_17629,N_18134);
nand U18920 (N_18920,N_18182,N_17750);
xor U18921 (N_18921,N_17801,N_17652);
nand U18922 (N_18922,N_18019,N_17948);
xor U18923 (N_18923,N_17800,N_18010);
xor U18924 (N_18924,N_18195,N_17863);
xnor U18925 (N_18925,N_17893,N_18232);
nor U18926 (N_18926,N_18120,N_18197);
and U18927 (N_18927,N_18137,N_17845);
and U18928 (N_18928,N_18254,N_18318);
xnor U18929 (N_18929,N_18228,N_17621);
and U18930 (N_18930,N_17726,N_17900);
and U18931 (N_18931,N_18387,N_17878);
nor U18932 (N_18932,N_18118,N_18110);
nand U18933 (N_18933,N_17987,N_18292);
or U18934 (N_18934,N_17670,N_18202);
and U18935 (N_18935,N_18395,N_18122);
or U18936 (N_18936,N_17995,N_17639);
or U18937 (N_18937,N_17606,N_18108);
nand U18938 (N_18938,N_18255,N_18241);
and U18939 (N_18939,N_17751,N_18194);
and U18940 (N_18940,N_17950,N_18329);
nor U18941 (N_18941,N_17797,N_17981);
and U18942 (N_18942,N_18041,N_18343);
and U18943 (N_18943,N_17872,N_17705);
nand U18944 (N_18944,N_17981,N_18310);
and U18945 (N_18945,N_18002,N_18365);
nor U18946 (N_18946,N_17716,N_17980);
nand U18947 (N_18947,N_17667,N_18040);
nor U18948 (N_18948,N_17827,N_18003);
nand U18949 (N_18949,N_17620,N_17622);
nor U18950 (N_18950,N_17855,N_18277);
nor U18951 (N_18951,N_18264,N_18164);
xnor U18952 (N_18952,N_17860,N_18211);
or U18953 (N_18953,N_17735,N_17717);
nor U18954 (N_18954,N_17862,N_17910);
xor U18955 (N_18955,N_17675,N_18140);
xnor U18956 (N_18956,N_18067,N_17816);
nor U18957 (N_18957,N_17876,N_17790);
nand U18958 (N_18958,N_17838,N_17822);
nor U18959 (N_18959,N_18359,N_18077);
nor U18960 (N_18960,N_17783,N_17777);
or U18961 (N_18961,N_18382,N_18226);
or U18962 (N_18962,N_17650,N_17963);
nand U18963 (N_18963,N_18101,N_18009);
and U18964 (N_18964,N_18149,N_17979);
xnor U18965 (N_18965,N_18290,N_17765);
nor U18966 (N_18966,N_17639,N_18314);
nand U18967 (N_18967,N_18081,N_18198);
nor U18968 (N_18968,N_18345,N_18033);
or U18969 (N_18969,N_18001,N_18380);
and U18970 (N_18970,N_17770,N_18297);
and U18971 (N_18971,N_18121,N_17844);
xnor U18972 (N_18972,N_18155,N_17760);
nand U18973 (N_18973,N_18024,N_18012);
nand U18974 (N_18974,N_17835,N_17931);
nor U18975 (N_18975,N_18324,N_18365);
nand U18976 (N_18976,N_17662,N_17671);
and U18977 (N_18977,N_18362,N_18299);
or U18978 (N_18978,N_17842,N_18167);
or U18979 (N_18979,N_17883,N_17810);
xnor U18980 (N_18980,N_18138,N_18103);
and U18981 (N_18981,N_17973,N_17814);
and U18982 (N_18982,N_18333,N_17660);
or U18983 (N_18983,N_18076,N_18198);
xor U18984 (N_18984,N_17744,N_17610);
and U18985 (N_18985,N_17624,N_17684);
nand U18986 (N_18986,N_18303,N_17840);
or U18987 (N_18987,N_18281,N_18283);
and U18988 (N_18988,N_18067,N_17963);
and U18989 (N_18989,N_17811,N_17937);
nand U18990 (N_18990,N_18249,N_17631);
nor U18991 (N_18991,N_17622,N_18064);
nand U18992 (N_18992,N_18010,N_17873);
nor U18993 (N_18993,N_17894,N_17618);
and U18994 (N_18994,N_17651,N_17771);
nand U18995 (N_18995,N_17761,N_17850);
xor U18996 (N_18996,N_18071,N_18098);
nand U18997 (N_18997,N_18338,N_18071);
xor U18998 (N_18998,N_18038,N_18071);
or U18999 (N_18999,N_17731,N_17848);
nand U19000 (N_19000,N_17832,N_17973);
xor U19001 (N_19001,N_18032,N_17948);
xnor U19002 (N_19002,N_18063,N_17949);
or U19003 (N_19003,N_17663,N_18372);
nor U19004 (N_19004,N_17669,N_18347);
nor U19005 (N_19005,N_18182,N_18108);
nor U19006 (N_19006,N_17847,N_18282);
xnor U19007 (N_19007,N_17815,N_18285);
or U19008 (N_19008,N_18375,N_17868);
nor U19009 (N_19009,N_18221,N_17700);
or U19010 (N_19010,N_17728,N_17914);
nor U19011 (N_19011,N_18054,N_17904);
nand U19012 (N_19012,N_17724,N_17685);
and U19013 (N_19013,N_18224,N_17612);
nand U19014 (N_19014,N_17879,N_18367);
nor U19015 (N_19015,N_17668,N_17674);
or U19016 (N_19016,N_17787,N_17802);
xor U19017 (N_19017,N_18024,N_18064);
and U19018 (N_19018,N_17780,N_17647);
and U19019 (N_19019,N_17896,N_18085);
and U19020 (N_19020,N_18054,N_18035);
nand U19021 (N_19021,N_17650,N_17961);
nor U19022 (N_19022,N_17847,N_18269);
and U19023 (N_19023,N_18141,N_17805);
and U19024 (N_19024,N_18018,N_17735);
nand U19025 (N_19025,N_18001,N_18387);
or U19026 (N_19026,N_18204,N_18036);
or U19027 (N_19027,N_17784,N_17842);
or U19028 (N_19028,N_18056,N_18297);
and U19029 (N_19029,N_17876,N_17696);
or U19030 (N_19030,N_18191,N_17869);
or U19031 (N_19031,N_17907,N_17638);
nor U19032 (N_19032,N_18048,N_18149);
nor U19033 (N_19033,N_18032,N_17850);
nor U19034 (N_19034,N_18180,N_18181);
nor U19035 (N_19035,N_17749,N_18086);
and U19036 (N_19036,N_17934,N_17989);
or U19037 (N_19037,N_17752,N_18247);
xnor U19038 (N_19038,N_17967,N_17976);
nor U19039 (N_19039,N_17995,N_18301);
nand U19040 (N_19040,N_17874,N_17678);
and U19041 (N_19041,N_18397,N_17898);
nand U19042 (N_19042,N_18392,N_18000);
nor U19043 (N_19043,N_18138,N_17968);
nand U19044 (N_19044,N_18223,N_18231);
and U19045 (N_19045,N_18350,N_17970);
xor U19046 (N_19046,N_18192,N_17849);
xor U19047 (N_19047,N_17890,N_18196);
nand U19048 (N_19048,N_17668,N_17788);
xor U19049 (N_19049,N_18220,N_17838);
nor U19050 (N_19050,N_17875,N_17843);
and U19051 (N_19051,N_18297,N_17924);
nand U19052 (N_19052,N_18314,N_18034);
nor U19053 (N_19053,N_18344,N_17873);
nor U19054 (N_19054,N_18142,N_18217);
xor U19055 (N_19055,N_18314,N_18346);
nor U19056 (N_19056,N_17975,N_18386);
nand U19057 (N_19057,N_18303,N_18052);
nor U19058 (N_19058,N_18309,N_18358);
xor U19059 (N_19059,N_18132,N_18276);
and U19060 (N_19060,N_17785,N_18163);
nor U19061 (N_19061,N_18335,N_18352);
nor U19062 (N_19062,N_18366,N_18168);
nand U19063 (N_19063,N_18209,N_17943);
xnor U19064 (N_19064,N_17973,N_18161);
nor U19065 (N_19065,N_18266,N_18230);
nand U19066 (N_19066,N_17753,N_18072);
xor U19067 (N_19067,N_17635,N_17614);
or U19068 (N_19068,N_18177,N_18170);
or U19069 (N_19069,N_17745,N_17804);
xnor U19070 (N_19070,N_17931,N_18150);
and U19071 (N_19071,N_17703,N_17639);
or U19072 (N_19072,N_17773,N_17697);
xor U19073 (N_19073,N_17866,N_17985);
and U19074 (N_19074,N_17974,N_18135);
nand U19075 (N_19075,N_17909,N_18392);
and U19076 (N_19076,N_17940,N_18001);
or U19077 (N_19077,N_18234,N_17950);
nor U19078 (N_19078,N_17628,N_17656);
or U19079 (N_19079,N_18366,N_18195);
or U19080 (N_19080,N_18252,N_17993);
or U19081 (N_19081,N_18177,N_17628);
xor U19082 (N_19082,N_18383,N_18090);
nor U19083 (N_19083,N_18297,N_17870);
xnor U19084 (N_19084,N_18137,N_17702);
nand U19085 (N_19085,N_17979,N_17950);
xnor U19086 (N_19086,N_17872,N_17949);
nand U19087 (N_19087,N_18304,N_17919);
and U19088 (N_19088,N_17735,N_18081);
and U19089 (N_19089,N_17850,N_18287);
nor U19090 (N_19090,N_17820,N_17781);
nor U19091 (N_19091,N_17721,N_18061);
xor U19092 (N_19092,N_17800,N_17891);
xnor U19093 (N_19093,N_17752,N_18078);
or U19094 (N_19094,N_18379,N_18104);
or U19095 (N_19095,N_17903,N_17736);
or U19096 (N_19096,N_18055,N_18284);
nand U19097 (N_19097,N_18254,N_18046);
or U19098 (N_19098,N_18252,N_18268);
and U19099 (N_19099,N_17870,N_18082);
xnor U19100 (N_19100,N_17761,N_17717);
and U19101 (N_19101,N_18193,N_18125);
nor U19102 (N_19102,N_18362,N_18004);
nor U19103 (N_19103,N_17699,N_17856);
nand U19104 (N_19104,N_18034,N_17806);
and U19105 (N_19105,N_18032,N_17760);
xnor U19106 (N_19106,N_18295,N_17629);
or U19107 (N_19107,N_18230,N_17619);
or U19108 (N_19108,N_17887,N_18220);
and U19109 (N_19109,N_17996,N_17677);
nor U19110 (N_19110,N_17644,N_18262);
or U19111 (N_19111,N_18291,N_17814);
nor U19112 (N_19112,N_18233,N_17655);
or U19113 (N_19113,N_17919,N_18344);
or U19114 (N_19114,N_18137,N_17900);
and U19115 (N_19115,N_18071,N_17802);
and U19116 (N_19116,N_18205,N_18143);
xor U19117 (N_19117,N_18159,N_17914);
or U19118 (N_19118,N_18399,N_18171);
nor U19119 (N_19119,N_17872,N_17697);
xor U19120 (N_19120,N_17784,N_17840);
or U19121 (N_19121,N_18389,N_17667);
and U19122 (N_19122,N_18369,N_18360);
and U19123 (N_19123,N_18316,N_18048);
or U19124 (N_19124,N_18047,N_17731);
nor U19125 (N_19125,N_17660,N_18380);
nor U19126 (N_19126,N_17861,N_18031);
xor U19127 (N_19127,N_17936,N_18188);
nor U19128 (N_19128,N_17913,N_18172);
or U19129 (N_19129,N_17842,N_17646);
nand U19130 (N_19130,N_18205,N_17810);
nor U19131 (N_19131,N_17878,N_17750);
nand U19132 (N_19132,N_17896,N_18378);
xnor U19133 (N_19133,N_18005,N_18334);
or U19134 (N_19134,N_17902,N_18270);
or U19135 (N_19135,N_18115,N_17924);
and U19136 (N_19136,N_17686,N_18183);
or U19137 (N_19137,N_17700,N_17897);
xor U19138 (N_19138,N_17860,N_18066);
nor U19139 (N_19139,N_18285,N_18343);
or U19140 (N_19140,N_18165,N_17735);
xnor U19141 (N_19141,N_18189,N_18350);
nand U19142 (N_19142,N_17735,N_18059);
xor U19143 (N_19143,N_17723,N_17646);
nor U19144 (N_19144,N_18033,N_18058);
nor U19145 (N_19145,N_18171,N_18249);
or U19146 (N_19146,N_18183,N_17946);
xnor U19147 (N_19147,N_18264,N_17864);
nor U19148 (N_19148,N_17710,N_18233);
nand U19149 (N_19149,N_17918,N_18075);
or U19150 (N_19150,N_17771,N_17874);
nor U19151 (N_19151,N_18020,N_18232);
or U19152 (N_19152,N_17710,N_18199);
or U19153 (N_19153,N_17755,N_17995);
nand U19154 (N_19154,N_18019,N_17619);
nand U19155 (N_19155,N_17896,N_18191);
nor U19156 (N_19156,N_17820,N_17893);
and U19157 (N_19157,N_17755,N_18211);
or U19158 (N_19158,N_18227,N_18276);
and U19159 (N_19159,N_17864,N_18239);
nand U19160 (N_19160,N_18389,N_17630);
or U19161 (N_19161,N_17999,N_18125);
xor U19162 (N_19162,N_17925,N_18271);
nor U19163 (N_19163,N_17701,N_18138);
nand U19164 (N_19164,N_18101,N_17838);
nor U19165 (N_19165,N_18268,N_18242);
nor U19166 (N_19166,N_17875,N_17691);
nand U19167 (N_19167,N_17605,N_17752);
or U19168 (N_19168,N_17700,N_18112);
or U19169 (N_19169,N_18115,N_17703);
xnor U19170 (N_19170,N_17939,N_18153);
and U19171 (N_19171,N_17837,N_17866);
and U19172 (N_19172,N_17879,N_18350);
nand U19173 (N_19173,N_17943,N_18248);
and U19174 (N_19174,N_17773,N_18365);
and U19175 (N_19175,N_17648,N_17909);
xor U19176 (N_19176,N_17880,N_18356);
and U19177 (N_19177,N_18052,N_18328);
xnor U19178 (N_19178,N_17748,N_17637);
nand U19179 (N_19179,N_18169,N_17706);
nand U19180 (N_19180,N_18157,N_17768);
nor U19181 (N_19181,N_17956,N_17837);
nor U19182 (N_19182,N_17762,N_17724);
nand U19183 (N_19183,N_17919,N_18397);
nand U19184 (N_19184,N_17972,N_18066);
or U19185 (N_19185,N_18322,N_18118);
nor U19186 (N_19186,N_18298,N_17685);
and U19187 (N_19187,N_17912,N_18323);
or U19188 (N_19188,N_18314,N_17646);
xnor U19189 (N_19189,N_17708,N_17654);
xor U19190 (N_19190,N_17603,N_18271);
xor U19191 (N_19191,N_18135,N_17944);
nand U19192 (N_19192,N_18131,N_18173);
xor U19193 (N_19193,N_18375,N_17887);
or U19194 (N_19194,N_18321,N_18259);
or U19195 (N_19195,N_17826,N_17701);
or U19196 (N_19196,N_18377,N_17897);
nor U19197 (N_19197,N_18296,N_18256);
nor U19198 (N_19198,N_17715,N_18295);
or U19199 (N_19199,N_18120,N_18103);
or U19200 (N_19200,N_19088,N_18408);
nand U19201 (N_19201,N_18919,N_18495);
and U19202 (N_19202,N_18897,N_19073);
and U19203 (N_19203,N_18908,N_18704);
nand U19204 (N_19204,N_18899,N_18861);
nor U19205 (N_19205,N_18541,N_19124);
or U19206 (N_19206,N_18810,N_18656);
nand U19207 (N_19207,N_18848,N_19009);
xnor U19208 (N_19208,N_19024,N_18869);
and U19209 (N_19209,N_18748,N_19185);
xor U19210 (N_19210,N_18996,N_18546);
and U19211 (N_19211,N_19065,N_18509);
nand U19212 (N_19212,N_18815,N_18809);
xnor U19213 (N_19213,N_18414,N_18781);
xor U19214 (N_19214,N_19197,N_18739);
or U19215 (N_19215,N_18792,N_18900);
xnor U19216 (N_19216,N_18597,N_19011);
nor U19217 (N_19217,N_18521,N_19178);
or U19218 (N_19218,N_18853,N_18641);
and U19219 (N_19219,N_19006,N_18403);
and U19220 (N_19220,N_19143,N_18516);
nor U19221 (N_19221,N_18494,N_18978);
or U19222 (N_19222,N_19007,N_18630);
nor U19223 (N_19223,N_18690,N_18746);
nand U19224 (N_19224,N_18984,N_18508);
and U19225 (N_19225,N_18967,N_18450);
or U19226 (N_19226,N_18581,N_19125);
nand U19227 (N_19227,N_18742,N_18816);
and U19228 (N_19228,N_19162,N_18913);
and U19229 (N_19229,N_19020,N_18895);
nor U19230 (N_19230,N_18664,N_19099);
and U19231 (N_19231,N_18653,N_18573);
and U19232 (N_19232,N_18836,N_19035);
nor U19233 (N_19233,N_18929,N_18717);
xnor U19234 (N_19234,N_18604,N_18842);
or U19235 (N_19235,N_18542,N_18587);
and U19236 (N_19236,N_18821,N_18472);
nor U19237 (N_19237,N_18938,N_18839);
and U19238 (N_19238,N_18902,N_18547);
or U19239 (N_19239,N_18773,N_18980);
xnor U19240 (N_19240,N_18402,N_18798);
nor U19241 (N_19241,N_19174,N_19087);
nand U19242 (N_19242,N_18598,N_18670);
nor U19243 (N_19243,N_19127,N_18669);
nand U19244 (N_19244,N_18496,N_18483);
nor U19245 (N_19245,N_18756,N_18813);
nor U19246 (N_19246,N_19026,N_18990);
or U19247 (N_19247,N_19091,N_18804);
nor U19248 (N_19248,N_19058,N_18763);
xnor U19249 (N_19249,N_19064,N_18624);
and U19250 (N_19250,N_18885,N_18643);
xor U19251 (N_19251,N_18966,N_18969);
xnor U19252 (N_19252,N_18805,N_18918);
nand U19253 (N_19253,N_19140,N_19031);
xnor U19254 (N_19254,N_18735,N_18401);
or U19255 (N_19255,N_18847,N_18903);
xor U19256 (N_19256,N_18826,N_18466);
nor U19257 (N_19257,N_18436,N_19160);
xor U19258 (N_19258,N_18762,N_18473);
xnor U19259 (N_19259,N_18979,N_18513);
nand U19260 (N_19260,N_18755,N_19086);
nand U19261 (N_19261,N_18820,N_18824);
or U19262 (N_19262,N_18727,N_18648);
or U19263 (N_19263,N_18993,N_19013);
and U19264 (N_19264,N_18831,N_19032);
nand U19265 (N_19265,N_19167,N_18437);
or U19266 (N_19266,N_18609,N_18991);
xor U19267 (N_19267,N_18960,N_18412);
nand U19268 (N_19268,N_18556,N_18856);
or U19269 (N_19269,N_19089,N_18439);
and U19270 (N_19270,N_18603,N_18877);
xnor U19271 (N_19271,N_18927,N_18775);
xnor U19272 (N_19272,N_19102,N_19153);
nand U19273 (N_19273,N_18757,N_18552);
xnor U19274 (N_19274,N_18779,N_18713);
and U19275 (N_19275,N_18997,N_18544);
or U19276 (N_19276,N_18693,N_18409);
xor U19277 (N_19277,N_18589,N_19095);
and U19278 (N_19278,N_19169,N_19199);
nand U19279 (N_19279,N_18873,N_18404);
or U19280 (N_19280,N_18768,N_18889);
nand U19281 (N_19281,N_18711,N_18553);
nand U19282 (N_19282,N_18788,N_18501);
xnor U19283 (N_19283,N_18539,N_18844);
nor U19284 (N_19284,N_18837,N_18658);
nor U19285 (N_19285,N_18920,N_18534);
nor U19286 (N_19286,N_18600,N_19093);
and U19287 (N_19287,N_19131,N_18857);
nand U19288 (N_19288,N_18745,N_18536);
nor U19289 (N_19289,N_18944,N_18417);
and U19290 (N_19290,N_18761,N_18968);
and U19291 (N_19291,N_18667,N_18550);
nor U19292 (N_19292,N_18945,N_19021);
nand U19293 (N_19293,N_19048,N_18580);
xor U19294 (N_19294,N_18794,N_18703);
and U19295 (N_19295,N_18500,N_18796);
and U19296 (N_19296,N_18965,N_18622);
nand U19297 (N_19297,N_18971,N_19076);
nand U19298 (N_19298,N_18679,N_18685);
nor U19299 (N_19299,N_18753,N_18435);
and U19300 (N_19300,N_18705,N_18935);
xnor U19301 (N_19301,N_18493,N_18766);
xnor U19302 (N_19302,N_18479,N_18531);
nor U19303 (N_19303,N_18645,N_18465);
nand U19304 (N_19304,N_18649,N_18486);
nand U19305 (N_19305,N_19193,N_18438);
xnor U19306 (N_19306,N_18497,N_19052);
nor U19307 (N_19307,N_18575,N_18511);
or U19308 (N_19308,N_18599,N_19106);
xor U19309 (N_19309,N_18429,N_19036);
nand U19310 (N_19310,N_19196,N_18778);
and U19311 (N_19311,N_18988,N_18817);
and U19312 (N_19312,N_18886,N_18750);
nand U19313 (N_19313,N_18563,N_18661);
xor U19314 (N_19314,N_18596,N_19018);
and U19315 (N_19315,N_18428,N_19016);
nand U19316 (N_19316,N_19156,N_18904);
nor U19317 (N_19317,N_18449,N_18852);
nand U19318 (N_19318,N_19141,N_18887);
or U19319 (N_19319,N_18652,N_18478);
nand U19320 (N_19320,N_19150,N_18623);
nand U19321 (N_19321,N_19175,N_18973);
xor U19322 (N_19322,N_18884,N_19038);
xnor U19323 (N_19323,N_18941,N_19066);
nor U19324 (N_19324,N_18448,N_19133);
or U19325 (N_19325,N_18456,N_18870);
and U19326 (N_19326,N_18601,N_19028);
nand U19327 (N_19327,N_19062,N_19115);
xor U19328 (N_19328,N_18865,N_18590);
xor U19329 (N_19329,N_19136,N_18424);
xor U19330 (N_19330,N_19050,N_18827);
nor U19331 (N_19331,N_19117,N_18504);
nor U19332 (N_19332,N_19148,N_19039);
nor U19333 (N_19333,N_18460,N_18636);
nor U19334 (N_19334,N_18795,N_18642);
or U19335 (N_19335,N_18738,N_19033);
xor U19336 (N_19336,N_19154,N_18832);
xnor U19337 (N_19337,N_18416,N_18663);
or U19338 (N_19338,N_18946,N_18540);
and U19339 (N_19339,N_18789,N_18606);
nand U19340 (N_19340,N_18673,N_18519);
xor U19341 (N_19341,N_18894,N_18771);
or U19342 (N_19342,N_19015,N_18505);
xnor U19343 (N_19343,N_19135,N_19166);
and U19344 (N_19344,N_18879,N_18999);
or U19345 (N_19345,N_18684,N_18480);
xor U19346 (N_19346,N_18744,N_18931);
or U19347 (N_19347,N_18660,N_18721);
and U19348 (N_19348,N_19137,N_19004);
xnor U19349 (N_19349,N_19054,N_18593);
and U19350 (N_19350,N_18605,N_18972);
nand U19351 (N_19351,N_19138,N_18706);
or U19352 (N_19352,N_18614,N_18625);
and U19353 (N_19353,N_18862,N_18440);
and U19354 (N_19354,N_18469,N_18898);
and U19355 (N_19355,N_18740,N_18595);
nor U19356 (N_19356,N_18674,N_18953);
nand U19357 (N_19357,N_18916,N_18492);
nor U19358 (N_19358,N_19030,N_18503);
or U19359 (N_19359,N_18621,N_18880);
and U19360 (N_19360,N_18883,N_19147);
nand U19361 (N_19361,N_18785,N_19134);
xor U19362 (N_19362,N_18634,N_19042);
and U19363 (N_19363,N_18797,N_18459);
xor U19364 (N_19364,N_18724,N_18940);
xnor U19365 (N_19365,N_19155,N_18400);
nor U19366 (N_19366,N_18627,N_18825);
nand U19367 (N_19367,N_19126,N_18992);
nand U19368 (N_19368,N_18567,N_18675);
and U19369 (N_19369,N_18640,N_18922);
xnor U19370 (N_19370,N_19025,N_18612);
or U19371 (N_19371,N_18850,N_19080);
and U19372 (N_19372,N_18561,N_18475);
or U19373 (N_19373,N_18720,N_19188);
or U19374 (N_19374,N_19023,N_18680);
and U19375 (N_19375,N_18729,N_19097);
xor U19376 (N_19376,N_18682,N_19128);
nor U19377 (N_19377,N_19149,N_18970);
or U19378 (N_19378,N_19075,N_18714);
xnor U19379 (N_19379,N_18422,N_18974);
nor U19380 (N_19380,N_18583,N_18780);
nand U19381 (N_19381,N_18989,N_19057);
nor U19382 (N_19382,N_18591,N_18770);
nor U19383 (N_19383,N_18543,N_18566);
xnor U19384 (N_19384,N_19053,N_19070);
xnor U19385 (N_19385,N_18558,N_18777);
nand U19386 (N_19386,N_18787,N_18925);
nand U19387 (N_19387,N_18823,N_19047);
and U19388 (N_19388,N_18602,N_19094);
and U19389 (N_19389,N_19130,N_18774);
and U19390 (N_19390,N_18526,N_18863);
or U19391 (N_19391,N_18607,N_19002);
nor U19392 (N_19392,N_18854,N_18515);
nand U19393 (N_19393,N_19179,N_18518);
or U19394 (N_19394,N_18951,N_18851);
and U19395 (N_19395,N_18699,N_19000);
nor U19396 (N_19396,N_19029,N_18876);
nor U19397 (N_19397,N_18843,N_19186);
or U19398 (N_19398,N_18783,N_18523);
nand U19399 (N_19399,N_19177,N_18845);
nor U19400 (N_19400,N_18741,N_18710);
and U19401 (N_19401,N_18822,N_18431);
nor U19402 (N_19402,N_18632,N_18864);
xnor U19403 (N_19403,N_18507,N_19017);
xor U19404 (N_19404,N_18426,N_18882);
xnor U19405 (N_19405,N_19192,N_18579);
nor U19406 (N_19406,N_18734,N_18678);
and U19407 (N_19407,N_18793,N_18430);
nor U19408 (N_19408,N_18712,N_19168);
xnor U19409 (N_19409,N_18709,N_18906);
nand U19410 (N_19410,N_18737,N_18538);
nor U19411 (N_19411,N_18617,N_18814);
nand U19412 (N_19412,N_18976,N_18432);
and U19413 (N_19413,N_18584,N_18671);
nor U19414 (N_19414,N_18665,N_18878);
and U19415 (N_19415,N_18828,N_19043);
nor U19416 (N_19416,N_18462,N_19119);
nand U19417 (N_19417,N_19181,N_19142);
and U19418 (N_19418,N_18803,N_18866);
nand U19419 (N_19419,N_19146,N_18517);
nand U19420 (N_19420,N_19012,N_19069);
and U19421 (N_19421,N_18835,N_18514);
xnor U19422 (N_19422,N_18691,N_18715);
nor U19423 (N_19423,N_18707,N_18405);
and U19424 (N_19424,N_19158,N_18421);
or U19425 (N_19425,N_18743,N_18926);
nor U19426 (N_19426,N_18985,N_18659);
or U19427 (N_19427,N_18957,N_19083);
xnor U19428 (N_19428,N_18427,N_18445);
nand U19429 (N_19429,N_18611,N_18628);
nand U19430 (N_19430,N_18719,N_18618);
nor U19431 (N_19431,N_19123,N_18451);
nor U19432 (N_19432,N_19191,N_18644);
nor U19433 (N_19433,N_19139,N_19040);
xor U19434 (N_19434,N_18728,N_18752);
xor U19435 (N_19435,N_18819,N_18891);
and U19436 (N_19436,N_18930,N_18535);
nand U19437 (N_19437,N_18829,N_19045);
or U19438 (N_19438,N_18463,N_18812);
xnor U19439 (N_19439,N_18950,N_18551);
and U19440 (N_19440,N_18694,N_18565);
xnor U19441 (N_19441,N_18754,N_18808);
or U19442 (N_19442,N_19046,N_18731);
xnor U19443 (N_19443,N_18681,N_18868);
nand U19444 (N_19444,N_18942,N_18568);
nand U19445 (N_19445,N_18616,N_19077);
xor U19446 (N_19446,N_18489,N_18470);
nor U19447 (N_19447,N_18646,N_18655);
xnor U19448 (N_19448,N_19090,N_18928);
nand U19449 (N_19449,N_19072,N_18994);
nor U19450 (N_19450,N_18423,N_18963);
nor U19451 (N_19451,N_19098,N_18910);
xor U19452 (N_19452,N_18716,N_18924);
nand U19453 (N_19453,N_18613,N_18441);
xor U19454 (N_19454,N_19085,N_18725);
nand U19455 (N_19455,N_18917,N_19116);
or U19456 (N_19456,N_19105,N_18830);
and U19457 (N_19457,N_18415,N_18672);
nand U19458 (N_19458,N_18764,N_18800);
nor U19459 (N_19459,N_18533,N_18477);
nor U19460 (N_19460,N_19060,N_18512);
nor U19461 (N_19461,N_18686,N_18801);
and U19462 (N_19462,N_19037,N_18776);
or U19463 (N_19463,N_18695,N_18954);
or U19464 (N_19464,N_19184,N_19172);
nor U19465 (N_19465,N_19055,N_19121);
nand U19466 (N_19466,N_18867,N_18859);
or U19467 (N_19467,N_19061,N_18406);
or U19468 (N_19468,N_19059,N_18442);
nand U19469 (N_19469,N_18912,N_18502);
nand U19470 (N_19470,N_18998,N_19014);
or U19471 (N_19471,N_19107,N_18932);
nor U19472 (N_19472,N_19129,N_18548);
and U19473 (N_19473,N_18697,N_18959);
nand U19474 (N_19474,N_18555,N_18615);
or U19475 (N_19475,N_18958,N_18807);
nand U19476 (N_19476,N_19152,N_18983);
nand U19477 (N_19477,N_18948,N_19079);
nor U19478 (N_19478,N_18549,N_18911);
or U19479 (N_19479,N_18443,N_18557);
xor U19480 (N_19480,N_18410,N_18901);
xnor U19481 (N_19481,N_18458,N_18767);
nand U19482 (N_19482,N_18708,N_19180);
nand U19483 (N_19483,N_19111,N_18446);
nor U19484 (N_19484,N_19161,N_18457);
nor U19485 (N_19485,N_18564,N_19071);
nor U19486 (N_19486,N_19078,N_19194);
nor U19487 (N_19487,N_18955,N_19103);
nand U19488 (N_19488,N_18524,N_18453);
and U19489 (N_19489,N_19051,N_18855);
nand U19490 (N_19490,N_18461,N_19092);
xor U19491 (N_19491,N_18425,N_18892);
or U19492 (N_19492,N_19034,N_18937);
xor U19493 (N_19493,N_18760,N_18571);
xnor U19494 (N_19494,N_18975,N_18841);
xnor U19495 (N_19495,N_19173,N_18818);
xor U19496 (N_19496,N_19001,N_19100);
nor U19497 (N_19497,N_19122,N_18482);
nand U19498 (N_19498,N_18806,N_18525);
and U19499 (N_19499,N_19108,N_18982);
nor U19500 (N_19500,N_18488,N_19190);
and U19501 (N_19501,N_19170,N_18939);
xnor U19502 (N_19502,N_19068,N_18576);
nand U19503 (N_19503,N_18474,N_18677);
or U19504 (N_19504,N_18981,N_19159);
or U19505 (N_19505,N_19198,N_19003);
nand U19506 (N_19506,N_18802,N_18582);
nor U19507 (N_19507,N_19164,N_18730);
and U19508 (N_19508,N_18858,N_18433);
and U19509 (N_19509,N_19104,N_19182);
nand U19510 (N_19510,N_18452,N_18657);
or U19511 (N_19511,N_18639,N_18620);
or U19512 (N_19512,N_18718,N_18545);
nor U19513 (N_19513,N_19157,N_18413);
nor U19514 (N_19514,N_18933,N_18529);
or U19515 (N_19515,N_19019,N_18949);
nand U19516 (N_19516,N_18875,N_18947);
nor U19517 (N_19517,N_18896,N_19084);
nor U19518 (N_19518,N_19110,N_18487);
nor U19519 (N_19519,N_18554,N_18676);
nor U19520 (N_19520,N_18633,N_18733);
and U19521 (N_19521,N_18471,N_18592);
nor U19522 (N_19522,N_18484,N_18419);
and U19523 (N_19523,N_18464,N_18528);
nor U19524 (N_19524,N_18995,N_18689);
nor U19525 (N_19525,N_18586,N_18881);
nor U19526 (N_19526,N_19176,N_18467);
and U19527 (N_19527,N_18476,N_18570);
nor U19528 (N_19528,N_18418,N_18687);
and U19529 (N_19529,N_18688,N_19010);
xor U19530 (N_19530,N_18594,N_18637);
xor U19531 (N_19531,N_19145,N_18700);
and U19532 (N_19532,N_18610,N_18987);
xnor U19533 (N_19533,N_18510,N_18562);
or U19534 (N_19534,N_18874,N_18838);
nor U19535 (N_19535,N_18654,N_18608);
nor U19536 (N_19536,N_18638,N_18769);
nand U19537 (N_19537,N_19005,N_18666);
and U19538 (N_19538,N_18647,N_18833);
nor U19539 (N_19539,N_18407,N_18702);
xor U19540 (N_19540,N_18444,N_18952);
or U19541 (N_19541,N_18499,N_18964);
nand U19542 (N_19542,N_18520,N_18668);
nor U19543 (N_19543,N_19044,N_18588);
and U19544 (N_19544,N_18698,N_19096);
and U19545 (N_19545,N_18651,N_19082);
nor U19546 (N_19546,N_18522,N_18572);
xor U19547 (N_19547,N_18751,N_19144);
xor U19548 (N_19548,N_18726,N_18786);
or U19549 (N_19549,N_18585,N_18915);
xnor U19550 (N_19550,N_19189,N_18732);
or U19551 (N_19551,N_18914,N_18956);
nand U19552 (N_19552,N_19049,N_19132);
nand U19553 (N_19553,N_18532,N_18559);
and U19554 (N_19554,N_18723,N_18888);
or U19555 (N_19555,N_19067,N_18890);
nand U19556 (N_19556,N_18447,N_18934);
xor U19557 (N_19557,N_18811,N_19113);
and U19558 (N_19558,N_18468,N_18790);
xnor U19559 (N_19559,N_18747,N_18683);
nand U19560 (N_19560,N_18782,N_18696);
xor U19561 (N_19561,N_19027,N_18635);
or U19562 (N_19562,N_18455,N_18420);
or U19563 (N_19563,N_18626,N_18560);
nand U19564 (N_19564,N_18784,N_18631);
and U19565 (N_19565,N_18871,N_19163);
and U19566 (N_19566,N_19008,N_18846);
and U19567 (N_19567,N_18569,N_18905);
nor U19568 (N_19568,N_18921,N_18577);
and U19569 (N_19569,N_18791,N_18527);
nand U19570 (N_19570,N_18961,N_19187);
nand U19571 (N_19571,N_19041,N_19112);
and U19572 (N_19572,N_18537,N_18943);
or U19573 (N_19573,N_18530,N_18434);
and U19574 (N_19574,N_18849,N_18619);
nand U19575 (N_19575,N_18772,N_18650);
and U19576 (N_19576,N_18701,N_18749);
nand U19577 (N_19577,N_19151,N_19109);
or U19578 (N_19578,N_18923,N_18977);
or U19579 (N_19579,N_19101,N_18872);
nand U19580 (N_19580,N_18907,N_18481);
nand U19581 (N_19581,N_18893,N_18986);
nand U19582 (N_19582,N_18758,N_18578);
or U19583 (N_19583,N_18491,N_18629);
or U19584 (N_19584,N_18936,N_18692);
nor U19585 (N_19585,N_18662,N_18498);
xor U19586 (N_19586,N_19081,N_18909);
nor U19587 (N_19587,N_18736,N_18840);
nor U19588 (N_19588,N_18490,N_18485);
or U19589 (N_19589,N_19165,N_18411);
nor U19590 (N_19590,N_19022,N_19120);
nand U19591 (N_19591,N_18722,N_18574);
or U19592 (N_19592,N_18759,N_18506);
and U19593 (N_19593,N_19063,N_18799);
nand U19594 (N_19594,N_19195,N_19056);
and U19595 (N_19595,N_19114,N_19183);
and U19596 (N_19596,N_18860,N_18962);
xnor U19597 (N_19597,N_18765,N_18454);
xnor U19598 (N_19598,N_19171,N_18834);
nor U19599 (N_19599,N_19074,N_19118);
nor U19600 (N_19600,N_18486,N_18688);
nor U19601 (N_19601,N_18549,N_18871);
or U19602 (N_19602,N_18827,N_18735);
xnor U19603 (N_19603,N_18622,N_18657);
nor U19604 (N_19604,N_19196,N_19016);
or U19605 (N_19605,N_18698,N_18949);
or U19606 (N_19606,N_18492,N_18775);
nor U19607 (N_19607,N_18959,N_18784);
nand U19608 (N_19608,N_19098,N_18489);
or U19609 (N_19609,N_18934,N_18433);
nor U19610 (N_19610,N_18762,N_19167);
nand U19611 (N_19611,N_18820,N_18621);
nand U19612 (N_19612,N_18548,N_18568);
or U19613 (N_19613,N_19197,N_18422);
or U19614 (N_19614,N_18457,N_18734);
or U19615 (N_19615,N_18672,N_18524);
nor U19616 (N_19616,N_19021,N_19159);
nand U19617 (N_19617,N_19137,N_18682);
xnor U19618 (N_19618,N_19052,N_18484);
and U19619 (N_19619,N_18752,N_18845);
and U19620 (N_19620,N_18835,N_18534);
xnor U19621 (N_19621,N_18724,N_18758);
nor U19622 (N_19622,N_19083,N_18610);
and U19623 (N_19623,N_18962,N_18445);
and U19624 (N_19624,N_18415,N_18556);
xor U19625 (N_19625,N_18801,N_19057);
xor U19626 (N_19626,N_18882,N_18888);
xor U19627 (N_19627,N_19172,N_19042);
nor U19628 (N_19628,N_19037,N_19048);
and U19629 (N_19629,N_19056,N_18766);
nor U19630 (N_19630,N_19128,N_18881);
nand U19631 (N_19631,N_19196,N_19153);
nand U19632 (N_19632,N_18711,N_18916);
nand U19633 (N_19633,N_18592,N_18823);
xnor U19634 (N_19634,N_18956,N_19139);
or U19635 (N_19635,N_18461,N_18453);
xnor U19636 (N_19636,N_19127,N_18792);
and U19637 (N_19637,N_18563,N_19088);
nand U19638 (N_19638,N_18411,N_18807);
or U19639 (N_19639,N_19100,N_19077);
nor U19640 (N_19640,N_19139,N_18546);
nand U19641 (N_19641,N_18691,N_19100);
and U19642 (N_19642,N_18456,N_18542);
nor U19643 (N_19643,N_18822,N_18970);
and U19644 (N_19644,N_18600,N_18923);
xnor U19645 (N_19645,N_18714,N_18476);
or U19646 (N_19646,N_18953,N_18449);
xor U19647 (N_19647,N_19077,N_18455);
nor U19648 (N_19648,N_18650,N_19195);
or U19649 (N_19649,N_18810,N_18764);
xor U19650 (N_19650,N_19141,N_18776);
and U19651 (N_19651,N_18528,N_18582);
or U19652 (N_19652,N_18433,N_19076);
nand U19653 (N_19653,N_18474,N_18495);
xnor U19654 (N_19654,N_18502,N_18783);
nand U19655 (N_19655,N_18578,N_19110);
nor U19656 (N_19656,N_18576,N_18801);
xnor U19657 (N_19657,N_19004,N_18840);
nor U19658 (N_19658,N_18867,N_18409);
and U19659 (N_19659,N_19060,N_18428);
nand U19660 (N_19660,N_18830,N_18626);
nand U19661 (N_19661,N_19044,N_18826);
nor U19662 (N_19662,N_18525,N_18565);
nor U19663 (N_19663,N_18588,N_18618);
nand U19664 (N_19664,N_18747,N_18534);
xor U19665 (N_19665,N_18522,N_19078);
xnor U19666 (N_19666,N_18868,N_19130);
nand U19667 (N_19667,N_18830,N_18424);
nand U19668 (N_19668,N_18875,N_18769);
nand U19669 (N_19669,N_18494,N_18403);
and U19670 (N_19670,N_18861,N_18508);
and U19671 (N_19671,N_18626,N_18617);
nand U19672 (N_19672,N_18988,N_18538);
and U19673 (N_19673,N_18855,N_19158);
nand U19674 (N_19674,N_18942,N_19131);
nand U19675 (N_19675,N_18535,N_18485);
nor U19676 (N_19676,N_19154,N_18497);
nor U19677 (N_19677,N_18796,N_19016);
and U19678 (N_19678,N_18839,N_18967);
nand U19679 (N_19679,N_18725,N_18467);
xnor U19680 (N_19680,N_19012,N_18680);
or U19681 (N_19681,N_19168,N_18724);
nand U19682 (N_19682,N_18757,N_19137);
nand U19683 (N_19683,N_18893,N_19052);
nand U19684 (N_19684,N_18794,N_19041);
xnor U19685 (N_19685,N_19177,N_18917);
or U19686 (N_19686,N_19016,N_18697);
nor U19687 (N_19687,N_18894,N_19133);
xor U19688 (N_19688,N_19179,N_18964);
nor U19689 (N_19689,N_19121,N_18575);
xor U19690 (N_19690,N_18546,N_19034);
nor U19691 (N_19691,N_18409,N_19173);
and U19692 (N_19692,N_18708,N_18514);
xor U19693 (N_19693,N_19161,N_18957);
nor U19694 (N_19694,N_18774,N_18423);
or U19695 (N_19695,N_18899,N_19190);
and U19696 (N_19696,N_18954,N_19158);
xnor U19697 (N_19697,N_19008,N_18588);
xnor U19698 (N_19698,N_18913,N_19182);
and U19699 (N_19699,N_18834,N_19188);
nand U19700 (N_19700,N_18933,N_19140);
nor U19701 (N_19701,N_18674,N_19135);
nand U19702 (N_19702,N_18981,N_19179);
or U19703 (N_19703,N_18493,N_18665);
and U19704 (N_19704,N_18795,N_19024);
xnor U19705 (N_19705,N_18514,N_18501);
nor U19706 (N_19706,N_18616,N_18943);
nor U19707 (N_19707,N_18568,N_18624);
and U19708 (N_19708,N_18763,N_18953);
or U19709 (N_19709,N_18717,N_18465);
nand U19710 (N_19710,N_18940,N_18832);
and U19711 (N_19711,N_18944,N_18404);
nand U19712 (N_19712,N_18667,N_18927);
nor U19713 (N_19713,N_19002,N_19125);
and U19714 (N_19714,N_19049,N_18402);
nand U19715 (N_19715,N_18707,N_18661);
nand U19716 (N_19716,N_19102,N_18512);
and U19717 (N_19717,N_18587,N_18676);
nor U19718 (N_19718,N_18441,N_18572);
and U19719 (N_19719,N_19142,N_18728);
nor U19720 (N_19720,N_18748,N_19113);
nand U19721 (N_19721,N_18663,N_18922);
or U19722 (N_19722,N_18516,N_18400);
and U19723 (N_19723,N_18639,N_19089);
nor U19724 (N_19724,N_18963,N_19082);
nor U19725 (N_19725,N_18800,N_19164);
and U19726 (N_19726,N_18966,N_18458);
nor U19727 (N_19727,N_19118,N_19032);
nand U19728 (N_19728,N_19101,N_18506);
nor U19729 (N_19729,N_18611,N_18507);
or U19730 (N_19730,N_18808,N_19042);
nor U19731 (N_19731,N_18492,N_19090);
or U19732 (N_19732,N_18624,N_18953);
and U19733 (N_19733,N_18894,N_19136);
nor U19734 (N_19734,N_18966,N_18666);
or U19735 (N_19735,N_18551,N_19015);
xnor U19736 (N_19736,N_19195,N_18681);
nor U19737 (N_19737,N_18608,N_18984);
or U19738 (N_19738,N_18984,N_18459);
nand U19739 (N_19739,N_18771,N_18919);
and U19740 (N_19740,N_18930,N_18587);
and U19741 (N_19741,N_18883,N_18415);
nor U19742 (N_19742,N_18642,N_19138);
or U19743 (N_19743,N_18995,N_18816);
xor U19744 (N_19744,N_18689,N_18727);
nand U19745 (N_19745,N_18863,N_19128);
and U19746 (N_19746,N_19150,N_19088);
xor U19747 (N_19747,N_18934,N_18571);
and U19748 (N_19748,N_18595,N_18714);
or U19749 (N_19749,N_18916,N_18601);
or U19750 (N_19750,N_18876,N_19093);
nor U19751 (N_19751,N_18788,N_18711);
nand U19752 (N_19752,N_18787,N_18680);
nor U19753 (N_19753,N_18873,N_18662);
xnor U19754 (N_19754,N_19176,N_18657);
nor U19755 (N_19755,N_18534,N_18656);
nand U19756 (N_19756,N_18468,N_18712);
xnor U19757 (N_19757,N_18530,N_18719);
and U19758 (N_19758,N_18501,N_19012);
and U19759 (N_19759,N_18738,N_19180);
nor U19760 (N_19760,N_18825,N_18705);
or U19761 (N_19761,N_18659,N_19002);
or U19762 (N_19762,N_18854,N_18878);
or U19763 (N_19763,N_18769,N_18923);
nor U19764 (N_19764,N_18489,N_18462);
or U19765 (N_19765,N_18820,N_18684);
nand U19766 (N_19766,N_18471,N_18681);
nor U19767 (N_19767,N_18658,N_18770);
nor U19768 (N_19768,N_18722,N_18427);
xor U19769 (N_19769,N_19021,N_18869);
xor U19770 (N_19770,N_18942,N_19099);
nand U19771 (N_19771,N_18511,N_18510);
nand U19772 (N_19772,N_18999,N_19007);
or U19773 (N_19773,N_18709,N_18593);
and U19774 (N_19774,N_19065,N_18690);
xnor U19775 (N_19775,N_18959,N_19118);
xor U19776 (N_19776,N_18602,N_18699);
xor U19777 (N_19777,N_18588,N_18971);
nand U19778 (N_19778,N_18969,N_18822);
or U19779 (N_19779,N_19183,N_19057);
or U19780 (N_19780,N_18898,N_18574);
xnor U19781 (N_19781,N_18502,N_18951);
nand U19782 (N_19782,N_19040,N_19037);
and U19783 (N_19783,N_19132,N_18886);
nand U19784 (N_19784,N_19127,N_18530);
nand U19785 (N_19785,N_18478,N_18948);
nand U19786 (N_19786,N_18740,N_18816);
nand U19787 (N_19787,N_18663,N_18802);
nor U19788 (N_19788,N_19049,N_18513);
nand U19789 (N_19789,N_18897,N_18821);
and U19790 (N_19790,N_18566,N_19171);
xor U19791 (N_19791,N_18499,N_19027);
nand U19792 (N_19792,N_18716,N_18522);
nor U19793 (N_19793,N_18907,N_19035);
and U19794 (N_19794,N_18516,N_18953);
and U19795 (N_19795,N_18922,N_18433);
nor U19796 (N_19796,N_18563,N_18744);
and U19797 (N_19797,N_18898,N_18778);
and U19798 (N_19798,N_18446,N_18518);
nor U19799 (N_19799,N_19131,N_19177);
xnor U19800 (N_19800,N_18602,N_19035);
and U19801 (N_19801,N_19081,N_18432);
and U19802 (N_19802,N_18792,N_18989);
xor U19803 (N_19803,N_18730,N_18480);
nand U19804 (N_19804,N_18464,N_18584);
xor U19805 (N_19805,N_18823,N_18764);
or U19806 (N_19806,N_18712,N_19127);
and U19807 (N_19807,N_18576,N_19116);
nor U19808 (N_19808,N_19033,N_18748);
and U19809 (N_19809,N_18490,N_18694);
nor U19810 (N_19810,N_19038,N_18492);
and U19811 (N_19811,N_18612,N_18850);
xor U19812 (N_19812,N_19004,N_19068);
xor U19813 (N_19813,N_18911,N_18610);
or U19814 (N_19814,N_18651,N_18572);
and U19815 (N_19815,N_19195,N_18470);
or U19816 (N_19816,N_18870,N_18794);
xnor U19817 (N_19817,N_18579,N_18972);
nand U19818 (N_19818,N_19064,N_18957);
or U19819 (N_19819,N_19132,N_18690);
and U19820 (N_19820,N_19059,N_18630);
or U19821 (N_19821,N_18546,N_18530);
xor U19822 (N_19822,N_18641,N_18580);
and U19823 (N_19823,N_18679,N_18964);
nand U19824 (N_19824,N_18419,N_18546);
xnor U19825 (N_19825,N_19188,N_18818);
and U19826 (N_19826,N_18832,N_19094);
and U19827 (N_19827,N_18405,N_18864);
and U19828 (N_19828,N_18964,N_18619);
and U19829 (N_19829,N_19098,N_18595);
and U19830 (N_19830,N_19116,N_19026);
xor U19831 (N_19831,N_18765,N_18517);
xnor U19832 (N_19832,N_18597,N_19156);
nor U19833 (N_19833,N_19016,N_18957);
nand U19834 (N_19834,N_18964,N_19151);
xnor U19835 (N_19835,N_18619,N_19115);
or U19836 (N_19836,N_18467,N_18517);
xnor U19837 (N_19837,N_19155,N_18870);
xnor U19838 (N_19838,N_18436,N_19171);
nor U19839 (N_19839,N_18427,N_18719);
or U19840 (N_19840,N_18619,N_19025);
xnor U19841 (N_19841,N_18572,N_18984);
and U19842 (N_19842,N_18687,N_18930);
nand U19843 (N_19843,N_18986,N_18611);
and U19844 (N_19844,N_19033,N_19170);
xor U19845 (N_19845,N_18541,N_18551);
and U19846 (N_19846,N_18988,N_18800);
nand U19847 (N_19847,N_18738,N_18860);
or U19848 (N_19848,N_19096,N_18910);
xor U19849 (N_19849,N_18413,N_18854);
or U19850 (N_19850,N_19127,N_18908);
nor U19851 (N_19851,N_18481,N_18580);
and U19852 (N_19852,N_18810,N_19184);
or U19853 (N_19853,N_18750,N_18556);
or U19854 (N_19854,N_18523,N_18528);
xnor U19855 (N_19855,N_18873,N_18535);
xor U19856 (N_19856,N_19065,N_19014);
nor U19857 (N_19857,N_18724,N_19101);
or U19858 (N_19858,N_18975,N_18811);
or U19859 (N_19859,N_18830,N_19189);
nand U19860 (N_19860,N_19184,N_18815);
nor U19861 (N_19861,N_18888,N_18540);
nand U19862 (N_19862,N_18658,N_18740);
and U19863 (N_19863,N_18965,N_19118);
nand U19864 (N_19864,N_18921,N_18870);
and U19865 (N_19865,N_18452,N_18676);
and U19866 (N_19866,N_18654,N_18656);
xnor U19867 (N_19867,N_18468,N_18570);
nor U19868 (N_19868,N_18481,N_18776);
nand U19869 (N_19869,N_18522,N_18954);
xor U19870 (N_19870,N_19182,N_18599);
or U19871 (N_19871,N_18631,N_18603);
nand U19872 (N_19872,N_19064,N_18606);
xnor U19873 (N_19873,N_19086,N_19031);
nand U19874 (N_19874,N_18615,N_18926);
or U19875 (N_19875,N_18747,N_18554);
or U19876 (N_19876,N_19138,N_18717);
xnor U19877 (N_19877,N_18612,N_18733);
or U19878 (N_19878,N_18883,N_18837);
nand U19879 (N_19879,N_18657,N_19140);
nand U19880 (N_19880,N_18777,N_18897);
xor U19881 (N_19881,N_18403,N_18718);
xnor U19882 (N_19882,N_18863,N_18691);
xnor U19883 (N_19883,N_18449,N_18530);
nor U19884 (N_19884,N_19127,N_18445);
nor U19885 (N_19885,N_18962,N_18939);
nand U19886 (N_19886,N_18661,N_18739);
nand U19887 (N_19887,N_19193,N_18641);
nand U19888 (N_19888,N_19184,N_18797);
nand U19889 (N_19889,N_18616,N_18442);
and U19890 (N_19890,N_19110,N_18775);
nand U19891 (N_19891,N_18509,N_18787);
xor U19892 (N_19892,N_19075,N_19175);
and U19893 (N_19893,N_18455,N_18453);
xor U19894 (N_19894,N_18669,N_18618);
nor U19895 (N_19895,N_19099,N_18768);
xnor U19896 (N_19896,N_18859,N_18968);
or U19897 (N_19897,N_18822,N_18634);
xor U19898 (N_19898,N_18923,N_18553);
xnor U19899 (N_19899,N_18639,N_18821);
or U19900 (N_19900,N_18789,N_18847);
and U19901 (N_19901,N_19034,N_19079);
nand U19902 (N_19902,N_18646,N_18549);
and U19903 (N_19903,N_19116,N_19110);
and U19904 (N_19904,N_18829,N_18538);
and U19905 (N_19905,N_19195,N_18687);
or U19906 (N_19906,N_18507,N_18736);
nand U19907 (N_19907,N_18502,N_18527);
or U19908 (N_19908,N_18927,N_18751);
xnor U19909 (N_19909,N_18652,N_19033);
or U19910 (N_19910,N_19111,N_18763);
xnor U19911 (N_19911,N_19199,N_18519);
and U19912 (N_19912,N_18983,N_18791);
nand U19913 (N_19913,N_18486,N_18592);
or U19914 (N_19914,N_18459,N_18538);
nand U19915 (N_19915,N_19196,N_18754);
or U19916 (N_19916,N_19153,N_18996);
nand U19917 (N_19917,N_19063,N_18578);
and U19918 (N_19918,N_18465,N_18767);
nand U19919 (N_19919,N_19035,N_18884);
xnor U19920 (N_19920,N_18677,N_18469);
nand U19921 (N_19921,N_18675,N_18906);
nand U19922 (N_19922,N_18630,N_19130);
or U19923 (N_19923,N_18839,N_18972);
nor U19924 (N_19924,N_18436,N_18999);
nand U19925 (N_19925,N_18999,N_18662);
and U19926 (N_19926,N_18673,N_18496);
xnor U19927 (N_19927,N_18954,N_18931);
nand U19928 (N_19928,N_19125,N_18896);
nand U19929 (N_19929,N_18546,N_18668);
nor U19930 (N_19930,N_18539,N_18410);
nand U19931 (N_19931,N_19050,N_18512);
xnor U19932 (N_19932,N_18560,N_18824);
and U19933 (N_19933,N_18494,N_19131);
nand U19934 (N_19934,N_18721,N_19066);
and U19935 (N_19935,N_18931,N_18901);
nand U19936 (N_19936,N_18715,N_19090);
xor U19937 (N_19937,N_18402,N_18673);
xor U19938 (N_19938,N_18904,N_18682);
and U19939 (N_19939,N_18829,N_18571);
nand U19940 (N_19940,N_18685,N_18558);
nor U19941 (N_19941,N_18511,N_18746);
nor U19942 (N_19942,N_18498,N_19195);
or U19943 (N_19943,N_19035,N_18454);
nand U19944 (N_19944,N_18735,N_18425);
nand U19945 (N_19945,N_18742,N_18867);
or U19946 (N_19946,N_19185,N_18691);
nand U19947 (N_19947,N_18475,N_18434);
and U19948 (N_19948,N_18777,N_18714);
and U19949 (N_19949,N_18949,N_18747);
xnor U19950 (N_19950,N_19092,N_18434);
xnor U19951 (N_19951,N_18814,N_18674);
nand U19952 (N_19952,N_18556,N_18784);
nor U19953 (N_19953,N_19140,N_19012);
nor U19954 (N_19954,N_18724,N_18503);
xor U19955 (N_19955,N_19109,N_18699);
nand U19956 (N_19956,N_18634,N_18440);
or U19957 (N_19957,N_18793,N_19045);
xnor U19958 (N_19958,N_18781,N_19075);
xor U19959 (N_19959,N_18789,N_18873);
and U19960 (N_19960,N_18972,N_18746);
and U19961 (N_19961,N_18993,N_18888);
xnor U19962 (N_19962,N_18993,N_18639);
and U19963 (N_19963,N_19127,N_18977);
and U19964 (N_19964,N_18449,N_19116);
and U19965 (N_19965,N_18673,N_18458);
xnor U19966 (N_19966,N_19124,N_18779);
or U19967 (N_19967,N_18976,N_18693);
nor U19968 (N_19968,N_18912,N_18964);
xor U19969 (N_19969,N_18982,N_18587);
and U19970 (N_19970,N_18902,N_19094);
xnor U19971 (N_19971,N_18503,N_18754);
or U19972 (N_19972,N_18493,N_18588);
and U19973 (N_19973,N_19096,N_18613);
or U19974 (N_19974,N_18867,N_19155);
or U19975 (N_19975,N_18857,N_18421);
nor U19976 (N_19976,N_18627,N_18774);
xor U19977 (N_19977,N_18471,N_19099);
xor U19978 (N_19978,N_18706,N_18923);
nand U19979 (N_19979,N_18513,N_19199);
and U19980 (N_19980,N_18931,N_18890);
nand U19981 (N_19981,N_19000,N_18954);
and U19982 (N_19982,N_19006,N_19107);
nand U19983 (N_19983,N_18424,N_18483);
or U19984 (N_19984,N_18745,N_18422);
nor U19985 (N_19985,N_18424,N_18850);
and U19986 (N_19986,N_18401,N_18493);
xor U19987 (N_19987,N_19147,N_18651);
and U19988 (N_19988,N_19106,N_18766);
xor U19989 (N_19989,N_18817,N_18702);
xor U19990 (N_19990,N_19156,N_18680);
and U19991 (N_19991,N_18496,N_18890);
xnor U19992 (N_19992,N_19059,N_18750);
or U19993 (N_19993,N_18972,N_19009);
nand U19994 (N_19994,N_18423,N_18653);
nor U19995 (N_19995,N_18951,N_19007);
and U19996 (N_19996,N_19041,N_19121);
xnor U19997 (N_19997,N_18949,N_19057);
nand U19998 (N_19998,N_18756,N_18494);
or U19999 (N_19999,N_19174,N_18790);
or UO_0 (O_0,N_19304,N_19436);
nand UO_1 (O_1,N_19967,N_19988);
and UO_2 (O_2,N_19995,N_19771);
nand UO_3 (O_3,N_19764,N_19628);
xor UO_4 (O_4,N_19239,N_19648);
nand UO_5 (O_5,N_19668,N_19241);
xor UO_6 (O_6,N_19641,N_19341);
nand UO_7 (O_7,N_19819,N_19428);
xnor UO_8 (O_8,N_19235,N_19607);
nor UO_9 (O_9,N_19937,N_19587);
nor UO_10 (O_10,N_19775,N_19841);
and UO_11 (O_11,N_19933,N_19281);
nor UO_12 (O_12,N_19792,N_19258);
nor UO_13 (O_13,N_19441,N_19635);
nor UO_14 (O_14,N_19808,N_19907);
nand UO_15 (O_15,N_19538,N_19362);
or UO_16 (O_16,N_19694,N_19813);
or UO_17 (O_17,N_19610,N_19577);
and UO_18 (O_18,N_19615,N_19274);
nor UO_19 (O_19,N_19499,N_19413);
xor UO_20 (O_20,N_19454,N_19971);
nand UO_21 (O_21,N_19493,N_19925);
nand UO_22 (O_22,N_19367,N_19226);
nor UO_23 (O_23,N_19541,N_19859);
nor UO_24 (O_24,N_19679,N_19714);
xor UO_25 (O_25,N_19581,N_19784);
nor UO_26 (O_26,N_19981,N_19748);
or UO_27 (O_27,N_19650,N_19715);
nand UO_28 (O_28,N_19705,N_19811);
and UO_29 (O_29,N_19488,N_19872);
nand UO_30 (O_30,N_19564,N_19254);
nor UO_31 (O_31,N_19291,N_19580);
xor UO_32 (O_32,N_19838,N_19217);
and UO_33 (O_33,N_19869,N_19334);
and UO_34 (O_34,N_19793,N_19930);
xor UO_35 (O_35,N_19985,N_19647);
nand UO_36 (O_36,N_19415,N_19721);
nor UO_37 (O_37,N_19213,N_19206);
or UO_38 (O_38,N_19251,N_19982);
or UO_39 (O_39,N_19884,N_19236);
xor UO_40 (O_40,N_19261,N_19826);
and UO_41 (O_41,N_19658,N_19565);
and UO_42 (O_42,N_19398,N_19309);
and UO_43 (O_43,N_19754,N_19680);
nor UO_44 (O_44,N_19944,N_19916);
or UO_45 (O_45,N_19856,N_19455);
xor UO_46 (O_46,N_19932,N_19588);
nor UO_47 (O_47,N_19876,N_19910);
or UO_48 (O_48,N_19660,N_19232);
xnor UO_49 (O_49,N_19388,N_19282);
and UO_50 (O_50,N_19257,N_19697);
and UO_51 (O_51,N_19358,N_19598);
or UO_52 (O_52,N_19529,N_19516);
and UO_53 (O_53,N_19256,N_19247);
xnor UO_54 (O_54,N_19221,N_19585);
and UO_55 (O_55,N_19459,N_19484);
and UO_56 (O_56,N_19339,N_19605);
or UO_57 (O_57,N_19702,N_19699);
nand UO_58 (O_58,N_19417,N_19552);
xnor UO_59 (O_59,N_19794,N_19314);
and UO_60 (O_60,N_19323,N_19534);
xor UO_61 (O_61,N_19750,N_19922);
and UO_62 (O_62,N_19940,N_19501);
or UO_63 (O_63,N_19224,N_19374);
nor UO_64 (O_64,N_19480,N_19543);
xor UO_65 (O_65,N_19200,N_19207);
nor UO_66 (O_66,N_19453,N_19521);
nor UO_67 (O_67,N_19861,N_19407);
nand UO_68 (O_68,N_19809,N_19810);
nor UO_69 (O_69,N_19812,N_19974);
or UO_70 (O_70,N_19498,N_19465);
nor UO_71 (O_71,N_19406,N_19209);
and UO_72 (O_72,N_19576,N_19346);
or UO_73 (O_73,N_19700,N_19980);
or UO_74 (O_74,N_19762,N_19586);
xor UO_75 (O_75,N_19503,N_19344);
or UO_76 (O_76,N_19905,N_19550);
nand UO_77 (O_77,N_19471,N_19849);
or UO_78 (O_78,N_19890,N_19763);
xor UO_79 (O_79,N_19487,N_19751);
xor UO_80 (O_80,N_19929,N_19693);
xnor UO_81 (O_81,N_19947,N_19926);
xnor UO_82 (O_82,N_19644,N_19682);
and UO_83 (O_83,N_19882,N_19765);
nor UO_84 (O_84,N_19228,N_19973);
nor UO_85 (O_85,N_19871,N_19776);
and UO_86 (O_86,N_19442,N_19215);
xor UO_87 (O_87,N_19683,N_19507);
nor UO_88 (O_88,N_19900,N_19593);
nor UO_89 (O_89,N_19955,N_19411);
or UO_90 (O_90,N_19796,N_19698);
nor UO_91 (O_91,N_19246,N_19681);
nand UO_92 (O_92,N_19512,N_19475);
nand UO_93 (O_93,N_19558,N_19865);
nand UO_94 (O_94,N_19238,N_19584);
and UO_95 (O_95,N_19338,N_19653);
nand UO_96 (O_96,N_19440,N_19991);
or UO_97 (O_97,N_19616,N_19275);
nand UO_98 (O_98,N_19877,N_19898);
nor UO_99 (O_99,N_19662,N_19460);
and UO_100 (O_100,N_19383,N_19335);
nor UO_101 (O_101,N_19695,N_19536);
nand UO_102 (O_102,N_19726,N_19544);
xor UO_103 (O_103,N_19677,N_19868);
and UO_104 (O_104,N_19302,N_19242);
nor UO_105 (O_105,N_19360,N_19920);
or UO_106 (O_106,N_19408,N_19836);
nand UO_107 (O_107,N_19456,N_19555);
xnor UO_108 (O_108,N_19825,N_19663);
xnor UO_109 (O_109,N_19761,N_19957);
or UO_110 (O_110,N_19404,N_19208);
nor UO_111 (O_111,N_19785,N_19773);
or UO_112 (O_112,N_19477,N_19692);
nor UO_113 (O_113,N_19359,N_19746);
xnor UO_114 (O_114,N_19831,N_19289);
xor UO_115 (O_115,N_19504,N_19918);
nand UO_116 (O_116,N_19457,N_19600);
or UO_117 (O_117,N_19685,N_19546);
or UO_118 (O_118,N_19523,N_19225);
or UO_119 (O_119,N_19294,N_19393);
nor UO_120 (O_120,N_19379,N_19963);
or UO_121 (O_121,N_19288,N_19655);
nor UO_122 (O_122,N_19840,N_19476);
xor UO_123 (O_123,N_19626,N_19672);
nor UO_124 (O_124,N_19828,N_19913);
and UO_125 (O_125,N_19848,N_19864);
xor UO_126 (O_126,N_19566,N_19827);
nor UO_127 (O_127,N_19621,N_19964);
nand UO_128 (O_128,N_19999,N_19327);
and UO_129 (O_129,N_19667,N_19328);
or UO_130 (O_130,N_19976,N_19752);
nand UO_131 (O_131,N_19496,N_19560);
and UO_132 (O_132,N_19899,N_19945);
nand UO_133 (O_133,N_19965,N_19342);
and UO_134 (O_134,N_19337,N_19203);
or UO_135 (O_135,N_19351,N_19462);
nor UO_136 (O_136,N_19422,N_19515);
nand UO_137 (O_137,N_19903,N_19285);
or UO_138 (O_138,N_19265,N_19956);
or UO_139 (O_139,N_19759,N_19734);
and UO_140 (O_140,N_19350,N_19755);
xnor UO_141 (O_141,N_19343,N_19718);
nand UO_142 (O_142,N_19286,N_19998);
nand UO_143 (O_143,N_19330,N_19527);
nor UO_144 (O_144,N_19347,N_19366);
or UO_145 (O_145,N_19969,N_19632);
nor UO_146 (O_146,N_19535,N_19572);
xnor UO_147 (O_147,N_19629,N_19329);
or UO_148 (O_148,N_19696,N_19263);
xor UO_149 (O_149,N_19799,N_19262);
nor UO_150 (O_150,N_19354,N_19514);
and UO_151 (O_151,N_19893,N_19452);
nand UO_152 (O_152,N_19519,N_19928);
or UO_153 (O_153,N_19279,N_19817);
nor UO_154 (O_154,N_19858,N_19887);
nand UO_155 (O_155,N_19387,N_19528);
nor UO_156 (O_156,N_19670,N_19997);
xnor UO_157 (O_157,N_19252,N_19896);
nand UO_158 (O_158,N_19741,N_19518);
nand UO_159 (O_159,N_19579,N_19297);
xor UO_160 (O_160,N_19287,N_19402);
nor UO_161 (O_161,N_19448,N_19352);
nor UO_162 (O_162,N_19391,N_19537);
xnor UO_163 (O_163,N_19949,N_19269);
xor UO_164 (O_164,N_19961,N_19481);
nor UO_165 (O_165,N_19300,N_19911);
nor UO_166 (O_166,N_19711,N_19375);
nand UO_167 (O_167,N_19712,N_19774);
or UO_168 (O_168,N_19397,N_19268);
or UO_169 (O_169,N_19492,N_19474);
xor UO_170 (O_170,N_19870,N_19533);
nand UO_171 (O_171,N_19385,N_19637);
nand UO_172 (O_172,N_19325,N_19332);
xor UO_173 (O_173,N_19218,N_19539);
and UO_174 (O_174,N_19790,N_19888);
or UO_175 (O_175,N_19993,N_19205);
and UO_176 (O_176,N_19201,N_19639);
nor UO_177 (O_177,N_19839,N_19701);
nand UO_178 (O_178,N_19760,N_19979);
nor UO_179 (O_179,N_19418,N_19376);
nand UO_180 (O_180,N_19311,N_19780);
xor UO_181 (O_181,N_19709,N_19889);
nor UO_182 (O_182,N_19227,N_19390);
nor UO_183 (O_183,N_19722,N_19652);
nand UO_184 (O_184,N_19449,N_19638);
and UO_185 (O_185,N_19284,N_19816);
xnor UO_186 (O_186,N_19972,N_19823);
or UO_187 (O_187,N_19571,N_19267);
nor UO_188 (O_188,N_19704,N_19767);
nor UO_189 (O_189,N_19283,N_19509);
or UO_190 (O_190,N_19483,N_19549);
or UO_191 (O_191,N_19249,N_19312);
and UO_192 (O_192,N_19691,N_19992);
nor UO_193 (O_193,N_19725,N_19219);
nand UO_194 (O_194,N_19835,N_19657);
xnor UO_195 (O_195,N_19707,N_19430);
and UO_196 (O_196,N_19664,N_19468);
or UO_197 (O_197,N_19622,N_19253);
nor UO_198 (O_198,N_19659,N_19747);
nand UO_199 (O_199,N_19603,N_19738);
and UO_200 (O_200,N_19936,N_19782);
nor UO_201 (O_201,N_19943,N_19744);
and UO_202 (O_202,N_19340,N_19906);
nand UO_203 (O_203,N_19651,N_19486);
and UO_204 (O_204,N_19815,N_19317);
and UO_205 (O_205,N_19666,N_19821);
nor UO_206 (O_206,N_19420,N_19333);
xnor UO_207 (O_207,N_19984,N_19954);
nand UO_208 (O_208,N_19909,N_19661);
and UO_209 (O_209,N_19290,N_19270);
xnor UO_210 (O_210,N_19434,N_19800);
and UO_211 (O_211,N_19608,N_19927);
xnor UO_212 (O_212,N_19319,N_19834);
and UO_213 (O_213,N_19688,N_19307);
and UO_214 (O_214,N_19904,N_19803);
xnor UO_215 (O_215,N_19931,N_19886);
nor UO_216 (O_216,N_19400,N_19820);
nand UO_217 (O_217,N_19551,N_19613);
or UO_218 (O_218,N_19386,N_19582);
nor UO_219 (O_219,N_19950,N_19273);
and UO_220 (O_220,N_19723,N_19464);
nand UO_221 (O_221,N_19645,N_19941);
xor UO_222 (O_222,N_19497,N_19601);
or UO_223 (O_223,N_19892,N_19237);
and UO_224 (O_224,N_19562,N_19673);
nand UO_225 (O_225,N_19495,N_19717);
nand UO_226 (O_226,N_19532,N_19426);
xnor UO_227 (O_227,N_19654,N_19299);
nand UO_228 (O_228,N_19489,N_19743);
nand UO_229 (O_229,N_19783,N_19570);
or UO_230 (O_230,N_19505,N_19953);
or UO_231 (O_231,N_19990,N_19806);
or UO_232 (O_232,N_19547,N_19389);
or UO_233 (O_233,N_19364,N_19623);
and UO_234 (O_234,N_19278,N_19409);
and UO_235 (O_235,N_19919,N_19636);
xnor UO_236 (O_236,N_19749,N_19575);
and UO_237 (O_237,N_19791,N_19234);
nor UO_238 (O_238,N_19727,N_19624);
and UO_239 (O_239,N_19240,N_19435);
and UO_240 (O_240,N_19914,N_19689);
nor UO_241 (O_241,N_19363,N_19322);
nand UO_242 (O_242,N_19960,N_19958);
xnor UO_243 (O_243,N_19934,N_19445);
xnor UO_244 (O_244,N_19573,N_19517);
nor UO_245 (O_245,N_19438,N_19804);
xnor UO_246 (O_246,N_19676,N_19733);
or UO_247 (O_247,N_19399,N_19378);
xnor UO_248 (O_248,N_19447,N_19852);
xor UO_249 (O_249,N_19729,N_19470);
or UO_250 (O_250,N_19482,N_19298);
xnor UO_251 (O_251,N_19766,N_19614);
nor UO_252 (O_252,N_19365,N_19305);
nand UO_253 (O_253,N_19271,N_19873);
nand UO_254 (O_254,N_19371,N_19951);
xor UO_255 (O_255,N_19781,N_19502);
or UO_256 (O_256,N_19917,N_19844);
nand UO_257 (O_257,N_19490,N_19370);
and UO_258 (O_258,N_19557,N_19837);
and UO_259 (O_259,N_19611,N_19842);
nor UO_260 (O_260,N_19461,N_19915);
or UO_261 (O_261,N_19901,N_19874);
xnor UO_262 (O_262,N_19912,N_19530);
nand UO_263 (O_263,N_19772,N_19604);
or UO_264 (O_264,N_19966,N_19211);
nor UO_265 (O_265,N_19935,N_19416);
xnor UO_266 (O_266,N_19862,N_19214);
nand UO_267 (O_267,N_19769,N_19789);
nor UO_268 (O_268,N_19778,N_19602);
or UO_269 (O_269,N_19845,N_19757);
and UO_270 (O_270,N_19567,N_19382);
xor UO_271 (O_271,N_19553,N_19627);
or UO_272 (O_272,N_19433,N_19634);
xor UO_273 (O_273,N_19710,N_19703);
nor UO_274 (O_274,N_19620,N_19318);
xnor UO_275 (O_275,N_19293,N_19807);
xnor UO_276 (O_276,N_19561,N_19414);
nand UO_277 (O_277,N_19938,N_19277);
xnor UO_278 (O_278,N_19822,N_19353);
and UO_279 (O_279,N_19625,N_19427);
and UO_280 (O_280,N_19511,N_19948);
nor UO_281 (O_281,N_19924,N_19316);
or UO_282 (O_282,N_19545,N_19403);
xor UO_283 (O_283,N_19805,N_19472);
and UO_284 (O_284,N_19569,N_19216);
or UO_285 (O_285,N_19473,N_19758);
nor UO_286 (O_286,N_19356,N_19212);
nand UO_287 (O_287,N_19591,N_19987);
and UO_288 (O_288,N_19939,N_19690);
nand UO_289 (O_289,N_19589,N_19590);
and UO_290 (O_290,N_19745,N_19578);
nor UO_291 (O_291,N_19878,N_19768);
nand UO_292 (O_292,N_19599,N_19424);
nand UO_293 (O_293,N_19233,N_19315);
nor UO_294 (O_294,N_19897,N_19731);
nand UO_295 (O_295,N_19770,N_19324);
nand UO_296 (O_296,N_19313,N_19419);
nand UO_297 (O_297,N_19372,N_19349);
and UO_298 (O_298,N_19260,N_19675);
nand UO_299 (O_299,N_19786,N_19824);
nor UO_300 (O_300,N_19439,N_19618);
xnor UO_301 (O_301,N_19272,N_19429);
or UO_302 (O_302,N_19526,N_19788);
or UO_303 (O_303,N_19735,N_19875);
and UO_304 (O_304,N_19850,N_19879);
and UO_305 (O_305,N_19345,N_19431);
nor UO_306 (O_306,N_19357,N_19630);
nor UO_307 (O_307,N_19479,N_19742);
nand UO_308 (O_308,N_19619,N_19996);
nand UO_309 (O_309,N_19500,N_19423);
nor UO_310 (O_310,N_19866,N_19377);
or UO_311 (O_311,N_19708,N_19853);
xnor UO_312 (O_312,N_19308,N_19656);
xnor UO_313 (O_313,N_19437,N_19520);
nand UO_314 (O_314,N_19478,N_19983);
nand UO_315 (O_315,N_19494,N_19245);
xnor UO_316 (O_316,N_19970,N_19306);
and UO_317 (O_317,N_19597,N_19994);
and UO_318 (O_318,N_19563,N_19394);
or UO_319 (O_319,N_19777,N_19202);
nand UO_320 (O_320,N_19881,N_19860);
and UO_321 (O_321,N_19451,N_19458);
nor UO_322 (O_322,N_19857,N_19463);
nand UO_323 (O_323,N_19851,N_19425);
and UO_324 (O_324,N_19466,N_19355);
xor UO_325 (O_325,N_19846,N_19908);
nor UO_326 (O_326,N_19421,N_19978);
nand UO_327 (O_327,N_19412,N_19814);
or UO_328 (O_328,N_19368,N_19432);
nor UO_329 (O_329,N_19331,N_19508);
or UO_330 (O_330,N_19229,N_19855);
xor UO_331 (O_331,N_19450,N_19867);
nor UO_332 (O_332,N_19280,N_19401);
xor UO_333 (O_333,N_19802,N_19326);
nor UO_334 (O_334,N_19556,N_19833);
or UO_335 (O_335,N_19923,N_19829);
nand UO_336 (O_336,N_19230,N_19392);
or UO_337 (O_337,N_19583,N_19303);
nand UO_338 (O_338,N_19231,N_19310);
nand UO_339 (O_339,N_19797,N_19885);
and UO_340 (O_340,N_19843,N_19381);
or UO_341 (O_341,N_19467,N_19609);
xnor UO_342 (O_342,N_19671,N_19292);
and UO_343 (O_343,N_19266,N_19491);
xor UO_344 (O_344,N_19646,N_19642);
or UO_345 (O_345,N_19739,N_19204);
and UO_346 (O_346,N_19730,N_19818);
and UO_347 (O_347,N_19832,N_19895);
nand UO_348 (O_348,N_19264,N_19525);
nand UO_349 (O_349,N_19801,N_19369);
nand UO_350 (O_350,N_19248,N_19687);
nor UO_351 (O_351,N_19276,N_19643);
or UO_352 (O_352,N_19295,N_19606);
xor UO_353 (O_353,N_19863,N_19720);
xnor UO_354 (O_354,N_19380,N_19740);
nor UO_355 (O_355,N_19395,N_19724);
nor UO_356 (O_356,N_19522,N_19223);
and UO_357 (O_357,N_19594,N_19942);
and UO_358 (O_358,N_19446,N_19716);
nand UO_359 (O_359,N_19959,N_19531);
or UO_360 (O_360,N_19250,N_19485);
nand UO_361 (O_361,N_19779,N_19296);
or UO_362 (O_362,N_19678,N_19548);
and UO_363 (O_363,N_19736,N_19612);
nand UO_364 (O_364,N_19921,N_19830);
nand UO_365 (O_365,N_19592,N_19719);
nor UO_366 (O_366,N_19244,N_19559);
nand UO_367 (O_367,N_19649,N_19902);
nand UO_368 (O_368,N_19222,N_19513);
xnor UO_369 (O_369,N_19946,N_19361);
nand UO_370 (O_370,N_19880,N_19210);
or UO_371 (O_371,N_19568,N_19259);
nand UO_372 (O_372,N_19542,N_19405);
xor UO_373 (O_373,N_19320,N_19674);
nor UO_374 (O_374,N_19986,N_19713);
and UO_375 (O_375,N_19384,N_19510);
nor UO_376 (O_376,N_19753,N_19574);
nand UO_377 (O_377,N_19396,N_19469);
nand UO_378 (O_378,N_19631,N_19795);
nor UO_379 (O_379,N_19506,N_19977);
and UO_380 (O_380,N_19373,N_19410);
xor UO_381 (O_381,N_19596,N_19595);
and UO_382 (O_382,N_19891,N_19686);
xnor UO_383 (O_383,N_19854,N_19952);
or UO_384 (O_384,N_19617,N_19706);
xnor UO_385 (O_385,N_19443,N_19989);
xor UO_386 (O_386,N_19444,N_19336);
nand UO_387 (O_387,N_19732,N_19348);
nor UO_388 (O_388,N_19798,N_19554);
xor UO_389 (O_389,N_19301,N_19756);
and UO_390 (O_390,N_19728,N_19684);
or UO_391 (O_391,N_19665,N_19633);
nor UO_392 (O_392,N_19737,N_19220);
nand UO_393 (O_393,N_19255,N_19243);
nand UO_394 (O_394,N_19968,N_19975);
nor UO_395 (O_395,N_19540,N_19894);
and UO_396 (O_396,N_19962,N_19524);
and UO_397 (O_397,N_19321,N_19787);
nor UO_398 (O_398,N_19669,N_19883);
or UO_399 (O_399,N_19847,N_19640);
and UO_400 (O_400,N_19307,N_19392);
and UO_401 (O_401,N_19408,N_19844);
nand UO_402 (O_402,N_19328,N_19821);
xor UO_403 (O_403,N_19319,N_19798);
or UO_404 (O_404,N_19843,N_19315);
nor UO_405 (O_405,N_19756,N_19331);
xor UO_406 (O_406,N_19267,N_19642);
nor UO_407 (O_407,N_19843,N_19688);
or UO_408 (O_408,N_19268,N_19920);
xnor UO_409 (O_409,N_19917,N_19871);
and UO_410 (O_410,N_19278,N_19951);
and UO_411 (O_411,N_19765,N_19351);
nand UO_412 (O_412,N_19465,N_19240);
nand UO_413 (O_413,N_19948,N_19504);
and UO_414 (O_414,N_19585,N_19616);
nand UO_415 (O_415,N_19889,N_19657);
nor UO_416 (O_416,N_19397,N_19311);
nor UO_417 (O_417,N_19758,N_19911);
or UO_418 (O_418,N_19217,N_19402);
xor UO_419 (O_419,N_19656,N_19575);
xnor UO_420 (O_420,N_19267,N_19406);
xor UO_421 (O_421,N_19216,N_19765);
and UO_422 (O_422,N_19570,N_19491);
or UO_423 (O_423,N_19290,N_19911);
nor UO_424 (O_424,N_19917,N_19534);
xnor UO_425 (O_425,N_19774,N_19234);
and UO_426 (O_426,N_19503,N_19316);
and UO_427 (O_427,N_19571,N_19393);
xnor UO_428 (O_428,N_19686,N_19317);
xor UO_429 (O_429,N_19854,N_19201);
nor UO_430 (O_430,N_19281,N_19229);
xnor UO_431 (O_431,N_19740,N_19700);
nand UO_432 (O_432,N_19733,N_19544);
xor UO_433 (O_433,N_19434,N_19997);
nor UO_434 (O_434,N_19833,N_19430);
xor UO_435 (O_435,N_19715,N_19976);
or UO_436 (O_436,N_19971,N_19710);
xnor UO_437 (O_437,N_19578,N_19738);
nand UO_438 (O_438,N_19271,N_19823);
nor UO_439 (O_439,N_19806,N_19208);
nand UO_440 (O_440,N_19625,N_19240);
xnor UO_441 (O_441,N_19887,N_19245);
nand UO_442 (O_442,N_19743,N_19371);
nor UO_443 (O_443,N_19942,N_19424);
xor UO_444 (O_444,N_19732,N_19499);
xnor UO_445 (O_445,N_19955,N_19357);
and UO_446 (O_446,N_19579,N_19657);
nor UO_447 (O_447,N_19473,N_19666);
nand UO_448 (O_448,N_19878,N_19518);
xnor UO_449 (O_449,N_19415,N_19955);
or UO_450 (O_450,N_19696,N_19269);
xnor UO_451 (O_451,N_19385,N_19491);
xor UO_452 (O_452,N_19879,N_19784);
nand UO_453 (O_453,N_19909,N_19626);
and UO_454 (O_454,N_19814,N_19912);
nor UO_455 (O_455,N_19684,N_19323);
nand UO_456 (O_456,N_19374,N_19803);
nor UO_457 (O_457,N_19405,N_19985);
nand UO_458 (O_458,N_19791,N_19937);
nand UO_459 (O_459,N_19807,N_19619);
nor UO_460 (O_460,N_19552,N_19659);
nand UO_461 (O_461,N_19503,N_19569);
or UO_462 (O_462,N_19385,N_19971);
nand UO_463 (O_463,N_19638,N_19636);
xnor UO_464 (O_464,N_19819,N_19488);
xor UO_465 (O_465,N_19442,N_19596);
nand UO_466 (O_466,N_19471,N_19415);
nand UO_467 (O_467,N_19624,N_19594);
xor UO_468 (O_468,N_19298,N_19729);
nor UO_469 (O_469,N_19903,N_19839);
and UO_470 (O_470,N_19967,N_19817);
nor UO_471 (O_471,N_19912,N_19612);
nor UO_472 (O_472,N_19500,N_19386);
xnor UO_473 (O_473,N_19297,N_19260);
or UO_474 (O_474,N_19217,N_19532);
nor UO_475 (O_475,N_19762,N_19675);
or UO_476 (O_476,N_19235,N_19509);
xnor UO_477 (O_477,N_19694,N_19651);
nand UO_478 (O_478,N_19379,N_19259);
and UO_479 (O_479,N_19365,N_19902);
xor UO_480 (O_480,N_19711,N_19575);
xor UO_481 (O_481,N_19312,N_19686);
xor UO_482 (O_482,N_19658,N_19477);
nor UO_483 (O_483,N_19534,N_19696);
or UO_484 (O_484,N_19722,N_19379);
xnor UO_485 (O_485,N_19562,N_19496);
or UO_486 (O_486,N_19636,N_19216);
and UO_487 (O_487,N_19555,N_19349);
nand UO_488 (O_488,N_19420,N_19845);
and UO_489 (O_489,N_19389,N_19414);
and UO_490 (O_490,N_19464,N_19741);
or UO_491 (O_491,N_19481,N_19877);
nand UO_492 (O_492,N_19579,N_19727);
nand UO_493 (O_493,N_19878,N_19497);
nor UO_494 (O_494,N_19813,N_19844);
nand UO_495 (O_495,N_19559,N_19491);
nand UO_496 (O_496,N_19822,N_19676);
nor UO_497 (O_497,N_19329,N_19866);
or UO_498 (O_498,N_19919,N_19961);
xor UO_499 (O_499,N_19222,N_19655);
nand UO_500 (O_500,N_19519,N_19797);
nor UO_501 (O_501,N_19480,N_19697);
nor UO_502 (O_502,N_19257,N_19860);
and UO_503 (O_503,N_19540,N_19906);
nor UO_504 (O_504,N_19657,N_19312);
or UO_505 (O_505,N_19504,N_19697);
nand UO_506 (O_506,N_19636,N_19364);
or UO_507 (O_507,N_19929,N_19205);
or UO_508 (O_508,N_19744,N_19307);
nor UO_509 (O_509,N_19277,N_19857);
nor UO_510 (O_510,N_19705,N_19561);
nand UO_511 (O_511,N_19703,N_19322);
nor UO_512 (O_512,N_19558,N_19478);
nand UO_513 (O_513,N_19846,N_19433);
nor UO_514 (O_514,N_19443,N_19851);
nor UO_515 (O_515,N_19388,N_19687);
xor UO_516 (O_516,N_19678,N_19991);
and UO_517 (O_517,N_19405,N_19554);
nor UO_518 (O_518,N_19448,N_19227);
nor UO_519 (O_519,N_19915,N_19716);
and UO_520 (O_520,N_19433,N_19866);
or UO_521 (O_521,N_19637,N_19827);
or UO_522 (O_522,N_19582,N_19803);
or UO_523 (O_523,N_19986,N_19202);
or UO_524 (O_524,N_19601,N_19757);
and UO_525 (O_525,N_19685,N_19422);
nand UO_526 (O_526,N_19377,N_19673);
and UO_527 (O_527,N_19496,N_19737);
nand UO_528 (O_528,N_19591,N_19429);
and UO_529 (O_529,N_19268,N_19759);
xnor UO_530 (O_530,N_19735,N_19407);
xor UO_531 (O_531,N_19948,N_19796);
nand UO_532 (O_532,N_19928,N_19415);
and UO_533 (O_533,N_19417,N_19805);
or UO_534 (O_534,N_19846,N_19563);
xnor UO_535 (O_535,N_19540,N_19833);
or UO_536 (O_536,N_19945,N_19515);
and UO_537 (O_537,N_19297,N_19721);
or UO_538 (O_538,N_19782,N_19788);
or UO_539 (O_539,N_19472,N_19528);
or UO_540 (O_540,N_19840,N_19838);
xnor UO_541 (O_541,N_19969,N_19679);
xor UO_542 (O_542,N_19824,N_19455);
and UO_543 (O_543,N_19874,N_19413);
nand UO_544 (O_544,N_19411,N_19422);
and UO_545 (O_545,N_19813,N_19743);
xor UO_546 (O_546,N_19228,N_19564);
nand UO_547 (O_547,N_19348,N_19381);
xnor UO_548 (O_548,N_19236,N_19770);
xnor UO_549 (O_549,N_19288,N_19686);
or UO_550 (O_550,N_19969,N_19628);
nor UO_551 (O_551,N_19905,N_19504);
xnor UO_552 (O_552,N_19384,N_19363);
nor UO_553 (O_553,N_19839,N_19228);
or UO_554 (O_554,N_19810,N_19892);
and UO_555 (O_555,N_19356,N_19501);
nor UO_556 (O_556,N_19332,N_19931);
xnor UO_557 (O_557,N_19336,N_19260);
and UO_558 (O_558,N_19857,N_19488);
and UO_559 (O_559,N_19867,N_19446);
and UO_560 (O_560,N_19771,N_19204);
and UO_561 (O_561,N_19894,N_19587);
nor UO_562 (O_562,N_19924,N_19766);
nand UO_563 (O_563,N_19765,N_19362);
xnor UO_564 (O_564,N_19878,N_19640);
or UO_565 (O_565,N_19401,N_19568);
nor UO_566 (O_566,N_19552,N_19614);
and UO_567 (O_567,N_19207,N_19694);
nand UO_568 (O_568,N_19725,N_19323);
xor UO_569 (O_569,N_19850,N_19508);
nand UO_570 (O_570,N_19851,N_19721);
or UO_571 (O_571,N_19958,N_19347);
nor UO_572 (O_572,N_19226,N_19236);
or UO_573 (O_573,N_19578,N_19939);
and UO_574 (O_574,N_19684,N_19992);
xor UO_575 (O_575,N_19759,N_19639);
xor UO_576 (O_576,N_19833,N_19622);
nor UO_577 (O_577,N_19594,N_19665);
and UO_578 (O_578,N_19992,N_19440);
nor UO_579 (O_579,N_19396,N_19549);
nor UO_580 (O_580,N_19902,N_19890);
nor UO_581 (O_581,N_19671,N_19622);
xnor UO_582 (O_582,N_19906,N_19207);
xor UO_583 (O_583,N_19443,N_19266);
nand UO_584 (O_584,N_19572,N_19208);
xnor UO_585 (O_585,N_19803,N_19822);
nand UO_586 (O_586,N_19837,N_19820);
xnor UO_587 (O_587,N_19919,N_19539);
xor UO_588 (O_588,N_19357,N_19806);
xnor UO_589 (O_589,N_19846,N_19477);
xor UO_590 (O_590,N_19252,N_19934);
and UO_591 (O_591,N_19506,N_19429);
or UO_592 (O_592,N_19521,N_19205);
nor UO_593 (O_593,N_19454,N_19344);
nand UO_594 (O_594,N_19467,N_19855);
xnor UO_595 (O_595,N_19835,N_19418);
nor UO_596 (O_596,N_19250,N_19204);
xnor UO_597 (O_597,N_19372,N_19524);
xor UO_598 (O_598,N_19626,N_19356);
or UO_599 (O_599,N_19604,N_19979);
and UO_600 (O_600,N_19929,N_19656);
or UO_601 (O_601,N_19801,N_19804);
nor UO_602 (O_602,N_19224,N_19244);
nor UO_603 (O_603,N_19648,N_19716);
or UO_604 (O_604,N_19523,N_19352);
nor UO_605 (O_605,N_19264,N_19574);
and UO_606 (O_606,N_19488,N_19503);
xnor UO_607 (O_607,N_19936,N_19752);
or UO_608 (O_608,N_19938,N_19726);
or UO_609 (O_609,N_19769,N_19341);
or UO_610 (O_610,N_19871,N_19310);
xnor UO_611 (O_611,N_19980,N_19329);
nor UO_612 (O_612,N_19491,N_19249);
and UO_613 (O_613,N_19404,N_19291);
nand UO_614 (O_614,N_19276,N_19445);
nand UO_615 (O_615,N_19950,N_19234);
nor UO_616 (O_616,N_19456,N_19233);
nor UO_617 (O_617,N_19743,N_19384);
and UO_618 (O_618,N_19913,N_19347);
nor UO_619 (O_619,N_19836,N_19845);
nor UO_620 (O_620,N_19589,N_19271);
nor UO_621 (O_621,N_19780,N_19802);
or UO_622 (O_622,N_19424,N_19416);
nor UO_623 (O_623,N_19883,N_19902);
and UO_624 (O_624,N_19614,N_19206);
and UO_625 (O_625,N_19814,N_19255);
xnor UO_626 (O_626,N_19823,N_19718);
or UO_627 (O_627,N_19610,N_19284);
and UO_628 (O_628,N_19880,N_19738);
nand UO_629 (O_629,N_19249,N_19914);
xnor UO_630 (O_630,N_19383,N_19656);
nor UO_631 (O_631,N_19803,N_19753);
nand UO_632 (O_632,N_19671,N_19326);
and UO_633 (O_633,N_19928,N_19317);
nor UO_634 (O_634,N_19373,N_19301);
nand UO_635 (O_635,N_19417,N_19462);
nand UO_636 (O_636,N_19961,N_19405);
nand UO_637 (O_637,N_19802,N_19303);
xor UO_638 (O_638,N_19712,N_19796);
or UO_639 (O_639,N_19867,N_19842);
xor UO_640 (O_640,N_19300,N_19858);
nand UO_641 (O_641,N_19713,N_19374);
xor UO_642 (O_642,N_19443,N_19601);
xnor UO_643 (O_643,N_19288,N_19587);
and UO_644 (O_644,N_19858,N_19658);
or UO_645 (O_645,N_19677,N_19795);
nor UO_646 (O_646,N_19877,N_19807);
nand UO_647 (O_647,N_19421,N_19356);
and UO_648 (O_648,N_19429,N_19659);
and UO_649 (O_649,N_19525,N_19763);
nor UO_650 (O_650,N_19684,N_19581);
nand UO_651 (O_651,N_19525,N_19777);
nor UO_652 (O_652,N_19830,N_19452);
nand UO_653 (O_653,N_19323,N_19257);
nor UO_654 (O_654,N_19311,N_19242);
nor UO_655 (O_655,N_19677,N_19444);
or UO_656 (O_656,N_19788,N_19501);
nand UO_657 (O_657,N_19321,N_19207);
or UO_658 (O_658,N_19908,N_19843);
and UO_659 (O_659,N_19584,N_19803);
nor UO_660 (O_660,N_19724,N_19833);
nand UO_661 (O_661,N_19813,N_19988);
nor UO_662 (O_662,N_19932,N_19243);
nor UO_663 (O_663,N_19669,N_19708);
nor UO_664 (O_664,N_19360,N_19379);
or UO_665 (O_665,N_19440,N_19428);
or UO_666 (O_666,N_19922,N_19292);
and UO_667 (O_667,N_19876,N_19816);
and UO_668 (O_668,N_19221,N_19880);
xor UO_669 (O_669,N_19387,N_19443);
nand UO_670 (O_670,N_19831,N_19417);
nor UO_671 (O_671,N_19587,N_19869);
xor UO_672 (O_672,N_19292,N_19817);
and UO_673 (O_673,N_19319,N_19607);
nor UO_674 (O_674,N_19332,N_19937);
nand UO_675 (O_675,N_19770,N_19345);
nor UO_676 (O_676,N_19739,N_19994);
xnor UO_677 (O_677,N_19415,N_19868);
nand UO_678 (O_678,N_19474,N_19946);
or UO_679 (O_679,N_19229,N_19402);
xnor UO_680 (O_680,N_19710,N_19841);
xnor UO_681 (O_681,N_19729,N_19366);
nor UO_682 (O_682,N_19985,N_19538);
xnor UO_683 (O_683,N_19294,N_19439);
or UO_684 (O_684,N_19716,N_19240);
xnor UO_685 (O_685,N_19800,N_19455);
nor UO_686 (O_686,N_19560,N_19888);
xnor UO_687 (O_687,N_19528,N_19835);
and UO_688 (O_688,N_19327,N_19716);
xor UO_689 (O_689,N_19785,N_19905);
and UO_690 (O_690,N_19615,N_19239);
or UO_691 (O_691,N_19794,N_19674);
and UO_692 (O_692,N_19938,N_19801);
xor UO_693 (O_693,N_19213,N_19767);
nor UO_694 (O_694,N_19750,N_19574);
and UO_695 (O_695,N_19783,N_19739);
and UO_696 (O_696,N_19457,N_19419);
and UO_697 (O_697,N_19815,N_19646);
nand UO_698 (O_698,N_19259,N_19427);
or UO_699 (O_699,N_19554,N_19631);
xor UO_700 (O_700,N_19988,N_19757);
xnor UO_701 (O_701,N_19807,N_19395);
and UO_702 (O_702,N_19697,N_19329);
and UO_703 (O_703,N_19406,N_19835);
and UO_704 (O_704,N_19640,N_19461);
nand UO_705 (O_705,N_19896,N_19998);
nand UO_706 (O_706,N_19406,N_19716);
xnor UO_707 (O_707,N_19544,N_19215);
and UO_708 (O_708,N_19723,N_19677);
nor UO_709 (O_709,N_19900,N_19508);
nand UO_710 (O_710,N_19909,N_19728);
or UO_711 (O_711,N_19327,N_19707);
or UO_712 (O_712,N_19223,N_19310);
or UO_713 (O_713,N_19409,N_19631);
or UO_714 (O_714,N_19865,N_19621);
nand UO_715 (O_715,N_19794,N_19784);
xor UO_716 (O_716,N_19232,N_19362);
xnor UO_717 (O_717,N_19430,N_19632);
or UO_718 (O_718,N_19903,N_19617);
and UO_719 (O_719,N_19391,N_19281);
nand UO_720 (O_720,N_19704,N_19593);
and UO_721 (O_721,N_19650,N_19877);
nand UO_722 (O_722,N_19462,N_19392);
and UO_723 (O_723,N_19689,N_19775);
nor UO_724 (O_724,N_19459,N_19895);
xnor UO_725 (O_725,N_19774,N_19609);
nor UO_726 (O_726,N_19865,N_19705);
nor UO_727 (O_727,N_19456,N_19759);
nand UO_728 (O_728,N_19256,N_19401);
nand UO_729 (O_729,N_19841,N_19926);
nand UO_730 (O_730,N_19807,N_19850);
or UO_731 (O_731,N_19818,N_19706);
and UO_732 (O_732,N_19691,N_19920);
and UO_733 (O_733,N_19601,N_19227);
and UO_734 (O_734,N_19456,N_19959);
or UO_735 (O_735,N_19346,N_19639);
xnor UO_736 (O_736,N_19275,N_19579);
or UO_737 (O_737,N_19269,N_19522);
and UO_738 (O_738,N_19898,N_19304);
and UO_739 (O_739,N_19710,N_19552);
and UO_740 (O_740,N_19208,N_19810);
nor UO_741 (O_741,N_19822,N_19377);
nor UO_742 (O_742,N_19525,N_19606);
and UO_743 (O_743,N_19350,N_19702);
and UO_744 (O_744,N_19322,N_19596);
nand UO_745 (O_745,N_19706,N_19863);
and UO_746 (O_746,N_19382,N_19359);
or UO_747 (O_747,N_19816,N_19841);
xnor UO_748 (O_748,N_19965,N_19200);
xor UO_749 (O_749,N_19440,N_19354);
nand UO_750 (O_750,N_19776,N_19957);
and UO_751 (O_751,N_19673,N_19320);
and UO_752 (O_752,N_19407,N_19236);
nor UO_753 (O_753,N_19696,N_19865);
or UO_754 (O_754,N_19284,N_19783);
nand UO_755 (O_755,N_19686,N_19784);
or UO_756 (O_756,N_19691,N_19356);
and UO_757 (O_757,N_19980,N_19687);
xnor UO_758 (O_758,N_19785,N_19622);
xor UO_759 (O_759,N_19589,N_19435);
xor UO_760 (O_760,N_19324,N_19539);
xor UO_761 (O_761,N_19515,N_19366);
or UO_762 (O_762,N_19419,N_19870);
and UO_763 (O_763,N_19598,N_19952);
and UO_764 (O_764,N_19754,N_19324);
nor UO_765 (O_765,N_19422,N_19212);
and UO_766 (O_766,N_19958,N_19452);
nand UO_767 (O_767,N_19647,N_19863);
nor UO_768 (O_768,N_19596,N_19320);
and UO_769 (O_769,N_19308,N_19768);
xor UO_770 (O_770,N_19668,N_19844);
xnor UO_771 (O_771,N_19414,N_19870);
xnor UO_772 (O_772,N_19873,N_19585);
and UO_773 (O_773,N_19742,N_19371);
nor UO_774 (O_774,N_19732,N_19419);
nand UO_775 (O_775,N_19797,N_19613);
nor UO_776 (O_776,N_19578,N_19574);
xnor UO_777 (O_777,N_19865,N_19443);
xor UO_778 (O_778,N_19552,N_19778);
nor UO_779 (O_779,N_19314,N_19387);
or UO_780 (O_780,N_19276,N_19498);
xnor UO_781 (O_781,N_19808,N_19621);
xor UO_782 (O_782,N_19695,N_19373);
and UO_783 (O_783,N_19211,N_19714);
nor UO_784 (O_784,N_19929,N_19291);
and UO_785 (O_785,N_19419,N_19775);
or UO_786 (O_786,N_19552,N_19611);
nor UO_787 (O_787,N_19603,N_19721);
nor UO_788 (O_788,N_19491,N_19802);
or UO_789 (O_789,N_19651,N_19577);
nor UO_790 (O_790,N_19464,N_19945);
or UO_791 (O_791,N_19299,N_19426);
nor UO_792 (O_792,N_19584,N_19372);
nand UO_793 (O_793,N_19861,N_19629);
or UO_794 (O_794,N_19883,N_19475);
nand UO_795 (O_795,N_19396,N_19789);
xor UO_796 (O_796,N_19799,N_19319);
xnor UO_797 (O_797,N_19887,N_19410);
and UO_798 (O_798,N_19655,N_19398);
and UO_799 (O_799,N_19294,N_19512);
nor UO_800 (O_800,N_19646,N_19224);
and UO_801 (O_801,N_19882,N_19503);
nand UO_802 (O_802,N_19634,N_19554);
and UO_803 (O_803,N_19433,N_19306);
and UO_804 (O_804,N_19608,N_19288);
and UO_805 (O_805,N_19591,N_19730);
nand UO_806 (O_806,N_19479,N_19873);
nand UO_807 (O_807,N_19372,N_19594);
nor UO_808 (O_808,N_19255,N_19434);
nor UO_809 (O_809,N_19923,N_19722);
or UO_810 (O_810,N_19271,N_19558);
nor UO_811 (O_811,N_19386,N_19295);
nor UO_812 (O_812,N_19481,N_19566);
xnor UO_813 (O_813,N_19688,N_19275);
or UO_814 (O_814,N_19344,N_19306);
nand UO_815 (O_815,N_19701,N_19620);
xnor UO_816 (O_816,N_19992,N_19786);
xor UO_817 (O_817,N_19730,N_19630);
nand UO_818 (O_818,N_19866,N_19683);
xor UO_819 (O_819,N_19680,N_19686);
and UO_820 (O_820,N_19965,N_19806);
nor UO_821 (O_821,N_19321,N_19518);
nor UO_822 (O_822,N_19246,N_19962);
nor UO_823 (O_823,N_19722,N_19497);
or UO_824 (O_824,N_19508,N_19979);
nand UO_825 (O_825,N_19205,N_19862);
and UO_826 (O_826,N_19658,N_19959);
xor UO_827 (O_827,N_19966,N_19281);
and UO_828 (O_828,N_19224,N_19586);
or UO_829 (O_829,N_19809,N_19488);
nor UO_830 (O_830,N_19352,N_19801);
or UO_831 (O_831,N_19755,N_19944);
and UO_832 (O_832,N_19712,N_19651);
nor UO_833 (O_833,N_19678,N_19525);
and UO_834 (O_834,N_19917,N_19449);
and UO_835 (O_835,N_19457,N_19346);
nor UO_836 (O_836,N_19254,N_19655);
xnor UO_837 (O_837,N_19458,N_19991);
nand UO_838 (O_838,N_19560,N_19472);
nand UO_839 (O_839,N_19885,N_19520);
nor UO_840 (O_840,N_19466,N_19928);
xor UO_841 (O_841,N_19726,N_19336);
or UO_842 (O_842,N_19488,N_19485);
nor UO_843 (O_843,N_19991,N_19964);
nand UO_844 (O_844,N_19733,N_19860);
nand UO_845 (O_845,N_19916,N_19504);
nor UO_846 (O_846,N_19212,N_19244);
nand UO_847 (O_847,N_19983,N_19331);
or UO_848 (O_848,N_19895,N_19214);
or UO_849 (O_849,N_19793,N_19618);
nor UO_850 (O_850,N_19765,N_19824);
and UO_851 (O_851,N_19750,N_19916);
nand UO_852 (O_852,N_19867,N_19870);
nor UO_853 (O_853,N_19760,N_19762);
or UO_854 (O_854,N_19357,N_19208);
or UO_855 (O_855,N_19503,N_19528);
nand UO_856 (O_856,N_19974,N_19328);
nand UO_857 (O_857,N_19249,N_19847);
xnor UO_858 (O_858,N_19876,N_19779);
xor UO_859 (O_859,N_19913,N_19720);
or UO_860 (O_860,N_19981,N_19468);
xnor UO_861 (O_861,N_19647,N_19234);
nand UO_862 (O_862,N_19752,N_19209);
xor UO_863 (O_863,N_19517,N_19780);
xnor UO_864 (O_864,N_19460,N_19588);
nor UO_865 (O_865,N_19909,N_19271);
xor UO_866 (O_866,N_19894,N_19882);
xnor UO_867 (O_867,N_19415,N_19730);
nand UO_868 (O_868,N_19910,N_19684);
and UO_869 (O_869,N_19439,N_19772);
or UO_870 (O_870,N_19407,N_19725);
and UO_871 (O_871,N_19615,N_19562);
and UO_872 (O_872,N_19248,N_19843);
nand UO_873 (O_873,N_19589,N_19319);
and UO_874 (O_874,N_19830,N_19728);
nor UO_875 (O_875,N_19554,N_19819);
and UO_876 (O_876,N_19371,N_19972);
and UO_877 (O_877,N_19670,N_19472);
xnor UO_878 (O_878,N_19956,N_19570);
nor UO_879 (O_879,N_19865,N_19953);
and UO_880 (O_880,N_19423,N_19458);
or UO_881 (O_881,N_19428,N_19295);
and UO_882 (O_882,N_19485,N_19962);
xor UO_883 (O_883,N_19794,N_19629);
or UO_884 (O_884,N_19720,N_19252);
xnor UO_885 (O_885,N_19462,N_19468);
nand UO_886 (O_886,N_19737,N_19859);
and UO_887 (O_887,N_19638,N_19352);
and UO_888 (O_888,N_19526,N_19758);
nand UO_889 (O_889,N_19503,N_19435);
and UO_890 (O_890,N_19364,N_19386);
nand UO_891 (O_891,N_19372,N_19741);
nand UO_892 (O_892,N_19507,N_19807);
xnor UO_893 (O_893,N_19574,N_19302);
and UO_894 (O_894,N_19481,N_19597);
xor UO_895 (O_895,N_19401,N_19580);
or UO_896 (O_896,N_19916,N_19662);
nand UO_897 (O_897,N_19575,N_19510);
or UO_898 (O_898,N_19459,N_19769);
nor UO_899 (O_899,N_19768,N_19348);
nand UO_900 (O_900,N_19687,N_19533);
and UO_901 (O_901,N_19560,N_19450);
and UO_902 (O_902,N_19361,N_19821);
nand UO_903 (O_903,N_19571,N_19599);
and UO_904 (O_904,N_19307,N_19797);
nand UO_905 (O_905,N_19871,N_19855);
nor UO_906 (O_906,N_19857,N_19847);
nand UO_907 (O_907,N_19868,N_19758);
and UO_908 (O_908,N_19626,N_19447);
or UO_909 (O_909,N_19352,N_19323);
and UO_910 (O_910,N_19567,N_19328);
or UO_911 (O_911,N_19902,N_19788);
xnor UO_912 (O_912,N_19655,N_19760);
nor UO_913 (O_913,N_19779,N_19881);
nand UO_914 (O_914,N_19929,N_19930);
and UO_915 (O_915,N_19825,N_19674);
nand UO_916 (O_916,N_19977,N_19399);
nand UO_917 (O_917,N_19964,N_19251);
nor UO_918 (O_918,N_19533,N_19726);
nor UO_919 (O_919,N_19681,N_19299);
or UO_920 (O_920,N_19662,N_19239);
and UO_921 (O_921,N_19832,N_19485);
and UO_922 (O_922,N_19245,N_19774);
and UO_923 (O_923,N_19693,N_19689);
nor UO_924 (O_924,N_19294,N_19598);
nand UO_925 (O_925,N_19833,N_19523);
nand UO_926 (O_926,N_19645,N_19581);
or UO_927 (O_927,N_19930,N_19603);
nor UO_928 (O_928,N_19832,N_19624);
and UO_929 (O_929,N_19557,N_19802);
xor UO_930 (O_930,N_19353,N_19964);
nor UO_931 (O_931,N_19305,N_19495);
nand UO_932 (O_932,N_19481,N_19651);
nand UO_933 (O_933,N_19425,N_19775);
nand UO_934 (O_934,N_19712,N_19273);
or UO_935 (O_935,N_19380,N_19838);
xor UO_936 (O_936,N_19210,N_19382);
xnor UO_937 (O_937,N_19725,N_19579);
and UO_938 (O_938,N_19236,N_19548);
nand UO_939 (O_939,N_19867,N_19743);
and UO_940 (O_940,N_19753,N_19590);
xor UO_941 (O_941,N_19771,N_19590);
nor UO_942 (O_942,N_19471,N_19798);
and UO_943 (O_943,N_19473,N_19358);
and UO_944 (O_944,N_19557,N_19567);
and UO_945 (O_945,N_19987,N_19981);
nor UO_946 (O_946,N_19423,N_19900);
nor UO_947 (O_947,N_19690,N_19368);
nor UO_948 (O_948,N_19262,N_19982);
nand UO_949 (O_949,N_19961,N_19450);
and UO_950 (O_950,N_19664,N_19805);
nor UO_951 (O_951,N_19748,N_19760);
nor UO_952 (O_952,N_19724,N_19821);
xnor UO_953 (O_953,N_19336,N_19616);
nor UO_954 (O_954,N_19734,N_19883);
or UO_955 (O_955,N_19799,N_19399);
xnor UO_956 (O_956,N_19492,N_19943);
and UO_957 (O_957,N_19848,N_19215);
and UO_958 (O_958,N_19919,N_19340);
or UO_959 (O_959,N_19668,N_19713);
or UO_960 (O_960,N_19982,N_19402);
and UO_961 (O_961,N_19680,N_19791);
and UO_962 (O_962,N_19454,N_19490);
and UO_963 (O_963,N_19838,N_19741);
nor UO_964 (O_964,N_19828,N_19452);
xor UO_965 (O_965,N_19535,N_19426);
or UO_966 (O_966,N_19963,N_19553);
xnor UO_967 (O_967,N_19254,N_19703);
xor UO_968 (O_968,N_19287,N_19712);
nand UO_969 (O_969,N_19240,N_19393);
or UO_970 (O_970,N_19987,N_19442);
or UO_971 (O_971,N_19423,N_19917);
and UO_972 (O_972,N_19938,N_19803);
nand UO_973 (O_973,N_19946,N_19364);
or UO_974 (O_974,N_19562,N_19683);
xnor UO_975 (O_975,N_19241,N_19265);
or UO_976 (O_976,N_19254,N_19653);
xor UO_977 (O_977,N_19517,N_19774);
and UO_978 (O_978,N_19745,N_19843);
nand UO_979 (O_979,N_19249,N_19423);
nor UO_980 (O_980,N_19855,N_19978);
or UO_981 (O_981,N_19954,N_19958);
or UO_982 (O_982,N_19570,N_19453);
xnor UO_983 (O_983,N_19791,N_19321);
nand UO_984 (O_984,N_19690,N_19869);
nand UO_985 (O_985,N_19928,N_19768);
nand UO_986 (O_986,N_19333,N_19551);
xor UO_987 (O_987,N_19422,N_19772);
xnor UO_988 (O_988,N_19408,N_19957);
and UO_989 (O_989,N_19864,N_19434);
nor UO_990 (O_990,N_19588,N_19207);
nor UO_991 (O_991,N_19228,N_19690);
and UO_992 (O_992,N_19638,N_19904);
or UO_993 (O_993,N_19467,N_19878);
nor UO_994 (O_994,N_19267,N_19348);
nor UO_995 (O_995,N_19203,N_19390);
or UO_996 (O_996,N_19454,N_19711);
nand UO_997 (O_997,N_19228,N_19472);
nand UO_998 (O_998,N_19930,N_19270);
and UO_999 (O_999,N_19326,N_19343);
and UO_1000 (O_1000,N_19985,N_19971);
and UO_1001 (O_1001,N_19597,N_19523);
nand UO_1002 (O_1002,N_19807,N_19433);
nor UO_1003 (O_1003,N_19608,N_19664);
nor UO_1004 (O_1004,N_19649,N_19678);
xor UO_1005 (O_1005,N_19256,N_19304);
or UO_1006 (O_1006,N_19745,N_19446);
or UO_1007 (O_1007,N_19564,N_19587);
nand UO_1008 (O_1008,N_19977,N_19391);
xor UO_1009 (O_1009,N_19410,N_19767);
nor UO_1010 (O_1010,N_19937,N_19233);
nand UO_1011 (O_1011,N_19964,N_19555);
nand UO_1012 (O_1012,N_19839,N_19410);
nand UO_1013 (O_1013,N_19982,N_19766);
and UO_1014 (O_1014,N_19886,N_19618);
xnor UO_1015 (O_1015,N_19965,N_19543);
nand UO_1016 (O_1016,N_19921,N_19726);
xor UO_1017 (O_1017,N_19200,N_19247);
or UO_1018 (O_1018,N_19578,N_19603);
nor UO_1019 (O_1019,N_19687,N_19851);
nand UO_1020 (O_1020,N_19805,N_19554);
nand UO_1021 (O_1021,N_19872,N_19455);
and UO_1022 (O_1022,N_19903,N_19493);
and UO_1023 (O_1023,N_19223,N_19744);
nand UO_1024 (O_1024,N_19526,N_19532);
and UO_1025 (O_1025,N_19344,N_19470);
nand UO_1026 (O_1026,N_19431,N_19901);
or UO_1027 (O_1027,N_19350,N_19410);
nor UO_1028 (O_1028,N_19925,N_19359);
nor UO_1029 (O_1029,N_19301,N_19329);
or UO_1030 (O_1030,N_19295,N_19987);
xor UO_1031 (O_1031,N_19990,N_19748);
or UO_1032 (O_1032,N_19275,N_19644);
nand UO_1033 (O_1033,N_19583,N_19800);
nor UO_1034 (O_1034,N_19953,N_19932);
or UO_1035 (O_1035,N_19929,N_19361);
or UO_1036 (O_1036,N_19681,N_19581);
or UO_1037 (O_1037,N_19340,N_19749);
and UO_1038 (O_1038,N_19646,N_19247);
or UO_1039 (O_1039,N_19759,N_19774);
or UO_1040 (O_1040,N_19547,N_19576);
xnor UO_1041 (O_1041,N_19621,N_19504);
nand UO_1042 (O_1042,N_19253,N_19615);
or UO_1043 (O_1043,N_19848,N_19536);
or UO_1044 (O_1044,N_19419,N_19388);
or UO_1045 (O_1045,N_19642,N_19282);
xnor UO_1046 (O_1046,N_19444,N_19566);
nand UO_1047 (O_1047,N_19631,N_19949);
or UO_1048 (O_1048,N_19938,N_19334);
nand UO_1049 (O_1049,N_19245,N_19575);
nor UO_1050 (O_1050,N_19899,N_19439);
or UO_1051 (O_1051,N_19526,N_19236);
nand UO_1052 (O_1052,N_19976,N_19364);
xor UO_1053 (O_1053,N_19774,N_19703);
or UO_1054 (O_1054,N_19989,N_19705);
xnor UO_1055 (O_1055,N_19304,N_19712);
xor UO_1056 (O_1056,N_19515,N_19318);
nand UO_1057 (O_1057,N_19786,N_19457);
or UO_1058 (O_1058,N_19337,N_19754);
xor UO_1059 (O_1059,N_19452,N_19827);
nor UO_1060 (O_1060,N_19253,N_19769);
or UO_1061 (O_1061,N_19446,N_19695);
and UO_1062 (O_1062,N_19674,N_19256);
or UO_1063 (O_1063,N_19412,N_19390);
and UO_1064 (O_1064,N_19436,N_19615);
and UO_1065 (O_1065,N_19951,N_19541);
or UO_1066 (O_1066,N_19419,N_19288);
xnor UO_1067 (O_1067,N_19945,N_19365);
nor UO_1068 (O_1068,N_19369,N_19758);
xor UO_1069 (O_1069,N_19806,N_19547);
nor UO_1070 (O_1070,N_19269,N_19894);
nor UO_1071 (O_1071,N_19597,N_19908);
or UO_1072 (O_1072,N_19247,N_19751);
nand UO_1073 (O_1073,N_19588,N_19403);
nand UO_1074 (O_1074,N_19286,N_19914);
nand UO_1075 (O_1075,N_19970,N_19680);
nand UO_1076 (O_1076,N_19525,N_19801);
nand UO_1077 (O_1077,N_19382,N_19808);
xor UO_1078 (O_1078,N_19355,N_19490);
nand UO_1079 (O_1079,N_19779,N_19272);
or UO_1080 (O_1080,N_19797,N_19843);
nor UO_1081 (O_1081,N_19954,N_19839);
or UO_1082 (O_1082,N_19820,N_19935);
nand UO_1083 (O_1083,N_19405,N_19612);
xor UO_1084 (O_1084,N_19949,N_19739);
xor UO_1085 (O_1085,N_19419,N_19222);
or UO_1086 (O_1086,N_19780,N_19266);
or UO_1087 (O_1087,N_19617,N_19450);
or UO_1088 (O_1088,N_19356,N_19349);
xnor UO_1089 (O_1089,N_19337,N_19476);
and UO_1090 (O_1090,N_19384,N_19959);
or UO_1091 (O_1091,N_19268,N_19270);
xor UO_1092 (O_1092,N_19988,N_19759);
nor UO_1093 (O_1093,N_19685,N_19370);
nand UO_1094 (O_1094,N_19576,N_19662);
or UO_1095 (O_1095,N_19212,N_19671);
nand UO_1096 (O_1096,N_19884,N_19279);
nand UO_1097 (O_1097,N_19880,N_19201);
or UO_1098 (O_1098,N_19219,N_19400);
xnor UO_1099 (O_1099,N_19505,N_19545);
nand UO_1100 (O_1100,N_19602,N_19871);
and UO_1101 (O_1101,N_19389,N_19516);
nor UO_1102 (O_1102,N_19341,N_19237);
and UO_1103 (O_1103,N_19691,N_19897);
nand UO_1104 (O_1104,N_19326,N_19502);
and UO_1105 (O_1105,N_19767,N_19530);
or UO_1106 (O_1106,N_19379,N_19862);
or UO_1107 (O_1107,N_19560,N_19729);
and UO_1108 (O_1108,N_19350,N_19673);
xor UO_1109 (O_1109,N_19568,N_19923);
nor UO_1110 (O_1110,N_19357,N_19309);
and UO_1111 (O_1111,N_19698,N_19609);
nor UO_1112 (O_1112,N_19310,N_19909);
or UO_1113 (O_1113,N_19659,N_19752);
or UO_1114 (O_1114,N_19321,N_19633);
nand UO_1115 (O_1115,N_19333,N_19808);
and UO_1116 (O_1116,N_19962,N_19510);
and UO_1117 (O_1117,N_19814,N_19971);
nor UO_1118 (O_1118,N_19563,N_19886);
and UO_1119 (O_1119,N_19472,N_19536);
and UO_1120 (O_1120,N_19992,N_19569);
or UO_1121 (O_1121,N_19552,N_19599);
or UO_1122 (O_1122,N_19929,N_19525);
nor UO_1123 (O_1123,N_19961,N_19540);
nand UO_1124 (O_1124,N_19521,N_19237);
or UO_1125 (O_1125,N_19542,N_19380);
nor UO_1126 (O_1126,N_19427,N_19725);
or UO_1127 (O_1127,N_19385,N_19541);
and UO_1128 (O_1128,N_19840,N_19785);
nand UO_1129 (O_1129,N_19464,N_19368);
and UO_1130 (O_1130,N_19388,N_19823);
or UO_1131 (O_1131,N_19274,N_19629);
xnor UO_1132 (O_1132,N_19568,N_19230);
xnor UO_1133 (O_1133,N_19951,N_19638);
nor UO_1134 (O_1134,N_19635,N_19378);
nor UO_1135 (O_1135,N_19518,N_19323);
nand UO_1136 (O_1136,N_19497,N_19535);
nand UO_1137 (O_1137,N_19863,N_19870);
or UO_1138 (O_1138,N_19775,N_19616);
xor UO_1139 (O_1139,N_19776,N_19450);
and UO_1140 (O_1140,N_19291,N_19534);
nand UO_1141 (O_1141,N_19369,N_19435);
xor UO_1142 (O_1142,N_19381,N_19708);
nand UO_1143 (O_1143,N_19300,N_19888);
xnor UO_1144 (O_1144,N_19823,N_19726);
nor UO_1145 (O_1145,N_19919,N_19467);
or UO_1146 (O_1146,N_19998,N_19791);
nand UO_1147 (O_1147,N_19261,N_19502);
nand UO_1148 (O_1148,N_19668,N_19956);
nor UO_1149 (O_1149,N_19503,N_19343);
xor UO_1150 (O_1150,N_19604,N_19788);
nor UO_1151 (O_1151,N_19432,N_19846);
or UO_1152 (O_1152,N_19503,N_19481);
xnor UO_1153 (O_1153,N_19872,N_19202);
and UO_1154 (O_1154,N_19884,N_19923);
nor UO_1155 (O_1155,N_19265,N_19895);
or UO_1156 (O_1156,N_19772,N_19577);
or UO_1157 (O_1157,N_19721,N_19403);
xor UO_1158 (O_1158,N_19331,N_19605);
and UO_1159 (O_1159,N_19223,N_19479);
and UO_1160 (O_1160,N_19762,N_19807);
nor UO_1161 (O_1161,N_19571,N_19624);
xnor UO_1162 (O_1162,N_19266,N_19209);
and UO_1163 (O_1163,N_19431,N_19917);
xor UO_1164 (O_1164,N_19777,N_19541);
and UO_1165 (O_1165,N_19756,N_19237);
and UO_1166 (O_1166,N_19225,N_19747);
or UO_1167 (O_1167,N_19242,N_19634);
or UO_1168 (O_1168,N_19395,N_19893);
and UO_1169 (O_1169,N_19930,N_19385);
nor UO_1170 (O_1170,N_19579,N_19923);
xor UO_1171 (O_1171,N_19331,N_19313);
nor UO_1172 (O_1172,N_19704,N_19826);
xor UO_1173 (O_1173,N_19725,N_19507);
nand UO_1174 (O_1174,N_19716,N_19659);
or UO_1175 (O_1175,N_19401,N_19772);
or UO_1176 (O_1176,N_19401,N_19779);
nand UO_1177 (O_1177,N_19499,N_19549);
and UO_1178 (O_1178,N_19279,N_19879);
nand UO_1179 (O_1179,N_19660,N_19894);
xnor UO_1180 (O_1180,N_19811,N_19392);
nand UO_1181 (O_1181,N_19265,N_19992);
nand UO_1182 (O_1182,N_19471,N_19433);
or UO_1183 (O_1183,N_19777,N_19262);
or UO_1184 (O_1184,N_19822,N_19221);
and UO_1185 (O_1185,N_19863,N_19593);
xor UO_1186 (O_1186,N_19544,N_19922);
or UO_1187 (O_1187,N_19470,N_19998);
nor UO_1188 (O_1188,N_19717,N_19647);
or UO_1189 (O_1189,N_19981,N_19660);
nand UO_1190 (O_1190,N_19563,N_19441);
nor UO_1191 (O_1191,N_19429,N_19896);
xnor UO_1192 (O_1192,N_19938,N_19459);
and UO_1193 (O_1193,N_19404,N_19870);
and UO_1194 (O_1194,N_19585,N_19295);
xor UO_1195 (O_1195,N_19306,N_19783);
or UO_1196 (O_1196,N_19669,N_19555);
or UO_1197 (O_1197,N_19325,N_19685);
nand UO_1198 (O_1198,N_19592,N_19295);
or UO_1199 (O_1199,N_19587,N_19263);
or UO_1200 (O_1200,N_19366,N_19573);
and UO_1201 (O_1201,N_19317,N_19650);
xnor UO_1202 (O_1202,N_19322,N_19469);
xor UO_1203 (O_1203,N_19345,N_19661);
or UO_1204 (O_1204,N_19983,N_19920);
xnor UO_1205 (O_1205,N_19404,N_19981);
xnor UO_1206 (O_1206,N_19562,N_19327);
or UO_1207 (O_1207,N_19910,N_19686);
or UO_1208 (O_1208,N_19349,N_19350);
xnor UO_1209 (O_1209,N_19794,N_19957);
nand UO_1210 (O_1210,N_19593,N_19321);
or UO_1211 (O_1211,N_19418,N_19671);
nand UO_1212 (O_1212,N_19460,N_19232);
xor UO_1213 (O_1213,N_19642,N_19917);
or UO_1214 (O_1214,N_19451,N_19752);
and UO_1215 (O_1215,N_19550,N_19925);
xor UO_1216 (O_1216,N_19237,N_19685);
or UO_1217 (O_1217,N_19223,N_19500);
xor UO_1218 (O_1218,N_19835,N_19779);
nand UO_1219 (O_1219,N_19356,N_19532);
xnor UO_1220 (O_1220,N_19868,N_19898);
nor UO_1221 (O_1221,N_19996,N_19405);
and UO_1222 (O_1222,N_19672,N_19559);
xnor UO_1223 (O_1223,N_19857,N_19722);
nor UO_1224 (O_1224,N_19915,N_19416);
xnor UO_1225 (O_1225,N_19741,N_19890);
nand UO_1226 (O_1226,N_19666,N_19656);
and UO_1227 (O_1227,N_19348,N_19607);
xor UO_1228 (O_1228,N_19395,N_19437);
or UO_1229 (O_1229,N_19509,N_19977);
and UO_1230 (O_1230,N_19991,N_19372);
xnor UO_1231 (O_1231,N_19230,N_19692);
nand UO_1232 (O_1232,N_19320,N_19560);
or UO_1233 (O_1233,N_19492,N_19785);
nand UO_1234 (O_1234,N_19573,N_19802);
nand UO_1235 (O_1235,N_19258,N_19511);
nand UO_1236 (O_1236,N_19449,N_19427);
and UO_1237 (O_1237,N_19362,N_19684);
and UO_1238 (O_1238,N_19733,N_19271);
and UO_1239 (O_1239,N_19602,N_19543);
or UO_1240 (O_1240,N_19745,N_19886);
nand UO_1241 (O_1241,N_19392,N_19414);
or UO_1242 (O_1242,N_19280,N_19778);
and UO_1243 (O_1243,N_19745,N_19275);
xnor UO_1244 (O_1244,N_19757,N_19299);
nand UO_1245 (O_1245,N_19898,N_19836);
nor UO_1246 (O_1246,N_19204,N_19585);
nand UO_1247 (O_1247,N_19351,N_19416);
or UO_1248 (O_1248,N_19753,N_19938);
nand UO_1249 (O_1249,N_19742,N_19981);
or UO_1250 (O_1250,N_19803,N_19426);
or UO_1251 (O_1251,N_19712,N_19636);
nor UO_1252 (O_1252,N_19213,N_19928);
nand UO_1253 (O_1253,N_19465,N_19733);
or UO_1254 (O_1254,N_19772,N_19780);
nand UO_1255 (O_1255,N_19287,N_19318);
xor UO_1256 (O_1256,N_19527,N_19676);
nor UO_1257 (O_1257,N_19787,N_19793);
or UO_1258 (O_1258,N_19414,N_19239);
and UO_1259 (O_1259,N_19349,N_19973);
nand UO_1260 (O_1260,N_19327,N_19844);
or UO_1261 (O_1261,N_19949,N_19955);
and UO_1262 (O_1262,N_19701,N_19691);
nor UO_1263 (O_1263,N_19851,N_19862);
nand UO_1264 (O_1264,N_19602,N_19621);
nand UO_1265 (O_1265,N_19539,N_19844);
nand UO_1266 (O_1266,N_19957,N_19511);
nor UO_1267 (O_1267,N_19216,N_19583);
nor UO_1268 (O_1268,N_19891,N_19451);
xnor UO_1269 (O_1269,N_19489,N_19673);
nand UO_1270 (O_1270,N_19965,N_19620);
or UO_1271 (O_1271,N_19663,N_19728);
or UO_1272 (O_1272,N_19580,N_19619);
and UO_1273 (O_1273,N_19502,N_19514);
nor UO_1274 (O_1274,N_19683,N_19555);
and UO_1275 (O_1275,N_19249,N_19326);
or UO_1276 (O_1276,N_19965,N_19702);
and UO_1277 (O_1277,N_19267,N_19650);
or UO_1278 (O_1278,N_19558,N_19830);
nand UO_1279 (O_1279,N_19930,N_19420);
or UO_1280 (O_1280,N_19976,N_19913);
and UO_1281 (O_1281,N_19211,N_19405);
xor UO_1282 (O_1282,N_19203,N_19923);
and UO_1283 (O_1283,N_19421,N_19707);
nand UO_1284 (O_1284,N_19250,N_19304);
nand UO_1285 (O_1285,N_19258,N_19491);
xor UO_1286 (O_1286,N_19376,N_19603);
and UO_1287 (O_1287,N_19494,N_19650);
and UO_1288 (O_1288,N_19809,N_19897);
and UO_1289 (O_1289,N_19794,N_19984);
nor UO_1290 (O_1290,N_19385,N_19556);
and UO_1291 (O_1291,N_19280,N_19709);
and UO_1292 (O_1292,N_19353,N_19233);
nand UO_1293 (O_1293,N_19820,N_19674);
or UO_1294 (O_1294,N_19893,N_19887);
nor UO_1295 (O_1295,N_19600,N_19858);
nor UO_1296 (O_1296,N_19768,N_19608);
and UO_1297 (O_1297,N_19411,N_19834);
and UO_1298 (O_1298,N_19982,N_19207);
or UO_1299 (O_1299,N_19760,N_19309);
nor UO_1300 (O_1300,N_19684,N_19926);
or UO_1301 (O_1301,N_19666,N_19240);
or UO_1302 (O_1302,N_19859,N_19724);
and UO_1303 (O_1303,N_19213,N_19797);
xor UO_1304 (O_1304,N_19972,N_19404);
or UO_1305 (O_1305,N_19926,N_19407);
and UO_1306 (O_1306,N_19643,N_19613);
nand UO_1307 (O_1307,N_19566,N_19707);
nand UO_1308 (O_1308,N_19220,N_19378);
and UO_1309 (O_1309,N_19646,N_19609);
and UO_1310 (O_1310,N_19733,N_19753);
nor UO_1311 (O_1311,N_19377,N_19801);
nand UO_1312 (O_1312,N_19743,N_19866);
xnor UO_1313 (O_1313,N_19758,N_19404);
xor UO_1314 (O_1314,N_19791,N_19508);
or UO_1315 (O_1315,N_19700,N_19320);
nand UO_1316 (O_1316,N_19604,N_19649);
nand UO_1317 (O_1317,N_19971,N_19895);
nand UO_1318 (O_1318,N_19275,N_19606);
nor UO_1319 (O_1319,N_19672,N_19565);
and UO_1320 (O_1320,N_19473,N_19820);
and UO_1321 (O_1321,N_19224,N_19483);
nor UO_1322 (O_1322,N_19228,N_19337);
or UO_1323 (O_1323,N_19654,N_19613);
xor UO_1324 (O_1324,N_19493,N_19948);
and UO_1325 (O_1325,N_19788,N_19950);
nor UO_1326 (O_1326,N_19978,N_19446);
xor UO_1327 (O_1327,N_19628,N_19941);
xnor UO_1328 (O_1328,N_19875,N_19957);
xnor UO_1329 (O_1329,N_19890,N_19412);
xnor UO_1330 (O_1330,N_19455,N_19957);
xor UO_1331 (O_1331,N_19394,N_19400);
nor UO_1332 (O_1332,N_19220,N_19766);
and UO_1333 (O_1333,N_19248,N_19924);
nor UO_1334 (O_1334,N_19917,N_19806);
nor UO_1335 (O_1335,N_19200,N_19647);
nor UO_1336 (O_1336,N_19998,N_19429);
or UO_1337 (O_1337,N_19400,N_19717);
xor UO_1338 (O_1338,N_19217,N_19726);
nor UO_1339 (O_1339,N_19782,N_19319);
and UO_1340 (O_1340,N_19250,N_19409);
nand UO_1341 (O_1341,N_19219,N_19208);
nand UO_1342 (O_1342,N_19685,N_19964);
nand UO_1343 (O_1343,N_19247,N_19889);
or UO_1344 (O_1344,N_19474,N_19609);
nor UO_1345 (O_1345,N_19530,N_19842);
or UO_1346 (O_1346,N_19770,N_19406);
and UO_1347 (O_1347,N_19807,N_19605);
and UO_1348 (O_1348,N_19244,N_19430);
and UO_1349 (O_1349,N_19278,N_19500);
and UO_1350 (O_1350,N_19523,N_19803);
nor UO_1351 (O_1351,N_19944,N_19680);
and UO_1352 (O_1352,N_19841,N_19579);
nand UO_1353 (O_1353,N_19819,N_19976);
and UO_1354 (O_1354,N_19262,N_19482);
or UO_1355 (O_1355,N_19695,N_19251);
nand UO_1356 (O_1356,N_19805,N_19422);
xnor UO_1357 (O_1357,N_19443,N_19563);
xnor UO_1358 (O_1358,N_19962,N_19473);
or UO_1359 (O_1359,N_19308,N_19253);
nor UO_1360 (O_1360,N_19477,N_19575);
xor UO_1361 (O_1361,N_19828,N_19987);
xnor UO_1362 (O_1362,N_19379,N_19335);
or UO_1363 (O_1363,N_19244,N_19257);
and UO_1364 (O_1364,N_19244,N_19808);
nand UO_1365 (O_1365,N_19736,N_19397);
and UO_1366 (O_1366,N_19917,N_19500);
or UO_1367 (O_1367,N_19665,N_19825);
or UO_1368 (O_1368,N_19446,N_19741);
and UO_1369 (O_1369,N_19438,N_19858);
xnor UO_1370 (O_1370,N_19947,N_19515);
xor UO_1371 (O_1371,N_19969,N_19359);
or UO_1372 (O_1372,N_19304,N_19687);
nor UO_1373 (O_1373,N_19974,N_19667);
xnor UO_1374 (O_1374,N_19649,N_19663);
nand UO_1375 (O_1375,N_19827,N_19482);
nor UO_1376 (O_1376,N_19342,N_19665);
and UO_1377 (O_1377,N_19355,N_19324);
or UO_1378 (O_1378,N_19744,N_19313);
nand UO_1379 (O_1379,N_19580,N_19926);
and UO_1380 (O_1380,N_19569,N_19582);
nand UO_1381 (O_1381,N_19964,N_19366);
nand UO_1382 (O_1382,N_19678,N_19788);
and UO_1383 (O_1383,N_19600,N_19387);
nand UO_1384 (O_1384,N_19217,N_19434);
nor UO_1385 (O_1385,N_19459,N_19892);
nand UO_1386 (O_1386,N_19401,N_19491);
xnor UO_1387 (O_1387,N_19897,N_19361);
nor UO_1388 (O_1388,N_19314,N_19339);
xor UO_1389 (O_1389,N_19256,N_19993);
nor UO_1390 (O_1390,N_19879,N_19623);
nor UO_1391 (O_1391,N_19705,N_19790);
nor UO_1392 (O_1392,N_19448,N_19277);
nand UO_1393 (O_1393,N_19208,N_19963);
or UO_1394 (O_1394,N_19517,N_19284);
or UO_1395 (O_1395,N_19295,N_19211);
xor UO_1396 (O_1396,N_19603,N_19910);
nand UO_1397 (O_1397,N_19887,N_19215);
nor UO_1398 (O_1398,N_19268,N_19865);
or UO_1399 (O_1399,N_19979,N_19718);
nand UO_1400 (O_1400,N_19728,N_19419);
xor UO_1401 (O_1401,N_19615,N_19865);
and UO_1402 (O_1402,N_19588,N_19527);
nand UO_1403 (O_1403,N_19501,N_19758);
nand UO_1404 (O_1404,N_19579,N_19992);
nor UO_1405 (O_1405,N_19537,N_19411);
nor UO_1406 (O_1406,N_19931,N_19799);
or UO_1407 (O_1407,N_19245,N_19281);
xnor UO_1408 (O_1408,N_19473,N_19388);
nor UO_1409 (O_1409,N_19314,N_19935);
or UO_1410 (O_1410,N_19869,N_19678);
nand UO_1411 (O_1411,N_19607,N_19664);
nand UO_1412 (O_1412,N_19946,N_19590);
nor UO_1413 (O_1413,N_19639,N_19368);
nor UO_1414 (O_1414,N_19320,N_19307);
xor UO_1415 (O_1415,N_19339,N_19656);
nor UO_1416 (O_1416,N_19988,N_19614);
or UO_1417 (O_1417,N_19690,N_19388);
and UO_1418 (O_1418,N_19853,N_19446);
nor UO_1419 (O_1419,N_19877,N_19795);
or UO_1420 (O_1420,N_19971,N_19369);
xor UO_1421 (O_1421,N_19549,N_19764);
nand UO_1422 (O_1422,N_19348,N_19230);
xor UO_1423 (O_1423,N_19783,N_19975);
xnor UO_1424 (O_1424,N_19831,N_19492);
nand UO_1425 (O_1425,N_19975,N_19902);
xor UO_1426 (O_1426,N_19800,N_19227);
xnor UO_1427 (O_1427,N_19343,N_19383);
or UO_1428 (O_1428,N_19621,N_19586);
nand UO_1429 (O_1429,N_19433,N_19402);
xor UO_1430 (O_1430,N_19829,N_19990);
nand UO_1431 (O_1431,N_19764,N_19208);
nand UO_1432 (O_1432,N_19462,N_19295);
xnor UO_1433 (O_1433,N_19439,N_19201);
nor UO_1434 (O_1434,N_19321,N_19318);
nand UO_1435 (O_1435,N_19976,N_19759);
nor UO_1436 (O_1436,N_19969,N_19921);
xnor UO_1437 (O_1437,N_19630,N_19566);
nor UO_1438 (O_1438,N_19697,N_19574);
xnor UO_1439 (O_1439,N_19265,N_19809);
and UO_1440 (O_1440,N_19908,N_19940);
or UO_1441 (O_1441,N_19555,N_19312);
and UO_1442 (O_1442,N_19808,N_19266);
nor UO_1443 (O_1443,N_19446,N_19713);
nand UO_1444 (O_1444,N_19257,N_19275);
and UO_1445 (O_1445,N_19725,N_19770);
nand UO_1446 (O_1446,N_19458,N_19497);
xnor UO_1447 (O_1447,N_19883,N_19693);
or UO_1448 (O_1448,N_19805,N_19309);
nand UO_1449 (O_1449,N_19497,N_19681);
and UO_1450 (O_1450,N_19491,N_19836);
and UO_1451 (O_1451,N_19672,N_19775);
or UO_1452 (O_1452,N_19281,N_19750);
nor UO_1453 (O_1453,N_19331,N_19821);
or UO_1454 (O_1454,N_19838,N_19697);
nand UO_1455 (O_1455,N_19963,N_19260);
or UO_1456 (O_1456,N_19224,N_19745);
and UO_1457 (O_1457,N_19537,N_19667);
nand UO_1458 (O_1458,N_19713,N_19244);
or UO_1459 (O_1459,N_19766,N_19964);
xor UO_1460 (O_1460,N_19331,N_19408);
or UO_1461 (O_1461,N_19992,N_19676);
nor UO_1462 (O_1462,N_19448,N_19800);
xnor UO_1463 (O_1463,N_19943,N_19984);
xnor UO_1464 (O_1464,N_19444,N_19760);
and UO_1465 (O_1465,N_19342,N_19707);
or UO_1466 (O_1466,N_19584,N_19853);
nor UO_1467 (O_1467,N_19440,N_19649);
nor UO_1468 (O_1468,N_19848,N_19447);
and UO_1469 (O_1469,N_19842,N_19205);
and UO_1470 (O_1470,N_19925,N_19445);
nor UO_1471 (O_1471,N_19606,N_19221);
xnor UO_1472 (O_1472,N_19570,N_19522);
nand UO_1473 (O_1473,N_19827,N_19862);
or UO_1474 (O_1474,N_19956,N_19855);
nor UO_1475 (O_1475,N_19222,N_19956);
and UO_1476 (O_1476,N_19478,N_19360);
nand UO_1477 (O_1477,N_19478,N_19598);
nand UO_1478 (O_1478,N_19855,N_19557);
and UO_1479 (O_1479,N_19203,N_19263);
nand UO_1480 (O_1480,N_19931,N_19451);
or UO_1481 (O_1481,N_19867,N_19497);
nand UO_1482 (O_1482,N_19893,N_19630);
and UO_1483 (O_1483,N_19285,N_19370);
xor UO_1484 (O_1484,N_19516,N_19270);
nor UO_1485 (O_1485,N_19464,N_19762);
nand UO_1486 (O_1486,N_19495,N_19848);
nand UO_1487 (O_1487,N_19551,N_19356);
or UO_1488 (O_1488,N_19644,N_19863);
nor UO_1489 (O_1489,N_19222,N_19414);
nand UO_1490 (O_1490,N_19455,N_19958);
and UO_1491 (O_1491,N_19273,N_19468);
nor UO_1492 (O_1492,N_19697,N_19459);
and UO_1493 (O_1493,N_19771,N_19402);
nor UO_1494 (O_1494,N_19726,N_19265);
nand UO_1495 (O_1495,N_19869,N_19248);
xor UO_1496 (O_1496,N_19683,N_19655);
nand UO_1497 (O_1497,N_19659,N_19800);
or UO_1498 (O_1498,N_19565,N_19358);
and UO_1499 (O_1499,N_19834,N_19397);
or UO_1500 (O_1500,N_19554,N_19767);
and UO_1501 (O_1501,N_19212,N_19563);
xor UO_1502 (O_1502,N_19724,N_19764);
or UO_1503 (O_1503,N_19625,N_19629);
or UO_1504 (O_1504,N_19556,N_19360);
xor UO_1505 (O_1505,N_19212,N_19809);
and UO_1506 (O_1506,N_19526,N_19949);
and UO_1507 (O_1507,N_19508,N_19476);
nand UO_1508 (O_1508,N_19993,N_19423);
or UO_1509 (O_1509,N_19286,N_19826);
and UO_1510 (O_1510,N_19606,N_19472);
nand UO_1511 (O_1511,N_19215,N_19761);
nor UO_1512 (O_1512,N_19521,N_19815);
or UO_1513 (O_1513,N_19382,N_19286);
nor UO_1514 (O_1514,N_19276,N_19684);
nor UO_1515 (O_1515,N_19921,N_19966);
nor UO_1516 (O_1516,N_19911,N_19550);
xnor UO_1517 (O_1517,N_19464,N_19291);
and UO_1518 (O_1518,N_19268,N_19512);
and UO_1519 (O_1519,N_19463,N_19698);
nor UO_1520 (O_1520,N_19212,N_19864);
nand UO_1521 (O_1521,N_19720,N_19518);
nand UO_1522 (O_1522,N_19542,N_19857);
nor UO_1523 (O_1523,N_19565,N_19267);
and UO_1524 (O_1524,N_19383,N_19267);
and UO_1525 (O_1525,N_19950,N_19388);
and UO_1526 (O_1526,N_19577,N_19827);
or UO_1527 (O_1527,N_19980,N_19506);
or UO_1528 (O_1528,N_19356,N_19869);
and UO_1529 (O_1529,N_19852,N_19773);
nand UO_1530 (O_1530,N_19771,N_19604);
nor UO_1531 (O_1531,N_19387,N_19594);
nor UO_1532 (O_1532,N_19555,N_19486);
nand UO_1533 (O_1533,N_19924,N_19414);
or UO_1534 (O_1534,N_19931,N_19325);
nand UO_1535 (O_1535,N_19841,N_19845);
xor UO_1536 (O_1536,N_19549,N_19953);
or UO_1537 (O_1537,N_19753,N_19697);
xor UO_1538 (O_1538,N_19282,N_19468);
nor UO_1539 (O_1539,N_19487,N_19245);
nor UO_1540 (O_1540,N_19536,N_19566);
nor UO_1541 (O_1541,N_19644,N_19756);
or UO_1542 (O_1542,N_19510,N_19283);
nand UO_1543 (O_1543,N_19665,N_19239);
and UO_1544 (O_1544,N_19353,N_19426);
nor UO_1545 (O_1545,N_19391,N_19720);
nand UO_1546 (O_1546,N_19762,N_19531);
xnor UO_1547 (O_1547,N_19437,N_19766);
nand UO_1548 (O_1548,N_19842,N_19657);
nor UO_1549 (O_1549,N_19706,N_19853);
nor UO_1550 (O_1550,N_19740,N_19482);
nor UO_1551 (O_1551,N_19483,N_19806);
xnor UO_1552 (O_1552,N_19605,N_19489);
or UO_1553 (O_1553,N_19787,N_19984);
nor UO_1554 (O_1554,N_19449,N_19794);
xor UO_1555 (O_1555,N_19525,N_19268);
nand UO_1556 (O_1556,N_19743,N_19900);
and UO_1557 (O_1557,N_19904,N_19780);
or UO_1558 (O_1558,N_19448,N_19357);
nor UO_1559 (O_1559,N_19376,N_19610);
or UO_1560 (O_1560,N_19854,N_19757);
or UO_1561 (O_1561,N_19571,N_19611);
or UO_1562 (O_1562,N_19632,N_19358);
xor UO_1563 (O_1563,N_19489,N_19338);
nor UO_1564 (O_1564,N_19405,N_19845);
nor UO_1565 (O_1565,N_19441,N_19620);
nand UO_1566 (O_1566,N_19260,N_19946);
xor UO_1567 (O_1567,N_19536,N_19526);
or UO_1568 (O_1568,N_19947,N_19677);
and UO_1569 (O_1569,N_19502,N_19384);
nand UO_1570 (O_1570,N_19507,N_19284);
or UO_1571 (O_1571,N_19740,N_19881);
nand UO_1572 (O_1572,N_19767,N_19504);
nand UO_1573 (O_1573,N_19204,N_19892);
xnor UO_1574 (O_1574,N_19910,N_19963);
or UO_1575 (O_1575,N_19588,N_19697);
and UO_1576 (O_1576,N_19410,N_19355);
nand UO_1577 (O_1577,N_19221,N_19230);
nand UO_1578 (O_1578,N_19880,N_19346);
nor UO_1579 (O_1579,N_19909,N_19370);
or UO_1580 (O_1580,N_19621,N_19975);
xor UO_1581 (O_1581,N_19209,N_19670);
nand UO_1582 (O_1582,N_19450,N_19602);
nor UO_1583 (O_1583,N_19935,N_19888);
and UO_1584 (O_1584,N_19822,N_19537);
or UO_1585 (O_1585,N_19782,N_19800);
or UO_1586 (O_1586,N_19488,N_19408);
nor UO_1587 (O_1587,N_19997,N_19623);
nand UO_1588 (O_1588,N_19867,N_19490);
nand UO_1589 (O_1589,N_19758,N_19308);
nand UO_1590 (O_1590,N_19213,N_19514);
nor UO_1591 (O_1591,N_19982,N_19522);
and UO_1592 (O_1592,N_19286,N_19769);
or UO_1593 (O_1593,N_19341,N_19847);
nor UO_1594 (O_1594,N_19987,N_19520);
or UO_1595 (O_1595,N_19253,N_19219);
nand UO_1596 (O_1596,N_19655,N_19685);
xor UO_1597 (O_1597,N_19923,N_19408);
nor UO_1598 (O_1598,N_19707,N_19733);
or UO_1599 (O_1599,N_19298,N_19872);
nand UO_1600 (O_1600,N_19213,N_19999);
nand UO_1601 (O_1601,N_19551,N_19542);
xor UO_1602 (O_1602,N_19564,N_19220);
xor UO_1603 (O_1603,N_19864,N_19511);
nand UO_1604 (O_1604,N_19906,N_19785);
nor UO_1605 (O_1605,N_19751,N_19828);
xnor UO_1606 (O_1606,N_19269,N_19866);
xor UO_1607 (O_1607,N_19260,N_19305);
and UO_1608 (O_1608,N_19352,N_19762);
nand UO_1609 (O_1609,N_19237,N_19858);
nor UO_1610 (O_1610,N_19907,N_19498);
nand UO_1611 (O_1611,N_19391,N_19234);
nand UO_1612 (O_1612,N_19325,N_19583);
and UO_1613 (O_1613,N_19397,N_19357);
nor UO_1614 (O_1614,N_19697,N_19777);
nor UO_1615 (O_1615,N_19897,N_19784);
nor UO_1616 (O_1616,N_19585,N_19315);
nand UO_1617 (O_1617,N_19719,N_19358);
nor UO_1618 (O_1618,N_19704,N_19856);
or UO_1619 (O_1619,N_19516,N_19256);
xor UO_1620 (O_1620,N_19552,N_19383);
nor UO_1621 (O_1621,N_19356,N_19387);
xnor UO_1622 (O_1622,N_19891,N_19476);
and UO_1623 (O_1623,N_19614,N_19246);
and UO_1624 (O_1624,N_19672,N_19673);
or UO_1625 (O_1625,N_19334,N_19467);
nand UO_1626 (O_1626,N_19213,N_19285);
and UO_1627 (O_1627,N_19666,N_19320);
or UO_1628 (O_1628,N_19827,N_19563);
xor UO_1629 (O_1629,N_19234,N_19825);
nand UO_1630 (O_1630,N_19676,N_19278);
and UO_1631 (O_1631,N_19419,N_19738);
xnor UO_1632 (O_1632,N_19230,N_19864);
and UO_1633 (O_1633,N_19961,N_19426);
and UO_1634 (O_1634,N_19563,N_19877);
and UO_1635 (O_1635,N_19504,N_19965);
or UO_1636 (O_1636,N_19277,N_19656);
and UO_1637 (O_1637,N_19984,N_19688);
nor UO_1638 (O_1638,N_19502,N_19821);
and UO_1639 (O_1639,N_19845,N_19895);
or UO_1640 (O_1640,N_19905,N_19348);
xnor UO_1641 (O_1641,N_19579,N_19928);
and UO_1642 (O_1642,N_19901,N_19272);
nor UO_1643 (O_1643,N_19486,N_19823);
and UO_1644 (O_1644,N_19322,N_19536);
nor UO_1645 (O_1645,N_19378,N_19795);
nor UO_1646 (O_1646,N_19819,N_19882);
nor UO_1647 (O_1647,N_19250,N_19654);
and UO_1648 (O_1648,N_19845,N_19710);
or UO_1649 (O_1649,N_19830,N_19223);
nand UO_1650 (O_1650,N_19220,N_19617);
nor UO_1651 (O_1651,N_19259,N_19455);
and UO_1652 (O_1652,N_19324,N_19953);
and UO_1653 (O_1653,N_19465,N_19224);
or UO_1654 (O_1654,N_19918,N_19235);
and UO_1655 (O_1655,N_19825,N_19556);
and UO_1656 (O_1656,N_19255,N_19262);
nand UO_1657 (O_1657,N_19251,N_19774);
xor UO_1658 (O_1658,N_19291,N_19773);
xor UO_1659 (O_1659,N_19290,N_19339);
and UO_1660 (O_1660,N_19610,N_19490);
nand UO_1661 (O_1661,N_19378,N_19248);
xnor UO_1662 (O_1662,N_19268,N_19342);
nor UO_1663 (O_1663,N_19509,N_19249);
nand UO_1664 (O_1664,N_19469,N_19373);
xor UO_1665 (O_1665,N_19622,N_19780);
nand UO_1666 (O_1666,N_19972,N_19919);
nand UO_1667 (O_1667,N_19988,N_19418);
or UO_1668 (O_1668,N_19384,N_19254);
or UO_1669 (O_1669,N_19938,N_19518);
xnor UO_1670 (O_1670,N_19854,N_19768);
nand UO_1671 (O_1671,N_19247,N_19551);
nor UO_1672 (O_1672,N_19896,N_19745);
nand UO_1673 (O_1673,N_19972,N_19362);
and UO_1674 (O_1674,N_19659,N_19409);
nor UO_1675 (O_1675,N_19789,N_19788);
nand UO_1676 (O_1676,N_19427,N_19916);
nor UO_1677 (O_1677,N_19964,N_19241);
nand UO_1678 (O_1678,N_19726,N_19770);
xnor UO_1679 (O_1679,N_19251,N_19341);
or UO_1680 (O_1680,N_19494,N_19636);
nor UO_1681 (O_1681,N_19630,N_19739);
and UO_1682 (O_1682,N_19417,N_19299);
or UO_1683 (O_1683,N_19616,N_19313);
nand UO_1684 (O_1684,N_19462,N_19348);
or UO_1685 (O_1685,N_19454,N_19809);
nand UO_1686 (O_1686,N_19367,N_19425);
nand UO_1687 (O_1687,N_19882,N_19674);
xor UO_1688 (O_1688,N_19723,N_19963);
and UO_1689 (O_1689,N_19547,N_19449);
or UO_1690 (O_1690,N_19864,N_19730);
nand UO_1691 (O_1691,N_19222,N_19578);
nand UO_1692 (O_1692,N_19541,N_19365);
or UO_1693 (O_1693,N_19290,N_19920);
xor UO_1694 (O_1694,N_19767,N_19233);
nand UO_1695 (O_1695,N_19389,N_19667);
and UO_1696 (O_1696,N_19291,N_19813);
or UO_1697 (O_1697,N_19912,N_19247);
and UO_1698 (O_1698,N_19644,N_19368);
and UO_1699 (O_1699,N_19413,N_19366);
and UO_1700 (O_1700,N_19393,N_19886);
xnor UO_1701 (O_1701,N_19930,N_19773);
nand UO_1702 (O_1702,N_19336,N_19902);
xor UO_1703 (O_1703,N_19203,N_19325);
or UO_1704 (O_1704,N_19859,N_19518);
or UO_1705 (O_1705,N_19273,N_19475);
nand UO_1706 (O_1706,N_19299,N_19737);
nand UO_1707 (O_1707,N_19891,N_19754);
and UO_1708 (O_1708,N_19564,N_19330);
or UO_1709 (O_1709,N_19754,N_19792);
xnor UO_1710 (O_1710,N_19600,N_19931);
nor UO_1711 (O_1711,N_19292,N_19421);
and UO_1712 (O_1712,N_19884,N_19806);
nor UO_1713 (O_1713,N_19384,N_19446);
nand UO_1714 (O_1714,N_19225,N_19495);
and UO_1715 (O_1715,N_19669,N_19738);
or UO_1716 (O_1716,N_19539,N_19578);
nor UO_1717 (O_1717,N_19724,N_19907);
and UO_1718 (O_1718,N_19265,N_19968);
or UO_1719 (O_1719,N_19684,N_19834);
xor UO_1720 (O_1720,N_19943,N_19441);
nand UO_1721 (O_1721,N_19638,N_19851);
nand UO_1722 (O_1722,N_19311,N_19795);
nor UO_1723 (O_1723,N_19548,N_19589);
nand UO_1724 (O_1724,N_19655,N_19472);
xnor UO_1725 (O_1725,N_19476,N_19925);
xnor UO_1726 (O_1726,N_19432,N_19929);
nor UO_1727 (O_1727,N_19965,N_19548);
and UO_1728 (O_1728,N_19971,N_19818);
and UO_1729 (O_1729,N_19474,N_19790);
nand UO_1730 (O_1730,N_19735,N_19587);
or UO_1731 (O_1731,N_19316,N_19283);
xor UO_1732 (O_1732,N_19747,N_19626);
nor UO_1733 (O_1733,N_19316,N_19899);
or UO_1734 (O_1734,N_19819,N_19469);
and UO_1735 (O_1735,N_19358,N_19797);
nand UO_1736 (O_1736,N_19502,N_19787);
or UO_1737 (O_1737,N_19865,N_19357);
and UO_1738 (O_1738,N_19915,N_19927);
xnor UO_1739 (O_1739,N_19444,N_19525);
xor UO_1740 (O_1740,N_19965,N_19474);
xor UO_1741 (O_1741,N_19897,N_19978);
and UO_1742 (O_1742,N_19947,N_19709);
nand UO_1743 (O_1743,N_19927,N_19867);
nor UO_1744 (O_1744,N_19755,N_19329);
and UO_1745 (O_1745,N_19969,N_19354);
nand UO_1746 (O_1746,N_19870,N_19230);
and UO_1747 (O_1747,N_19445,N_19704);
nand UO_1748 (O_1748,N_19263,N_19233);
xor UO_1749 (O_1749,N_19994,N_19665);
or UO_1750 (O_1750,N_19311,N_19949);
nor UO_1751 (O_1751,N_19229,N_19570);
and UO_1752 (O_1752,N_19460,N_19716);
xnor UO_1753 (O_1753,N_19373,N_19971);
nor UO_1754 (O_1754,N_19879,N_19351);
nor UO_1755 (O_1755,N_19866,N_19438);
or UO_1756 (O_1756,N_19587,N_19619);
and UO_1757 (O_1757,N_19772,N_19419);
xor UO_1758 (O_1758,N_19407,N_19704);
and UO_1759 (O_1759,N_19557,N_19884);
and UO_1760 (O_1760,N_19880,N_19981);
nor UO_1761 (O_1761,N_19692,N_19375);
xnor UO_1762 (O_1762,N_19936,N_19802);
nor UO_1763 (O_1763,N_19301,N_19328);
nor UO_1764 (O_1764,N_19548,N_19997);
xor UO_1765 (O_1765,N_19845,N_19218);
xor UO_1766 (O_1766,N_19680,N_19782);
and UO_1767 (O_1767,N_19687,N_19861);
and UO_1768 (O_1768,N_19569,N_19869);
or UO_1769 (O_1769,N_19425,N_19733);
nor UO_1770 (O_1770,N_19411,N_19602);
nand UO_1771 (O_1771,N_19508,N_19396);
or UO_1772 (O_1772,N_19758,N_19871);
and UO_1773 (O_1773,N_19302,N_19977);
xnor UO_1774 (O_1774,N_19661,N_19334);
nor UO_1775 (O_1775,N_19573,N_19562);
or UO_1776 (O_1776,N_19400,N_19586);
nor UO_1777 (O_1777,N_19674,N_19684);
nand UO_1778 (O_1778,N_19970,N_19289);
xnor UO_1779 (O_1779,N_19773,N_19469);
nand UO_1780 (O_1780,N_19885,N_19656);
xnor UO_1781 (O_1781,N_19682,N_19241);
xor UO_1782 (O_1782,N_19555,N_19630);
or UO_1783 (O_1783,N_19654,N_19811);
nor UO_1784 (O_1784,N_19889,N_19321);
nor UO_1785 (O_1785,N_19879,N_19413);
nand UO_1786 (O_1786,N_19692,N_19768);
nand UO_1787 (O_1787,N_19574,N_19639);
xor UO_1788 (O_1788,N_19373,N_19858);
nor UO_1789 (O_1789,N_19537,N_19285);
nand UO_1790 (O_1790,N_19504,N_19370);
nand UO_1791 (O_1791,N_19941,N_19622);
xor UO_1792 (O_1792,N_19790,N_19851);
xor UO_1793 (O_1793,N_19407,N_19481);
or UO_1794 (O_1794,N_19986,N_19459);
xnor UO_1795 (O_1795,N_19441,N_19456);
and UO_1796 (O_1796,N_19250,N_19251);
nor UO_1797 (O_1797,N_19921,N_19458);
nand UO_1798 (O_1798,N_19923,N_19685);
nor UO_1799 (O_1799,N_19247,N_19466);
xnor UO_1800 (O_1800,N_19687,N_19612);
and UO_1801 (O_1801,N_19352,N_19282);
nor UO_1802 (O_1802,N_19384,N_19260);
or UO_1803 (O_1803,N_19971,N_19419);
nand UO_1804 (O_1804,N_19648,N_19951);
nor UO_1805 (O_1805,N_19652,N_19826);
or UO_1806 (O_1806,N_19898,N_19583);
or UO_1807 (O_1807,N_19523,N_19331);
xor UO_1808 (O_1808,N_19444,N_19939);
and UO_1809 (O_1809,N_19236,N_19249);
or UO_1810 (O_1810,N_19522,N_19763);
and UO_1811 (O_1811,N_19959,N_19244);
nor UO_1812 (O_1812,N_19245,N_19698);
nor UO_1813 (O_1813,N_19896,N_19631);
nand UO_1814 (O_1814,N_19654,N_19565);
or UO_1815 (O_1815,N_19267,N_19213);
nand UO_1816 (O_1816,N_19975,N_19970);
nand UO_1817 (O_1817,N_19253,N_19563);
and UO_1818 (O_1818,N_19277,N_19722);
nand UO_1819 (O_1819,N_19570,N_19285);
nor UO_1820 (O_1820,N_19555,N_19984);
nor UO_1821 (O_1821,N_19952,N_19835);
and UO_1822 (O_1822,N_19986,N_19297);
nand UO_1823 (O_1823,N_19398,N_19459);
or UO_1824 (O_1824,N_19590,N_19480);
and UO_1825 (O_1825,N_19400,N_19802);
and UO_1826 (O_1826,N_19839,N_19847);
and UO_1827 (O_1827,N_19260,N_19572);
nand UO_1828 (O_1828,N_19933,N_19719);
or UO_1829 (O_1829,N_19306,N_19700);
nor UO_1830 (O_1830,N_19246,N_19652);
or UO_1831 (O_1831,N_19509,N_19687);
xnor UO_1832 (O_1832,N_19639,N_19895);
or UO_1833 (O_1833,N_19569,N_19393);
nand UO_1834 (O_1834,N_19368,N_19752);
and UO_1835 (O_1835,N_19514,N_19946);
and UO_1836 (O_1836,N_19614,N_19708);
nor UO_1837 (O_1837,N_19510,N_19294);
nand UO_1838 (O_1838,N_19409,N_19774);
xnor UO_1839 (O_1839,N_19778,N_19903);
nand UO_1840 (O_1840,N_19897,N_19655);
nor UO_1841 (O_1841,N_19383,N_19462);
or UO_1842 (O_1842,N_19819,N_19393);
nor UO_1843 (O_1843,N_19530,N_19329);
or UO_1844 (O_1844,N_19354,N_19875);
or UO_1845 (O_1845,N_19989,N_19340);
and UO_1846 (O_1846,N_19237,N_19522);
nand UO_1847 (O_1847,N_19253,N_19236);
xor UO_1848 (O_1848,N_19952,N_19652);
and UO_1849 (O_1849,N_19475,N_19666);
xor UO_1850 (O_1850,N_19610,N_19484);
and UO_1851 (O_1851,N_19385,N_19571);
nor UO_1852 (O_1852,N_19503,N_19474);
or UO_1853 (O_1853,N_19623,N_19474);
nand UO_1854 (O_1854,N_19727,N_19902);
xor UO_1855 (O_1855,N_19289,N_19273);
nor UO_1856 (O_1856,N_19345,N_19285);
nand UO_1857 (O_1857,N_19294,N_19715);
xor UO_1858 (O_1858,N_19353,N_19425);
nand UO_1859 (O_1859,N_19414,N_19796);
and UO_1860 (O_1860,N_19893,N_19762);
or UO_1861 (O_1861,N_19996,N_19690);
xnor UO_1862 (O_1862,N_19540,N_19271);
xnor UO_1863 (O_1863,N_19245,N_19530);
nand UO_1864 (O_1864,N_19516,N_19662);
or UO_1865 (O_1865,N_19364,N_19688);
nor UO_1866 (O_1866,N_19682,N_19899);
and UO_1867 (O_1867,N_19895,N_19490);
xnor UO_1868 (O_1868,N_19308,N_19616);
nor UO_1869 (O_1869,N_19441,N_19377);
nor UO_1870 (O_1870,N_19518,N_19654);
xor UO_1871 (O_1871,N_19271,N_19444);
nand UO_1872 (O_1872,N_19431,N_19914);
xnor UO_1873 (O_1873,N_19432,N_19376);
xor UO_1874 (O_1874,N_19687,N_19893);
nand UO_1875 (O_1875,N_19829,N_19405);
xor UO_1876 (O_1876,N_19864,N_19301);
nand UO_1877 (O_1877,N_19838,N_19232);
or UO_1878 (O_1878,N_19843,N_19514);
nor UO_1879 (O_1879,N_19739,N_19704);
or UO_1880 (O_1880,N_19517,N_19490);
or UO_1881 (O_1881,N_19488,N_19614);
and UO_1882 (O_1882,N_19540,N_19992);
nand UO_1883 (O_1883,N_19980,N_19485);
xnor UO_1884 (O_1884,N_19497,N_19728);
xnor UO_1885 (O_1885,N_19697,N_19740);
xor UO_1886 (O_1886,N_19289,N_19592);
nor UO_1887 (O_1887,N_19600,N_19489);
nand UO_1888 (O_1888,N_19442,N_19724);
nor UO_1889 (O_1889,N_19459,N_19489);
nand UO_1890 (O_1890,N_19902,N_19408);
xnor UO_1891 (O_1891,N_19387,N_19896);
or UO_1892 (O_1892,N_19418,N_19228);
or UO_1893 (O_1893,N_19584,N_19307);
and UO_1894 (O_1894,N_19295,N_19210);
nand UO_1895 (O_1895,N_19476,N_19498);
nand UO_1896 (O_1896,N_19334,N_19399);
nand UO_1897 (O_1897,N_19906,N_19485);
and UO_1898 (O_1898,N_19984,N_19382);
nand UO_1899 (O_1899,N_19756,N_19958);
or UO_1900 (O_1900,N_19998,N_19389);
and UO_1901 (O_1901,N_19665,N_19330);
nor UO_1902 (O_1902,N_19645,N_19478);
nor UO_1903 (O_1903,N_19564,N_19941);
or UO_1904 (O_1904,N_19551,N_19447);
or UO_1905 (O_1905,N_19424,N_19482);
and UO_1906 (O_1906,N_19254,N_19934);
xor UO_1907 (O_1907,N_19700,N_19218);
nor UO_1908 (O_1908,N_19906,N_19967);
nor UO_1909 (O_1909,N_19535,N_19399);
nor UO_1910 (O_1910,N_19962,N_19360);
or UO_1911 (O_1911,N_19816,N_19491);
nor UO_1912 (O_1912,N_19777,N_19362);
xor UO_1913 (O_1913,N_19518,N_19641);
nand UO_1914 (O_1914,N_19767,N_19744);
or UO_1915 (O_1915,N_19854,N_19861);
or UO_1916 (O_1916,N_19429,N_19498);
or UO_1917 (O_1917,N_19974,N_19715);
or UO_1918 (O_1918,N_19491,N_19885);
nand UO_1919 (O_1919,N_19354,N_19884);
and UO_1920 (O_1920,N_19683,N_19704);
xor UO_1921 (O_1921,N_19590,N_19288);
xor UO_1922 (O_1922,N_19523,N_19811);
or UO_1923 (O_1923,N_19668,N_19450);
nor UO_1924 (O_1924,N_19877,N_19833);
xnor UO_1925 (O_1925,N_19429,N_19796);
or UO_1926 (O_1926,N_19534,N_19621);
nand UO_1927 (O_1927,N_19900,N_19402);
nand UO_1928 (O_1928,N_19385,N_19917);
nand UO_1929 (O_1929,N_19584,N_19261);
nor UO_1930 (O_1930,N_19867,N_19658);
nor UO_1931 (O_1931,N_19303,N_19301);
or UO_1932 (O_1932,N_19464,N_19396);
or UO_1933 (O_1933,N_19541,N_19439);
or UO_1934 (O_1934,N_19257,N_19529);
nor UO_1935 (O_1935,N_19546,N_19584);
and UO_1936 (O_1936,N_19671,N_19981);
nand UO_1937 (O_1937,N_19373,N_19627);
or UO_1938 (O_1938,N_19719,N_19786);
and UO_1939 (O_1939,N_19293,N_19892);
or UO_1940 (O_1940,N_19426,N_19522);
nand UO_1941 (O_1941,N_19228,N_19641);
nand UO_1942 (O_1942,N_19481,N_19482);
nor UO_1943 (O_1943,N_19311,N_19875);
nand UO_1944 (O_1944,N_19647,N_19330);
nor UO_1945 (O_1945,N_19830,N_19903);
or UO_1946 (O_1946,N_19206,N_19550);
xnor UO_1947 (O_1947,N_19793,N_19525);
or UO_1948 (O_1948,N_19363,N_19504);
or UO_1949 (O_1949,N_19857,N_19452);
or UO_1950 (O_1950,N_19913,N_19934);
nand UO_1951 (O_1951,N_19943,N_19979);
nand UO_1952 (O_1952,N_19407,N_19284);
nor UO_1953 (O_1953,N_19783,N_19592);
nand UO_1954 (O_1954,N_19741,N_19319);
nor UO_1955 (O_1955,N_19863,N_19767);
or UO_1956 (O_1956,N_19990,N_19342);
nor UO_1957 (O_1957,N_19977,N_19797);
xnor UO_1958 (O_1958,N_19249,N_19648);
xnor UO_1959 (O_1959,N_19297,N_19557);
or UO_1960 (O_1960,N_19584,N_19854);
nor UO_1961 (O_1961,N_19245,N_19734);
nand UO_1962 (O_1962,N_19358,N_19583);
nor UO_1963 (O_1963,N_19613,N_19631);
nor UO_1964 (O_1964,N_19386,N_19583);
nand UO_1965 (O_1965,N_19335,N_19975);
and UO_1966 (O_1966,N_19364,N_19938);
or UO_1967 (O_1967,N_19324,N_19484);
xor UO_1968 (O_1968,N_19869,N_19645);
and UO_1969 (O_1969,N_19394,N_19613);
nor UO_1970 (O_1970,N_19665,N_19766);
and UO_1971 (O_1971,N_19217,N_19313);
nand UO_1972 (O_1972,N_19564,N_19804);
and UO_1973 (O_1973,N_19392,N_19831);
and UO_1974 (O_1974,N_19542,N_19735);
nor UO_1975 (O_1975,N_19767,N_19226);
and UO_1976 (O_1976,N_19314,N_19779);
xnor UO_1977 (O_1977,N_19947,N_19582);
nand UO_1978 (O_1978,N_19694,N_19740);
or UO_1979 (O_1979,N_19531,N_19859);
nor UO_1980 (O_1980,N_19505,N_19259);
nor UO_1981 (O_1981,N_19795,N_19960);
and UO_1982 (O_1982,N_19731,N_19650);
nor UO_1983 (O_1983,N_19512,N_19473);
and UO_1984 (O_1984,N_19608,N_19343);
or UO_1985 (O_1985,N_19300,N_19576);
nand UO_1986 (O_1986,N_19338,N_19862);
nor UO_1987 (O_1987,N_19597,N_19455);
xor UO_1988 (O_1988,N_19506,N_19513);
or UO_1989 (O_1989,N_19644,N_19591);
or UO_1990 (O_1990,N_19293,N_19903);
nor UO_1991 (O_1991,N_19218,N_19314);
nand UO_1992 (O_1992,N_19221,N_19406);
or UO_1993 (O_1993,N_19351,N_19741);
nand UO_1994 (O_1994,N_19684,N_19991);
and UO_1995 (O_1995,N_19782,N_19551);
nand UO_1996 (O_1996,N_19429,N_19616);
or UO_1997 (O_1997,N_19831,N_19916);
nand UO_1998 (O_1998,N_19923,N_19339);
nand UO_1999 (O_1999,N_19593,N_19661);
and UO_2000 (O_2000,N_19412,N_19256);
nand UO_2001 (O_2001,N_19244,N_19795);
nor UO_2002 (O_2002,N_19737,N_19440);
or UO_2003 (O_2003,N_19745,N_19858);
xnor UO_2004 (O_2004,N_19603,N_19353);
nor UO_2005 (O_2005,N_19410,N_19774);
nor UO_2006 (O_2006,N_19548,N_19495);
nor UO_2007 (O_2007,N_19455,N_19849);
xor UO_2008 (O_2008,N_19801,N_19269);
or UO_2009 (O_2009,N_19626,N_19715);
and UO_2010 (O_2010,N_19246,N_19979);
or UO_2011 (O_2011,N_19277,N_19525);
xnor UO_2012 (O_2012,N_19543,N_19850);
nor UO_2013 (O_2013,N_19294,N_19406);
nand UO_2014 (O_2014,N_19469,N_19308);
xnor UO_2015 (O_2015,N_19884,N_19398);
nor UO_2016 (O_2016,N_19393,N_19492);
and UO_2017 (O_2017,N_19750,N_19997);
nand UO_2018 (O_2018,N_19415,N_19803);
nor UO_2019 (O_2019,N_19927,N_19661);
nand UO_2020 (O_2020,N_19915,N_19578);
and UO_2021 (O_2021,N_19386,N_19508);
and UO_2022 (O_2022,N_19409,N_19987);
and UO_2023 (O_2023,N_19952,N_19749);
nand UO_2024 (O_2024,N_19850,N_19921);
or UO_2025 (O_2025,N_19936,N_19529);
and UO_2026 (O_2026,N_19313,N_19533);
nand UO_2027 (O_2027,N_19743,N_19871);
and UO_2028 (O_2028,N_19903,N_19444);
nand UO_2029 (O_2029,N_19732,N_19478);
nand UO_2030 (O_2030,N_19889,N_19997);
and UO_2031 (O_2031,N_19299,N_19864);
nor UO_2032 (O_2032,N_19823,N_19317);
or UO_2033 (O_2033,N_19225,N_19852);
or UO_2034 (O_2034,N_19718,N_19612);
nand UO_2035 (O_2035,N_19930,N_19332);
and UO_2036 (O_2036,N_19730,N_19663);
or UO_2037 (O_2037,N_19939,N_19524);
nor UO_2038 (O_2038,N_19807,N_19586);
nand UO_2039 (O_2039,N_19900,N_19921);
nand UO_2040 (O_2040,N_19501,N_19867);
and UO_2041 (O_2041,N_19289,N_19568);
or UO_2042 (O_2042,N_19742,N_19469);
and UO_2043 (O_2043,N_19917,N_19548);
nand UO_2044 (O_2044,N_19618,N_19872);
or UO_2045 (O_2045,N_19764,N_19745);
or UO_2046 (O_2046,N_19311,N_19856);
xor UO_2047 (O_2047,N_19885,N_19908);
or UO_2048 (O_2048,N_19676,N_19301);
nor UO_2049 (O_2049,N_19412,N_19720);
or UO_2050 (O_2050,N_19344,N_19375);
and UO_2051 (O_2051,N_19298,N_19276);
nand UO_2052 (O_2052,N_19652,N_19252);
nor UO_2053 (O_2053,N_19758,N_19288);
and UO_2054 (O_2054,N_19760,N_19534);
and UO_2055 (O_2055,N_19696,N_19344);
nand UO_2056 (O_2056,N_19264,N_19573);
and UO_2057 (O_2057,N_19370,N_19286);
nand UO_2058 (O_2058,N_19916,N_19970);
nand UO_2059 (O_2059,N_19252,N_19857);
nand UO_2060 (O_2060,N_19776,N_19426);
and UO_2061 (O_2061,N_19944,N_19208);
nand UO_2062 (O_2062,N_19301,N_19476);
nor UO_2063 (O_2063,N_19302,N_19346);
nand UO_2064 (O_2064,N_19891,N_19532);
nor UO_2065 (O_2065,N_19627,N_19230);
or UO_2066 (O_2066,N_19717,N_19579);
and UO_2067 (O_2067,N_19675,N_19853);
nand UO_2068 (O_2068,N_19348,N_19529);
or UO_2069 (O_2069,N_19649,N_19822);
nand UO_2070 (O_2070,N_19336,N_19317);
nand UO_2071 (O_2071,N_19585,N_19695);
nor UO_2072 (O_2072,N_19530,N_19671);
nor UO_2073 (O_2073,N_19321,N_19528);
nand UO_2074 (O_2074,N_19371,N_19511);
or UO_2075 (O_2075,N_19642,N_19323);
xor UO_2076 (O_2076,N_19722,N_19284);
and UO_2077 (O_2077,N_19689,N_19547);
or UO_2078 (O_2078,N_19733,N_19799);
or UO_2079 (O_2079,N_19904,N_19781);
and UO_2080 (O_2080,N_19855,N_19462);
nor UO_2081 (O_2081,N_19933,N_19391);
nor UO_2082 (O_2082,N_19965,N_19460);
nor UO_2083 (O_2083,N_19557,N_19747);
nor UO_2084 (O_2084,N_19323,N_19415);
xor UO_2085 (O_2085,N_19300,N_19740);
nor UO_2086 (O_2086,N_19457,N_19790);
or UO_2087 (O_2087,N_19242,N_19276);
nand UO_2088 (O_2088,N_19790,N_19967);
or UO_2089 (O_2089,N_19245,N_19857);
or UO_2090 (O_2090,N_19853,N_19225);
nor UO_2091 (O_2091,N_19835,N_19758);
or UO_2092 (O_2092,N_19545,N_19574);
or UO_2093 (O_2093,N_19583,N_19396);
or UO_2094 (O_2094,N_19505,N_19327);
and UO_2095 (O_2095,N_19542,N_19697);
xnor UO_2096 (O_2096,N_19274,N_19533);
nand UO_2097 (O_2097,N_19258,N_19496);
and UO_2098 (O_2098,N_19461,N_19408);
xnor UO_2099 (O_2099,N_19756,N_19546);
and UO_2100 (O_2100,N_19820,N_19940);
and UO_2101 (O_2101,N_19392,N_19424);
or UO_2102 (O_2102,N_19290,N_19865);
and UO_2103 (O_2103,N_19734,N_19384);
nor UO_2104 (O_2104,N_19427,N_19726);
nor UO_2105 (O_2105,N_19863,N_19807);
or UO_2106 (O_2106,N_19963,N_19900);
nand UO_2107 (O_2107,N_19566,N_19863);
or UO_2108 (O_2108,N_19538,N_19744);
xor UO_2109 (O_2109,N_19658,N_19779);
and UO_2110 (O_2110,N_19496,N_19279);
and UO_2111 (O_2111,N_19297,N_19448);
xor UO_2112 (O_2112,N_19650,N_19829);
or UO_2113 (O_2113,N_19408,N_19672);
and UO_2114 (O_2114,N_19550,N_19774);
xnor UO_2115 (O_2115,N_19340,N_19270);
xor UO_2116 (O_2116,N_19396,N_19604);
or UO_2117 (O_2117,N_19434,N_19801);
nand UO_2118 (O_2118,N_19892,N_19873);
nor UO_2119 (O_2119,N_19430,N_19301);
nor UO_2120 (O_2120,N_19957,N_19733);
nor UO_2121 (O_2121,N_19711,N_19749);
xor UO_2122 (O_2122,N_19628,N_19289);
nor UO_2123 (O_2123,N_19276,N_19993);
nor UO_2124 (O_2124,N_19458,N_19963);
nor UO_2125 (O_2125,N_19928,N_19451);
and UO_2126 (O_2126,N_19509,N_19472);
nand UO_2127 (O_2127,N_19457,N_19233);
or UO_2128 (O_2128,N_19946,N_19509);
and UO_2129 (O_2129,N_19493,N_19737);
nand UO_2130 (O_2130,N_19252,N_19911);
xor UO_2131 (O_2131,N_19789,N_19966);
nand UO_2132 (O_2132,N_19513,N_19643);
or UO_2133 (O_2133,N_19542,N_19703);
nand UO_2134 (O_2134,N_19730,N_19265);
and UO_2135 (O_2135,N_19864,N_19225);
xor UO_2136 (O_2136,N_19668,N_19822);
or UO_2137 (O_2137,N_19582,N_19333);
nor UO_2138 (O_2138,N_19348,N_19819);
nand UO_2139 (O_2139,N_19859,N_19662);
and UO_2140 (O_2140,N_19865,N_19526);
nand UO_2141 (O_2141,N_19553,N_19315);
nand UO_2142 (O_2142,N_19563,N_19477);
or UO_2143 (O_2143,N_19924,N_19242);
nand UO_2144 (O_2144,N_19791,N_19900);
nand UO_2145 (O_2145,N_19610,N_19347);
and UO_2146 (O_2146,N_19795,N_19932);
nor UO_2147 (O_2147,N_19984,N_19640);
xor UO_2148 (O_2148,N_19455,N_19932);
nor UO_2149 (O_2149,N_19903,N_19886);
nor UO_2150 (O_2150,N_19302,N_19361);
xor UO_2151 (O_2151,N_19931,N_19398);
xor UO_2152 (O_2152,N_19485,N_19810);
and UO_2153 (O_2153,N_19480,N_19420);
nor UO_2154 (O_2154,N_19932,N_19707);
or UO_2155 (O_2155,N_19292,N_19995);
xor UO_2156 (O_2156,N_19471,N_19813);
nand UO_2157 (O_2157,N_19408,N_19494);
nor UO_2158 (O_2158,N_19923,N_19839);
and UO_2159 (O_2159,N_19926,N_19757);
nand UO_2160 (O_2160,N_19567,N_19816);
and UO_2161 (O_2161,N_19681,N_19338);
xor UO_2162 (O_2162,N_19440,N_19641);
and UO_2163 (O_2163,N_19680,N_19574);
and UO_2164 (O_2164,N_19663,N_19612);
or UO_2165 (O_2165,N_19238,N_19965);
nand UO_2166 (O_2166,N_19637,N_19870);
or UO_2167 (O_2167,N_19676,N_19850);
xnor UO_2168 (O_2168,N_19289,N_19271);
nor UO_2169 (O_2169,N_19737,N_19984);
nor UO_2170 (O_2170,N_19383,N_19278);
nand UO_2171 (O_2171,N_19260,N_19247);
nand UO_2172 (O_2172,N_19349,N_19235);
and UO_2173 (O_2173,N_19932,N_19336);
or UO_2174 (O_2174,N_19473,N_19500);
and UO_2175 (O_2175,N_19506,N_19982);
and UO_2176 (O_2176,N_19285,N_19830);
nand UO_2177 (O_2177,N_19900,N_19510);
or UO_2178 (O_2178,N_19609,N_19588);
nand UO_2179 (O_2179,N_19456,N_19778);
and UO_2180 (O_2180,N_19438,N_19580);
xnor UO_2181 (O_2181,N_19591,N_19342);
or UO_2182 (O_2182,N_19594,N_19470);
xnor UO_2183 (O_2183,N_19753,N_19426);
or UO_2184 (O_2184,N_19467,N_19522);
nor UO_2185 (O_2185,N_19613,N_19717);
and UO_2186 (O_2186,N_19543,N_19899);
nor UO_2187 (O_2187,N_19896,N_19304);
nor UO_2188 (O_2188,N_19275,N_19676);
nand UO_2189 (O_2189,N_19506,N_19675);
or UO_2190 (O_2190,N_19869,N_19729);
and UO_2191 (O_2191,N_19617,N_19695);
and UO_2192 (O_2192,N_19661,N_19539);
and UO_2193 (O_2193,N_19315,N_19656);
nand UO_2194 (O_2194,N_19716,N_19612);
or UO_2195 (O_2195,N_19403,N_19846);
and UO_2196 (O_2196,N_19880,N_19202);
and UO_2197 (O_2197,N_19643,N_19367);
nor UO_2198 (O_2198,N_19300,N_19823);
or UO_2199 (O_2199,N_19350,N_19725);
and UO_2200 (O_2200,N_19393,N_19277);
nor UO_2201 (O_2201,N_19773,N_19954);
xnor UO_2202 (O_2202,N_19967,N_19891);
nand UO_2203 (O_2203,N_19303,N_19443);
and UO_2204 (O_2204,N_19418,N_19283);
or UO_2205 (O_2205,N_19404,N_19904);
nor UO_2206 (O_2206,N_19268,N_19984);
or UO_2207 (O_2207,N_19559,N_19373);
nand UO_2208 (O_2208,N_19731,N_19765);
xnor UO_2209 (O_2209,N_19284,N_19812);
or UO_2210 (O_2210,N_19495,N_19739);
or UO_2211 (O_2211,N_19466,N_19715);
or UO_2212 (O_2212,N_19911,N_19270);
and UO_2213 (O_2213,N_19258,N_19912);
or UO_2214 (O_2214,N_19957,N_19401);
and UO_2215 (O_2215,N_19927,N_19724);
nand UO_2216 (O_2216,N_19668,N_19528);
nand UO_2217 (O_2217,N_19630,N_19210);
xor UO_2218 (O_2218,N_19307,N_19975);
and UO_2219 (O_2219,N_19923,N_19398);
nor UO_2220 (O_2220,N_19259,N_19492);
nor UO_2221 (O_2221,N_19398,N_19475);
xnor UO_2222 (O_2222,N_19738,N_19926);
or UO_2223 (O_2223,N_19757,N_19400);
xnor UO_2224 (O_2224,N_19373,N_19309);
xor UO_2225 (O_2225,N_19414,N_19559);
or UO_2226 (O_2226,N_19800,N_19817);
and UO_2227 (O_2227,N_19247,N_19714);
nor UO_2228 (O_2228,N_19553,N_19486);
nor UO_2229 (O_2229,N_19957,N_19627);
nor UO_2230 (O_2230,N_19827,N_19301);
nor UO_2231 (O_2231,N_19660,N_19898);
or UO_2232 (O_2232,N_19345,N_19942);
nand UO_2233 (O_2233,N_19781,N_19975);
and UO_2234 (O_2234,N_19576,N_19478);
nand UO_2235 (O_2235,N_19630,N_19286);
nor UO_2236 (O_2236,N_19892,N_19398);
nand UO_2237 (O_2237,N_19582,N_19860);
nand UO_2238 (O_2238,N_19908,N_19279);
or UO_2239 (O_2239,N_19412,N_19554);
xnor UO_2240 (O_2240,N_19551,N_19749);
or UO_2241 (O_2241,N_19299,N_19639);
or UO_2242 (O_2242,N_19784,N_19683);
nand UO_2243 (O_2243,N_19432,N_19775);
nand UO_2244 (O_2244,N_19492,N_19250);
nand UO_2245 (O_2245,N_19598,N_19717);
or UO_2246 (O_2246,N_19295,N_19333);
xnor UO_2247 (O_2247,N_19362,N_19427);
nor UO_2248 (O_2248,N_19935,N_19725);
nand UO_2249 (O_2249,N_19828,N_19581);
and UO_2250 (O_2250,N_19453,N_19598);
or UO_2251 (O_2251,N_19920,N_19323);
or UO_2252 (O_2252,N_19847,N_19854);
xnor UO_2253 (O_2253,N_19649,N_19963);
and UO_2254 (O_2254,N_19395,N_19993);
nand UO_2255 (O_2255,N_19755,N_19736);
nand UO_2256 (O_2256,N_19467,N_19896);
nand UO_2257 (O_2257,N_19544,N_19440);
or UO_2258 (O_2258,N_19642,N_19488);
nor UO_2259 (O_2259,N_19319,N_19936);
or UO_2260 (O_2260,N_19989,N_19750);
or UO_2261 (O_2261,N_19323,N_19329);
or UO_2262 (O_2262,N_19558,N_19356);
xor UO_2263 (O_2263,N_19341,N_19657);
nor UO_2264 (O_2264,N_19909,N_19376);
nor UO_2265 (O_2265,N_19648,N_19354);
or UO_2266 (O_2266,N_19419,N_19761);
or UO_2267 (O_2267,N_19722,N_19520);
nand UO_2268 (O_2268,N_19541,N_19747);
nor UO_2269 (O_2269,N_19493,N_19845);
nor UO_2270 (O_2270,N_19787,N_19768);
nor UO_2271 (O_2271,N_19349,N_19473);
xnor UO_2272 (O_2272,N_19854,N_19652);
xor UO_2273 (O_2273,N_19449,N_19970);
nand UO_2274 (O_2274,N_19230,N_19562);
nand UO_2275 (O_2275,N_19470,N_19779);
nor UO_2276 (O_2276,N_19810,N_19689);
nor UO_2277 (O_2277,N_19897,N_19225);
nand UO_2278 (O_2278,N_19994,N_19869);
or UO_2279 (O_2279,N_19494,N_19248);
xnor UO_2280 (O_2280,N_19277,N_19960);
or UO_2281 (O_2281,N_19299,N_19495);
and UO_2282 (O_2282,N_19655,N_19387);
nor UO_2283 (O_2283,N_19380,N_19297);
xnor UO_2284 (O_2284,N_19700,N_19502);
nand UO_2285 (O_2285,N_19876,N_19820);
nor UO_2286 (O_2286,N_19924,N_19548);
and UO_2287 (O_2287,N_19859,N_19571);
nand UO_2288 (O_2288,N_19456,N_19368);
xnor UO_2289 (O_2289,N_19543,N_19311);
and UO_2290 (O_2290,N_19747,N_19837);
nand UO_2291 (O_2291,N_19748,N_19428);
and UO_2292 (O_2292,N_19948,N_19878);
nor UO_2293 (O_2293,N_19790,N_19787);
nor UO_2294 (O_2294,N_19901,N_19700);
or UO_2295 (O_2295,N_19418,N_19845);
nor UO_2296 (O_2296,N_19508,N_19682);
and UO_2297 (O_2297,N_19448,N_19644);
nor UO_2298 (O_2298,N_19911,N_19609);
nor UO_2299 (O_2299,N_19214,N_19344);
nand UO_2300 (O_2300,N_19290,N_19729);
xnor UO_2301 (O_2301,N_19568,N_19391);
xnor UO_2302 (O_2302,N_19577,N_19414);
nor UO_2303 (O_2303,N_19346,N_19895);
nor UO_2304 (O_2304,N_19651,N_19335);
nand UO_2305 (O_2305,N_19344,N_19578);
xnor UO_2306 (O_2306,N_19209,N_19583);
or UO_2307 (O_2307,N_19930,N_19275);
nand UO_2308 (O_2308,N_19990,N_19464);
nand UO_2309 (O_2309,N_19970,N_19529);
or UO_2310 (O_2310,N_19714,N_19472);
nor UO_2311 (O_2311,N_19202,N_19370);
or UO_2312 (O_2312,N_19381,N_19355);
nor UO_2313 (O_2313,N_19487,N_19214);
and UO_2314 (O_2314,N_19750,N_19732);
nor UO_2315 (O_2315,N_19927,N_19900);
and UO_2316 (O_2316,N_19526,N_19591);
nand UO_2317 (O_2317,N_19333,N_19807);
or UO_2318 (O_2318,N_19215,N_19822);
or UO_2319 (O_2319,N_19934,N_19917);
or UO_2320 (O_2320,N_19736,N_19413);
nand UO_2321 (O_2321,N_19390,N_19525);
xor UO_2322 (O_2322,N_19271,N_19646);
or UO_2323 (O_2323,N_19464,N_19416);
and UO_2324 (O_2324,N_19661,N_19229);
and UO_2325 (O_2325,N_19614,N_19865);
and UO_2326 (O_2326,N_19247,N_19707);
and UO_2327 (O_2327,N_19821,N_19612);
nor UO_2328 (O_2328,N_19902,N_19302);
and UO_2329 (O_2329,N_19957,N_19302);
and UO_2330 (O_2330,N_19902,N_19262);
nor UO_2331 (O_2331,N_19543,N_19418);
xnor UO_2332 (O_2332,N_19788,N_19571);
nor UO_2333 (O_2333,N_19931,N_19476);
nor UO_2334 (O_2334,N_19805,N_19641);
nor UO_2335 (O_2335,N_19475,N_19817);
nand UO_2336 (O_2336,N_19434,N_19699);
nand UO_2337 (O_2337,N_19551,N_19524);
or UO_2338 (O_2338,N_19230,N_19468);
nor UO_2339 (O_2339,N_19238,N_19349);
or UO_2340 (O_2340,N_19946,N_19644);
and UO_2341 (O_2341,N_19729,N_19279);
and UO_2342 (O_2342,N_19342,N_19698);
or UO_2343 (O_2343,N_19219,N_19944);
nand UO_2344 (O_2344,N_19507,N_19990);
nand UO_2345 (O_2345,N_19951,N_19470);
and UO_2346 (O_2346,N_19523,N_19233);
nand UO_2347 (O_2347,N_19936,N_19557);
nand UO_2348 (O_2348,N_19303,N_19374);
nand UO_2349 (O_2349,N_19824,N_19775);
xor UO_2350 (O_2350,N_19794,N_19404);
nor UO_2351 (O_2351,N_19715,N_19892);
xnor UO_2352 (O_2352,N_19904,N_19443);
or UO_2353 (O_2353,N_19710,N_19653);
or UO_2354 (O_2354,N_19502,N_19720);
xor UO_2355 (O_2355,N_19416,N_19465);
nor UO_2356 (O_2356,N_19355,N_19942);
and UO_2357 (O_2357,N_19426,N_19997);
or UO_2358 (O_2358,N_19969,N_19890);
nand UO_2359 (O_2359,N_19640,N_19487);
nor UO_2360 (O_2360,N_19415,N_19841);
or UO_2361 (O_2361,N_19552,N_19852);
nor UO_2362 (O_2362,N_19558,N_19740);
nand UO_2363 (O_2363,N_19798,N_19780);
nand UO_2364 (O_2364,N_19905,N_19834);
xnor UO_2365 (O_2365,N_19678,N_19431);
and UO_2366 (O_2366,N_19554,N_19413);
or UO_2367 (O_2367,N_19301,N_19808);
nor UO_2368 (O_2368,N_19245,N_19681);
xor UO_2369 (O_2369,N_19395,N_19947);
nor UO_2370 (O_2370,N_19567,N_19450);
nor UO_2371 (O_2371,N_19537,N_19440);
nand UO_2372 (O_2372,N_19788,N_19944);
nor UO_2373 (O_2373,N_19709,N_19434);
nor UO_2374 (O_2374,N_19243,N_19849);
or UO_2375 (O_2375,N_19968,N_19330);
and UO_2376 (O_2376,N_19594,N_19851);
nand UO_2377 (O_2377,N_19453,N_19482);
and UO_2378 (O_2378,N_19850,N_19421);
xor UO_2379 (O_2379,N_19815,N_19905);
nand UO_2380 (O_2380,N_19744,N_19609);
or UO_2381 (O_2381,N_19381,N_19296);
nor UO_2382 (O_2382,N_19926,N_19899);
or UO_2383 (O_2383,N_19838,N_19875);
nor UO_2384 (O_2384,N_19883,N_19673);
xor UO_2385 (O_2385,N_19292,N_19335);
or UO_2386 (O_2386,N_19757,N_19632);
and UO_2387 (O_2387,N_19755,N_19307);
nor UO_2388 (O_2388,N_19762,N_19871);
nand UO_2389 (O_2389,N_19923,N_19467);
or UO_2390 (O_2390,N_19587,N_19526);
nand UO_2391 (O_2391,N_19932,N_19803);
or UO_2392 (O_2392,N_19474,N_19894);
and UO_2393 (O_2393,N_19901,N_19323);
xnor UO_2394 (O_2394,N_19977,N_19316);
or UO_2395 (O_2395,N_19630,N_19387);
nand UO_2396 (O_2396,N_19688,N_19643);
or UO_2397 (O_2397,N_19671,N_19486);
nor UO_2398 (O_2398,N_19684,N_19953);
xnor UO_2399 (O_2399,N_19779,N_19369);
and UO_2400 (O_2400,N_19832,N_19363);
or UO_2401 (O_2401,N_19340,N_19854);
or UO_2402 (O_2402,N_19482,N_19794);
xor UO_2403 (O_2403,N_19361,N_19828);
and UO_2404 (O_2404,N_19272,N_19963);
nand UO_2405 (O_2405,N_19459,N_19297);
and UO_2406 (O_2406,N_19262,N_19565);
and UO_2407 (O_2407,N_19212,N_19787);
nand UO_2408 (O_2408,N_19357,N_19374);
and UO_2409 (O_2409,N_19414,N_19257);
xor UO_2410 (O_2410,N_19596,N_19711);
or UO_2411 (O_2411,N_19993,N_19200);
nor UO_2412 (O_2412,N_19409,N_19869);
xnor UO_2413 (O_2413,N_19518,N_19934);
or UO_2414 (O_2414,N_19472,N_19748);
nand UO_2415 (O_2415,N_19598,N_19232);
nor UO_2416 (O_2416,N_19858,N_19851);
or UO_2417 (O_2417,N_19953,N_19433);
or UO_2418 (O_2418,N_19763,N_19455);
and UO_2419 (O_2419,N_19347,N_19504);
nand UO_2420 (O_2420,N_19234,N_19287);
nor UO_2421 (O_2421,N_19997,N_19867);
nand UO_2422 (O_2422,N_19331,N_19532);
nor UO_2423 (O_2423,N_19291,N_19541);
and UO_2424 (O_2424,N_19830,N_19380);
nor UO_2425 (O_2425,N_19569,N_19530);
nand UO_2426 (O_2426,N_19594,N_19563);
nor UO_2427 (O_2427,N_19275,N_19329);
nand UO_2428 (O_2428,N_19984,N_19247);
and UO_2429 (O_2429,N_19937,N_19693);
nand UO_2430 (O_2430,N_19779,N_19663);
nand UO_2431 (O_2431,N_19250,N_19383);
and UO_2432 (O_2432,N_19416,N_19943);
nor UO_2433 (O_2433,N_19877,N_19401);
and UO_2434 (O_2434,N_19543,N_19767);
xor UO_2435 (O_2435,N_19529,N_19469);
nor UO_2436 (O_2436,N_19689,N_19694);
nor UO_2437 (O_2437,N_19350,N_19656);
xor UO_2438 (O_2438,N_19984,N_19448);
xor UO_2439 (O_2439,N_19345,N_19507);
or UO_2440 (O_2440,N_19997,N_19492);
xor UO_2441 (O_2441,N_19642,N_19720);
xnor UO_2442 (O_2442,N_19922,N_19582);
and UO_2443 (O_2443,N_19614,N_19409);
and UO_2444 (O_2444,N_19713,N_19747);
nor UO_2445 (O_2445,N_19269,N_19962);
or UO_2446 (O_2446,N_19739,N_19767);
or UO_2447 (O_2447,N_19719,N_19682);
or UO_2448 (O_2448,N_19350,N_19880);
nor UO_2449 (O_2449,N_19421,N_19798);
nor UO_2450 (O_2450,N_19560,N_19342);
nor UO_2451 (O_2451,N_19434,N_19799);
nor UO_2452 (O_2452,N_19303,N_19988);
or UO_2453 (O_2453,N_19909,N_19778);
or UO_2454 (O_2454,N_19719,N_19940);
nand UO_2455 (O_2455,N_19292,N_19337);
and UO_2456 (O_2456,N_19386,N_19944);
nand UO_2457 (O_2457,N_19965,N_19994);
nand UO_2458 (O_2458,N_19504,N_19724);
xnor UO_2459 (O_2459,N_19735,N_19630);
xor UO_2460 (O_2460,N_19239,N_19623);
xor UO_2461 (O_2461,N_19518,N_19834);
or UO_2462 (O_2462,N_19383,N_19452);
and UO_2463 (O_2463,N_19458,N_19804);
or UO_2464 (O_2464,N_19675,N_19283);
or UO_2465 (O_2465,N_19955,N_19238);
nand UO_2466 (O_2466,N_19574,N_19381);
and UO_2467 (O_2467,N_19906,N_19662);
and UO_2468 (O_2468,N_19502,N_19611);
and UO_2469 (O_2469,N_19456,N_19886);
and UO_2470 (O_2470,N_19324,N_19360);
nor UO_2471 (O_2471,N_19280,N_19394);
nor UO_2472 (O_2472,N_19517,N_19773);
and UO_2473 (O_2473,N_19500,N_19924);
nor UO_2474 (O_2474,N_19471,N_19388);
xor UO_2475 (O_2475,N_19822,N_19707);
xnor UO_2476 (O_2476,N_19423,N_19207);
and UO_2477 (O_2477,N_19934,N_19394);
nor UO_2478 (O_2478,N_19634,N_19928);
and UO_2479 (O_2479,N_19672,N_19298);
nor UO_2480 (O_2480,N_19637,N_19293);
and UO_2481 (O_2481,N_19285,N_19472);
xnor UO_2482 (O_2482,N_19648,N_19399);
or UO_2483 (O_2483,N_19316,N_19833);
nand UO_2484 (O_2484,N_19924,N_19914);
nand UO_2485 (O_2485,N_19994,N_19318);
nand UO_2486 (O_2486,N_19992,N_19631);
nor UO_2487 (O_2487,N_19639,N_19793);
and UO_2488 (O_2488,N_19872,N_19720);
or UO_2489 (O_2489,N_19538,N_19816);
or UO_2490 (O_2490,N_19587,N_19430);
or UO_2491 (O_2491,N_19325,N_19747);
or UO_2492 (O_2492,N_19395,N_19797);
nand UO_2493 (O_2493,N_19900,N_19749);
nor UO_2494 (O_2494,N_19614,N_19454);
nor UO_2495 (O_2495,N_19263,N_19540);
nor UO_2496 (O_2496,N_19217,N_19510);
nor UO_2497 (O_2497,N_19902,N_19395);
or UO_2498 (O_2498,N_19760,N_19903);
or UO_2499 (O_2499,N_19984,N_19507);
endmodule